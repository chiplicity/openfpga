magic
tech sky130A
magscale 1 2
timestamp 1605004037
<< locali >>
rect 949 15963 983 16609
rect 949 13175 983 15929
rect 3065 15351 3099 15453
rect 20453 14807 20487 14909
rect 949 12835 983 13141
rect 949 10999 983 12801
rect 17417 12699 17451 12937
rect 1501 11611 1535 11849
rect 12081 11543 12115 11781
<< viali >>
rect 1593 23817 1627 23851
rect 22661 23817 22695 23851
rect 24777 23817 24811 23851
rect 1409 23613 1443 23647
rect 1961 23613 1995 23647
rect 22477 23613 22511 23647
rect 23029 23613 23063 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 1593 23273 1627 23307
rect 19809 23205 19843 23239
rect 1409 23137 1443 23171
rect 19533 23137 19567 23171
rect 1869 22593 1903 22627
rect 1685 22525 1719 22559
rect 2513 22389 2547 22423
rect 19533 22389 19567 22423
rect 1409 22049 1443 22083
rect 1593 21913 1627 21947
rect 2053 21845 2087 21879
rect 1593 21641 1627 21675
rect 24777 21641 24811 21675
rect 1409 21437 1443 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 2053 21301 2087 21335
rect 2421 21301 2455 21335
rect 1593 21097 1627 21131
rect 4629 21097 4663 21131
rect 23949 21029 23983 21063
rect 1409 20961 1443 20995
rect 4445 20961 4479 20995
rect 23673 20961 23707 20995
rect 1593 20553 1627 20587
rect 24777 20553 24811 20587
rect 4537 20417 4571 20451
rect 5365 20417 5399 20451
rect 1409 20349 1443 20383
rect 2053 20349 2087 20383
rect 5181 20349 5215 20383
rect 24593 20349 24627 20383
rect 25145 20349 25179 20383
rect 2421 20213 2455 20247
rect 6009 20213 6043 20247
rect 23857 20213 23891 20247
rect 1593 20009 1627 20043
rect 2697 20009 2731 20043
rect 24777 20009 24811 20043
rect 1409 19873 1443 19907
rect 2513 19873 2547 19907
rect 24593 19873 24627 19907
rect 23581 19805 23615 19839
rect 1961 19669 1995 19703
rect 1409 19261 1443 19295
rect 2513 19261 2547 19295
rect 3065 19261 3099 19295
rect 18153 19261 18187 19295
rect 18705 19261 18739 19295
rect 24593 19261 24627 19295
rect 25145 19261 25179 19295
rect 1593 19125 1627 19159
rect 2053 19125 2087 19159
rect 2421 19125 2455 19159
rect 2697 19125 2731 19159
rect 18337 19125 18371 19159
rect 22569 19125 22603 19159
rect 24409 19125 24443 19159
rect 24777 19125 24811 19159
rect 4261 18921 4295 18955
rect 24777 18921 24811 18955
rect 17417 18853 17451 18887
rect 1501 18785 1535 18819
rect 2789 18785 2823 18819
rect 4077 18785 4111 18819
rect 17141 18785 17175 18819
rect 22385 18785 22419 18819
rect 23489 18785 23523 18819
rect 24593 18785 24627 18819
rect 1777 18717 1811 18751
rect 22569 18649 22603 18683
rect 2605 18581 2639 18615
rect 2973 18581 3007 18615
rect 23673 18581 23707 18615
rect 24869 18377 24903 18411
rect 1685 18241 1719 18275
rect 2881 18241 2915 18275
rect 3985 18241 4019 18275
rect 4445 18241 4479 18275
rect 1409 18173 1443 18207
rect 3709 18173 3743 18207
rect 21373 18173 21407 18207
rect 21925 18173 21959 18207
rect 22293 18173 22327 18207
rect 22477 18173 22511 18207
rect 24317 18173 24351 18207
rect 25421 18173 25455 18207
rect 2513 18105 2547 18139
rect 23121 18105 23155 18139
rect 2145 18037 2179 18071
rect 3617 18037 3651 18071
rect 17141 18037 17175 18071
rect 19625 18037 19659 18071
rect 21557 18037 21591 18071
rect 22661 18037 22695 18071
rect 23489 18037 23523 18071
rect 24133 18037 24167 18071
rect 24501 18037 24535 18071
rect 25605 18037 25639 18071
rect 26065 18037 26099 18071
rect 5365 17833 5399 17867
rect 24777 17833 24811 17867
rect 1961 17765 1995 17799
rect 1869 17697 1903 17731
rect 4077 17697 4111 17731
rect 5181 17697 5215 17731
rect 19625 17697 19659 17731
rect 21281 17697 21315 17731
rect 22385 17697 22419 17731
rect 23489 17697 23523 17731
rect 24593 17697 24627 17731
rect 2145 17629 2179 17663
rect 17417 17629 17451 17663
rect 19717 17629 19751 17663
rect 19901 17629 19935 17663
rect 4629 17561 4663 17595
rect 21465 17561 21499 17595
rect 22569 17561 22603 17595
rect 1501 17493 1535 17527
rect 2513 17493 2547 17527
rect 2973 17493 3007 17527
rect 3341 17493 3375 17527
rect 3709 17493 3743 17527
rect 4261 17493 4295 17527
rect 19073 17493 19107 17527
rect 19257 17493 19291 17527
rect 20361 17493 20395 17527
rect 20637 17493 20671 17527
rect 21925 17493 21959 17527
rect 23673 17493 23707 17527
rect 2789 17289 2823 17323
rect 3985 17289 4019 17323
rect 16037 17289 16071 17323
rect 18797 17289 18831 17323
rect 21281 17289 21315 17323
rect 24777 17289 24811 17323
rect 19717 17221 19751 17255
rect 2053 17153 2087 17187
rect 3525 17153 3559 17187
rect 20453 17153 20487 17187
rect 21925 17153 21959 17187
rect 22017 17153 22051 17187
rect 1777 17085 1811 17119
rect 4537 17085 4571 17119
rect 4813 17085 4847 17119
rect 15853 17085 15887 17119
rect 16405 17085 16439 17119
rect 19349 17085 19383 17119
rect 20269 17085 20303 17119
rect 24593 17085 24627 17119
rect 3433 17017 3467 17051
rect 24409 17017 24443 17051
rect 1409 16949 1443 16983
rect 1869 16949 1903 16983
rect 2513 16949 2547 16983
rect 2973 16949 3007 16983
rect 3341 16949 3375 16983
rect 4353 16949 4387 16983
rect 5273 16949 5307 16983
rect 16957 16949 16991 16983
rect 18889 16949 18923 16983
rect 19901 16949 19935 16983
rect 20361 16949 20395 16983
rect 20913 16949 20947 16983
rect 21465 16949 21499 16983
rect 21833 16949 21867 16983
rect 22569 16949 22603 16983
rect 23857 16949 23891 16983
rect 25145 16949 25179 16983
rect 2605 16745 2639 16779
rect 3249 16745 3283 16779
rect 5549 16745 5583 16779
rect 6929 16745 6963 16779
rect 7941 16745 7975 16779
rect 17417 16745 17451 16779
rect 18613 16745 18647 16779
rect 19257 16745 19291 16779
rect 20913 16745 20947 16779
rect 21925 16745 21959 16779
rect 22477 16745 22511 16779
rect 23765 16745 23799 16779
rect 25513 16745 25547 16779
rect 6469 16677 6503 16711
rect 7389 16677 7423 16711
rect 16282 16677 16316 16711
rect 22293 16677 22327 16711
rect 24317 16677 24351 16711
rect 949 16609 983 16643
rect 1869 16609 1903 16643
rect 1961 16609 1995 16643
rect 3617 16609 3651 16643
rect 4077 16609 4111 16643
rect 4353 16609 4387 16643
rect 5365 16609 5399 16643
rect 6837 16609 6871 16643
rect 7297 16609 7331 16643
rect 13277 16609 13311 16643
rect 19625 16609 19659 16643
rect 20361 16609 20395 16643
rect 21281 16609 21315 16643
rect 21373 16609 21407 16643
rect 22845 16609 22879 16643
rect 24041 16609 24075 16643
rect 24777 16609 24811 16643
rect 25329 16609 25363 16643
rect 2053 16541 2087 16575
rect 2881 16541 2915 16575
rect 7573 16541 7607 16575
rect 16037 16541 16071 16575
rect 19717 16541 19751 16575
rect 19901 16541 19935 16575
rect 21465 16541 21499 16575
rect 22937 16541 22971 16575
rect 23029 16541 23063 16575
rect 4813 16473 4847 16507
rect 1501 16405 1535 16439
rect 5181 16405 5215 16439
rect 5917 16405 5951 16439
rect 18245 16405 18279 16439
rect 19165 16405 19199 16439
rect 20637 16405 20671 16439
rect 2421 16201 2455 16235
rect 5365 16201 5399 16235
rect 5825 16201 5859 16235
rect 7113 16201 7147 16235
rect 9045 16201 9079 16235
rect 16129 16201 16163 16235
rect 22385 16201 22419 16235
rect 22661 16201 22695 16235
rect 23673 16201 23707 16235
rect 25421 16201 25455 16235
rect 1409 16133 1443 16167
rect 1961 16065 1995 16099
rect 7665 16065 7699 16099
rect 13737 16065 13771 16099
rect 15209 16065 15243 16099
rect 18797 16065 18831 16099
rect 19717 16065 19751 16099
rect 21649 16065 21683 16099
rect 24225 16065 24259 16099
rect 24685 16065 24719 16099
rect 1777 15997 1811 16031
rect 3157 15997 3191 16031
rect 5641 15997 5675 16031
rect 13093 15997 13127 16031
rect 14933 15997 14967 16031
rect 15669 15997 15703 16031
rect 17509 15997 17543 16031
rect 18613 15997 18647 16031
rect 22477 15997 22511 16031
rect 23029 15997 23063 16031
rect 24133 15997 24167 16031
rect 25237 15997 25271 16031
rect 949 15929 983 15963
rect 2789 15929 2823 15963
rect 3424 15929 3458 15963
rect 7481 15929 7515 15963
rect 7910 15929 7944 15963
rect 13645 15929 13679 15963
rect 18521 15929 18555 15963
rect 19984 15929 20018 15963
rect 23489 15929 23523 15963
rect 24041 15929 24075 15963
rect 1869 15861 1903 15895
rect 4537 15861 4571 15895
rect 6285 15861 6319 15895
rect 6653 15861 6687 15895
rect 11069 15861 11103 15895
rect 12725 15861 12759 15895
rect 13185 15861 13219 15895
rect 13553 15861 13587 15895
rect 14289 15861 14323 15895
rect 16497 15861 16531 15895
rect 17049 15861 17083 15895
rect 17785 15861 17819 15895
rect 18153 15861 18187 15895
rect 19349 15861 19383 15895
rect 21097 15861 21131 15895
rect 25053 15861 25087 15895
rect 25789 15861 25823 15895
rect 3617 15657 3651 15691
rect 4353 15657 4387 15691
rect 4997 15657 5031 15691
rect 6285 15657 6319 15691
rect 6653 15657 6687 15691
rect 6837 15657 6871 15691
rect 8217 15657 8251 15691
rect 8861 15657 8895 15691
rect 9229 15657 9263 15691
rect 19901 15657 19935 15691
rect 20729 15657 20763 15691
rect 22569 15657 22603 15691
rect 7297 15589 7331 15623
rect 13553 15589 13587 15623
rect 15577 15589 15611 15623
rect 23918 15589 23952 15623
rect 1869 15521 1903 15555
rect 1961 15521 1995 15555
rect 4905 15521 4939 15555
rect 5549 15521 5583 15555
rect 7205 15521 7239 15555
rect 8401 15521 8435 15555
rect 10968 15521 11002 15555
rect 13093 15521 13127 15555
rect 15301 15521 15335 15555
rect 17305 15521 17339 15555
rect 19717 15521 19751 15555
rect 21189 15521 21223 15555
rect 21445 15521 21479 15555
rect 2053 15453 2087 15487
rect 3065 15453 3099 15487
rect 5181 15453 5215 15487
rect 7389 15453 7423 15487
rect 9689 15453 9723 15487
rect 10701 15453 10735 15487
rect 13645 15453 13679 15487
rect 13829 15453 13863 15487
rect 17049 15453 17083 15487
rect 23673 15453 23707 15487
rect 2973 15385 3007 15419
rect 5917 15385 5951 15419
rect 7849 15385 7883 15419
rect 13185 15385 13219 15419
rect 1501 15317 1535 15351
rect 2605 15317 2639 15351
rect 3065 15317 3099 15351
rect 3341 15317 3375 15351
rect 4537 15317 4571 15351
rect 10149 15317 10183 15351
rect 10517 15317 10551 15351
rect 12081 15317 12115 15351
rect 12633 15317 12667 15351
rect 14289 15317 14323 15351
rect 14657 15317 14691 15351
rect 15025 15317 15059 15351
rect 16037 15317 16071 15351
rect 16865 15317 16899 15351
rect 18429 15317 18463 15351
rect 19349 15317 19383 15351
rect 20269 15317 20303 15351
rect 23121 15317 23155 15351
rect 23581 15317 23615 15351
rect 25053 15317 25087 15351
rect 1593 15113 1627 15147
rect 2513 15113 2547 15147
rect 3709 15113 3743 15147
rect 6193 15113 6227 15147
rect 6653 15113 6687 15147
rect 7021 15113 7055 15147
rect 16221 15113 16255 15147
rect 19625 15045 19659 15079
rect 23673 15045 23707 15079
rect 2053 14977 2087 15011
rect 3157 14977 3191 15011
rect 8033 14977 8067 15011
rect 10609 14977 10643 15011
rect 11253 14977 11287 15011
rect 11437 14977 11471 15011
rect 13001 14977 13035 15011
rect 18245 14977 18279 15011
rect 21465 14977 21499 15011
rect 22477 14977 22511 15011
rect 22661 14977 22695 15011
rect 24225 14977 24259 15011
rect 24685 14977 24719 15011
rect 25053 14977 25087 15011
rect 25421 14977 25455 15011
rect 1409 14909 1443 14943
rect 4261 14909 4295 14943
rect 4517 14909 4551 14943
rect 6837 14909 6871 14943
rect 10333 14909 10367 14943
rect 11161 14909 11195 14943
rect 12817 14909 12851 14943
rect 14289 14909 14323 14943
rect 16865 14909 16899 14943
rect 18512 14909 18546 14943
rect 20453 14909 20487 14943
rect 20729 14909 20763 14943
rect 23397 14909 23431 14943
rect 24133 14909 24167 14943
rect 25237 14909 25271 14943
rect 25973 14909 26007 14943
rect 2329 14841 2363 14875
rect 8278 14841 8312 14875
rect 11805 14841 11839 14875
rect 12909 14841 12943 14875
rect 14556 14841 14590 14875
rect 17877 14841 17911 14875
rect 21005 14841 21039 14875
rect 21925 14841 21959 14875
rect 22385 14841 22419 14875
rect 23121 14841 23155 14875
rect 24041 14841 24075 14875
rect 2881 14773 2915 14807
rect 2973 14773 3007 14807
rect 4169 14773 4203 14807
rect 5641 14773 5675 14807
rect 7481 14773 7515 14807
rect 7941 14773 7975 14807
rect 9413 14773 9447 14807
rect 10793 14773 10827 14807
rect 12173 14773 12207 14807
rect 12449 14773 12483 14807
rect 13461 14773 13495 14807
rect 13921 14773 13955 14807
rect 15669 14773 15703 14807
rect 16681 14773 16715 14807
rect 17049 14773 17083 14807
rect 17417 14773 17451 14807
rect 20269 14773 20303 14807
rect 20453 14773 20487 14807
rect 20545 14773 20579 14807
rect 22017 14773 22051 14807
rect 2605 14569 2639 14603
rect 4077 14569 4111 14603
rect 4445 14569 4479 14603
rect 5917 14569 5951 14603
rect 9045 14569 9079 14603
rect 9413 14569 9447 14603
rect 19257 14569 19291 14603
rect 21373 14569 21407 14603
rect 22477 14569 22511 14603
rect 25421 14569 25455 14603
rect 5181 14501 5215 14535
rect 12440 14501 12474 14535
rect 15761 14501 15795 14535
rect 17693 14501 17727 14535
rect 18613 14501 18647 14535
rect 20361 14501 20395 14535
rect 24685 14501 24719 14535
rect 25053 14501 25087 14535
rect 3617 14433 3651 14467
rect 6285 14433 6319 14467
rect 6377 14433 6411 14467
rect 8401 14433 8435 14467
rect 8493 14433 8527 14467
rect 9689 14433 9723 14467
rect 9956 14433 9990 14467
rect 15669 14433 15703 14467
rect 17601 14433 17635 14467
rect 19165 14433 19199 14467
rect 19625 14433 19659 14467
rect 21281 14433 21315 14467
rect 22109 14433 22143 14467
rect 23020 14433 23054 14467
rect 25237 14433 25271 14467
rect 1685 14365 1719 14399
rect 2053 14365 2087 14399
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 5825 14365 5859 14399
rect 6469 14365 6503 14399
rect 7573 14365 7607 14399
rect 8585 14365 8619 14399
rect 12173 14365 12207 14399
rect 14381 14365 14415 14399
rect 15945 14365 15979 14399
rect 17877 14365 17911 14399
rect 19717 14365 19751 14399
rect 19901 14365 19935 14399
rect 21557 14365 21591 14399
rect 22753 14365 22787 14399
rect 17141 14297 17175 14331
rect 20913 14297 20947 14331
rect 2237 14229 2271 14263
rect 3249 14229 3283 14263
rect 7021 14229 7055 14263
rect 7941 14229 7975 14263
rect 8033 14229 8067 14263
rect 11069 14229 11103 14263
rect 11713 14229 11747 14263
rect 11989 14229 12023 14263
rect 13553 14229 13587 14263
rect 14749 14229 14783 14263
rect 15025 14229 15059 14263
rect 15301 14229 15335 14263
rect 16497 14229 16531 14263
rect 17233 14229 17267 14263
rect 18245 14229 18279 14263
rect 20729 14229 20763 14263
rect 24133 14229 24167 14263
rect 7757 14025 7791 14059
rect 9321 14025 9355 14059
rect 12173 14025 12207 14059
rect 16405 14025 16439 14059
rect 17417 14025 17451 14059
rect 18061 14025 18095 14059
rect 19165 14025 19199 14059
rect 19625 14025 19659 14059
rect 20913 14025 20947 14059
rect 21373 14025 21407 14059
rect 21649 14025 21683 14059
rect 23029 14025 23063 14059
rect 23489 14025 23523 14059
rect 24777 14025 24811 14059
rect 5181 13957 5215 13991
rect 10793 13957 10827 13991
rect 17877 13957 17911 13991
rect 25973 13957 26007 13991
rect 5641 13889 5675 13923
rect 5733 13889 5767 13923
rect 6285 13889 6319 13923
rect 7481 13889 7515 13923
rect 10333 13889 10367 13923
rect 11345 13889 11379 13923
rect 17049 13889 17083 13923
rect 18613 13889 18647 13923
rect 20269 13889 20303 13923
rect 22661 13889 22695 13923
rect 24317 13889 24351 13923
rect 25421 13889 25455 13923
rect 2053 13821 2087 13855
rect 4721 13821 4755 13855
rect 6653 13821 6687 13855
rect 7941 13821 7975 13855
rect 8197 13821 8231 13855
rect 9873 13821 9907 13855
rect 10701 13821 10735 13855
rect 11253 13821 11287 13855
rect 13185 13821 13219 13855
rect 13277 13821 13311 13855
rect 13533 13821 13567 13855
rect 15301 13821 15335 13855
rect 15669 13821 15703 13855
rect 16865 13821 16899 13855
rect 18521 13821 18555 13855
rect 20085 13821 20119 13855
rect 25053 13821 25087 13855
rect 25237 13821 25271 13855
rect 2298 13753 2332 13787
rect 5089 13753 5123 13787
rect 5549 13753 5583 13787
rect 18429 13753 18463 13787
rect 19993 13753 20027 13787
rect 22385 13753 22419 13787
rect 24041 13753 24075 13787
rect 24133 13753 24167 13787
rect 1961 13685 1995 13719
rect 3433 13685 3467 13719
rect 4077 13685 4111 13719
rect 6929 13685 6963 13719
rect 11161 13685 11195 13719
rect 11897 13685 11931 13719
rect 12633 13685 12667 13719
rect 14657 13685 14691 13719
rect 16313 13685 16347 13719
rect 16773 13685 16807 13719
rect 19441 13685 19475 13719
rect 22017 13685 22051 13719
rect 22477 13685 22511 13719
rect 23673 13685 23707 13719
rect 1869 13481 1903 13515
rect 4353 13481 4387 13515
rect 4721 13481 4755 13515
rect 6285 13481 6319 13515
rect 7757 13481 7791 13515
rect 8493 13481 8527 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 11621 13481 11655 13515
rect 11713 13481 11747 13515
rect 13185 13481 13219 13515
rect 14013 13481 14047 13515
rect 15301 13481 15335 13515
rect 16497 13481 16531 13515
rect 18797 13481 18831 13515
rect 19257 13481 19291 13515
rect 20085 13481 20119 13515
rect 20913 13481 20947 13515
rect 22109 13481 22143 13515
rect 23305 13481 23339 13515
rect 23673 13481 23707 13515
rect 5172 13413 5206 13447
rect 9413 13413 9447 13447
rect 21281 13413 21315 13447
rect 24032 13413 24066 13447
rect 2237 13345 2271 13379
rect 6837 13345 6871 13379
rect 7481 13345 7515 13379
rect 8401 13345 8435 13379
rect 10057 13345 10091 13379
rect 15025 13345 15059 13379
rect 15669 13345 15703 13379
rect 17132 13345 17166 13379
rect 19349 13345 19383 13379
rect 22477 13345 22511 13379
rect 2329 13277 2363 13311
rect 2421 13277 2455 13311
rect 4905 13277 4939 13311
rect 8677 13277 8711 13311
rect 10241 13277 10275 13311
rect 11897 13277 11931 13311
rect 12725 13277 12759 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15761 13277 15795 13311
rect 15853 13277 15887 13311
rect 16865 13277 16899 13311
rect 19625 13277 19659 13311
rect 20729 13277 20763 13311
rect 21373 13277 21407 13311
rect 21557 13277 21591 13311
rect 22661 13277 22695 13311
rect 23765 13277 23799 13311
rect 8033 13209 8067 13243
rect 13645 13209 13679 13243
rect 18245 13209 18279 13243
rect 949 13141 983 13175
rect 1593 13141 1627 13175
rect 2973 13141 3007 13175
rect 3249 13141 3283 13175
rect 3709 13141 3743 13175
rect 10793 13141 10827 13175
rect 11253 13141 11287 13175
rect 12265 13141 12299 13175
rect 13461 13141 13495 13175
rect 14657 13141 14691 13175
rect 25145 13141 25179 13175
rect 4537 12937 4571 12971
rect 5181 12937 5215 12971
rect 5825 12937 5859 12971
rect 7757 12937 7791 12971
rect 8769 12937 8803 12971
rect 9137 12937 9171 12971
rect 10701 12937 10735 12971
rect 11897 12937 11931 12971
rect 12265 12937 12299 12971
rect 13645 12937 13679 12971
rect 17141 12937 17175 12971
rect 17417 12937 17451 12971
rect 17693 12937 17727 12971
rect 19441 12937 19475 12971
rect 19901 12937 19935 12971
rect 22661 12937 22695 12971
rect 23029 12937 23063 12971
rect 23489 12937 23523 12971
rect 1593 12869 1627 12903
rect 7297 12869 7331 12903
rect 13553 12869 13587 12903
rect 16589 12869 16623 12903
rect 949 12801 983 12835
rect 2053 12801 2087 12835
rect 2145 12801 2179 12835
rect 5549 12801 5583 12835
rect 8217 12801 8251 12835
rect 8309 12801 8343 12835
rect 9873 12801 9907 12835
rect 13185 12801 13219 12835
rect 14197 12801 14231 12835
rect 14657 12801 14691 12835
rect 15117 12801 15151 12835
rect 3157 12733 3191 12767
rect 5641 12733 5675 12767
rect 6193 12733 6227 12767
rect 7573 12733 7607 12767
rect 8125 12733 8159 12767
rect 11069 12733 11103 12767
rect 14013 12733 14047 12767
rect 15209 12733 15243 12767
rect 15476 12733 15510 12767
rect 18613 12801 18647 12835
rect 19073 12801 19107 12835
rect 20361 12801 20395 12835
rect 24225 12801 24259 12835
rect 24869 12801 24903 12835
rect 25053 12801 25087 12835
rect 25421 12801 25455 12835
rect 17509 12733 17543 12767
rect 17877 12733 17911 12767
rect 20085 12733 20119 12767
rect 20617 12733 20651 12767
rect 2605 12665 2639 12699
rect 3402 12665 3436 12699
rect 9689 12665 9723 12699
rect 10425 12665 10459 12699
rect 11345 12665 11379 12699
rect 17417 12665 17451 12699
rect 18429 12665 18463 12699
rect 23949 12665 23983 12699
rect 24777 12665 24811 12699
rect 1961 12597 1995 12631
rect 2973 12597 3007 12631
rect 6653 12597 6687 12631
rect 9321 12597 9355 12631
rect 9781 12597 9815 12631
rect 12633 12597 12667 12631
rect 14105 12597 14139 12631
rect 18061 12597 18095 12631
rect 18521 12597 18555 12631
rect 21741 12597 21775 12631
rect 22293 12597 22327 12631
rect 24409 12597 24443 12631
rect 25881 12597 25915 12631
rect 26157 12597 26191 12631
rect 1685 12393 1719 12427
rect 3525 12393 3559 12427
rect 4261 12393 4295 12427
rect 4445 12393 4479 12427
rect 6009 12393 6043 12427
rect 8769 12393 8803 12427
rect 12265 12393 12299 12427
rect 13185 12393 13219 12427
rect 15117 12393 15151 12427
rect 15301 12393 15335 12427
rect 17417 12393 17451 12427
rect 19349 12393 19383 12427
rect 20453 12393 20487 12427
rect 20913 12393 20947 12427
rect 21925 12393 21959 12427
rect 24869 12393 24903 12427
rect 4905 12325 4939 12359
rect 10600 12325 10634 12359
rect 14749 12325 14783 12359
rect 2053 12257 2087 12291
rect 2145 12257 2179 12291
rect 3801 12257 3835 12291
rect 4813 12257 4847 12291
rect 6193 12257 6227 12291
rect 6469 12257 6503 12291
rect 7104 12257 7138 12291
rect 9505 12257 9539 12291
rect 14013 12257 14047 12291
rect 15669 12257 15703 12291
rect 16865 12257 16899 12291
rect 17969 12257 18003 12291
rect 18236 12257 18270 12291
rect 19993 12257 20027 12291
rect 21281 12257 21315 12291
rect 23213 12257 23247 12291
rect 24777 12257 24811 12291
rect 2329 12189 2363 12223
rect 3157 12189 3191 12223
rect 5089 12189 5123 12223
rect 6837 12189 6871 12223
rect 10333 12189 10367 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 21373 12189 21407 12223
rect 21465 12189 21499 12223
rect 23305 12189 23339 12223
rect 23489 12189 23523 12223
rect 24225 12189 24259 12223
rect 25053 12189 25087 12223
rect 5917 12121 5951 12155
rect 9321 12121 9355 12155
rect 13645 12121 13679 12155
rect 22753 12121 22787 12155
rect 2697 12053 2731 12087
rect 5457 12053 5491 12087
rect 8217 12053 8251 12087
rect 9137 12053 9171 12087
rect 9965 12053 9999 12087
rect 11713 12053 11747 12087
rect 12725 12053 12759 12087
rect 13553 12053 13587 12087
rect 16405 12053 16439 12087
rect 16773 12053 16807 12087
rect 17049 12053 17083 12087
rect 17785 12053 17819 12087
rect 22385 12053 22419 12087
rect 22845 12053 22879 12087
rect 24409 12053 24443 12087
rect 25513 12053 25547 12087
rect 1501 11849 1535 11883
rect 3709 11849 3743 11883
rect 4169 11849 4203 11883
rect 7665 11849 7699 11883
rect 10793 11849 10827 11883
rect 14381 11849 14415 11883
rect 15853 11849 15887 11883
rect 17049 11849 17083 11883
rect 17601 11849 17635 11883
rect 18613 11849 18647 11883
rect 19257 11849 19291 11883
rect 20729 11849 20763 11883
rect 21281 11849 21315 11883
rect 23305 11849 23339 11883
rect 23949 11849 23983 11883
rect 5917 11781 5951 11815
rect 9137 11781 9171 11815
rect 12081 11781 12115 11815
rect 12173 11781 12207 11815
rect 16037 11781 16071 11815
rect 17693 11781 17727 11815
rect 21741 11781 21775 11815
rect 1777 11713 1811 11747
rect 5365 11713 5399 11747
rect 5549 11713 5583 11747
rect 7573 11713 7607 11747
rect 8217 11713 8251 11747
rect 9781 11713 9815 11747
rect 11437 11713 11471 11747
rect 2033 11645 2067 11679
rect 8125 11645 8159 11679
rect 9689 11645 9723 11679
rect 1501 11577 1535 11611
rect 1685 11577 1719 11611
rect 4537 11577 4571 11611
rect 6653 11577 6687 11611
rect 8033 11577 8067 11611
rect 10609 11577 10643 11611
rect 11253 11577 11287 11611
rect 16589 11713 16623 11747
rect 22477 11713 22511 11747
rect 12449 11645 12483 11679
rect 12705 11645 12739 11679
rect 14933 11645 14967 11679
rect 16405 11645 16439 11679
rect 17877 11645 17911 11679
rect 18061 11645 18095 11679
rect 19349 11645 19383 11679
rect 19605 11645 19639 11679
rect 22293 11645 22327 11679
rect 24133 11645 24167 11679
rect 14841 11577 14875 11611
rect 24400 11577 24434 11611
rect 3157 11509 3191 11543
rect 4905 11509 4939 11543
rect 5273 11509 5307 11543
rect 7113 11509 7147 11543
rect 8677 11509 8711 11543
rect 9229 11509 9263 11543
rect 9597 11509 9631 11543
rect 10241 11509 10275 11543
rect 11161 11509 11195 11543
rect 11805 11509 11839 11543
rect 12081 11509 12115 11543
rect 13829 11509 13863 11543
rect 15117 11509 15151 11543
rect 15485 11509 15519 11543
rect 16497 11509 16531 11543
rect 18245 11509 18279 11543
rect 21925 11509 21959 11543
rect 22385 11509 22419 11543
rect 22937 11509 22971 11543
rect 25513 11509 25547 11543
rect 26065 11509 26099 11543
rect 1593 11305 1627 11339
rect 2053 11305 2087 11339
rect 3341 11305 3375 11339
rect 4537 11305 4571 11339
rect 6101 11305 6135 11339
rect 8309 11305 8343 11339
rect 8585 11305 8619 11339
rect 8769 11305 8803 11339
rect 14197 11305 14231 11339
rect 14565 11305 14599 11339
rect 15485 11305 15519 11339
rect 16405 11305 16439 11339
rect 16773 11305 16807 11339
rect 19073 11305 19107 11339
rect 20729 11305 20763 11339
rect 21281 11305 21315 11339
rect 22017 11305 22051 11339
rect 24317 11305 24351 11339
rect 24869 11305 24903 11339
rect 25237 11305 25271 11339
rect 2697 11237 2731 11271
rect 4966 11237 5000 11271
rect 7573 11237 7607 11271
rect 9321 11237 9355 11271
rect 10149 11237 10183 11271
rect 13553 11237 13587 11271
rect 16221 11237 16255 11271
rect 17509 11237 17543 11271
rect 19441 11237 19475 11271
rect 22845 11237 22879 11271
rect 1961 11169 1995 11203
rect 3709 11169 3743 11203
rect 6745 11169 6779 11203
rect 7113 11169 7147 11203
rect 8953 11169 8987 11203
rect 10497 11169 10531 11203
rect 15301 11169 15335 11203
rect 18337 11169 18371 11203
rect 19533 11169 19567 11203
rect 22937 11169 22971 11203
rect 23204 11169 23238 11203
rect 2145 11101 2179 11135
rect 4721 11101 4755 11135
rect 7665 11101 7699 11135
rect 7849 11101 7883 11135
rect 10241 11101 10275 11135
rect 12541 11101 12575 11135
rect 13645 11101 13679 11135
rect 13737 11101 13771 11135
rect 15945 11101 15979 11135
rect 16865 11101 16899 11135
rect 16957 11101 16991 11135
rect 18429 11101 18463 11135
rect 18613 11101 18647 11135
rect 20177 11101 20211 11135
rect 21373 11101 21407 11135
rect 21465 11101 21499 11135
rect 25421 11101 25455 11135
rect 7205 11033 7239 11067
rect 12173 11033 12207 11067
rect 13093 11033 13127 11067
rect 14933 11033 14967 11067
rect 17877 11033 17911 11067
rect 17969 11033 18003 11067
rect 19717 11033 19751 11067
rect 20913 11033 20947 11067
rect 949 10965 983 10999
rect 2973 10965 3007 10999
rect 11621 10965 11655 10999
rect 13185 10965 13219 10999
rect 22385 10965 22419 10999
rect 4445 10761 4479 10795
rect 5549 10761 5583 10795
rect 6561 10761 6595 10795
rect 11529 10761 11563 10795
rect 14933 10761 14967 10795
rect 16865 10761 16899 10795
rect 20085 10761 20119 10795
rect 20453 10761 20487 10795
rect 22293 10761 22327 10795
rect 24225 10761 24259 10795
rect 25881 10761 25915 10795
rect 10149 10693 10183 10727
rect 17417 10693 17451 10727
rect 25421 10693 25455 10727
rect 1685 10625 1719 10659
rect 3985 10625 4019 10659
rect 4905 10625 4939 10659
rect 4997 10625 5031 10659
rect 6837 10625 6871 10659
rect 10057 10625 10091 10659
rect 10701 10625 10735 10659
rect 21741 10625 21775 10659
rect 21925 10625 21959 10659
rect 24869 10625 24903 10659
rect 25053 10625 25087 10659
rect 1952 10557 1986 10591
rect 4353 10557 4387 10591
rect 9321 10557 9355 10591
rect 10609 10557 10643 10591
rect 13001 10557 13035 10591
rect 15485 10557 15519 10591
rect 18061 10557 18095 10591
rect 4813 10489 4847 10523
rect 5825 10489 5859 10523
rect 7082 10489 7116 10523
rect 9689 10489 9723 10523
rect 10517 10489 10551 10523
rect 11161 10489 11195 10523
rect 12265 10489 12299 10523
rect 13268 10489 13302 10523
rect 15393 10489 15427 10523
rect 15752 10489 15786 10523
rect 18306 10489 18340 10523
rect 21097 10489 21131 10523
rect 21649 10489 21683 10523
rect 24777 10489 24811 10523
rect 3065 10421 3099 10455
rect 6193 10421 6227 10455
rect 8217 10421 8251 10455
rect 8769 10421 8803 10455
rect 12909 10421 12943 10455
rect 14381 10421 14415 10455
rect 17785 10421 17819 10455
rect 19441 10421 19475 10455
rect 20821 10421 20855 10455
rect 21281 10421 21315 10455
rect 23029 10421 23063 10455
rect 23397 10421 23431 10455
rect 23949 10421 23983 10455
rect 24409 10421 24443 10455
rect 1409 10217 1443 10251
rect 2789 10217 2823 10251
rect 3433 10217 3467 10251
rect 6285 10217 6319 10251
rect 6837 10217 6871 10251
rect 7297 10217 7331 10251
rect 8401 10217 8435 10251
rect 11437 10217 11471 10251
rect 11989 10217 12023 10251
rect 12633 10217 12667 10251
rect 13461 10217 13495 10251
rect 14473 10217 14507 10251
rect 15117 10217 15151 10251
rect 15301 10217 15335 10251
rect 15761 10217 15795 10251
rect 17693 10217 17727 10251
rect 18245 10217 18279 10251
rect 18613 10217 18647 10251
rect 19717 10217 19751 10251
rect 21925 10217 21959 10251
rect 22661 10217 22695 10251
rect 23121 10217 23155 10251
rect 24225 10217 24259 10251
rect 2329 10149 2363 10183
rect 4261 10149 4295 10183
rect 5172 10149 5206 10183
rect 8493 10149 8527 10183
rect 10302 10149 10336 10183
rect 16580 10149 16614 10183
rect 19625 10149 19659 10183
rect 21373 10149 21407 10183
rect 25421 10149 25455 10183
rect 1961 10081 1995 10115
rect 4905 10081 4939 10115
rect 14105 10081 14139 10115
rect 16313 10081 16347 10115
rect 21281 10081 21315 10115
rect 23029 10081 23063 10115
rect 24777 10081 24811 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 8677 10013 8711 10047
rect 10057 10013 10091 10047
rect 13001 10013 13035 10047
rect 13553 10013 13587 10047
rect 13645 10013 13679 10047
rect 19809 10013 19843 10047
rect 20361 10013 20395 10047
rect 20637 10013 20671 10047
rect 21557 10013 21591 10047
rect 23213 10013 23247 10047
rect 24869 10013 24903 10047
rect 24961 10013 24995 10047
rect 2421 9945 2455 9979
rect 9137 9945 9171 9979
rect 16129 9945 16163 9979
rect 3893 9877 3927 9911
rect 4721 9877 4755 9911
rect 7849 9877 7883 9911
rect 8033 9877 8067 9911
rect 9413 9877 9447 9911
rect 9965 9877 9999 9911
rect 13093 9877 13127 9911
rect 19073 9877 19107 9911
rect 19257 9877 19291 9911
rect 20913 9877 20947 9911
rect 22385 9877 22419 9911
rect 23765 9877 23799 9911
rect 24409 9877 24443 9911
rect 2881 9673 2915 9707
rect 4629 9673 4663 9707
rect 9689 9673 9723 9707
rect 10057 9673 10091 9707
rect 10241 9673 10275 9707
rect 16865 9673 16899 9707
rect 17785 9673 17819 9707
rect 19349 9673 19383 9707
rect 22385 9673 22419 9707
rect 24041 9673 24075 9707
rect 1409 9605 1443 9639
rect 2513 9605 2547 9639
rect 3065 9605 3099 9639
rect 4537 9605 4571 9639
rect 5641 9605 5675 9639
rect 7297 9605 7331 9639
rect 9137 9605 9171 9639
rect 11989 9605 12023 9639
rect 13001 9605 13035 9639
rect 15853 9605 15887 9639
rect 18061 9605 18095 9639
rect 22661 9605 22695 9639
rect 1961 9537 1995 9571
rect 3709 9537 3743 9571
rect 5181 9537 5215 9571
rect 7573 9537 7607 9571
rect 10793 9537 10827 9571
rect 16405 9537 16439 9571
rect 17509 9537 17543 9571
rect 18521 9537 18555 9571
rect 18613 9537 18647 9571
rect 24133 9537 24167 9571
rect 1869 9469 1903 9503
rect 3525 9469 3559 9503
rect 4169 9469 4203 9503
rect 7757 9469 7791 9503
rect 10609 9469 10643 9503
rect 11621 9469 11655 9503
rect 13185 9469 13219 9503
rect 16221 9469 16255 9503
rect 18429 9469 18463 9503
rect 19625 9469 19659 9503
rect 22477 9469 22511 9503
rect 23029 9469 23063 9503
rect 24389 9469 24423 9503
rect 26065 9469 26099 9503
rect 1777 9401 1811 9435
rect 4997 9401 5031 9435
rect 8002 9401 8036 9435
rect 12725 9401 12759 9435
rect 14933 9401 14967 9435
rect 16313 9401 16347 9435
rect 19892 9401 19926 9435
rect 3433 9333 3467 9367
rect 5089 9333 5123 9367
rect 6193 9333 6227 9367
rect 6561 9333 6595 9367
rect 10701 9333 10735 9367
rect 11253 9333 11287 9367
rect 15301 9333 15335 9367
rect 15669 9333 15703 9367
rect 21005 9333 21039 9367
rect 21557 9333 21591 9367
rect 21925 9333 21959 9367
rect 23489 9333 23523 9367
rect 25513 9333 25547 9367
rect 1409 9129 1443 9163
rect 1961 9129 1995 9163
rect 2421 9129 2455 9163
rect 5549 9129 5583 9163
rect 8493 9129 8527 9163
rect 10425 9129 10459 9163
rect 17141 9129 17175 9163
rect 17601 9129 17635 9163
rect 18705 9129 18739 9163
rect 19257 9129 19291 9163
rect 20269 9129 20303 9163
rect 21281 9129 21315 9163
rect 22753 9129 22787 9163
rect 24501 9129 24535 9163
rect 2789 9061 2823 9095
rect 6009 9061 6043 9095
rect 7380 9061 7414 9095
rect 10333 9061 10367 9095
rect 12449 9061 12483 9095
rect 18061 9061 18095 9095
rect 18153 9061 18187 9095
rect 19073 9061 19107 9095
rect 25421 9061 25455 9095
rect 2329 8993 2363 9027
rect 5917 8993 5951 9027
rect 9045 8993 9079 9027
rect 9965 8993 9999 9027
rect 10793 8993 10827 9027
rect 12357 8993 12391 9027
rect 13636 8993 13670 9027
rect 16497 8993 16531 9027
rect 19625 8993 19659 9027
rect 23121 8993 23155 9027
rect 23388 8993 23422 9027
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 4353 8925 4387 8959
rect 4537 8925 4571 8959
rect 6101 8925 6135 8959
rect 7113 8925 7147 8959
rect 10885 8925 10919 8959
rect 10977 8925 11011 8959
rect 12541 8925 12575 8959
rect 13369 8925 13403 8959
rect 16589 8925 16623 8959
rect 16681 8925 16715 8959
rect 18337 8925 18371 8959
rect 19717 8925 19751 8959
rect 19901 8925 19935 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 3801 8857 3835 8891
rect 11989 8857 12023 8891
rect 17693 8857 17727 8891
rect 20913 8857 20947 8891
rect 22293 8857 22327 8891
rect 3433 8789 3467 8823
rect 4997 8789 5031 8823
rect 5365 8789 5399 8823
rect 6929 8789 6963 8823
rect 9413 8789 9447 8823
rect 11529 8789 11563 8823
rect 11897 8789 11931 8823
rect 13277 8789 13311 8823
rect 14749 8789 14783 8823
rect 15485 8789 15519 8823
rect 15945 8789 15979 8823
rect 16129 8789 16163 8823
rect 20729 8789 20763 8823
rect 21925 8789 21959 8823
rect 25053 8789 25087 8823
rect 1777 8585 1811 8619
rect 3801 8585 3835 8619
rect 5641 8585 5675 8619
rect 9229 8585 9263 8619
rect 9965 8585 9999 8619
rect 10425 8585 10459 8619
rect 12449 8585 12483 8619
rect 13553 8585 13587 8619
rect 15393 8585 15427 8619
rect 15853 8585 15887 8619
rect 17785 8585 17819 8619
rect 18245 8585 18279 8619
rect 18613 8585 18647 8619
rect 20361 8585 20395 8619
rect 25605 8585 25639 8619
rect 3249 8517 3283 8551
rect 4353 8517 4387 8551
rect 8401 8517 8435 8551
rect 14381 8517 14415 8551
rect 21465 8517 21499 8551
rect 4905 8449 4939 8483
rect 7021 8449 7055 8483
rect 9597 8449 9631 8483
rect 10977 8449 11011 8483
rect 13001 8449 13035 8483
rect 14105 8449 14139 8483
rect 14933 8449 14967 8483
rect 16957 8449 16991 8483
rect 18981 8449 19015 8483
rect 22017 8449 22051 8483
rect 23673 8449 23707 8483
rect 1869 8381 1903 8415
rect 2136 8381 2170 8415
rect 4261 8381 4295 8415
rect 4721 8381 4755 8415
rect 6653 8381 6687 8415
rect 7288 8381 7322 8415
rect 10241 8381 10275 8415
rect 14013 8381 14047 8415
rect 14749 8381 14783 8415
rect 16773 8381 16807 8415
rect 16865 8381 16899 8415
rect 19237 8381 19271 8415
rect 21005 8381 21039 8415
rect 21833 8381 21867 8415
rect 4813 8313 4847 8347
rect 10793 8313 10827 8347
rect 10885 8313 10919 8347
rect 11713 8313 11747 8347
rect 12909 8313 12943 8347
rect 13921 8313 13955 8347
rect 16129 8313 16163 8347
rect 21373 8313 21407 8347
rect 21925 8313 21959 8347
rect 23918 8313 23952 8347
rect 6285 8245 6319 8279
rect 11989 8245 12023 8279
rect 12817 8245 12851 8279
rect 14841 8245 14875 8279
rect 16405 8245 16439 8279
rect 22753 8245 22787 8279
rect 23213 8245 23247 8279
rect 25053 8245 25087 8279
rect 1961 8041 1995 8075
rect 2237 8041 2271 8075
rect 2421 8041 2455 8075
rect 3893 8041 3927 8075
rect 4905 8041 4939 8075
rect 5549 8041 5583 8075
rect 5917 8041 5951 8075
rect 6837 8041 6871 8075
rect 7849 8041 7883 8075
rect 10425 8041 10459 8075
rect 10885 8041 10919 8075
rect 12357 8041 12391 8075
rect 13369 8041 13403 8075
rect 14473 8041 14507 8075
rect 15301 8041 15335 8075
rect 16129 8041 16163 8075
rect 17693 8041 17727 8075
rect 19073 8041 19107 8075
rect 19441 8041 19475 8075
rect 20177 8041 20211 8075
rect 20545 8041 20579 8075
rect 21097 8041 21131 8075
rect 21925 8041 21959 8075
rect 22937 8041 22971 8075
rect 23121 8041 23155 8075
rect 25053 8041 25087 8075
rect 4353 7973 4387 8007
rect 7573 7973 7607 8007
rect 11222 7973 11256 8007
rect 14841 7973 14875 8007
rect 18337 7973 18371 8007
rect 1409 7905 1443 7939
rect 2789 7905 2823 7939
rect 3525 7905 3559 7939
rect 8401 7905 8435 7939
rect 9689 7905 9723 7939
rect 10977 7905 11011 7939
rect 13829 7905 13863 7939
rect 13921 7905 13955 7939
rect 16569 7905 16603 7939
rect 18981 7905 19015 7939
rect 22661 7905 22695 7939
rect 23489 7905 23523 7939
rect 24133 7905 24167 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 6929 7837 6963 7871
rect 7113 7837 7147 7871
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 9965 7837 9999 7871
rect 14013 7837 14047 7871
rect 16313 7837 16347 7871
rect 19533 7837 19567 7871
rect 19625 7837 19659 7871
rect 22017 7837 22051 7871
rect 22109 7837 22143 7871
rect 23581 7837 23615 7871
rect 23673 7837 23707 7871
rect 25145 7837 25179 7871
rect 25329 7837 25363 7871
rect 4537 7769 4571 7803
rect 6469 7769 6503 7803
rect 18613 7769 18647 7803
rect 24685 7769 24719 7803
rect 6285 7701 6319 7735
rect 8033 7701 8067 7735
rect 9045 7701 9079 7735
rect 9505 7701 9539 7735
rect 12909 7701 12943 7735
rect 13461 7701 13495 7735
rect 15853 7701 15887 7735
rect 18797 7701 18831 7735
rect 21557 7701 21591 7735
rect 24501 7701 24535 7735
rect 1593 7497 1627 7531
rect 3617 7497 3651 7531
rect 5181 7497 5215 7531
rect 6837 7497 6871 7531
rect 9597 7497 9631 7531
rect 11897 7497 11931 7531
rect 12265 7497 12299 7531
rect 13277 7497 13311 7531
rect 15577 7497 15611 7531
rect 19165 7497 19199 7531
rect 19809 7497 19843 7531
rect 20821 7497 20855 7531
rect 21373 7497 21407 7531
rect 21833 7497 21867 7531
rect 22017 7497 22051 7531
rect 23213 7497 23247 7531
rect 24041 7497 24075 7531
rect 25605 7497 25639 7531
rect 25973 7497 26007 7531
rect 6653 7429 6687 7463
rect 8585 7429 8619 7463
rect 16313 7429 16347 7463
rect 21189 7429 21223 7463
rect 26341 7429 26375 7463
rect 2053 7361 2087 7395
rect 2145 7361 2179 7395
rect 4169 7361 4203 7395
rect 5733 7361 5767 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 9229 7361 9263 7395
rect 10793 7361 10827 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 18521 7361 18555 7395
rect 18613 7361 18647 7395
rect 20453 7361 20487 7395
rect 22661 7361 22695 7395
rect 25145 7361 25179 7395
rect 2697 7293 2731 7327
rect 4721 7293 4755 7327
rect 5641 7293 5675 7327
rect 8401 7293 8435 7327
rect 10517 7293 10551 7327
rect 13369 7293 13403 7327
rect 13636 7293 13670 7327
rect 16773 7293 16807 7327
rect 18429 7293 18463 7327
rect 20269 7293 20303 7327
rect 21557 7293 21591 7327
rect 25053 7293 25087 7327
rect 3525 7225 3559 7259
rect 4077 7225 4111 7259
rect 5089 7225 5123 7259
rect 5549 7225 5583 7259
rect 17417 7225 17451 7259
rect 20177 7225 20211 7259
rect 22385 7225 22419 7259
rect 24501 7225 24535 7259
rect 1961 7157 1995 7191
rect 2973 7157 3007 7191
rect 3985 7157 4019 7191
rect 6193 7157 6227 7191
rect 7205 7157 7239 7191
rect 8033 7157 8067 7191
rect 8953 7157 8987 7191
rect 9045 7157 9079 7191
rect 10057 7157 10091 7191
rect 10149 7157 10183 7191
rect 10609 7157 10643 7191
rect 11161 7157 11195 7191
rect 12909 7157 12943 7191
rect 14749 7157 14783 7191
rect 15945 7157 15979 7191
rect 16405 7157 16439 7191
rect 17785 7157 17819 7191
rect 18061 7157 18095 7191
rect 19441 7157 19475 7191
rect 22477 7157 22511 7191
rect 24593 7157 24627 7191
rect 24961 7157 24995 7191
rect 4629 6953 4663 6987
rect 5641 6953 5675 6987
rect 5825 6953 5859 6987
rect 7757 6953 7791 6987
rect 9413 6953 9447 6987
rect 11989 6953 12023 6987
rect 12633 6953 12667 6987
rect 14105 6953 14139 6987
rect 17509 6953 17543 6987
rect 20269 6953 20303 6987
rect 20729 6953 20763 6987
rect 22937 6953 22971 6987
rect 25789 6953 25823 6987
rect 2789 6885 2823 6919
rect 8585 6885 8619 6919
rect 13001 6885 13035 6919
rect 19533 6885 19567 6919
rect 1409 6817 1443 6851
rect 2329 6817 2363 6851
rect 4721 6817 4755 6851
rect 6193 6817 6227 6851
rect 9137 6817 9171 6851
rect 10517 6817 10551 6851
rect 10865 6817 10899 6851
rect 13461 6817 13495 6851
rect 14841 6817 14875 6851
rect 15577 6817 15611 6851
rect 16037 6817 16071 6851
rect 16396 6817 16430 6851
rect 18797 6817 18831 6851
rect 20913 6817 20947 6851
rect 21169 6817 21203 6851
rect 23305 6817 23339 6851
rect 23664 6817 23698 6851
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 4813 6749 4847 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 7849 6749 7883 6783
rect 8033 6749 8067 6783
rect 10609 6749 10643 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 16129 6749 16163 6783
rect 18521 6749 18555 6783
rect 19625 6749 19659 6783
rect 19809 6749 19843 6783
rect 23397 6749 23431 6783
rect 5365 6681 5399 6715
rect 10149 6681 10183 6715
rect 13093 6681 13127 6715
rect 24777 6681 24811 6715
rect 1961 6613 1995 6647
rect 2421 6613 2455 6647
rect 3617 6613 3651 6647
rect 4261 6613 4295 6647
rect 7021 6613 7055 6647
rect 7389 6613 7423 6647
rect 8953 6613 8987 6647
rect 14473 6613 14507 6647
rect 18061 6613 18095 6647
rect 18613 6613 18647 6647
rect 19165 6613 19199 6647
rect 22293 6613 22327 6647
rect 25329 6613 25363 6647
rect 1961 6409 1995 6443
rect 3801 6409 3835 6443
rect 4445 6409 4479 6443
rect 4721 6409 4755 6443
rect 5089 6409 5123 6443
rect 7941 6409 7975 6443
rect 13921 6409 13955 6443
rect 18613 6409 18647 6443
rect 21005 6409 21039 6443
rect 21557 6409 21591 6443
rect 22569 6409 22603 6443
rect 23673 6409 23707 6443
rect 26341 6409 26375 6443
rect 6653 6341 6687 6375
rect 11897 6341 11931 6375
rect 19073 6341 19107 6375
rect 2421 6273 2455 6307
rect 5549 6273 5583 6307
rect 5641 6273 5675 6307
rect 7573 6273 7607 6307
rect 9689 6273 9723 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 18061 6273 18095 6307
rect 19717 6273 19751 6307
rect 22017 6273 22051 6307
rect 22201 6273 22235 6307
rect 23489 6273 23523 6307
rect 24225 6273 24259 6307
rect 25421 6273 25455 6307
rect 8585 6205 8619 6239
rect 9873 6205 9907 6239
rect 10140 6205 10174 6239
rect 12173 6205 12207 6239
rect 14105 6205 14139 6239
rect 16589 6205 16623 6239
rect 17325 6205 17359 6239
rect 18889 6205 18923 6239
rect 21925 6205 21959 6239
rect 23121 6205 23155 6239
rect 24133 6205 24167 6239
rect 25237 6205 25271 6239
rect 25973 6205 26007 6239
rect 2237 6137 2271 6171
rect 2688 6137 2722 6171
rect 8861 6137 8895 6171
rect 12817 6137 12851 6171
rect 14350 6137 14384 6171
rect 16865 6137 16899 6171
rect 17877 6137 17911 6171
rect 19533 6137 19567 6171
rect 21465 6137 21499 6171
rect 24041 6137 24075 6171
rect 24685 6137 24719 6171
rect 1409 6069 1443 6103
rect 5457 6069 5491 6103
rect 6101 6069 6135 6103
rect 6929 6069 6963 6103
rect 7297 6069 7331 6103
rect 7389 6069 7423 6103
rect 8401 6069 8435 6103
rect 9413 6069 9447 6103
rect 11253 6069 11287 6103
rect 12449 6069 12483 6103
rect 13461 6069 13495 6103
rect 15485 6069 15519 6103
rect 16129 6069 16163 6103
rect 19441 6069 19475 6103
rect 20085 6069 20119 6103
rect 20545 6069 20579 6103
rect 25053 6069 25087 6103
rect 3893 5865 3927 5899
rect 5733 5865 5767 5899
rect 6653 5865 6687 5899
rect 9045 5865 9079 5899
rect 10517 5865 10551 5899
rect 13185 5865 13219 5899
rect 16773 5865 16807 5899
rect 17877 5865 17911 5899
rect 18245 5865 18279 5899
rect 20913 5865 20947 5899
rect 21925 5865 21959 5899
rect 22385 5865 22419 5899
rect 23949 5865 23983 5899
rect 24317 5865 24351 5899
rect 24961 5865 24995 5899
rect 25329 5865 25363 5899
rect 25697 5865 25731 5899
rect 4598 5797 4632 5831
rect 6285 5797 6319 5831
rect 10425 5797 10459 5831
rect 13093 5797 13127 5831
rect 17325 5797 17359 5831
rect 20269 5797 20303 5831
rect 22753 5797 22787 5831
rect 23765 5797 23799 5831
rect 1501 5729 1535 5763
rect 1768 5729 1802 5763
rect 7021 5729 7055 5763
rect 7380 5729 7414 5763
rect 10885 5729 10919 5763
rect 10977 5729 11011 5763
rect 11529 5729 11563 5763
rect 11897 5729 11931 5763
rect 12081 5729 12115 5763
rect 13553 5729 13587 5763
rect 13645 5729 13679 5763
rect 15649 5729 15683 5763
rect 18593 5729 18627 5763
rect 21281 5729 21315 5763
rect 22477 5729 22511 5763
rect 23213 5729 23247 5763
rect 24409 5729 24443 5763
rect 4353 5661 4387 5695
rect 7113 5661 7147 5695
rect 11069 5661 11103 5695
rect 13737 5661 13771 5695
rect 15393 5661 15427 5695
rect 18337 5661 18371 5695
rect 20729 5661 20763 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 24501 5661 24535 5695
rect 6837 5593 6871 5627
rect 8493 5593 8527 5627
rect 2881 5525 2915 5559
rect 3433 5525 3467 5559
rect 9413 5525 9447 5559
rect 10057 5525 10091 5559
rect 12265 5525 12299 5559
rect 12633 5525 12667 5559
rect 14289 5525 14323 5559
rect 14565 5525 14599 5559
rect 15025 5525 15059 5559
rect 19717 5525 19751 5559
rect 1501 5321 1535 5355
rect 3065 5321 3099 5355
rect 4353 5321 4387 5355
rect 6193 5321 6227 5355
rect 7849 5321 7883 5355
rect 8953 5321 8987 5355
rect 10425 5321 10459 5355
rect 10517 5321 10551 5355
rect 11897 5321 11931 5355
rect 14933 5321 14967 5355
rect 17233 5321 17267 5355
rect 17601 5321 17635 5355
rect 21373 5321 21407 5355
rect 23489 5321 23523 5355
rect 25605 5321 25639 5355
rect 25973 5321 26007 5355
rect 26341 5321 26375 5355
rect 2973 5253 3007 5287
rect 6653 5253 6687 5287
rect 10057 5253 10091 5287
rect 13921 5253 13955 5287
rect 16497 5253 16531 5287
rect 25053 5253 25087 5287
rect 2053 5185 2087 5219
rect 3617 5185 3651 5219
rect 4997 5185 5031 5219
rect 5733 5185 5767 5219
rect 6837 5185 6871 5219
rect 7389 5185 7423 5219
rect 8401 5185 8435 5219
rect 10977 5185 11011 5219
rect 11069 5185 11103 5219
rect 14473 5185 14507 5219
rect 15945 5185 15979 5219
rect 16037 5185 16071 5219
rect 18429 5185 18463 5219
rect 21925 5185 21959 5219
rect 23673 5185 23707 5219
rect 1869 5117 1903 5151
rect 3525 5117 3559 5151
rect 5549 5117 5583 5151
rect 9321 5117 9355 5151
rect 9413 5117 9447 5151
rect 10885 5117 10919 5151
rect 12265 5117 12299 5151
rect 12633 5117 12667 5151
rect 14381 5117 14415 5151
rect 15393 5117 15427 5151
rect 18889 5117 18923 5151
rect 23929 5117 23963 5151
rect 8309 5049 8343 5083
rect 12909 5049 12943 5083
rect 13829 5049 13863 5083
rect 14289 5049 14323 5083
rect 18797 5049 18831 5083
rect 19156 5049 19190 5083
rect 20913 5049 20947 5083
rect 21741 5049 21775 5083
rect 22385 5049 22419 5083
rect 23121 5049 23155 5083
rect 1961 4981 1995 5015
rect 2513 4981 2547 5015
rect 3433 4981 3467 5015
rect 5089 4981 5123 5015
rect 5457 4981 5491 5015
rect 7757 4981 7791 5015
rect 8217 4981 8251 5015
rect 9597 4981 9631 5015
rect 13461 4981 13495 5015
rect 15485 4981 15519 5015
rect 15853 4981 15887 5015
rect 16865 4981 16899 5015
rect 20269 4981 20303 5015
rect 21281 4981 21315 5015
rect 21833 4981 21867 5015
rect 1409 4777 1443 4811
rect 1777 4777 1811 4811
rect 1869 4777 1903 4811
rect 2421 4777 2455 4811
rect 6745 4777 6779 4811
rect 7389 4777 7423 4811
rect 9137 4777 9171 4811
rect 11161 4777 11195 4811
rect 11713 4777 11747 4811
rect 12357 4777 12391 4811
rect 12909 4777 12943 4811
rect 13001 4777 13035 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15853 4777 15887 4811
rect 17601 4777 17635 4811
rect 18245 4777 18279 4811
rect 19349 4777 19383 4811
rect 20729 4777 20763 4811
rect 21281 4777 21315 4811
rect 23489 4777 23523 4811
rect 24041 4777 24075 4811
rect 24501 4777 24535 4811
rect 25053 4777 25087 4811
rect 25421 4777 25455 4811
rect 3801 4709 3835 4743
rect 5610 4709 5644 4743
rect 8493 4709 8527 4743
rect 22017 4709 22051 4743
rect 22845 4709 22879 4743
rect 23949 4709 23983 4743
rect 4261 4641 4295 4675
rect 5365 4641 5399 4675
rect 8401 4641 8435 4675
rect 10048 4641 10082 4675
rect 14105 4641 14139 4675
rect 14657 4641 14691 4675
rect 16221 4641 16255 4675
rect 16488 4641 16522 4675
rect 19257 4641 19291 4675
rect 22385 4641 22419 4675
rect 22937 4641 22971 4675
rect 24409 4641 24443 4675
rect 1961 4573 1995 4607
rect 7941 4573 7975 4607
rect 8585 4573 8619 4607
rect 9781 4573 9815 4607
rect 13185 4573 13219 4607
rect 19441 4573 19475 4607
rect 21373 4573 21407 4607
rect 21465 4573 21499 4607
rect 23029 4573 23063 4607
rect 24685 4573 24719 4607
rect 3065 4505 3099 4539
rect 4905 4505 4939 4539
rect 3433 4437 3467 4471
rect 4445 4437 4479 4471
rect 8033 4437 8067 4471
rect 9505 4437 9539 4471
rect 12541 4437 12575 4471
rect 14289 4437 14323 4471
rect 15025 4437 15059 4471
rect 15577 4437 15611 4471
rect 18797 4437 18831 4471
rect 18889 4437 18923 4471
rect 19901 4437 19935 4471
rect 20269 4437 20303 4471
rect 20913 4437 20947 4471
rect 22477 4437 22511 4471
rect 1685 4233 1719 4267
rect 2053 4233 2087 4267
rect 4353 4233 4387 4267
rect 6285 4233 6319 4267
rect 9413 4233 9447 4267
rect 10793 4233 10827 4267
rect 15025 4233 15059 4267
rect 15485 4233 15519 4267
rect 16497 4233 16531 4267
rect 19073 4233 19107 4267
rect 20913 4233 20947 4267
rect 23029 4233 23063 4267
rect 25605 4233 25639 4267
rect 25973 4233 26007 4267
rect 26341 4233 26375 4267
rect 18061 4165 18095 4199
rect 2421 4097 2455 4131
rect 5457 4097 5491 4131
rect 7389 4097 7423 4131
rect 8125 4097 8159 4131
rect 8953 4097 8987 4131
rect 11345 4097 11379 4131
rect 12265 4097 12299 4131
rect 12725 4097 12759 4131
rect 15945 4097 15979 4131
rect 16037 4097 16071 4131
rect 16865 4097 16899 4131
rect 17233 4097 17267 4131
rect 18613 4097 18647 4131
rect 21005 4097 21039 4131
rect 23673 4097 23707 4131
rect 4813 4029 4847 4063
rect 8861 4029 8895 4063
rect 10241 4029 10275 4063
rect 11161 4029 11195 4063
rect 12992 4029 13026 4063
rect 15393 4029 15427 4063
rect 15853 4029 15887 4063
rect 19625 4029 19659 4063
rect 21272 4029 21306 4063
rect 2688 3961 2722 3995
rect 5273 3961 5307 3995
rect 6653 3961 6687 3995
rect 10701 3961 10735 3995
rect 11253 3961 11287 3995
rect 11805 3961 11839 3995
rect 18429 3961 18463 3995
rect 19901 3961 19935 3995
rect 23489 3961 23523 3995
rect 23918 3961 23952 3995
rect 3801 3893 3835 3927
rect 4905 3893 4939 3927
rect 5365 3893 5399 3927
rect 6837 3893 6871 3927
rect 7205 3893 7239 3927
rect 7297 3893 7331 3927
rect 8401 3893 8435 3927
rect 8769 3893 8803 3927
rect 9873 3893 9907 3927
rect 14105 3893 14139 3927
rect 17785 3893 17819 3927
rect 18521 3893 18555 3927
rect 19441 3893 19475 3927
rect 20453 3893 20487 3927
rect 22385 3893 22419 3927
rect 25053 3893 25087 3927
rect 1409 3689 1443 3723
rect 2421 3689 2455 3723
rect 4077 3689 4111 3723
rect 5089 3689 5123 3723
rect 5641 3689 5675 3723
rect 5825 3689 5859 3723
rect 6193 3689 6227 3723
rect 7389 3689 7423 3723
rect 9413 3689 9447 3723
rect 11069 3689 11103 3723
rect 11621 3689 11655 3723
rect 13001 3689 13035 3723
rect 13093 3689 13127 3723
rect 15301 3689 15335 3723
rect 15669 3689 15703 3723
rect 16865 3689 16899 3723
rect 17325 3689 17359 3723
rect 18153 3689 18187 3723
rect 19073 3689 19107 3723
rect 19165 3689 19199 3723
rect 20545 3689 20579 3723
rect 21189 3689 21223 3723
rect 23029 3689 23063 3723
rect 24133 3689 24167 3723
rect 24593 3689 24627 3723
rect 25145 3689 25179 3723
rect 25605 3689 25639 3723
rect 1869 3621 1903 3655
rect 4537 3621 4571 3655
rect 8401 3621 8435 3655
rect 9934 3621 9968 3655
rect 14197 3621 14231 3655
rect 14749 3621 14783 3655
rect 17233 3621 17267 3655
rect 1777 3553 1811 3587
rect 2973 3553 3007 3587
rect 4445 3553 4479 3587
rect 7757 3553 7791 3587
rect 7849 3553 7883 3587
rect 9137 3553 9171 3587
rect 12541 3553 12575 3587
rect 21649 3553 21683 3587
rect 21916 3553 21950 3587
rect 24501 3553 24535 3587
rect 2053 3485 2087 3519
rect 4721 3485 4755 3519
rect 6285 3485 6319 3519
rect 6377 3485 6411 3519
rect 7941 3485 7975 3519
rect 8861 3485 8895 3519
rect 9689 3485 9723 3519
rect 13277 3485 13311 3519
rect 13645 3485 13679 3519
rect 15025 3485 15059 3519
rect 15761 3485 15795 3519
rect 15945 3485 15979 3519
rect 17417 3485 17451 3519
rect 19349 3485 19383 3519
rect 24041 3485 24075 3519
rect 24685 3485 24719 3519
rect 3525 3417 3559 3451
rect 3893 3417 3927 3451
rect 6837 3417 6871 3451
rect 12173 3417 12207 3451
rect 16313 3417 16347 3451
rect 19717 3417 19751 3451
rect 21465 3417 21499 3451
rect 2881 3349 2915 3383
rect 7205 3349 7239 3383
rect 8953 3349 8987 3383
rect 12633 3349 12667 3383
rect 14013 3349 14047 3383
rect 16773 3349 16807 3383
rect 18521 3349 18555 3383
rect 18705 3349 18739 3383
rect 20177 3349 20211 3383
rect 23581 3349 23615 3383
rect 3433 3145 3467 3179
rect 5273 3145 5307 3179
rect 6561 3145 6595 3179
rect 8125 3145 8159 3179
rect 10793 3145 10827 3179
rect 12265 3145 12299 3179
rect 14105 3145 14139 3179
rect 16221 3145 16255 3179
rect 16681 3145 16715 3179
rect 19625 3145 19659 3179
rect 20361 3145 20395 3179
rect 20821 3145 20855 3179
rect 22293 3145 22327 3179
rect 23029 3145 23063 3179
rect 23673 3145 23707 3179
rect 26341 3145 26375 3179
rect 3709 3077 3743 3111
rect 16957 3077 16991 3111
rect 17693 3077 17727 3111
rect 3893 3009 3927 3043
rect 8309 3009 8343 3043
rect 10333 3009 10367 3043
rect 10609 3009 10643 3043
rect 11345 3009 11379 3043
rect 12725 3009 12759 3043
rect 15117 3009 15151 3043
rect 15669 3009 15703 3043
rect 15853 3009 15887 3043
rect 17325 3009 17359 3043
rect 24225 3009 24259 3043
rect 25421 3009 25455 3043
rect 1409 2941 1443 2975
rect 1676 2941 1710 2975
rect 4160 2941 4194 2975
rect 7021 2941 7055 2975
rect 8576 2941 8610 2975
rect 11897 2941 11931 2975
rect 12992 2941 13026 2975
rect 16773 2941 16807 2975
rect 18245 2941 18279 2975
rect 18512 2941 18546 2975
rect 20913 2941 20947 2975
rect 24133 2941 24167 2975
rect 25237 2941 25271 2975
rect 25973 2941 26007 2975
rect 5825 2873 5859 2907
rect 7297 2873 7331 2907
rect 14749 2873 14783 2907
rect 15577 2873 15611 2907
rect 21158 2873 21192 2907
rect 24777 2873 24811 2907
rect 2789 2805 2823 2839
rect 6193 2805 6227 2839
rect 7849 2805 7883 2839
rect 9689 2805 9723 2839
rect 11161 2805 11195 2839
rect 11253 2805 11287 2839
rect 15209 2805 15243 2839
rect 23489 2805 23523 2839
rect 24041 2805 24075 2839
rect 25145 2805 25179 2839
rect 1869 2601 1903 2635
rect 2237 2601 2271 2635
rect 2421 2601 2455 2635
rect 2881 2601 2915 2635
rect 4077 2601 4111 2635
rect 8401 2601 8435 2635
rect 10149 2601 10183 2635
rect 11161 2601 11195 2635
rect 12081 2601 12115 2635
rect 19901 2601 19935 2635
rect 20637 2601 20671 2635
rect 21281 2601 21315 2635
rect 21649 2601 21683 2635
rect 22293 2601 22327 2635
rect 22661 2601 22695 2635
rect 24041 2601 24075 2635
rect 24409 2601 24443 2635
rect 25513 2601 25547 2635
rect 3433 2533 3467 2567
rect 4445 2533 4479 2567
rect 7297 2533 7331 2567
rect 10241 2533 10275 2567
rect 12449 2533 12483 2567
rect 12878 2533 12912 2567
rect 19993 2533 20027 2567
rect 24501 2533 24535 2567
rect 25145 2533 25179 2567
rect 1409 2465 1443 2499
rect 2789 2465 2823 2499
rect 5733 2465 5767 2499
rect 7389 2465 7423 2499
rect 8585 2465 8619 2499
rect 10793 2465 10827 2499
rect 11437 2465 11471 2499
rect 12633 2465 12667 2499
rect 14841 2465 14875 2499
rect 15853 2465 15887 2499
rect 17049 2465 17083 2499
rect 17601 2465 17635 2499
rect 21005 2465 21039 2499
rect 25605 2465 25639 2499
rect 3065 2397 3099 2431
rect 4537 2397 4571 2431
rect 4721 2397 4755 2431
rect 5549 2397 5583 2431
rect 6745 2397 6779 2431
rect 7573 2397 7607 2431
rect 7941 2397 7975 2431
rect 9229 2397 9263 2431
rect 9597 2397 9631 2431
rect 10333 2397 10367 2431
rect 15209 2397 15243 2431
rect 15945 2397 15979 2431
rect 16037 2397 16071 2431
rect 16497 2397 16531 2431
rect 16865 2397 16899 2431
rect 19073 2397 19107 2431
rect 19441 2397 19475 2431
rect 20177 2397 20211 2431
rect 21741 2397 21775 2431
rect 21925 2397 21959 2431
rect 24685 2397 24719 2431
rect 5089 2329 5123 2363
rect 5917 2329 5951 2363
rect 9781 2329 9815 2363
rect 17233 2329 17267 2363
rect 19533 2329 19567 2363
rect 3801 2261 3835 2295
rect 6285 2261 6319 2295
rect 6929 2261 6963 2295
rect 8769 2261 8803 2295
rect 11621 2261 11655 2295
rect 14013 2261 14047 2295
rect 15485 2261 15519 2295
rect 17969 2261 18003 2295
rect 18613 2261 18647 2295
rect 23029 2261 23063 2295
rect 23673 2261 23707 2295
<< metal1 >>
rect 4062 26256 4068 26308
rect 4120 26296 4126 26308
rect 22462 26296 22468 26308
rect 4120 26268 22468 26296
rect 4120 26256 4126 26268
rect 22462 26256 22468 26268
rect 22520 26256 22526 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 3326 24828 3332 24880
rect 3384 24868 3390 24880
rect 7006 24868 7012 24880
rect 3384 24840 7012 24868
rect 3384 24828 3390 24840
rect 7006 24828 7012 24840
rect 7064 24828 7070 24880
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 22646 23848 22652 23860
rect 22607 23820 22652 23848
rect 22646 23808 22652 23820
rect 22704 23808 22710 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 1854 23644 1860 23656
rect 1443 23616 1860 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 1854 23604 1860 23616
rect 1912 23644 1918 23656
rect 1949 23647 2007 23653
rect 1949 23644 1961 23647
rect 1912 23616 1961 23644
rect 1912 23604 1918 23616
rect 1949 23613 1961 23616
rect 1995 23613 2007 23647
rect 22462 23644 22468 23656
rect 22423 23616 22468 23644
rect 1949 23607 2007 23613
rect 22462 23604 22468 23616
rect 22520 23644 22526 23656
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22520 23616 23029 23644
rect 22520 23604 22526 23616
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 24578 23644 24584 23656
rect 24539 23616 24584 23644
rect 23017 23607 23075 23613
rect 24578 23604 24584 23616
rect 24636 23644 24642 23656
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24636 23616 25145 23644
rect 24636 23604 24642 23616
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1486 23264 1492 23316
rect 1544 23304 1550 23316
rect 1581 23307 1639 23313
rect 1581 23304 1593 23307
rect 1544 23276 1593 23304
rect 1544 23264 1550 23276
rect 1581 23273 1593 23276
rect 1627 23273 1639 23307
rect 1581 23267 1639 23273
rect 19797 23239 19855 23245
rect 19797 23205 19809 23239
rect 19843 23236 19855 23239
rect 20622 23236 20628 23248
rect 19843 23208 20628 23236
rect 19843 23205 19855 23208
rect 19797 23199 19855 23205
rect 20622 23196 20628 23208
rect 20680 23196 20686 23248
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2498 23168 2504 23180
rect 1443 23140 2504 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2498 23128 2504 23140
rect 2556 23128 2562 23180
rect 19518 23168 19524 23180
rect 19479 23140 19524 23168
rect 19518 23128 19524 23140
rect 19576 23128 19582 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 1673 22559 1731 22565
rect 1673 22525 1685 22559
rect 1719 22556 1731 22559
rect 2222 22556 2228 22568
rect 1719 22528 2228 22556
rect 1719 22525 1731 22528
rect 1673 22519 1731 22525
rect 2222 22516 2228 22528
rect 2280 22516 2286 22568
rect 2498 22420 2504 22432
rect 2459 22392 2504 22420
rect 2498 22380 2504 22392
rect 2556 22380 2562 22432
rect 19518 22420 19524 22432
rect 19479 22392 19524 22420
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1397 22083 1455 22089
rect 1397 22049 1409 22083
rect 1443 22080 1455 22083
rect 2406 22080 2412 22092
rect 1443 22052 2412 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 2406 22040 2412 22052
rect 2464 22040 2470 22092
rect 1394 21904 1400 21956
rect 1452 21944 1458 21956
rect 1581 21947 1639 21953
rect 1581 21944 1593 21947
rect 1452 21916 1593 21944
rect 1452 21904 1458 21916
rect 1581 21913 1593 21916
rect 1627 21913 1639 21947
rect 1581 21907 1639 21913
rect 2041 21879 2099 21885
rect 2041 21845 2053 21879
rect 2087 21876 2099 21879
rect 2222 21876 2228 21888
rect 2087 21848 2228 21876
rect 2087 21845 2099 21848
rect 2041 21839 2099 21845
rect 2222 21836 2228 21848
rect 2280 21836 2286 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 1443 21440 2084 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2056 21344 2084 21440
rect 23934 21428 23940 21480
rect 23992 21468 23998 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 23992 21440 24593 21468
rect 23992 21428 23998 21440
rect 24581 21437 24593 21440
rect 24627 21468 24639 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24627 21440 25145 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 2038 21332 2044 21344
rect 1999 21304 2044 21332
rect 2038 21292 2044 21304
rect 2096 21292 2102 21344
rect 2406 21332 2412 21344
rect 2367 21304 2412 21332
rect 2406 21292 2412 21304
rect 2464 21292 2470 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1486 21088 1492 21140
rect 1544 21128 1550 21140
rect 1581 21131 1639 21137
rect 1581 21128 1593 21131
rect 1544 21100 1593 21128
rect 1544 21088 1550 21100
rect 1581 21097 1593 21100
rect 1627 21097 1639 21131
rect 4614 21128 4620 21140
rect 4575 21100 4620 21128
rect 1581 21091 1639 21097
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 23934 21060 23940 21072
rect 23895 21032 23940 21060
rect 23934 21020 23940 21032
rect 23992 21020 23998 21072
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 2314 20992 2320 21004
rect 1443 20964 2320 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 2314 20952 2320 20964
rect 2372 20952 2378 21004
rect 4430 20992 4436 21004
rect 4391 20964 4436 20992
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 23661 20995 23719 21001
rect 23661 20961 23673 20995
rect 23707 20992 23719 20995
rect 23842 20992 23848 21004
rect 23707 20964 23848 20992
rect 23707 20961 23719 20964
rect 23661 20955 23719 20961
rect 23842 20952 23848 20964
rect 23900 20952 23906 21004
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 24670 20544 24676 20596
rect 24728 20584 24734 20596
rect 24765 20587 24823 20593
rect 24765 20584 24777 20587
rect 24728 20556 24777 20584
rect 24728 20544 24734 20556
rect 24765 20553 24777 20556
rect 24811 20553 24823 20587
rect 24765 20547 24823 20553
rect 4430 20408 4436 20460
rect 4488 20448 4494 20460
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 4488 20420 4537 20448
rect 4488 20408 4494 20420
rect 4525 20417 4537 20420
rect 4571 20448 4583 20451
rect 5353 20451 5411 20457
rect 5353 20448 5365 20451
rect 4571 20420 5365 20448
rect 4571 20417 4583 20420
rect 4525 20411 4583 20417
rect 5353 20417 5365 20420
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20349 1455 20383
rect 1397 20343 1455 20349
rect 2041 20383 2099 20389
rect 2041 20349 2053 20383
rect 2087 20380 2099 20383
rect 2314 20380 2320 20392
rect 2087 20352 2320 20380
rect 2087 20349 2099 20352
rect 2041 20343 2099 20349
rect 1412 20312 1440 20343
rect 2314 20340 2320 20352
rect 2372 20340 2378 20392
rect 5169 20383 5227 20389
rect 5169 20349 5181 20383
rect 5215 20380 5227 20383
rect 24578 20380 24584 20392
rect 5215 20352 6040 20380
rect 24539 20352 24584 20380
rect 5215 20349 5227 20352
rect 5169 20343 5227 20349
rect 1412 20284 2452 20312
rect 2424 20256 2452 20284
rect 2406 20244 2412 20256
rect 2367 20216 2412 20244
rect 2406 20204 2412 20216
rect 2464 20204 2470 20256
rect 6012 20253 6040 20352
rect 24578 20340 24584 20352
rect 24636 20380 24642 20392
rect 25133 20383 25191 20389
rect 25133 20380 25145 20383
rect 24636 20352 25145 20380
rect 24636 20340 24642 20352
rect 25133 20349 25145 20352
rect 25179 20349 25191 20383
rect 25133 20343 25191 20349
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6086 20244 6092 20256
rect 6043 20216 6092 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6086 20204 6092 20216
rect 6144 20204 6150 20256
rect 23842 20244 23848 20256
rect 23803 20216 23848 20244
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 2682 20040 2688 20052
rect 2643 20012 2688 20040
rect 2682 20000 2688 20012
rect 2740 20000 2746 20052
rect 24762 20040 24768 20052
rect 24723 20012 24768 20040
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2406 19904 2412 19916
rect 1443 19876 2412 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2406 19864 2412 19876
rect 2464 19864 2470 19916
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19904 2559 19907
rect 2682 19904 2688 19916
rect 2547 19876 2688 19904
rect 2547 19873 2559 19876
rect 2501 19867 2559 19873
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 24581 19907 24639 19913
rect 24581 19873 24593 19907
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19836 23627 19839
rect 23934 19836 23940 19848
rect 23615 19808 23940 19836
rect 23615 19805 23627 19808
rect 23569 19799 23627 19805
rect 23934 19796 23940 19808
rect 23992 19796 23998 19848
rect 23842 19728 23848 19780
rect 23900 19768 23906 19780
rect 24596 19768 24624 19867
rect 23900 19740 24624 19768
rect 23900 19728 23906 19740
rect 1946 19700 1952 19712
rect 1907 19672 1952 19700
rect 1946 19660 1952 19672
rect 2004 19660 2010 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 2498 19292 2504 19304
rect 1443 19264 2084 19292
rect 2459 19264 2504 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 2056 19168 2084 19264
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 2682 19252 2688 19304
rect 2740 19292 2746 19304
rect 3053 19295 3111 19301
rect 3053 19292 3065 19295
rect 2740 19264 3065 19292
rect 2740 19252 2746 19264
rect 3053 19261 3065 19264
rect 3099 19292 3111 19295
rect 9214 19292 9220 19304
rect 3099 19264 9220 19292
rect 3099 19261 3111 19264
rect 3053 19255 3111 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 17402 19252 17408 19304
rect 17460 19292 17466 19304
rect 18141 19295 18199 19301
rect 18141 19292 18153 19295
rect 17460 19264 18153 19292
rect 17460 19252 17466 19264
rect 18141 19261 18153 19264
rect 18187 19292 18199 19295
rect 18693 19295 18751 19301
rect 18693 19292 18705 19295
rect 18187 19264 18705 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 18693 19261 18705 19264
rect 18739 19261 18751 19295
rect 24578 19292 24584 19304
rect 24539 19264 24584 19292
rect 18693 19255 18751 19261
rect 24578 19252 24584 19264
rect 24636 19292 24642 19304
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24636 19264 25145 19292
rect 24636 19252 24642 19264
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 2038 19156 2044 19168
rect 1999 19128 2044 19156
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 2406 19156 2412 19168
rect 2367 19128 2412 19156
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 2590 19116 2596 19168
rect 2648 19156 2654 19168
rect 2685 19159 2743 19165
rect 2685 19156 2697 19159
rect 2648 19128 2697 19156
rect 2648 19116 2654 19128
rect 2685 19125 2697 19128
rect 2731 19125 2743 19159
rect 18322 19156 18328 19168
rect 18283 19128 18328 19156
rect 2685 19119 2743 19125
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 22557 19159 22615 19165
rect 22557 19125 22569 19159
rect 22603 19156 22615 19159
rect 23014 19156 23020 19168
rect 22603 19128 23020 19156
rect 22603 19125 22615 19128
rect 22557 19119 22615 19125
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 23842 19116 23848 19168
rect 23900 19156 23906 19168
rect 24397 19159 24455 19165
rect 24397 19156 24409 19159
rect 23900 19128 24409 19156
rect 23900 19116 23906 19128
rect 24397 19125 24409 19128
rect 24443 19125 24455 19159
rect 24762 19156 24768 19168
rect 24723 19128 24768 19156
rect 24397 19119 24455 19125
rect 24762 19116 24768 19128
rect 24820 19116 24826 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 4246 18952 4252 18964
rect 4207 18924 4252 18952
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 24670 18912 24676 18964
rect 24728 18952 24734 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 24728 18924 24777 18952
rect 24728 18912 24734 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 17402 18884 17408 18896
rect 17363 18856 17408 18884
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 1489 18819 1547 18825
rect 1489 18785 1501 18819
rect 1535 18816 1547 18819
rect 1670 18816 1676 18828
rect 1535 18788 1676 18816
rect 1535 18785 1547 18788
rect 1489 18779 1547 18785
rect 1670 18776 1676 18788
rect 1728 18776 1734 18828
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 4062 18816 4068 18828
rect 2832 18788 2877 18816
rect 4023 18788 4068 18816
rect 2832 18776 2838 18788
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 17126 18816 17132 18828
rect 17087 18788 17132 18816
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 22370 18816 22376 18828
rect 22331 18788 22376 18816
rect 22370 18776 22376 18788
rect 22428 18776 22434 18828
rect 23474 18816 23480 18828
rect 23435 18788 23480 18816
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 24578 18816 24584 18828
rect 24539 18788 24584 18816
rect 24578 18776 24584 18788
rect 24636 18776 24642 18828
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 2866 18748 2872 18760
rect 1811 18720 2872 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 22557 18683 22615 18689
rect 22557 18649 22569 18683
rect 22603 18680 22615 18683
rect 25958 18680 25964 18692
rect 22603 18652 25964 18680
rect 22603 18649 22615 18652
rect 22557 18643 22615 18649
rect 25958 18640 25964 18652
rect 26016 18640 26022 18692
rect 2590 18612 2596 18624
rect 2551 18584 2596 18612
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 23661 18615 23719 18621
rect 23661 18581 23673 18615
rect 23707 18612 23719 18615
rect 24762 18612 24768 18624
rect 23707 18584 24768 18612
rect 23707 18581 23719 18584
rect 23661 18575 23719 18581
rect 24762 18572 24768 18584
rect 24820 18572 24826 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 24670 18368 24676 18420
rect 24728 18408 24734 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 24728 18380 24869 18408
rect 24728 18368 24734 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 24857 18371 24915 18377
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 2774 18272 2780 18284
rect 1719 18244 2780 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 2774 18232 2780 18244
rect 2832 18272 2838 18284
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2832 18244 2881 18272
rect 2832 18232 2838 18244
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 3973 18275 4031 18281
rect 3973 18241 3985 18275
rect 4019 18272 4031 18275
rect 4062 18272 4068 18284
rect 4019 18244 4068 18272
rect 4019 18241 4031 18244
rect 3973 18235 4031 18241
rect 4062 18232 4068 18244
rect 4120 18272 4126 18284
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4120 18244 4445 18272
rect 4120 18232 4126 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 23842 18232 23848 18284
rect 23900 18272 23906 18284
rect 24670 18272 24676 18284
rect 23900 18244 24676 18272
rect 23900 18232 23906 18244
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 1394 18204 1400 18216
rect 1307 18176 1400 18204
rect 1394 18164 1400 18176
rect 1452 18204 1458 18216
rect 1946 18204 1952 18216
rect 1452 18176 1952 18204
rect 1452 18164 1458 18176
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 3697 18207 3755 18213
rect 3697 18173 3709 18207
rect 3743 18173 3755 18207
rect 3697 18167 3755 18173
rect 1670 18096 1676 18148
rect 1728 18136 1734 18148
rect 2501 18139 2559 18145
rect 2501 18136 2513 18139
rect 1728 18108 2513 18136
rect 1728 18096 1734 18108
rect 2501 18105 2513 18108
rect 2547 18105 2559 18139
rect 2501 18099 2559 18105
rect 2130 18068 2136 18080
rect 2091 18040 2136 18068
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 3712 18068 3740 18167
rect 20714 18164 20720 18216
rect 20772 18204 20778 18216
rect 21361 18207 21419 18213
rect 21361 18204 21373 18207
rect 20772 18176 21373 18204
rect 20772 18164 20778 18176
rect 21361 18173 21373 18176
rect 21407 18204 21419 18207
rect 21913 18207 21971 18213
rect 21913 18204 21925 18207
rect 21407 18176 21925 18204
rect 21407 18173 21419 18176
rect 21361 18167 21419 18173
rect 21913 18173 21925 18176
rect 21959 18173 21971 18207
rect 21913 18167 21971 18173
rect 22281 18207 22339 18213
rect 22281 18173 22293 18207
rect 22327 18204 22339 18207
rect 22465 18207 22523 18213
rect 22465 18204 22477 18207
rect 22327 18176 22477 18204
rect 22327 18173 22339 18176
rect 22281 18167 22339 18173
rect 22465 18173 22477 18176
rect 22511 18204 22523 18207
rect 22922 18204 22928 18216
rect 22511 18176 22928 18204
rect 22511 18173 22523 18176
rect 22465 18167 22523 18173
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 24305 18207 24363 18213
rect 24305 18204 24317 18207
rect 24136 18176 24317 18204
rect 22370 18096 22376 18148
rect 22428 18136 22434 18148
rect 23109 18139 23167 18145
rect 23109 18136 23121 18139
rect 22428 18108 23121 18136
rect 22428 18096 22434 18108
rect 23109 18105 23121 18108
rect 23155 18136 23167 18139
rect 23382 18136 23388 18148
rect 23155 18108 23388 18136
rect 23155 18105 23167 18108
rect 23109 18099 23167 18105
rect 23382 18096 23388 18108
rect 23440 18096 23446 18148
rect 4062 18068 4068 18080
rect 3651 18040 4068 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 17126 18068 17132 18080
rect 16356 18040 17132 18068
rect 16356 18028 16362 18040
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19484 18040 19625 18068
rect 19484 18028 19490 18040
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 21542 18068 21548 18080
rect 21503 18040 21548 18068
rect 19613 18031 19671 18037
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 22646 18068 22652 18080
rect 22607 18040 22652 18068
rect 22646 18028 22652 18040
rect 22704 18028 22710 18080
rect 23474 18068 23480 18080
rect 23435 18040 23480 18068
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 23842 18028 23848 18080
rect 23900 18068 23906 18080
rect 24136 18077 24164 18176
rect 24305 18173 24317 18176
rect 24351 18173 24363 18207
rect 24305 18167 24363 18173
rect 25409 18207 25467 18213
rect 25409 18173 25421 18207
rect 25455 18204 25467 18207
rect 25455 18176 26096 18204
rect 25455 18173 25467 18176
rect 25409 18167 25467 18173
rect 24121 18071 24179 18077
rect 24121 18068 24133 18071
rect 23900 18040 24133 18068
rect 23900 18028 23906 18040
rect 24121 18037 24133 18040
rect 24167 18037 24179 18071
rect 24486 18068 24492 18080
rect 24447 18040 24492 18068
rect 24121 18031 24179 18037
rect 24486 18028 24492 18040
rect 24544 18028 24550 18080
rect 25590 18068 25596 18080
rect 25551 18040 25596 18068
rect 25590 18028 25596 18040
rect 25648 18028 25654 18080
rect 26068 18077 26096 18176
rect 26053 18071 26111 18077
rect 26053 18037 26065 18071
rect 26099 18068 26111 18071
rect 26142 18068 26148 18080
rect 26099 18040 26148 18068
rect 26099 18037 26111 18040
rect 26053 18031 26111 18037
rect 26142 18028 26148 18040
rect 26200 18028 26206 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 5353 17867 5411 17873
rect 5353 17864 5365 17867
rect 4212 17836 5365 17864
rect 4212 17824 4218 17836
rect 5353 17833 5365 17836
rect 5399 17833 5411 17867
rect 5353 17827 5411 17833
rect 23750 17824 23756 17876
rect 23808 17864 23814 17876
rect 24765 17867 24823 17873
rect 24765 17864 24777 17867
rect 23808 17836 24777 17864
rect 23808 17824 23814 17836
rect 24765 17833 24777 17836
rect 24811 17833 24823 17867
rect 24765 17827 24823 17833
rect 1949 17799 2007 17805
rect 1949 17765 1961 17799
rect 1995 17796 2007 17799
rect 2498 17796 2504 17808
rect 1995 17768 2504 17796
rect 1995 17765 2007 17768
rect 1949 17759 2007 17765
rect 2498 17756 2504 17768
rect 2556 17756 2562 17808
rect 19518 17756 19524 17808
rect 19576 17796 19582 17808
rect 20622 17796 20628 17808
rect 19576 17768 20628 17796
rect 19576 17756 19582 17768
rect 20622 17756 20628 17768
rect 20680 17756 20686 17808
rect 1854 17728 1860 17740
rect 1767 17700 1860 17728
rect 1854 17688 1860 17700
rect 1912 17728 1918 17740
rect 2774 17728 2780 17740
rect 1912 17700 2780 17728
rect 1912 17688 1918 17700
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 2866 17688 2872 17740
rect 2924 17728 2930 17740
rect 3970 17728 3976 17740
rect 2924 17700 3976 17728
rect 2924 17688 2930 17700
rect 3970 17688 3976 17700
rect 4028 17728 4034 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 4028 17700 4077 17728
rect 4028 17688 4034 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4982 17688 4988 17740
rect 5040 17728 5046 17740
rect 5169 17731 5227 17737
rect 5169 17728 5181 17731
rect 5040 17700 5181 17728
rect 5040 17688 5046 17700
rect 5169 17697 5181 17700
rect 5215 17697 5227 17731
rect 5169 17691 5227 17697
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 19613 17731 19671 17737
rect 19613 17728 19625 17731
rect 19392 17700 19625 17728
rect 19392 17688 19398 17700
rect 19613 17697 19625 17700
rect 19659 17697 19671 17731
rect 21266 17728 21272 17740
rect 21227 17700 21272 17728
rect 19613 17691 19671 17697
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 22373 17731 22431 17737
rect 22373 17697 22385 17731
rect 22419 17728 22431 17731
rect 22462 17728 22468 17740
rect 22419 17700 22468 17728
rect 22419 17697 22431 17700
rect 22373 17691 22431 17697
rect 22462 17688 22468 17700
rect 22520 17688 22526 17740
rect 23477 17731 23535 17737
rect 23477 17697 23489 17731
rect 23523 17728 23535 17731
rect 23566 17728 23572 17740
rect 23523 17700 23572 17728
rect 23523 17697 23535 17700
rect 23477 17691 23535 17697
rect 23566 17688 23572 17700
rect 23624 17688 23630 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 25130 17728 25136 17740
rect 24627 17700 25136 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 25130 17688 25136 17700
rect 25188 17688 25194 17740
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 17402 17660 17408 17672
rect 17363 17632 17408 17660
rect 17402 17620 17408 17632
rect 17460 17620 17466 17672
rect 19702 17660 19708 17672
rect 19663 17632 19708 17660
rect 19702 17620 19708 17632
rect 19760 17620 19766 17672
rect 19886 17660 19892 17672
rect 19847 17632 19892 17660
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 26510 17660 26516 17672
rect 21468 17632 26516 17660
rect 21468 17601 21496 17632
rect 26510 17620 26516 17632
rect 26568 17620 26574 17672
rect 4617 17595 4675 17601
rect 4617 17592 4629 17595
rect 3712 17564 4629 17592
rect 3712 17536 3740 17564
rect 4617 17561 4629 17564
rect 4663 17561 4675 17595
rect 4617 17555 4675 17561
rect 21453 17595 21511 17601
rect 21453 17561 21465 17595
rect 21499 17561 21511 17595
rect 22554 17592 22560 17604
rect 22515 17564 22560 17592
rect 21453 17555 21511 17561
rect 22554 17552 22560 17564
rect 22612 17552 22618 17604
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 2406 17524 2412 17536
rect 1820 17496 2412 17524
rect 1820 17484 1826 17496
rect 2406 17484 2412 17496
rect 2464 17524 2470 17536
rect 2501 17527 2559 17533
rect 2501 17524 2513 17527
rect 2464 17496 2513 17524
rect 2464 17484 2470 17496
rect 2501 17493 2513 17496
rect 2547 17493 2559 17527
rect 2501 17487 2559 17493
rect 2866 17484 2872 17536
rect 2924 17524 2930 17536
rect 2961 17527 3019 17533
rect 2961 17524 2973 17527
rect 2924 17496 2973 17524
rect 2924 17484 2930 17496
rect 2961 17493 2973 17496
rect 3007 17493 3019 17527
rect 3326 17524 3332 17536
rect 3287 17496 3332 17524
rect 2961 17487 3019 17493
rect 3326 17484 3332 17496
rect 3384 17484 3390 17536
rect 3694 17524 3700 17536
rect 3655 17496 3700 17524
rect 3694 17484 3700 17496
rect 3752 17484 3758 17536
rect 4246 17524 4252 17536
rect 4207 17496 4252 17524
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 19058 17524 19064 17536
rect 19019 17496 19064 17524
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 19242 17524 19248 17536
rect 19203 17496 19248 17524
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 20346 17524 20352 17536
rect 20307 17496 20352 17524
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20622 17524 20628 17536
rect 20583 17496 20628 17524
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 21910 17524 21916 17536
rect 21871 17496 21916 17524
rect 21910 17484 21916 17496
rect 21968 17484 21974 17536
rect 23661 17527 23719 17533
rect 23661 17493 23673 17527
rect 23707 17524 23719 17527
rect 23842 17524 23848 17536
rect 23707 17496 23848 17524
rect 23707 17493 23719 17496
rect 23661 17487 23719 17493
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 3970 17320 3976 17332
rect 2832 17292 2877 17320
rect 3931 17292 3976 17320
rect 2832 17280 2838 17292
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 16022 17320 16028 17332
rect 15983 17292 16028 17320
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 18598 17320 18604 17332
rect 17552 17292 18604 17320
rect 17552 17280 17558 17292
rect 18598 17280 18604 17292
rect 18656 17320 18662 17332
rect 18785 17323 18843 17329
rect 18785 17320 18797 17323
rect 18656 17292 18797 17320
rect 18656 17280 18662 17292
rect 18785 17289 18797 17292
rect 18831 17320 18843 17323
rect 19886 17320 19892 17332
rect 18831 17292 19892 17320
rect 18831 17289 18843 17292
rect 18785 17283 18843 17289
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 21266 17320 21272 17332
rect 21227 17292 21272 17320
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 24118 17280 24124 17332
rect 24176 17320 24182 17332
rect 24765 17323 24823 17329
rect 24765 17320 24777 17323
rect 24176 17292 24777 17320
rect 24176 17280 24182 17292
rect 24765 17289 24777 17292
rect 24811 17289 24823 17323
rect 24765 17283 24823 17289
rect 19702 17252 19708 17264
rect 19663 17224 19708 17252
rect 19702 17212 19708 17224
rect 19760 17252 19766 17264
rect 20530 17252 20536 17264
rect 19760 17224 20536 17252
rect 19760 17212 19766 17224
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 2041 17187 2099 17193
rect 2041 17153 2053 17187
rect 2087 17184 2099 17187
rect 2130 17184 2136 17196
rect 2087 17156 2136 17184
rect 2087 17153 2099 17156
rect 2041 17147 2099 17153
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3513 17187 3571 17193
rect 3513 17184 3525 17187
rect 2924 17156 3525 17184
rect 2924 17144 2930 17156
rect 3513 17153 3525 17156
rect 3559 17153 3571 17187
rect 20438 17184 20444 17196
rect 20399 17156 20444 17184
rect 3513 17147 3571 17153
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 21910 17184 21916 17196
rect 21871 17156 21916 17184
rect 21910 17144 21916 17156
rect 21968 17144 21974 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 4525 17119 4583 17125
rect 4525 17116 4537 17119
rect 4356 17088 4537 17116
rect 1946 17048 1952 17060
rect 1412 17020 1952 17048
rect 1412 16989 1440 17020
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 3421 17051 3479 17057
rect 3421 17048 3433 17051
rect 3200 17020 3433 17048
rect 3200 17008 3206 17020
rect 3421 17017 3433 17020
rect 3467 17017 3479 17051
rect 3421 17011 3479 17017
rect 4356 16992 4384 17088
rect 4525 17085 4537 17088
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 5258 17116 5264 17128
rect 4847 17088 5264 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 15838 17116 15844 17128
rect 15799 17088 15844 17116
rect 15838 17076 15844 17088
rect 15896 17116 15902 17128
rect 16393 17119 16451 17125
rect 16393 17116 16405 17119
rect 15896 17088 16405 17116
rect 15896 17076 15902 17088
rect 16393 17085 16405 17088
rect 16439 17085 16451 17119
rect 19334 17116 19340 17128
rect 19295 17088 19340 17116
rect 16393 17079 16451 17085
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 20257 17119 20315 17125
rect 20257 17085 20269 17119
rect 20303 17116 20315 17119
rect 20622 17116 20628 17128
rect 20303 17088 20628 17116
rect 20303 17085 20315 17088
rect 20257 17079 20315 17085
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 22020 17116 22048 17147
rect 20916 17088 22048 17116
rect 24581 17119 24639 17125
rect 20916 16992 20944 17088
rect 24581 17085 24593 17119
rect 24627 17085 24639 17119
rect 24581 17079 24639 17085
rect 20990 17008 20996 17060
rect 21048 17048 21054 17060
rect 24397 17051 24455 17057
rect 24397 17048 24409 17051
rect 21048 17020 24409 17048
rect 21048 17008 21054 17020
rect 24397 17017 24409 17020
rect 24443 17048 24455 17051
rect 24596 17048 24624 17079
rect 24443 17020 24624 17048
rect 24443 17017 24455 17020
rect 24397 17011 24455 17017
rect 1397 16983 1455 16989
rect 1397 16949 1409 16983
rect 1443 16949 1455 16983
rect 1397 16943 1455 16949
rect 1857 16983 1915 16989
rect 1857 16949 1869 16983
rect 1903 16980 1915 16983
rect 2314 16980 2320 16992
rect 1903 16952 2320 16980
rect 1903 16949 1915 16952
rect 1857 16943 1915 16949
rect 2314 16940 2320 16952
rect 2372 16940 2378 16992
rect 2498 16980 2504 16992
rect 2459 16952 2504 16980
rect 2498 16940 2504 16952
rect 2556 16940 2562 16992
rect 2958 16980 2964 16992
rect 2919 16952 2964 16980
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 3326 16980 3332 16992
rect 3287 16952 3332 16980
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 4338 16980 4344 16992
rect 4299 16952 4344 16980
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 5261 16983 5319 16989
rect 5261 16980 5273 16983
rect 5040 16952 5273 16980
rect 5040 16940 5046 16952
rect 5261 16949 5273 16952
rect 5307 16949 5319 16983
rect 5261 16943 5319 16949
rect 16758 16940 16764 16992
rect 16816 16980 16822 16992
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16816 16952 16957 16980
rect 16816 16940 16822 16952
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 18874 16980 18880 16992
rect 18835 16952 18880 16980
rect 16945 16943 17003 16949
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 19889 16983 19947 16989
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20162 16980 20168 16992
rect 19935 16952 20168 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 20898 16980 20904 16992
rect 20859 16952 20904 16980
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 21358 16940 21364 16992
rect 21416 16980 21422 16992
rect 21453 16983 21511 16989
rect 21453 16980 21465 16983
rect 21416 16952 21465 16980
rect 21416 16940 21422 16952
rect 21453 16949 21465 16952
rect 21499 16949 21511 16983
rect 21818 16980 21824 16992
rect 21779 16952 21824 16980
rect 21453 16943 21511 16949
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 22554 16980 22560 16992
rect 22515 16952 22560 16980
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 23566 16940 23572 16992
rect 23624 16980 23630 16992
rect 23845 16983 23903 16989
rect 23845 16980 23857 16983
rect 23624 16952 23857 16980
rect 23624 16940 23630 16952
rect 23845 16949 23857 16952
rect 23891 16949 23903 16983
rect 25130 16980 25136 16992
rect 25091 16952 25136 16980
rect 23845 16943 23903 16949
rect 25130 16940 25136 16952
rect 25188 16940 25194 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1946 16736 1952 16788
rect 2004 16776 2010 16788
rect 2130 16776 2136 16788
rect 2004 16748 2136 16776
rect 2004 16736 2010 16748
rect 2130 16736 2136 16748
rect 2188 16736 2194 16788
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 2593 16779 2651 16785
rect 2593 16776 2605 16779
rect 2372 16748 2605 16776
rect 2372 16736 2378 16748
rect 2593 16745 2605 16748
rect 2639 16776 2651 16779
rect 2639 16748 3096 16776
rect 2639 16745 2651 16748
rect 2593 16739 2651 16745
rect 2148 16708 2176 16736
rect 3068 16708 3096 16748
rect 3142 16736 3148 16788
rect 3200 16776 3206 16788
rect 3237 16779 3295 16785
rect 3237 16776 3249 16779
rect 3200 16748 3249 16776
rect 3200 16736 3206 16748
rect 3237 16745 3249 16748
rect 3283 16745 3295 16779
rect 5534 16776 5540 16788
rect 5495 16748 5540 16776
rect 3237 16739 3295 16745
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 7650 16776 7656 16788
rect 7116 16748 7656 16776
rect 5166 16708 5172 16720
rect 2148 16680 2636 16708
rect 3068 16680 5172 16708
rect 937 16643 995 16649
rect 937 16609 949 16643
rect 983 16640 995 16643
rect 1857 16643 1915 16649
rect 1857 16640 1869 16643
rect 983 16612 1869 16640
rect 983 16609 995 16612
rect 937 16603 995 16609
rect 1857 16609 1869 16612
rect 1903 16609 1915 16643
rect 1857 16603 1915 16609
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2314 16640 2320 16652
rect 1995 16612 2320 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 2608 16640 2636 16680
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 6457 16711 6515 16717
rect 6457 16677 6469 16711
rect 6503 16708 6515 16711
rect 7116 16708 7144 16748
rect 7650 16736 7656 16748
rect 7708 16776 7714 16788
rect 7929 16779 7987 16785
rect 7929 16776 7941 16779
rect 7708 16748 7941 16776
rect 7708 16736 7714 16748
rect 7929 16745 7941 16748
rect 7975 16745 7987 16779
rect 7929 16739 7987 16745
rect 17405 16779 17463 16785
rect 17405 16745 17417 16779
rect 17451 16776 17463 16779
rect 17494 16776 17500 16788
rect 17451 16748 17500 16776
rect 17451 16745 17463 16748
rect 17405 16739 17463 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16776 18659 16779
rect 19058 16776 19064 16788
rect 18647 16748 19064 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 19058 16736 19064 16748
rect 19116 16736 19122 16788
rect 19245 16779 19303 16785
rect 19245 16745 19257 16779
rect 19291 16776 19303 16779
rect 20346 16776 20352 16788
rect 19291 16748 20352 16776
rect 19291 16745 19303 16748
rect 19245 16739 19303 16745
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 20901 16779 20959 16785
rect 20901 16776 20913 16779
rect 20680 16748 20913 16776
rect 20680 16736 20686 16748
rect 20901 16745 20913 16748
rect 20947 16745 20959 16779
rect 20901 16739 20959 16745
rect 21818 16736 21824 16788
rect 21876 16776 21882 16788
rect 21913 16779 21971 16785
rect 21913 16776 21925 16779
rect 21876 16748 21925 16776
rect 21876 16736 21882 16748
rect 21913 16745 21925 16748
rect 21959 16776 21971 16779
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 21959 16748 22477 16776
rect 21959 16745 21971 16748
rect 21913 16739 21971 16745
rect 22465 16745 22477 16748
rect 22511 16745 22523 16779
rect 22465 16739 22523 16745
rect 23753 16779 23811 16785
rect 23753 16745 23765 16779
rect 23799 16776 23811 16779
rect 24026 16776 24032 16788
rect 23799 16748 24032 16776
rect 23799 16745 23811 16748
rect 23753 16739 23811 16745
rect 24026 16736 24032 16748
rect 24084 16736 24090 16788
rect 25501 16779 25559 16785
rect 25501 16745 25513 16779
rect 25547 16776 25559 16779
rect 25682 16776 25688 16788
rect 25547 16748 25688 16776
rect 25547 16745 25559 16748
rect 25501 16739 25559 16745
rect 25682 16736 25688 16748
rect 25740 16736 25746 16788
rect 6503 16680 7144 16708
rect 6503 16677 6515 16680
rect 6457 16671 6515 16677
rect 7190 16668 7196 16720
rect 7248 16708 7254 16720
rect 7377 16711 7435 16717
rect 7377 16708 7389 16711
rect 7248 16680 7389 16708
rect 7248 16668 7254 16680
rect 7377 16677 7389 16680
rect 7423 16677 7435 16711
rect 7377 16671 7435 16677
rect 16206 16668 16212 16720
rect 16264 16717 16270 16720
rect 16264 16711 16328 16717
rect 16264 16677 16282 16711
rect 16316 16677 16328 16711
rect 22278 16708 22284 16720
rect 22239 16680 22284 16708
rect 16264 16671 16328 16677
rect 16264 16668 16270 16671
rect 22278 16668 22284 16680
rect 22336 16668 22342 16720
rect 22554 16668 22560 16720
rect 22612 16708 22618 16720
rect 24305 16711 24363 16717
rect 24305 16708 24317 16711
rect 22612 16680 24317 16708
rect 22612 16668 22618 16680
rect 24305 16677 24317 16680
rect 24351 16677 24363 16711
rect 24305 16671 24363 16677
rect 3605 16643 3663 16649
rect 3605 16640 3617 16643
rect 2608 16612 3617 16640
rect 3605 16609 3617 16612
rect 3651 16609 3663 16643
rect 3605 16603 3663 16609
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4341 16643 4399 16649
rect 4341 16609 4353 16643
rect 4387 16640 4399 16643
rect 5350 16640 5356 16652
rect 4387 16612 5356 16640
rect 4387 16609 4399 16612
rect 4341 16603 4399 16609
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16572 2102 16584
rect 2682 16572 2688 16584
rect 2096 16544 2688 16572
rect 2096 16532 2102 16544
rect 2682 16532 2688 16544
rect 2740 16572 2746 16584
rect 2869 16575 2927 16581
rect 2869 16572 2881 16575
rect 2740 16544 2881 16572
rect 2740 16532 2746 16544
rect 2869 16541 2881 16544
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 4080 16504 4108 16603
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 6822 16640 6828 16652
rect 6735 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16640 6886 16652
rect 7285 16643 7343 16649
rect 7285 16640 7297 16643
rect 6880 16612 7297 16640
rect 6880 16600 6886 16612
rect 7285 16609 7297 16612
rect 7331 16609 7343 16643
rect 7285 16603 7343 16609
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13354 16640 13360 16652
rect 13311 16612 13360 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 19613 16643 19671 16649
rect 19613 16640 19625 16643
rect 19576 16612 19625 16640
rect 19576 16600 19582 16612
rect 19613 16609 19625 16612
rect 19659 16609 19671 16643
rect 19613 16603 19671 16609
rect 20349 16643 20407 16649
rect 20349 16609 20361 16643
rect 20395 16640 20407 16643
rect 20438 16640 20444 16652
rect 20395 16612 20444 16640
rect 20395 16609 20407 16612
rect 20349 16603 20407 16609
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 21266 16640 21272 16652
rect 21227 16612 21272 16640
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21361 16643 21419 16649
rect 21361 16609 21373 16643
rect 21407 16640 21419 16643
rect 21542 16640 21548 16652
rect 21407 16612 21548 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 22830 16640 22836 16652
rect 22791 16612 22836 16640
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 24029 16643 24087 16649
rect 24029 16609 24041 16643
rect 24075 16640 24087 16643
rect 24118 16640 24124 16652
rect 24075 16612 24124 16640
rect 24075 16609 24087 16612
rect 24029 16603 24087 16609
rect 24118 16600 24124 16612
rect 24176 16640 24182 16652
rect 24765 16643 24823 16649
rect 24765 16640 24777 16643
rect 24176 16612 24777 16640
rect 24176 16600 24182 16612
rect 24765 16609 24777 16612
rect 24811 16609 24823 16643
rect 24765 16603 24823 16609
rect 25317 16643 25375 16649
rect 25317 16609 25329 16643
rect 25363 16640 25375 16643
rect 25774 16640 25780 16652
rect 25363 16612 25780 16640
rect 25363 16609 25375 16612
rect 25317 16603 25375 16609
rect 25774 16600 25780 16612
rect 25832 16600 25838 16652
rect 7558 16572 7564 16584
rect 7471 16544 7564 16572
rect 7558 16532 7564 16544
rect 7616 16572 7622 16584
rect 9030 16572 9036 16584
rect 7616 16544 9036 16572
rect 7616 16532 7622 16544
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 16022 16572 16028 16584
rect 15983 16544 16028 16572
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 19334 16532 19340 16584
rect 19392 16572 19398 16584
rect 19705 16575 19763 16581
rect 19705 16572 19717 16575
rect 19392 16544 19717 16572
rect 19392 16532 19398 16544
rect 19705 16541 19717 16544
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 4801 16507 4859 16513
rect 4801 16504 4813 16507
rect 2648 16476 4813 16504
rect 2648 16464 2654 16476
rect 4801 16473 4813 16476
rect 4847 16473 4859 16507
rect 4801 16467 4859 16473
rect 1489 16439 1547 16445
rect 1489 16405 1501 16439
rect 1535 16436 1547 16439
rect 1946 16436 1952 16448
rect 1535 16408 1952 16436
rect 1535 16405 1547 16408
rect 1489 16399 1547 16405
rect 1946 16396 1952 16408
rect 2004 16396 2010 16448
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3694 16436 3700 16448
rect 3292 16408 3700 16436
rect 3292 16396 3298 16408
rect 3694 16396 3700 16408
rect 3752 16436 3758 16448
rect 5169 16439 5227 16445
rect 5169 16436 5181 16439
rect 3752 16408 5181 16436
rect 3752 16396 3758 16408
rect 5169 16405 5181 16408
rect 5215 16436 5227 16439
rect 5905 16439 5963 16445
rect 5905 16436 5917 16439
rect 5215 16408 5917 16436
rect 5215 16405 5227 16408
rect 5169 16399 5227 16405
rect 5905 16405 5917 16408
rect 5951 16436 5963 16439
rect 6270 16436 6276 16448
rect 5951 16408 6276 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16436 18291 16439
rect 18782 16436 18788 16448
rect 18279 16408 18788 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 18782 16396 18788 16408
rect 18840 16436 18846 16448
rect 19153 16439 19211 16445
rect 19153 16436 19165 16439
rect 18840 16408 19165 16436
rect 18840 16396 18846 16408
rect 19153 16405 19165 16408
rect 19199 16436 19211 16439
rect 19904 16436 19932 16535
rect 20898 16532 20904 16584
rect 20956 16572 20962 16584
rect 21453 16575 21511 16581
rect 21453 16572 21465 16575
rect 20956 16544 21465 16572
rect 20956 16532 20962 16544
rect 21453 16541 21465 16544
rect 21499 16541 21511 16575
rect 21453 16535 21511 16541
rect 22370 16532 22376 16584
rect 22428 16572 22434 16584
rect 22925 16575 22983 16581
rect 22925 16572 22937 16575
rect 22428 16544 22937 16572
rect 22428 16532 22434 16544
rect 22925 16541 22937 16544
rect 22971 16541 22983 16575
rect 22925 16535 22983 16541
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16541 23075 16575
rect 23017 16535 23075 16541
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 23032 16504 23060 16535
rect 24210 16504 24216 16516
rect 22336 16476 24216 16504
rect 22336 16464 22342 16476
rect 24210 16464 24216 16476
rect 24268 16464 24274 16516
rect 19978 16436 19984 16448
rect 19199 16408 19984 16436
rect 19199 16405 19211 16408
rect 19153 16399 19211 16405
rect 19978 16396 19984 16408
rect 20036 16436 20042 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20036 16408 20637 16436
rect 20036 16396 20042 16408
rect 20625 16405 20637 16408
rect 20671 16436 20683 16439
rect 20898 16436 20904 16448
rect 20671 16408 20904 16436
rect 20671 16405 20683 16408
rect 20625 16399 20683 16405
rect 20898 16396 20904 16408
rect 20956 16396 20962 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2409 16235 2467 16241
rect 2409 16232 2421 16235
rect 2372 16204 2421 16232
rect 2372 16192 2378 16204
rect 2409 16201 2421 16204
rect 2455 16232 2467 16235
rect 3418 16232 3424 16244
rect 2455 16204 3424 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 5350 16232 5356 16244
rect 5311 16204 5356 16232
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 5813 16235 5871 16241
rect 5813 16201 5825 16235
rect 5859 16232 5871 16235
rect 5994 16232 6000 16244
rect 5859 16204 6000 16232
rect 5859 16201 5871 16204
rect 5813 16195 5871 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 7558 16232 7564 16244
rect 7147 16204 7564 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 9030 16232 9036 16244
rect 8991 16204 9036 16232
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 16117 16235 16175 16241
rect 16117 16201 16129 16235
rect 16163 16232 16175 16235
rect 16206 16232 16212 16244
rect 16163 16204 16212 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16206 16192 16212 16204
rect 16264 16192 16270 16244
rect 22370 16232 22376 16244
rect 22331 16204 22376 16232
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 22649 16235 22707 16241
rect 22649 16201 22661 16235
rect 22695 16232 22707 16235
rect 22738 16232 22744 16244
rect 22695 16204 22744 16232
rect 22695 16201 22707 16204
rect 22649 16195 22707 16201
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 23658 16232 23664 16244
rect 23619 16204 23664 16232
rect 23658 16192 23664 16204
rect 23716 16192 23722 16244
rect 25406 16232 25412 16244
rect 25367 16204 25412 16232
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 1397 16167 1455 16173
rect 1397 16133 1409 16167
rect 1443 16164 1455 16167
rect 2038 16164 2044 16176
rect 1443 16136 2044 16164
rect 1443 16133 1455 16136
rect 1397 16127 1455 16133
rect 2038 16124 2044 16136
rect 2096 16124 2102 16176
rect 1854 16096 1860 16108
rect 1688 16068 1860 16096
rect 1688 16040 1716 16068
rect 1854 16056 1860 16068
rect 1912 16056 1918 16108
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16096 2007 16099
rect 2314 16096 2320 16108
rect 1995 16068 2320 16096
rect 1995 16065 2007 16068
rect 1949 16059 2007 16065
rect 2314 16056 2320 16068
rect 2372 16096 2378 16108
rect 2866 16096 2872 16108
rect 2372 16068 2872 16096
rect 2372 16056 2378 16068
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 7650 16096 7656 16108
rect 7611 16068 7656 16096
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 14274 16096 14280 16108
rect 13771 16068 14280 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 15197 16099 15255 16105
rect 15197 16065 15209 16099
rect 15243 16096 15255 16099
rect 15838 16096 15844 16108
rect 15243 16068 15844 16096
rect 15243 16065 15255 16068
rect 15197 16059 15255 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 18782 16096 18788 16108
rect 18743 16068 18788 16096
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 19058 16056 19064 16108
rect 19116 16096 19122 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19116 16068 19717 16096
rect 19116 16056 19122 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 1670 15988 1676 16040
rect 1728 15988 1734 16040
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 2130 16028 2136 16040
rect 1811 16000 2136 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 2130 15988 2136 16000
rect 2188 15988 2194 16040
rect 3145 16031 3203 16037
rect 3145 15997 3157 16031
rect 3191 16028 3203 16031
rect 3234 16028 3240 16040
rect 3191 16000 3240 16028
rect 3191 15997 3203 16000
rect 3145 15991 3203 15997
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 13081 16031 13139 16037
rect 5675 16000 6316 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 937 15963 995 15969
rect 937 15929 949 15963
rect 983 15960 995 15963
rect 2777 15963 2835 15969
rect 2777 15960 2789 15963
rect 983 15932 2789 15960
rect 983 15929 995 15932
rect 937 15923 995 15929
rect 2777 15929 2789 15932
rect 2823 15929 2835 15963
rect 2777 15923 2835 15929
rect 3412 15963 3470 15969
rect 3412 15929 3424 15963
rect 3458 15960 3470 15963
rect 3510 15960 3516 15972
rect 3458 15932 3516 15960
rect 3458 15929 3470 15932
rect 3412 15923 3470 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 1486 15852 1492 15904
rect 1544 15892 1550 15904
rect 1854 15892 1860 15904
rect 1544 15864 1860 15892
rect 1544 15852 1550 15864
rect 1854 15852 1860 15864
rect 1912 15852 1918 15904
rect 2130 15852 2136 15904
rect 2188 15892 2194 15904
rect 2498 15892 2504 15904
rect 2188 15864 2504 15892
rect 2188 15852 2194 15864
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 4338 15852 4344 15904
rect 4396 15892 4402 15904
rect 6288 15901 6316 16000
rect 13081 15997 13093 16031
rect 13127 16028 13139 16031
rect 13538 16028 13544 16040
rect 13127 16000 13544 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 13872 16000 14933 16028
rect 13872 15988 13878 16000
rect 14921 15997 14933 16000
rect 14967 16028 14979 16031
rect 15657 16031 15715 16037
rect 15657 16028 15669 16031
rect 14967 16000 15669 16028
rect 14967 15997 14979 16000
rect 14921 15991 14979 15997
rect 15657 15997 15669 16000
rect 15703 15997 15715 16031
rect 15657 15991 15715 15997
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 16028 17555 16031
rect 18601 16031 18659 16037
rect 18601 16028 18613 16031
rect 17543 16000 18613 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 18601 15997 18613 16000
rect 18647 16028 18659 16031
rect 19242 16028 19248 16040
rect 18647 16000 19248 16028
rect 18647 15997 18659 16000
rect 18601 15991 18659 15997
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 19720 16028 19748 16059
rect 21542 16056 21548 16108
rect 21600 16096 21606 16108
rect 21637 16099 21695 16105
rect 21637 16096 21649 16099
rect 21600 16068 21649 16096
rect 21600 16056 21606 16068
rect 21637 16065 21649 16068
rect 21683 16096 21695 16099
rect 21683 16068 22508 16096
rect 21683 16065 21695 16068
rect 21637 16059 21695 16065
rect 21082 16028 21088 16040
rect 19720 16000 21088 16028
rect 21082 15988 21088 16000
rect 21140 15988 21146 16040
rect 22480 16037 22508 16068
rect 24026 16056 24032 16108
rect 24084 16056 24090 16108
rect 24210 16096 24216 16108
rect 24171 16068 24216 16096
rect 24210 16056 24216 16068
rect 24268 16096 24274 16108
rect 24673 16099 24731 16105
rect 24673 16096 24685 16099
rect 24268 16068 24685 16096
rect 24268 16056 24274 16068
rect 24673 16065 24685 16068
rect 24719 16065 24731 16099
rect 24673 16059 24731 16065
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 16028 22523 16031
rect 23017 16031 23075 16037
rect 23017 16028 23029 16031
rect 22511 16000 23029 16028
rect 22511 15997 22523 16000
rect 22465 15991 22523 15997
rect 23017 15997 23029 16000
rect 23063 15997 23075 16031
rect 24044 16028 24072 16056
rect 24121 16031 24179 16037
rect 24121 16028 24133 16031
rect 24044 16000 24133 16028
rect 23017 15991 23075 15997
rect 24121 15997 24133 16000
rect 24167 15997 24179 16031
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 24121 15991 24179 15997
rect 25056 16000 25237 16028
rect 7098 15920 7104 15972
rect 7156 15960 7162 15972
rect 7469 15963 7527 15969
rect 7469 15960 7481 15963
rect 7156 15932 7481 15960
rect 7156 15920 7162 15932
rect 7469 15929 7481 15932
rect 7515 15960 7527 15963
rect 7898 15963 7956 15969
rect 7898 15960 7910 15963
rect 7515 15932 7910 15960
rect 7515 15929 7527 15932
rect 7469 15923 7527 15929
rect 7898 15929 7910 15932
rect 7944 15929 7956 15963
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 7898 15923 7956 15929
rect 12728 15932 13645 15960
rect 12728 15904 12756 15932
rect 13633 15929 13645 15932
rect 13679 15929 13691 15963
rect 18509 15963 18567 15969
rect 18509 15960 18521 15963
rect 13633 15923 13691 15929
rect 17788 15932 18521 15960
rect 17788 15904 17816 15932
rect 18509 15929 18521 15932
rect 18555 15929 18567 15963
rect 18509 15923 18567 15929
rect 19972 15963 20030 15969
rect 19972 15929 19984 15963
rect 20018 15960 20030 15963
rect 20254 15960 20260 15972
rect 20018 15932 20260 15960
rect 20018 15929 20030 15932
rect 19972 15923 20030 15929
rect 20254 15920 20260 15932
rect 20312 15920 20318 15972
rect 23477 15963 23535 15969
rect 23477 15929 23489 15963
rect 23523 15960 23535 15963
rect 24029 15963 24087 15969
rect 24029 15960 24041 15963
rect 23523 15932 24041 15960
rect 23523 15929 23535 15932
rect 23477 15923 23535 15929
rect 24029 15929 24041 15932
rect 24075 15960 24087 15963
rect 24670 15960 24676 15972
rect 24075 15932 24676 15960
rect 24075 15929 24087 15932
rect 24029 15923 24087 15929
rect 24670 15920 24676 15932
rect 24728 15920 24734 15972
rect 4525 15895 4583 15901
rect 4525 15892 4537 15895
rect 4396 15864 4537 15892
rect 4396 15852 4402 15864
rect 4525 15861 4537 15864
rect 4571 15861 4583 15895
rect 4525 15855 4583 15861
rect 6273 15895 6331 15901
rect 6273 15861 6285 15895
rect 6319 15892 6331 15895
rect 6362 15892 6368 15904
rect 6319 15864 6368 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7190 15892 7196 15904
rect 6687 15864 7196 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 11054 15892 11060 15904
rect 11015 15864 11060 15892
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 12710 15892 12716 15904
rect 12671 15864 12716 15892
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 13173 15895 13231 15901
rect 13173 15861 13185 15895
rect 13219 15892 13231 15895
rect 13262 15892 13268 15904
rect 13219 15864 13268 15892
rect 13219 15861 13231 15864
rect 13173 15855 13231 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 13538 15892 13544 15904
rect 13499 15864 13544 15892
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 14274 15892 14280 15904
rect 14235 15864 14280 15892
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 16485 15895 16543 15901
rect 16485 15892 16497 15895
rect 16264 15864 16497 15892
rect 16264 15852 16270 15864
rect 16485 15861 16497 15864
rect 16531 15861 16543 15895
rect 17034 15892 17040 15904
rect 16995 15864 17040 15892
rect 16485 15855 16543 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 17770 15892 17776 15904
rect 17731 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 18141 15895 18199 15901
rect 18141 15861 18153 15895
rect 18187 15892 18199 15895
rect 19150 15892 19156 15904
rect 18187 15864 19156 15892
rect 18187 15861 18199 15864
rect 18141 15855 18199 15861
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 19337 15895 19395 15901
rect 19337 15861 19349 15895
rect 19383 15892 19395 15895
rect 19518 15892 19524 15904
rect 19383 15864 19524 15892
rect 19383 15861 19395 15864
rect 19337 15855 19395 15861
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 21085 15895 21143 15901
rect 21085 15861 21097 15895
rect 21131 15892 21143 15895
rect 21174 15892 21180 15904
rect 21131 15864 21180 15892
rect 21131 15861 21143 15864
rect 21085 15855 21143 15861
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 24946 15852 24952 15904
rect 25004 15892 25010 15904
rect 25056 15901 25084 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 25041 15895 25099 15901
rect 25041 15892 25053 15895
rect 25004 15864 25053 15892
rect 25004 15852 25010 15864
rect 25041 15861 25053 15864
rect 25087 15861 25099 15895
rect 25774 15892 25780 15904
rect 25735 15864 25780 15892
rect 25041 15855 25099 15861
rect 25774 15852 25780 15864
rect 25832 15852 25838 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 3605 15691 3663 15697
rect 3605 15688 3617 15691
rect 1912 15660 3617 15688
rect 1912 15648 1918 15660
rect 3605 15657 3617 15660
rect 3651 15657 3663 15691
rect 4338 15688 4344 15700
rect 4299 15660 4344 15688
rect 3605 15651 3663 15657
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 4985 15691 5043 15697
rect 4985 15657 4997 15691
rect 5031 15688 5043 15691
rect 5074 15688 5080 15700
rect 5031 15660 5080 15688
rect 5031 15657 5043 15660
rect 4985 15651 5043 15657
rect 2682 15580 2688 15632
rect 2740 15620 2746 15632
rect 2740 15592 3004 15620
rect 2740 15580 2746 15592
rect 1854 15552 1860 15564
rect 1815 15524 1860 15552
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 1946 15512 1952 15564
rect 2004 15552 2010 15564
rect 2774 15552 2780 15564
rect 2004 15524 2780 15552
rect 2004 15512 2010 15524
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2314 15484 2320 15496
rect 2087 15456 2320 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 1946 15376 1952 15428
rect 2004 15416 2010 15428
rect 2056 15416 2084 15447
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 2976 15425 3004 15592
rect 3694 15580 3700 15632
rect 3752 15620 3758 15632
rect 5000 15620 5028 15651
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 6270 15688 6276 15700
rect 6231 15660 6276 15688
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 6638 15688 6644 15700
rect 6599 15660 6644 15688
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 6822 15688 6828 15700
rect 6783 15660 6828 15688
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7650 15648 7656 15700
rect 7708 15688 7714 15700
rect 8205 15691 8263 15697
rect 8205 15688 8217 15691
rect 7708 15660 8217 15688
rect 7708 15648 7714 15660
rect 8205 15657 8217 15660
rect 8251 15688 8263 15691
rect 8849 15691 8907 15697
rect 8849 15688 8861 15691
rect 8251 15660 8861 15688
rect 8251 15657 8263 15660
rect 8205 15651 8263 15657
rect 8849 15657 8861 15660
rect 8895 15688 8907 15691
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 8895 15660 9229 15688
rect 8895 15657 8907 15660
rect 8849 15651 8907 15657
rect 9217 15657 9229 15660
rect 9263 15688 9275 15691
rect 10134 15688 10140 15700
rect 9263 15660 10140 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 19889 15691 19947 15697
rect 12584 15660 15608 15688
rect 12584 15648 12590 15660
rect 3752 15592 5028 15620
rect 6656 15620 6684 15648
rect 7285 15623 7343 15629
rect 7285 15620 7297 15623
rect 6656 15592 7297 15620
rect 3752 15580 3758 15592
rect 7285 15589 7297 15592
rect 7331 15589 7343 15623
rect 7285 15583 7343 15589
rect 13541 15623 13599 15629
rect 13541 15589 13553 15623
rect 13587 15620 13599 15623
rect 13722 15620 13728 15632
rect 13587 15592 13728 15620
rect 13587 15589 13599 15592
rect 13541 15583 13599 15589
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 15580 15629 15608 15660
rect 19889 15657 19901 15691
rect 19935 15688 19947 15691
rect 20070 15688 20076 15700
rect 19935 15660 20076 15688
rect 19935 15657 19947 15660
rect 19889 15651 19947 15657
rect 20070 15648 20076 15660
rect 20128 15648 20134 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 21266 15688 21272 15700
rect 20763 15660 21272 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 22557 15691 22615 15697
rect 22557 15657 22569 15691
rect 22603 15657 22615 15691
rect 22557 15651 22615 15657
rect 15565 15623 15623 15629
rect 15565 15589 15577 15623
rect 15611 15589 15623 15623
rect 22572 15620 22600 15651
rect 23906 15623 23964 15629
rect 23906 15620 23918 15623
rect 22572 15592 23918 15620
rect 15565 15583 15623 15589
rect 23906 15589 23918 15592
rect 23952 15620 23964 15623
rect 24210 15620 24216 15632
rect 23952 15592 24216 15620
rect 23952 15589 23964 15592
rect 23906 15583 23964 15589
rect 24210 15580 24216 15592
rect 24268 15580 24274 15632
rect 4893 15555 4951 15561
rect 4893 15521 4905 15555
rect 4939 15552 4951 15555
rect 5074 15552 5080 15564
rect 4939 15524 5080 15552
rect 4939 15521 4951 15524
rect 4893 15515 4951 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 5534 15552 5540 15564
rect 5495 15524 5540 15552
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 6822 15512 6828 15564
rect 6880 15552 6886 15564
rect 10962 15561 10968 15564
rect 7193 15555 7251 15561
rect 7193 15552 7205 15555
rect 6880 15524 7205 15552
rect 6880 15512 6886 15524
rect 7193 15521 7205 15524
rect 7239 15552 7251 15555
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 7239 15524 8401 15552
rect 7239 15521 7251 15524
rect 7193 15515 7251 15521
rect 8389 15521 8401 15524
rect 8435 15521 8447 15555
rect 10956 15552 10968 15561
rect 10923 15524 10968 15552
rect 8389 15515 8447 15521
rect 10956 15515 10968 15524
rect 10962 15512 10968 15515
rect 11020 15512 11026 15564
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 15286 15552 15292 15564
rect 13127 15524 13860 15552
rect 15247 15524 15292 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 5169 15487 5227 15493
rect 3099 15456 3740 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 2004 15388 2084 15416
rect 2961 15419 3019 15425
rect 2004 15376 2010 15388
rect 2961 15385 2973 15419
rect 3007 15416 3019 15419
rect 3602 15416 3608 15428
rect 3007 15388 3608 15416
rect 3007 15385 3019 15388
rect 2961 15379 3019 15385
rect 3602 15376 3608 15388
rect 3660 15376 3666 15428
rect 3712 15416 3740 15456
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5442 15484 5448 15496
rect 5215 15456 5448 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7377 15487 7435 15493
rect 7377 15484 7389 15487
rect 7156 15456 7389 15484
rect 7156 15444 7162 15456
rect 7377 15453 7389 15456
rect 7423 15453 7435 15487
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 7377 15447 7435 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10520 15456 10701 15484
rect 5905 15419 5963 15425
rect 5905 15416 5917 15419
rect 3712 15388 5917 15416
rect 5905 15385 5917 15388
rect 5951 15385 5963 15419
rect 5905 15379 5963 15385
rect 6270 15376 6276 15428
rect 6328 15416 6334 15428
rect 7837 15419 7895 15425
rect 7837 15416 7849 15419
rect 6328 15388 7849 15416
rect 6328 15376 6334 15388
rect 7837 15385 7849 15388
rect 7883 15416 7895 15419
rect 9030 15416 9036 15428
rect 7883 15388 9036 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 9030 15376 9036 15388
rect 9088 15376 9094 15428
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 2593 15351 2651 15357
rect 2593 15317 2605 15351
rect 2639 15348 2651 15351
rect 2682 15348 2688 15360
rect 2639 15320 2688 15348
rect 2639 15317 2651 15320
rect 2593 15311 2651 15317
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 3053 15351 3111 15357
rect 3053 15348 3065 15351
rect 2924 15320 3065 15348
rect 2924 15308 2930 15320
rect 3053 15317 3065 15320
rect 3099 15317 3111 15351
rect 3053 15311 3111 15317
rect 3329 15351 3387 15357
rect 3329 15317 3341 15351
rect 3375 15348 3387 15351
rect 3510 15348 3516 15360
rect 3375 15320 3516 15348
rect 3375 15317 3387 15320
rect 3329 15311 3387 15317
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 4525 15351 4583 15357
rect 4525 15348 4537 15351
rect 4396 15320 4537 15348
rect 4396 15308 4402 15320
rect 4525 15317 4537 15320
rect 4571 15317 4583 15351
rect 10134 15348 10140 15360
rect 10095 15320 10140 15348
rect 4525 15311 4583 15317
rect 10134 15308 10140 15320
rect 10192 15348 10198 15360
rect 10520 15357 10548 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 13446 15444 13452 15496
rect 13504 15484 13510 15496
rect 13832 15493 13860 15524
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 17293 15555 17351 15561
rect 17293 15552 17305 15555
rect 16724 15524 17305 15552
rect 16724 15512 16730 15524
rect 17293 15521 17305 15524
rect 17339 15521 17351 15555
rect 17293 15515 17351 15521
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 20346 15552 20352 15564
rect 19751 15524 20352 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 20346 15512 20352 15524
rect 20404 15512 20410 15564
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21177 15555 21235 15561
rect 21177 15552 21189 15555
rect 21140 15524 21189 15552
rect 21140 15512 21146 15524
rect 21177 15521 21189 15524
rect 21223 15521 21235 15555
rect 21177 15515 21235 15521
rect 21266 15512 21272 15564
rect 21324 15552 21330 15564
rect 21433 15555 21491 15561
rect 21433 15552 21445 15555
rect 21324 15524 21445 15552
rect 21324 15512 21330 15524
rect 21433 15521 21445 15524
rect 21479 15521 21491 15555
rect 21433 15515 21491 15521
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13504 15456 13645 15484
rect 13504 15444 13510 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13817 15487 13875 15493
rect 13817 15453 13829 15487
rect 13863 15484 13875 15487
rect 14274 15484 14280 15496
rect 13863 15456 14280 15484
rect 13863 15453 13875 15456
rect 13817 15447 13875 15453
rect 14274 15444 14280 15456
rect 14332 15444 14338 15496
rect 17034 15484 17040 15496
rect 16868 15456 17040 15484
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 13173 15419 13231 15425
rect 13173 15416 13185 15419
rect 12308 15388 13185 15416
rect 12308 15376 12314 15388
rect 13173 15385 13185 15388
rect 13219 15385 13231 15419
rect 13173 15379 13231 15385
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 10192 15320 10517 15348
rect 10192 15308 10198 15320
rect 10505 15317 10517 15320
rect 10551 15317 10563 15351
rect 10505 15311 10563 15317
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 12434 15348 12440 15360
rect 12115 15320 12440 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 12434 15308 12440 15320
rect 12492 15348 12498 15360
rect 12621 15351 12679 15357
rect 12621 15348 12633 15351
rect 12492 15320 12633 15348
rect 12492 15308 12498 15320
rect 12621 15317 12633 15320
rect 12667 15317 12679 15351
rect 12621 15311 12679 15317
rect 14277 15351 14335 15357
rect 14277 15317 14289 15351
rect 14323 15348 14335 15351
rect 14645 15351 14703 15357
rect 14645 15348 14657 15351
rect 14323 15320 14657 15348
rect 14323 15317 14335 15320
rect 14277 15311 14335 15317
rect 14645 15317 14657 15320
rect 14691 15348 14703 15351
rect 14826 15348 14832 15360
rect 14691 15320 14832 15348
rect 14691 15317 14703 15320
rect 14645 15311 14703 15317
rect 14826 15308 14832 15320
rect 14884 15348 14890 15360
rect 15013 15351 15071 15357
rect 15013 15348 15025 15351
rect 14884 15320 15025 15348
rect 14884 15308 14890 15320
rect 15013 15317 15025 15320
rect 15059 15348 15071 15351
rect 16022 15348 16028 15360
rect 15059 15320 16028 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 16022 15308 16028 15320
rect 16080 15348 16086 15360
rect 16868 15357 16896 15456
rect 17034 15444 17040 15456
rect 17092 15444 17098 15496
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 23676 15360 23704 15447
rect 16853 15351 16911 15357
rect 16853 15348 16865 15351
rect 16080 15320 16865 15348
rect 16080 15308 16086 15320
rect 16853 15317 16865 15320
rect 16899 15317 16911 15351
rect 16853 15311 16911 15317
rect 18417 15351 18475 15357
rect 18417 15317 18429 15351
rect 18463 15348 18475 15351
rect 18506 15348 18512 15360
rect 18463 15320 18512 15348
rect 18463 15317 18475 15320
rect 18417 15311 18475 15317
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 19334 15348 19340 15360
rect 19295 15320 19340 15348
rect 19334 15308 19340 15320
rect 19392 15308 19398 15360
rect 20254 15348 20260 15360
rect 20215 15320 20260 15348
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 22094 15308 22100 15360
rect 22152 15348 22158 15360
rect 22830 15348 22836 15360
rect 22152 15320 22836 15348
rect 22152 15308 22158 15320
rect 22830 15308 22836 15320
rect 22888 15348 22894 15360
rect 23109 15351 23167 15357
rect 23109 15348 23121 15351
rect 22888 15320 23121 15348
rect 22888 15308 22894 15320
rect 23109 15317 23121 15320
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 23569 15351 23627 15357
rect 23569 15317 23581 15351
rect 23615 15348 23627 15351
rect 23658 15348 23664 15360
rect 23615 15320 23664 15348
rect 23615 15317 23627 15320
rect 23569 15311 23627 15317
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 24854 15308 24860 15360
rect 24912 15348 24918 15360
rect 25041 15351 25099 15357
rect 25041 15348 25053 15351
rect 24912 15320 25053 15348
rect 24912 15308 24918 15320
rect 25041 15317 25053 15320
rect 25087 15317 25099 15351
rect 25041 15311 25099 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1578 15144 1584 15156
rect 1539 15116 1584 15144
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2590 15144 2596 15156
rect 2547 15116 2596 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2590 15104 2596 15116
rect 2648 15104 2654 15156
rect 3694 15144 3700 15156
rect 3655 15116 3700 15144
rect 3694 15104 3700 15116
rect 3752 15104 3758 15156
rect 5442 15104 5448 15156
rect 5500 15144 5506 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 5500 15116 6193 15144
rect 5500 15104 5506 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 6181 15107 6239 15113
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 6822 15144 6828 15156
rect 6687 15116 6828 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7006 15144 7012 15156
rect 6967 15116 7012 15144
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 16209 15147 16267 15153
rect 16209 15144 16221 15147
rect 15344 15116 16221 15144
rect 15344 15104 15350 15116
rect 16209 15113 16221 15116
rect 16255 15113 16267 15147
rect 18966 15144 18972 15156
rect 16209 15107 16267 15113
rect 18248 15116 18972 15144
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2314 15008 2320 15020
rect 2087 14980 2320 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 2056 14940 2084 14971
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 2682 14968 2688 15020
rect 2740 15008 2746 15020
rect 3145 15011 3203 15017
rect 3145 15008 3157 15011
rect 2740 14980 3157 15008
rect 2740 14968 2746 14980
rect 3145 14977 3157 14980
rect 3191 15008 3203 15011
rect 3191 14980 4384 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 4356 14952 4384 14980
rect 7650 14968 7656 15020
rect 7708 15008 7714 15020
rect 8021 15011 8079 15017
rect 8021 15008 8033 15011
rect 7708 14980 8033 15008
rect 7708 14968 7714 14980
rect 8021 14977 8033 14980
rect 8067 14977 8079 15011
rect 10594 15008 10600 15020
rect 10555 14980 10600 15008
rect 8021 14971 8079 14977
rect 10594 14968 10600 14980
rect 10652 15008 10658 15020
rect 11241 15011 11299 15017
rect 11241 15008 11253 15011
rect 10652 14980 11253 15008
rect 10652 14968 10658 14980
rect 11241 14977 11253 14980
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 11425 15011 11483 15017
rect 11425 14977 11437 15011
rect 11471 15008 11483 15011
rect 12434 15008 12440 15020
rect 11471 14980 12440 15008
rect 11471 14977 11483 14980
rect 11425 14971 11483 14977
rect 12434 14968 12440 14980
rect 12492 15008 12498 15020
rect 18248 15017 18276 15116
rect 18966 15104 18972 15116
rect 19024 15144 19030 15156
rect 19518 15144 19524 15156
rect 19024 15116 19524 15144
rect 19024 15104 19030 15116
rect 19518 15104 19524 15116
rect 19576 15104 19582 15156
rect 19613 15079 19671 15085
rect 19613 15045 19625 15079
rect 19659 15076 19671 15079
rect 20254 15076 20260 15088
rect 19659 15048 20260 15076
rect 19659 15045 19671 15048
rect 19613 15039 19671 15045
rect 20254 15036 20260 15048
rect 20312 15036 20318 15088
rect 23661 15079 23719 15085
rect 23661 15076 23673 15079
rect 22480 15048 23673 15076
rect 22480 15020 22508 15048
rect 23661 15045 23673 15048
rect 23707 15045 23719 15079
rect 23661 15039 23719 15045
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12492 14980 13001 15008
rect 12492 14968 12498 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 21266 15008 21272 15020
rect 20128 14980 21272 15008
rect 20128 14968 20134 14980
rect 21266 14968 21272 14980
rect 21324 15008 21330 15020
rect 21453 15011 21511 15017
rect 21453 15008 21465 15011
rect 21324 14980 21465 15008
rect 21324 14968 21330 14980
rect 21453 14977 21465 14980
rect 21499 14977 21511 15011
rect 22462 15008 22468 15020
rect 22375 14980 22468 15008
rect 21453 14971 21511 14977
rect 22462 14968 22468 14980
rect 22520 14968 22526 15020
rect 22646 15008 22652 15020
rect 22607 14980 22652 15008
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 24210 15008 24216 15020
rect 24171 14980 24216 15008
rect 24210 14968 24216 14980
rect 24268 15008 24274 15020
rect 24673 15011 24731 15017
rect 24673 15008 24685 15011
rect 24268 14980 24685 15008
rect 24268 14968 24274 14980
rect 24673 14977 24685 14980
rect 24719 15008 24731 15011
rect 25041 15011 25099 15017
rect 25041 15008 25053 15011
rect 24719 14980 25053 15008
rect 24719 14977 24731 14980
rect 24673 14971 24731 14977
rect 25041 14977 25053 14980
rect 25087 14977 25099 15011
rect 25406 15008 25412 15020
rect 25367 14980 25412 15008
rect 25041 14971 25099 14977
rect 25406 14968 25412 14980
rect 25464 14968 25470 15020
rect 1443 14912 2084 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 2866 14900 2872 14952
rect 2924 14900 2930 14952
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3694 14940 3700 14952
rect 3292 14912 3700 14940
rect 3292 14900 3298 14912
rect 3694 14900 3700 14912
rect 3752 14940 3758 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 3752 14912 4261 14940
rect 3752 14900 3758 14912
rect 4249 14909 4261 14912
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 4505 14943 4563 14949
rect 4505 14940 4517 14943
rect 4396 14912 4517 14940
rect 4396 14900 4402 14912
rect 4505 14909 4517 14912
rect 4551 14909 4563 14943
rect 4505 14903 4563 14909
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 5132 14912 6837 14940
rect 5132 14900 5138 14912
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 10321 14943 10379 14949
rect 6871 14912 7512 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 1854 14832 1860 14884
rect 1912 14872 1918 14884
rect 2317 14875 2375 14881
rect 2317 14872 2329 14875
rect 1912 14844 2329 14872
rect 1912 14832 1918 14844
rect 2317 14841 2329 14844
rect 2363 14841 2375 14875
rect 2317 14835 2375 14841
rect 2590 14764 2596 14816
rect 2648 14804 2654 14816
rect 2884 14813 2912 14900
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 2648 14776 2881 14804
rect 2648 14764 2654 14776
rect 2869 14773 2881 14776
rect 2915 14773 2927 14807
rect 2869 14767 2927 14773
rect 2961 14807 3019 14813
rect 2961 14773 2973 14807
rect 3007 14804 3019 14807
rect 4062 14804 4068 14816
rect 3007 14776 4068 14804
rect 3007 14773 3019 14776
rect 2961 14767 3019 14773
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4157 14807 4215 14813
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 5092 14804 5120 14900
rect 7484 14816 7512 14912
rect 10321 14909 10333 14943
rect 10367 14940 10379 14943
rect 11054 14940 11060 14952
rect 10367 14912 11060 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 11054 14900 11060 14912
rect 11112 14940 11118 14952
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 11112 14912 11161 14940
rect 11112 14900 11118 14912
rect 11149 14909 11161 14912
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 12802 14940 12808 14952
rect 12124 14912 12808 14940
rect 12124 14900 12130 14912
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 14277 14943 14335 14949
rect 14277 14909 14289 14943
rect 14323 14940 14335 14943
rect 14826 14940 14832 14952
rect 14323 14912 14832 14940
rect 14323 14909 14335 14912
rect 14277 14903 14335 14909
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 18506 14949 18512 14952
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 18500 14940 18512 14949
rect 16899 14912 17356 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 8266 14875 8324 14881
rect 8266 14872 8278 14875
rect 7944 14844 8278 14872
rect 7944 14816 7972 14844
rect 8266 14841 8278 14844
rect 8312 14841 8324 14875
rect 11793 14875 11851 14881
rect 11793 14872 11805 14875
rect 8266 14835 8324 14841
rect 11072 14844 11805 14872
rect 11072 14816 11100 14844
rect 11793 14841 11805 14844
rect 11839 14841 11851 14875
rect 11793 14835 11851 14841
rect 11974 14832 11980 14884
rect 12032 14872 12038 14884
rect 12897 14875 12955 14881
rect 12897 14872 12909 14875
rect 12032 14844 12909 14872
rect 12032 14832 12038 14844
rect 12897 14841 12909 14844
rect 12943 14841 12955 14875
rect 12897 14835 12955 14841
rect 14544 14875 14602 14881
rect 14544 14841 14556 14875
rect 14590 14872 14602 14875
rect 14642 14872 14648 14884
rect 14590 14844 14648 14872
rect 14590 14841 14602 14844
rect 14544 14835 14602 14841
rect 14642 14832 14648 14844
rect 14700 14832 14706 14884
rect 17328 14816 17356 14912
rect 18340 14912 18512 14940
rect 17862 14872 17868 14884
rect 17775 14844 17868 14872
rect 17862 14832 17868 14844
rect 17920 14872 17926 14884
rect 18340 14872 18368 14912
rect 18500 14903 18512 14912
rect 18506 14900 18512 14903
rect 18564 14900 18570 14952
rect 20441 14943 20499 14949
rect 20441 14909 20453 14943
rect 20487 14940 20499 14943
rect 20717 14943 20775 14949
rect 20717 14940 20729 14943
rect 20487 14912 20729 14940
rect 20487 14909 20499 14912
rect 20441 14903 20499 14909
rect 20717 14909 20729 14912
rect 20763 14909 20775 14943
rect 20717 14903 20775 14909
rect 23198 14900 23204 14952
rect 23256 14940 23262 14952
rect 23385 14943 23443 14949
rect 23385 14940 23397 14943
rect 23256 14912 23397 14940
rect 23256 14900 23262 14912
rect 23385 14909 23397 14912
rect 23431 14940 23443 14943
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23431 14912 24133 14940
rect 23431 14909 23443 14912
rect 23385 14903 23443 14909
rect 24121 14909 24133 14912
rect 24167 14940 24179 14943
rect 24762 14940 24768 14952
rect 24167 14912 24768 14940
rect 24167 14909 24179 14912
rect 24121 14903 24179 14909
rect 24762 14900 24768 14912
rect 24820 14900 24826 14952
rect 25225 14943 25283 14949
rect 25225 14909 25237 14943
rect 25271 14940 25283 14943
rect 25314 14940 25320 14952
rect 25271 14912 25320 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25314 14900 25320 14912
rect 25372 14940 25378 14952
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25372 14912 25973 14940
rect 25372 14900 25378 14912
rect 25961 14909 25973 14912
rect 26007 14909 26019 14943
rect 25961 14903 26019 14909
rect 17920 14844 18368 14872
rect 17920 14832 17926 14844
rect 19058 14832 19064 14884
rect 19116 14872 19122 14884
rect 20990 14872 20996 14884
rect 19116 14844 20668 14872
rect 20951 14844 20996 14872
rect 19116 14832 19122 14844
rect 4203 14776 5120 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5500 14776 5641 14804
rect 5500 14764 5506 14776
rect 5629 14773 5641 14776
rect 5675 14773 5687 14807
rect 7466 14804 7472 14816
rect 7427 14776 7472 14804
rect 5629 14767 5687 14773
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 7926 14804 7932 14816
rect 7887 14776 7932 14804
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14804 9459 14807
rect 9950 14804 9956 14816
rect 9447 14776 9956 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10781 14807 10839 14813
rect 10781 14773 10793 14807
rect 10827 14804 10839 14807
rect 10870 14804 10876 14816
rect 10827 14776 10876 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 11054 14764 11060 14816
rect 11112 14764 11118 14816
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 12124 14776 12173 14804
rect 12124 14764 12130 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12161 14767 12219 14773
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12400 14776 12449 14804
rect 12400 14764 12406 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 13446 14804 13452 14816
rect 13407 14776 13452 14804
rect 12437 14767 12495 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 13909 14807 13967 14813
rect 13909 14804 13921 14807
rect 13872 14776 13921 14804
rect 13872 14764 13878 14776
rect 13909 14773 13921 14776
rect 13955 14804 13967 14807
rect 14734 14804 14740 14816
rect 13955 14776 14740 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 15470 14764 15476 14816
rect 15528 14804 15534 14816
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15528 14776 15669 14804
rect 15528 14764 15534 14776
rect 15657 14773 15669 14776
rect 15703 14773 15715 14807
rect 15657 14767 15715 14773
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 16666 14804 16672 14816
rect 16540 14776 16672 14804
rect 16540 14764 16546 14776
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 17034 14804 17040 14816
rect 16995 14776 17040 14804
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 17310 14764 17316 14816
rect 17368 14804 17374 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 17368 14776 17417 14804
rect 17368 14764 17374 14776
rect 17405 14773 17417 14776
rect 17451 14773 17463 14807
rect 17405 14767 17463 14773
rect 20257 14807 20315 14813
rect 20257 14773 20269 14807
rect 20303 14804 20315 14807
rect 20346 14804 20352 14816
rect 20303 14776 20352 14804
rect 20303 14773 20315 14776
rect 20257 14767 20315 14773
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 20441 14807 20499 14813
rect 20441 14773 20453 14807
rect 20487 14804 20499 14807
rect 20530 14804 20536 14816
rect 20487 14776 20536 14804
rect 20487 14773 20499 14776
rect 20441 14767 20499 14773
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 20640 14804 20668 14844
rect 20990 14832 20996 14844
rect 21048 14832 21054 14884
rect 21910 14872 21916 14884
rect 21823 14844 21916 14872
rect 21910 14832 21916 14844
rect 21968 14872 21974 14884
rect 22373 14875 22431 14881
rect 22373 14872 22385 14875
rect 21968 14844 22385 14872
rect 21968 14832 21974 14844
rect 22373 14841 22385 14844
rect 22419 14841 22431 14875
rect 22373 14835 22431 14841
rect 23109 14875 23167 14881
rect 23109 14841 23121 14875
rect 23155 14872 23167 14875
rect 24026 14872 24032 14884
rect 23155 14844 24032 14872
rect 23155 14841 23167 14844
rect 23109 14835 23167 14841
rect 24026 14832 24032 14844
rect 24084 14832 24090 14884
rect 21450 14804 21456 14816
rect 20640 14776 21456 14804
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 22002 14804 22008 14816
rect 21963 14776 22008 14804
rect 22002 14764 22008 14776
rect 22060 14764 22066 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1578 14560 1584 14612
rect 1636 14600 1642 14612
rect 2406 14600 2412 14612
rect 1636 14572 2412 14600
rect 1636 14560 1642 14572
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 2593 14603 2651 14609
rect 2593 14569 2605 14603
rect 2639 14600 2651 14603
rect 2866 14600 2872 14612
rect 2639 14572 2872 14600
rect 2639 14569 2651 14572
rect 2593 14563 2651 14569
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 4062 14600 4068 14612
rect 4023 14572 4068 14600
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 4706 14600 4712 14612
rect 4479 14572 4712 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 4706 14560 4712 14572
rect 4764 14600 4770 14612
rect 5905 14603 5963 14609
rect 5905 14600 5917 14603
rect 4764 14572 5917 14600
rect 4764 14560 4770 14572
rect 5905 14569 5917 14572
rect 5951 14569 5963 14603
rect 9030 14600 9036 14612
rect 8991 14572 9036 14600
rect 5905 14563 5963 14569
rect 9030 14560 9036 14572
rect 9088 14600 9094 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 9088 14572 9413 14600
rect 9088 14560 9094 14572
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 14918 14600 14924 14612
rect 12860 14572 14924 14600
rect 12860 14560 12866 14572
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 19245 14603 19303 14609
rect 19245 14569 19257 14603
rect 19291 14600 19303 14603
rect 20530 14600 20536 14612
rect 19291 14572 20536 14600
rect 19291 14569 19303 14572
rect 19245 14563 19303 14569
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 21361 14603 21419 14609
rect 21361 14569 21373 14603
rect 21407 14600 21419 14603
rect 21450 14600 21456 14612
rect 21407 14572 21456 14600
rect 21407 14569 21419 14572
rect 21361 14563 21419 14569
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 22462 14600 22468 14612
rect 22423 14572 22468 14600
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 23474 14560 23480 14612
rect 23532 14600 23538 14612
rect 23934 14600 23940 14612
rect 23532 14572 23940 14600
rect 23532 14560 23538 14572
rect 23934 14560 23940 14572
rect 23992 14560 23998 14612
rect 25409 14603 25467 14609
rect 25409 14569 25421 14603
rect 25455 14600 25467 14603
rect 25498 14600 25504 14612
rect 25455 14572 25504 14600
rect 25455 14569 25467 14572
rect 25409 14563 25467 14569
rect 25498 14560 25504 14572
rect 25556 14560 25562 14612
rect 1946 14424 1952 14476
rect 2004 14424 2010 14476
rect 2884 14464 2912 14560
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 4614 14532 4620 14544
rect 3752 14504 4620 14532
rect 3752 14492 3758 14504
rect 4614 14492 4620 14504
rect 4672 14492 4678 14544
rect 4798 14492 4804 14544
rect 4856 14532 4862 14544
rect 5169 14535 5227 14541
rect 5169 14532 5181 14535
rect 4856 14504 5181 14532
rect 4856 14492 4862 14504
rect 5169 14501 5181 14504
rect 5215 14501 5227 14535
rect 10134 14532 10140 14544
rect 5169 14495 5227 14501
rect 9692 14504 10140 14532
rect 3605 14467 3663 14473
rect 3605 14464 3617 14467
rect 2884 14436 3617 14464
rect 3605 14433 3617 14436
rect 3651 14433 3663 14467
rect 6270 14464 6276 14476
rect 6231 14436 6276 14464
rect 3605 14427 3663 14433
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 6365 14467 6423 14473
rect 6365 14433 6377 14467
rect 6411 14464 6423 14467
rect 6730 14464 6736 14476
rect 6411 14436 6736 14464
rect 6411 14433 6423 14436
rect 6365 14427 6423 14433
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 8386 14464 8392 14476
rect 7800 14436 8392 14464
rect 7800 14424 7806 14436
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 9582 14464 9588 14476
rect 8527 14436 9588 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1964 14396 1992 14424
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 1719 14368 2053 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2041 14365 2053 14368
rect 2087 14396 2099 14399
rect 2406 14396 2412 14408
rect 2087 14368 2412 14396
rect 2087 14365 2099 14368
rect 2041 14359 2099 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2682 14396 2688 14408
rect 2643 14368 2688 14396
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 4522 14396 4528 14408
rect 4483 14368 4528 14396
rect 2869 14359 2927 14365
rect 2314 14288 2320 14340
rect 2372 14328 2378 14340
rect 2884 14328 2912 14359
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14396 5871 14399
rect 6178 14396 6184 14408
rect 5859 14368 6184 14396
rect 5859 14365 5871 14368
rect 5813 14359 5871 14365
rect 2372 14300 2912 14328
rect 2372 14288 2378 14300
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 4632 14328 4660 14359
rect 6178 14356 6184 14368
rect 6236 14396 6242 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6236 14368 6469 14396
rect 6236 14356 6242 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14396 7619 14399
rect 8496 14396 8524 14427
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 9692 14473 9720 14504
rect 9950 14473 9956 14476
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14433 9735 14467
rect 9944 14464 9956 14473
rect 9911 14436 9956 14464
rect 9677 14427 9735 14433
rect 9944 14427 9956 14436
rect 9950 14424 9956 14427
rect 10008 14424 10014 14476
rect 10060 14464 10088 14504
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 11698 14492 11704 14544
rect 11756 14532 11762 14544
rect 12434 14541 12440 14544
rect 12428 14532 12440 14541
rect 11756 14504 12440 14532
rect 11756 14492 11762 14504
rect 12428 14495 12440 14504
rect 12492 14532 12498 14544
rect 12492 14504 12576 14532
rect 12434 14492 12440 14495
rect 12492 14492 12498 14504
rect 15286 14492 15292 14544
rect 15344 14532 15350 14544
rect 15749 14535 15807 14541
rect 15749 14532 15761 14535
rect 15344 14504 15761 14532
rect 15344 14492 15350 14504
rect 15749 14501 15761 14504
rect 15795 14501 15807 14535
rect 15749 14495 15807 14501
rect 16390 14492 16396 14544
rect 16448 14532 16454 14544
rect 17681 14535 17739 14541
rect 17681 14532 17693 14535
rect 16448 14504 17693 14532
rect 16448 14492 16454 14504
rect 17681 14501 17693 14504
rect 17727 14532 17739 14535
rect 18601 14535 18659 14541
rect 18601 14532 18613 14535
rect 17727 14504 18613 14532
rect 17727 14501 17739 14504
rect 17681 14495 17739 14501
rect 18601 14501 18613 14504
rect 18647 14501 18659 14535
rect 18601 14495 18659 14501
rect 20254 14492 20260 14544
rect 20312 14532 20318 14544
rect 20349 14535 20407 14541
rect 20349 14532 20361 14535
rect 20312 14504 20361 14532
rect 20312 14492 20318 14504
rect 20349 14501 20361 14504
rect 20395 14532 20407 14535
rect 20395 14504 21588 14532
rect 20395 14501 20407 14504
rect 20349 14495 20407 14501
rect 15654 14464 15660 14476
rect 10060 14436 12204 14464
rect 15615 14436 15660 14464
rect 12176 14408 12204 14436
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14464 17647 14467
rect 18046 14464 18052 14476
rect 17635 14436 18052 14464
rect 17635 14433 17647 14436
rect 17589 14427 17647 14433
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 19153 14467 19211 14473
rect 19153 14433 19165 14467
rect 19199 14464 19211 14467
rect 19610 14464 19616 14476
rect 19199 14436 19616 14464
rect 19199 14433 19211 14436
rect 19153 14427 19211 14433
rect 19610 14424 19616 14436
rect 19668 14424 19674 14476
rect 20898 14424 20904 14476
rect 20956 14464 20962 14476
rect 21269 14467 21327 14473
rect 21269 14464 21281 14467
rect 20956 14436 21281 14464
rect 20956 14424 20962 14436
rect 21269 14433 21281 14436
rect 21315 14433 21327 14467
rect 21269 14427 21327 14433
rect 7607 14368 8524 14396
rect 8573 14399 8631 14405
rect 7607 14365 7619 14368
rect 7561 14359 7619 14365
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 12158 14396 12164 14408
rect 12119 14368 12164 14396
rect 8573 14359 8631 14365
rect 8588 14328 8616 14359
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14396 14427 14399
rect 14642 14396 14648 14408
rect 14415 14368 14648 14396
rect 14415 14365 14427 14368
rect 14369 14359 14427 14365
rect 14642 14356 14648 14368
rect 14700 14356 14706 14408
rect 15746 14356 15752 14408
rect 15804 14396 15810 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15804 14368 15945 14396
rect 15804 14356 15810 14368
rect 15933 14365 15945 14368
rect 15979 14365 15991 14399
rect 17862 14396 17868 14408
rect 17823 14368 17868 14396
rect 15933 14359 15991 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20070 14396 20076 14408
rect 19935 14368 20076 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 9306 14328 9312 14340
rect 4120 14300 4660 14328
rect 7944 14300 9312 14328
rect 4120 14288 4126 14300
rect 7944 14272 7972 14300
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 17129 14331 17187 14337
rect 17129 14297 17141 14331
rect 17175 14328 17187 14331
rect 17880 14328 17908 14356
rect 17175 14300 17908 14328
rect 17175 14297 17187 14300
rect 17129 14291 17187 14297
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19720 14328 19748 14359
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 21560 14405 21588 14504
rect 22738 14492 22744 14544
rect 22796 14532 22802 14544
rect 23658 14532 23664 14544
rect 22796 14504 23664 14532
rect 22796 14492 22802 14504
rect 23658 14492 23664 14504
rect 23716 14532 23722 14544
rect 24673 14535 24731 14541
rect 24673 14532 24685 14535
rect 23716 14504 24685 14532
rect 23716 14492 23722 14504
rect 24673 14501 24685 14504
rect 24719 14532 24731 14535
rect 25041 14535 25099 14541
rect 25041 14532 25053 14535
rect 24719 14504 25053 14532
rect 24719 14501 24731 14504
rect 24673 14495 24731 14501
rect 25041 14501 25053 14504
rect 25087 14501 25099 14535
rect 25041 14495 25099 14501
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 22646 14464 22652 14476
rect 22143 14436 22652 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 22646 14424 22652 14436
rect 22704 14464 22710 14476
rect 23008 14467 23066 14473
rect 23008 14464 23020 14467
rect 22704 14436 23020 14464
rect 22704 14424 22710 14436
rect 23008 14433 23020 14436
rect 23054 14464 23066 14467
rect 23382 14464 23388 14476
rect 23054 14436 23388 14464
rect 23054 14433 23066 14436
rect 23008 14427 23066 14433
rect 23382 14424 23388 14436
rect 23440 14464 23446 14476
rect 24762 14464 24768 14476
rect 23440 14436 24768 14464
rect 23440 14424 23446 14436
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 25222 14464 25228 14476
rect 25183 14436 25228 14464
rect 25222 14424 25228 14436
rect 25280 14424 25286 14476
rect 21545 14399 21603 14405
rect 21545 14365 21557 14399
rect 21591 14396 21603 14399
rect 21634 14396 21640 14408
rect 21591 14368 21640 14396
rect 21591 14365 21603 14368
rect 21545 14359 21603 14365
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 22738 14396 22744 14408
rect 22699 14368 22744 14396
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 20901 14331 20959 14337
rect 20901 14328 20913 14331
rect 19392 14300 20913 14328
rect 19392 14288 19398 14300
rect 20901 14297 20913 14300
rect 20947 14297 20959 14331
rect 20901 14291 20959 14297
rect 2038 14220 2044 14272
rect 2096 14260 2102 14272
rect 2225 14263 2283 14269
rect 2225 14260 2237 14263
rect 2096 14232 2237 14260
rect 2096 14220 2102 14232
rect 2225 14229 2237 14232
rect 2271 14229 2283 14263
rect 2225 14223 2283 14229
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3237 14263 3295 14269
rect 3237 14260 3249 14263
rect 2832 14232 3249 14260
rect 2832 14220 2838 14232
rect 3237 14229 3249 14232
rect 3283 14229 3295 14263
rect 7006 14260 7012 14272
rect 6967 14232 7012 14260
rect 3237 14223 3295 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7926 14260 7932 14272
rect 7887 14232 7932 14260
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 8021 14263 8079 14269
rect 8021 14229 8033 14263
rect 8067 14260 8079 14263
rect 8294 14260 8300 14272
rect 8067 14232 8300 14260
rect 8067 14229 8079 14232
rect 8021 14223 8079 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 11054 14260 11060 14272
rect 11015 14232 11060 14260
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 11698 14260 11704 14272
rect 11659 14232 11704 14260
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 11974 14260 11980 14272
rect 11935 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 13541 14263 13599 14269
rect 13541 14260 13553 14263
rect 12492 14232 13553 14260
rect 12492 14220 12498 14232
rect 13541 14229 13553 14232
rect 13587 14229 13599 14263
rect 13541 14223 13599 14229
rect 14737 14263 14795 14269
rect 14737 14229 14749 14263
rect 14783 14260 14795 14263
rect 14826 14260 14832 14272
rect 14783 14232 14832 14260
rect 14783 14229 14795 14232
rect 14737 14223 14795 14229
rect 14826 14220 14832 14232
rect 14884 14260 14890 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14884 14232 15025 14260
rect 14884 14220 14890 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 15562 14260 15568 14272
rect 15335 14232 15568 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15562 14220 15568 14232
rect 15620 14220 15626 14272
rect 16482 14260 16488 14272
rect 16443 14232 16488 14260
rect 16482 14220 16488 14232
rect 16540 14220 16546 14272
rect 17218 14260 17224 14272
rect 17179 14232 17224 14260
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 18230 14260 18236 14272
rect 18191 14232 18236 14260
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 20714 14260 20720 14272
rect 20675 14232 20720 14260
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 24118 14260 24124 14272
rect 24079 14232 24124 14260
rect 24118 14220 24124 14232
rect 24176 14220 24182 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2406 14016 2412 14068
rect 2464 14056 2470 14068
rect 2774 14056 2780 14068
rect 2464 14028 2780 14056
rect 2464 14016 2470 14028
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 7742 14056 7748 14068
rect 3108 14028 7748 14056
rect 3108 14016 3114 14028
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 9306 14056 9312 14068
rect 9267 14028 9312 14056
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11756 14028 12173 14056
rect 11756 14016 11762 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 16390 14056 16396 14068
rect 16351 14028 16396 14056
rect 12161 14019 12219 14025
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 18046 14056 18052 14068
rect 18007 14028 18052 14056
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14056 19211 14059
rect 19242 14056 19248 14068
rect 19199 14028 19248 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 19610 14056 19616 14068
rect 19571 14028 19616 14056
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 20898 14056 20904 14068
rect 20859 14028 20904 14056
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21361 14059 21419 14065
rect 21361 14025 21373 14059
rect 21407 14056 21419 14059
rect 21450 14056 21456 14068
rect 21407 14028 21456 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 21450 14016 21456 14028
rect 21508 14016 21514 14068
rect 21634 14056 21640 14068
rect 21595 14028 21640 14056
rect 21634 14016 21640 14028
rect 21692 14016 21698 14068
rect 23014 14056 23020 14068
rect 22975 14028 23020 14056
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 23474 14056 23480 14068
rect 23435 14028 23480 14056
rect 23474 14016 23480 14028
rect 23532 14056 23538 14068
rect 24762 14056 24768 14068
rect 23532 14028 24256 14056
rect 24723 14028 24768 14056
rect 23532 14016 23538 14028
rect 4798 13948 4804 14000
rect 4856 13948 4862 14000
rect 5074 13948 5080 14000
rect 5132 13988 5138 14000
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 5132 13960 5181 13988
rect 5132 13948 5138 13960
rect 5169 13957 5181 13960
rect 5215 13957 5227 13991
rect 5169 13951 5227 13957
rect 10781 13991 10839 13997
rect 10781 13957 10793 13991
rect 10827 13988 10839 13991
rect 11974 13988 11980 14000
rect 10827 13960 11980 13988
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 11974 13948 11980 13960
rect 12032 13948 12038 14000
rect 15194 13948 15200 14000
rect 15252 13988 15258 14000
rect 15746 13988 15752 14000
rect 15252 13960 15752 13988
rect 15252 13948 15258 13960
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 17862 13988 17868 14000
rect 17775 13960 17868 13988
rect 17862 13948 17868 13960
rect 17920 13988 17926 14000
rect 18506 13988 18512 14000
rect 17920 13960 18512 13988
rect 17920 13948 17926 13960
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 4816 13920 4844 13948
rect 5626 13920 5632 13932
rect 4816 13892 5632 13920
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 6270 13920 6276 13932
rect 6183 13892 6276 13920
rect 5721 13883 5779 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 4709 13855 4767 13861
rect 2740 13824 2820 13852
rect 2740 13812 2746 13824
rect 2222 13744 2228 13796
rect 2280 13793 2286 13796
rect 2280 13787 2344 13793
rect 2280 13753 2298 13787
rect 2332 13753 2344 13787
rect 2792 13784 2820 13824
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4798 13852 4804 13864
rect 4755 13824 4804 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 4798 13812 4804 13824
rect 4856 13852 4862 13864
rect 5442 13852 5448 13864
rect 4856 13824 5448 13852
rect 4856 13812 4862 13824
rect 5442 13812 5448 13824
rect 5500 13852 5506 13864
rect 5736 13852 5764 13883
rect 6270 13880 6276 13892
rect 6328 13920 6334 13932
rect 7282 13920 7288 13932
rect 6328 13892 7288 13920
rect 6328 13880 6334 13892
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 10321 13923 10379 13929
rect 7515 13892 8064 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 5500 13824 5764 13852
rect 6641 13855 6699 13861
rect 5500 13812 5506 13824
rect 6641 13821 6653 13855
rect 6687 13852 6699 13855
rect 6730 13852 6736 13864
rect 6687 13824 6736 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 7929 13855 7987 13861
rect 7929 13852 7941 13855
rect 7708 13824 7941 13852
rect 7708 13812 7714 13824
rect 7929 13821 7941 13824
rect 7975 13821 7987 13855
rect 8036 13852 8064 13892
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 11054 13920 11060 13932
rect 10367 13892 11060 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 11054 13880 11060 13892
rect 11112 13920 11118 13932
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 11112 13892 11345 13920
rect 11112 13880 11118 13892
rect 11333 13889 11345 13892
rect 11379 13889 11391 13923
rect 11333 13883 11391 13889
rect 13188 13892 13400 13920
rect 13188 13864 13216 13892
rect 8202 13861 8208 13864
rect 8185 13855 8208 13861
rect 8185 13852 8197 13855
rect 8036 13824 8197 13852
rect 7929 13815 7987 13821
rect 8185 13821 8197 13824
rect 8260 13852 8266 13864
rect 8260 13824 8333 13852
rect 8185 13815 8208 13821
rect 8202 13812 8208 13815
rect 8260 13812 8266 13824
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 8812 13824 9873 13852
rect 8812 13812 8818 13824
rect 9861 13821 9873 13824
rect 9907 13852 9919 13855
rect 9950 13852 9956 13864
rect 9907 13824 9956 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 11241 13855 11299 13861
rect 10735 13824 11100 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 3694 13784 3700 13796
rect 2792 13756 3700 13784
rect 2280 13747 2344 13753
rect 2280 13744 2286 13747
rect 3694 13744 3700 13756
rect 3752 13744 3758 13796
rect 4982 13744 4988 13796
rect 5040 13784 5046 13796
rect 5077 13787 5135 13793
rect 5077 13784 5089 13787
rect 5040 13756 5089 13784
rect 5040 13744 5046 13756
rect 5077 13753 5089 13756
rect 5123 13784 5135 13787
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5123 13756 5549 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 5537 13753 5549 13756
rect 5583 13784 5595 13787
rect 5994 13784 6000 13796
rect 5583 13756 6000 13784
rect 5583 13753 5595 13756
rect 5537 13747 5595 13753
rect 5994 13744 6000 13756
rect 6052 13744 6058 13796
rect 11072 13784 11100 13824
rect 11241 13821 11253 13855
rect 11287 13852 11299 13855
rect 11422 13852 11428 13864
rect 11287 13824 11428 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 13170 13852 13176 13864
rect 13131 13824 13176 13852
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13821 13323 13855
rect 13372 13852 13400 13892
rect 16482 13880 16488 13932
rect 16540 13920 16546 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16540 13892 17049 13920
rect 16540 13880 16546 13892
rect 17037 13889 17049 13892
rect 17083 13920 17095 13923
rect 18230 13920 18236 13932
rect 17083 13892 18236 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 18230 13880 18236 13892
rect 18288 13920 18294 13932
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18288 13892 18613 13920
rect 18288 13880 18294 13892
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 20254 13920 20260 13932
rect 20215 13892 20260 13920
rect 18601 13883 18659 13889
rect 20254 13880 20260 13892
rect 20312 13880 20318 13932
rect 22002 13880 22008 13932
rect 22060 13920 22066 13932
rect 22462 13920 22468 13932
rect 22060 13892 22468 13920
rect 22060 13880 22066 13892
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22646 13920 22652 13932
rect 22559 13892 22652 13920
rect 22646 13880 22652 13892
rect 22704 13920 22710 13932
rect 24118 13920 24124 13932
rect 22704 13892 24124 13920
rect 22704 13880 22710 13892
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 13521 13855 13579 13861
rect 13521 13852 13533 13855
rect 13372 13824 13533 13852
rect 13265 13815 13323 13821
rect 13521 13821 13533 13824
rect 13567 13821 13579 13855
rect 14826 13852 14832 13864
rect 13521 13815 13579 13821
rect 13648 13824 14832 13852
rect 13280 13784 13308 13815
rect 13648 13784 13676 13824
rect 14826 13812 14832 13824
rect 14884 13852 14890 13864
rect 15286 13852 15292 13864
rect 14884 13824 15148 13852
rect 15247 13824 15292 13852
rect 14884 13812 14890 13824
rect 11072 13756 11192 13784
rect 13280 13756 13676 13784
rect 15120 13784 15148 13824
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15654 13852 15660 13864
rect 15615 13824 15660 13852
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 16850 13852 16856 13864
rect 16724 13824 16856 13852
rect 16724 13812 16730 13824
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17402 13812 17408 13864
rect 17460 13852 17466 13864
rect 18506 13852 18512 13864
rect 17460 13824 17908 13852
rect 18467 13824 18512 13852
rect 17460 13812 17466 13824
rect 16390 13784 16396 13796
rect 15120 13756 16396 13784
rect 11164 13728 11192 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 17880 13784 17908 13824
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 19242 13812 19248 13864
rect 19300 13812 19306 13864
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19484 13824 20085 13852
rect 19484 13812 19490 13824
rect 20073 13821 20085 13824
rect 20119 13852 20131 13855
rect 20530 13852 20536 13864
rect 20119 13824 20536 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 23014 13812 23020 13864
rect 23072 13852 23078 13864
rect 24228 13852 24256 14028
rect 24762 14016 24768 14028
rect 24820 14016 24826 14068
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13920 24363 13923
rect 24780 13920 24808 14016
rect 25222 13948 25228 14000
rect 25280 13988 25286 14000
rect 25961 13991 26019 13997
rect 25961 13988 25973 13991
rect 25280 13960 25973 13988
rect 25280 13948 25286 13960
rect 25961 13957 25973 13960
rect 26007 13957 26019 13991
rect 25961 13951 26019 13957
rect 24351 13892 24808 13920
rect 24351 13889 24363 13892
rect 24305 13883 24363 13889
rect 25130 13880 25136 13932
rect 25188 13920 25194 13932
rect 25409 13923 25467 13929
rect 25409 13920 25421 13923
rect 25188 13892 25421 13920
rect 25188 13880 25194 13892
rect 25409 13889 25421 13892
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 24854 13852 24860 13864
rect 23072 13824 23796 13852
rect 23072 13812 23078 13824
rect 18417 13787 18475 13793
rect 18417 13784 18429 13787
rect 17880 13756 18429 13784
rect 18417 13753 18429 13756
rect 18463 13753 18475 13787
rect 19260 13784 19288 13812
rect 19981 13787 20039 13793
rect 19981 13784 19993 13787
rect 19260 13756 19993 13784
rect 18417 13747 18475 13753
rect 19981 13753 19993 13756
rect 20027 13753 20039 13787
rect 19981 13747 20039 13753
rect 22373 13787 22431 13793
rect 22373 13753 22385 13787
rect 22419 13784 22431 13787
rect 23768 13784 23796 13824
rect 24136 13824 24860 13852
rect 24136 13793 24164 13824
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25038 13852 25044 13864
rect 24999 13824 25044 13852
rect 25038 13812 25044 13824
rect 25096 13852 25102 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 25096 13824 25237 13852
rect 25096 13812 25102 13824
rect 25225 13821 25237 13824
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 24029 13787 24087 13793
rect 24029 13784 24041 13787
rect 22419 13756 23704 13784
rect 23768 13756 24041 13784
rect 22419 13753 22431 13756
rect 22373 13747 22431 13753
rect 23676 13728 23704 13756
rect 24029 13753 24041 13756
rect 24075 13753 24087 13787
rect 24029 13747 24087 13753
rect 24121 13787 24179 13793
rect 24121 13753 24133 13787
rect 24167 13753 24179 13787
rect 24121 13747 24179 13753
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2406 13716 2412 13728
rect 1995 13688 2412 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2406 13676 2412 13688
rect 2464 13676 2470 13728
rect 3421 13719 3479 13725
rect 3421 13685 3433 13719
rect 3467 13716 3479 13719
rect 3510 13716 3516 13728
rect 3467 13688 3516 13716
rect 3467 13685 3479 13688
rect 3421 13679 3479 13685
rect 3510 13676 3516 13688
rect 3568 13716 3574 13728
rect 4062 13716 4068 13728
rect 3568 13688 4068 13716
rect 3568 13676 3574 13688
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 11146 13716 11152 13728
rect 11107 13688 11152 13716
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11885 13719 11943 13725
rect 11885 13685 11897 13719
rect 11931 13716 11943 13719
rect 12158 13716 12164 13728
rect 11931 13688 12164 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 12158 13676 12164 13688
rect 12216 13716 12222 13728
rect 12618 13716 12624 13728
rect 12216 13688 12624 13716
rect 12216 13676 12222 13688
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 14642 13716 14648 13728
rect 14603 13688 14648 13716
rect 14642 13676 14648 13688
rect 14700 13676 14706 13728
rect 16301 13719 16359 13725
rect 16301 13685 16313 13719
rect 16347 13716 16359 13719
rect 16761 13719 16819 13725
rect 16761 13716 16773 13719
rect 16347 13688 16773 13716
rect 16347 13685 16359 13688
rect 16301 13679 16359 13685
rect 16761 13685 16773 13688
rect 16807 13716 16819 13719
rect 17126 13716 17132 13728
rect 16807 13688 17132 13716
rect 16807 13685 16819 13688
rect 16761 13679 16819 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 18322 13676 18328 13728
rect 18380 13716 18386 13728
rect 19426 13716 19432 13728
rect 18380 13688 19432 13716
rect 18380 13676 18386 13688
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 22005 13719 22063 13725
rect 22005 13685 22017 13719
rect 22051 13716 22063 13719
rect 22278 13716 22284 13728
rect 22051 13688 22284 13716
rect 22051 13685 22063 13688
rect 22005 13679 22063 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 22462 13716 22468 13728
rect 22423 13688 22468 13716
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 23658 13716 23664 13728
rect 23571 13688 23664 13716
rect 23658 13676 23664 13688
rect 23716 13676 23722 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1857 13515 1915 13521
rect 1857 13481 1869 13515
rect 1903 13512 1915 13515
rect 2590 13512 2596 13524
rect 1903 13484 2596 13512
rect 1903 13481 1915 13484
rect 1857 13475 1915 13481
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4522 13512 4528 13524
rect 4387 13484 4528 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 4522 13472 4528 13484
rect 4580 13472 4586 13524
rect 4706 13512 4712 13524
rect 4667 13484 4712 13512
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 6178 13512 6184 13524
rect 5500 13484 6184 13512
rect 5500 13472 5506 13484
rect 6178 13472 6184 13484
rect 6236 13512 6242 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6236 13484 6285 13512
rect 6236 13472 6242 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6273 13475 6331 13481
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 6972 13484 7757 13512
rect 6972 13472 6978 13484
rect 7745 13481 7757 13484
rect 7791 13512 7803 13515
rect 8110 13512 8116 13524
rect 7791 13484 8116 13512
rect 7791 13481 7803 13484
rect 7745 13475 7803 13481
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8481 13515 8539 13521
rect 8481 13512 8493 13515
rect 8352 13484 8493 13512
rect 8352 13472 8358 13484
rect 8481 13481 8493 13484
rect 8527 13481 8539 13515
rect 8481 13475 8539 13481
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9640 13484 9689 13512
rect 9640 13472 9646 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 10100 13484 10149 13512
rect 10100 13472 10106 13484
rect 10137 13481 10149 13484
rect 10183 13481 10195 13515
rect 10137 13475 10195 13481
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 11606 13512 11612 13524
rect 11112 13484 11612 13512
rect 11112 13472 11118 13484
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 11701 13515 11759 13521
rect 11701 13481 11713 13515
rect 11747 13512 11759 13515
rect 12342 13512 12348 13524
rect 11747 13484 12348 13512
rect 11747 13481 11759 13484
rect 11701 13475 11759 13481
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 13173 13515 13231 13521
rect 13173 13481 13185 13515
rect 13219 13512 13231 13515
rect 14001 13515 14059 13521
rect 14001 13512 14013 13515
rect 13219 13484 14013 13512
rect 13219 13481 13231 13484
rect 13173 13475 13231 13481
rect 14001 13481 14013 13484
rect 14047 13512 14059 13515
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 14047 13484 15301 13512
rect 14047 13481 14059 13484
rect 14001 13475 14059 13481
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 16482 13512 16488 13524
rect 16443 13484 16488 13512
rect 15289 13475 15347 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 18785 13515 18843 13521
rect 18785 13512 18797 13515
rect 18104 13484 18797 13512
rect 18104 13472 18110 13484
rect 18785 13481 18797 13484
rect 18831 13481 18843 13515
rect 19242 13512 19248 13524
rect 19203 13484 19248 13512
rect 18785 13475 18843 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 20070 13512 20076 13524
rect 20031 13484 20076 13512
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20898 13512 20904 13524
rect 20859 13484 20904 13512
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 22097 13515 22155 13521
rect 22097 13481 22109 13515
rect 22143 13512 22155 13515
rect 22646 13512 22652 13524
rect 22143 13484 22652 13512
rect 22143 13481 22155 13484
rect 22097 13475 22155 13481
rect 22646 13472 22652 13484
rect 22704 13472 22710 13524
rect 23293 13515 23351 13521
rect 23293 13481 23305 13515
rect 23339 13512 23351 13515
rect 23382 13512 23388 13524
rect 23339 13484 23388 13512
rect 23339 13481 23351 13484
rect 23293 13475 23351 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 23658 13512 23664 13524
rect 23619 13484 23664 13512
rect 23658 13472 23664 13484
rect 23716 13472 23722 13524
rect 3510 13444 3516 13456
rect 2424 13416 3516 13444
rect 2222 13376 2228 13388
rect 2183 13348 2228 13376
rect 2222 13336 2228 13348
rect 2280 13336 2286 13388
rect 1210 13268 1216 13320
rect 1268 13308 1274 13320
rect 2424 13317 2452 13416
rect 3510 13404 3516 13416
rect 3568 13404 3574 13456
rect 5160 13447 5218 13453
rect 5160 13413 5172 13447
rect 5206 13444 5218 13447
rect 5350 13444 5356 13456
rect 5206 13416 5356 13444
rect 5206 13413 5218 13416
rect 5160 13407 5218 13413
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 9401 13447 9459 13453
rect 9401 13413 9413 13447
rect 9447 13444 9459 13447
rect 9858 13444 9864 13456
rect 9447 13416 9864 13444
rect 9447 13413 9459 13416
rect 9401 13407 9459 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 14642 13404 14648 13456
rect 14700 13444 14706 13456
rect 14700 13416 15884 13444
rect 14700 13404 14706 13416
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 4908 13348 6837 13376
rect 2317 13311 2375 13317
rect 2317 13308 2329 13311
rect 1268 13280 2329 13308
rect 1268 13268 1274 13280
rect 2317 13277 2329 13280
rect 2363 13277 2375 13311
rect 2317 13271 2375 13277
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 4908 13317 4936 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6825 13339 6883 13345
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13376 7527 13379
rect 7742 13376 7748 13388
rect 7515 13348 7748 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7742 13336 7748 13348
rect 7800 13376 7806 13388
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 7800 13348 8401 13376
rect 7800 13336 7806 13348
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 10042 13376 10048 13388
rect 10003 13348 10048 13376
rect 8389 13339 8447 13345
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 15013 13379 15071 13385
rect 15013 13376 15025 13379
rect 14424 13348 15025 13376
rect 14424 13336 14430 13348
rect 15013 13345 15025 13348
rect 15059 13376 15071 13379
rect 15102 13376 15108 13388
rect 15059 13348 15108 13376
rect 15059 13345 15071 13348
rect 15013 13339 15071 13345
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15344 13348 15669 13376
rect 15344 13336 15350 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4764 13280 4905 13308
rect 4764 13268 4770 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8754 13308 8760 13320
rect 8711 13280 8760 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 11882 13308 11888 13320
rect 10284 13280 10329 13308
rect 11795 13280 11888 13308
rect 10284 13268 10290 13280
rect 11882 13268 11888 13280
rect 11940 13308 11946 13320
rect 12434 13308 12440 13320
rect 11940 13280 12440 13308
rect 11940 13268 11946 13280
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12676 13280 12725 13308
rect 12676 13268 12682 13280
rect 12713 13277 12725 13280
rect 12759 13308 12771 13311
rect 14090 13308 14096 13320
rect 12759 13280 13768 13308
rect 14051 13280 14096 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 8018 13240 8024 13252
rect 7979 13212 8024 13240
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 13630 13240 13636 13252
rect 13591 13212 13636 13240
rect 13630 13200 13636 13212
rect 13688 13200 13694 13252
rect 937 13175 995 13181
rect 937 13141 949 13175
rect 983 13172 995 13175
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 983 13144 1593 13172
rect 983 13141 995 13144
rect 937 13135 995 13141
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13172 3019 13175
rect 3234 13172 3240 13184
rect 3007 13144 3240 13172
rect 3007 13141 3019 13144
rect 2961 13135 3019 13141
rect 3234 13132 3240 13144
rect 3292 13132 3298 13184
rect 3694 13172 3700 13184
rect 3655 13144 3700 13172
rect 3694 13132 3700 13144
rect 3752 13132 3758 13184
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 9398 13172 9404 13184
rect 4672 13144 9404 13172
rect 4672 13132 4678 13144
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 10781 13175 10839 13181
rect 10781 13172 10793 13175
rect 10744 13144 10793 13172
rect 10744 13132 10750 13144
rect 10781 13141 10793 13144
rect 10827 13141 10839 13175
rect 10781 13135 10839 13141
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11241 13175 11299 13181
rect 11241 13172 11253 13175
rect 11112 13144 11253 13172
rect 11112 13132 11118 13144
rect 11241 13141 11253 13144
rect 11287 13172 11299 13175
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 11287 13144 12265 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 12253 13141 12265 13144
rect 12299 13141 12311 13175
rect 13446 13172 13452 13184
rect 13407 13144 13452 13172
rect 12253 13135 12311 13141
rect 13446 13132 13452 13144
rect 13504 13132 13510 13184
rect 13740 13172 13768 13280
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 15470 13308 15476 13320
rect 14323 13280 15476 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 15746 13308 15752 13320
rect 15707 13280 15752 13308
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 15856 13317 15884 13416
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19978 13444 19984 13456
rect 19484 13416 19984 13444
rect 19484 13404 19490 13416
rect 19978 13404 19984 13416
rect 20036 13404 20042 13456
rect 20162 13404 20168 13456
rect 20220 13444 20226 13456
rect 21269 13447 21327 13453
rect 21269 13444 21281 13447
rect 20220 13416 21281 13444
rect 20220 13404 20226 13416
rect 21269 13413 21281 13416
rect 21315 13444 21327 13447
rect 21910 13444 21916 13456
rect 21315 13416 21916 13444
rect 21315 13413 21327 13416
rect 21269 13407 21327 13413
rect 21910 13404 21916 13416
rect 21968 13404 21974 13456
rect 24020 13447 24078 13453
rect 24020 13413 24032 13447
rect 24066 13444 24078 13447
rect 24118 13444 24124 13456
rect 24066 13416 24124 13444
rect 24066 13413 24078 13416
rect 24020 13407 24078 13413
rect 24118 13404 24124 13416
rect 24176 13404 24182 13456
rect 17120 13379 17178 13385
rect 17120 13345 17132 13379
rect 17166 13376 17178 13379
rect 17402 13376 17408 13388
rect 17166 13348 17408 13376
rect 17166 13345 17178 13348
rect 17120 13339 17178 13345
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 19334 13376 19340 13388
rect 19295 13348 19340 13376
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 22278 13336 22284 13388
rect 22336 13376 22342 13388
rect 22465 13379 22523 13385
rect 22465 13376 22477 13379
rect 22336 13348 22477 13376
rect 22336 13336 22342 13348
rect 22465 13345 22477 13348
rect 22511 13376 22523 13379
rect 23014 13376 23020 13388
rect 22511 13348 23020 13376
rect 22511 13345 22523 13348
rect 22465 13339 22523 13345
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 20162 13308 20168 13320
rect 19659 13280 20168 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 14550 13172 14556 13184
rect 13740 13144 14556 13172
rect 14550 13132 14556 13144
rect 14608 13172 14614 13184
rect 14645 13175 14703 13181
rect 14645 13172 14657 13175
rect 14608 13144 14657 13172
rect 14608 13132 14614 13144
rect 14645 13141 14657 13144
rect 14691 13141 14703 13175
rect 14645 13135 14703 13141
rect 16390 13132 16396 13184
rect 16448 13172 16454 13184
rect 16868 13172 16896 13271
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 20898 13308 20904 13320
rect 20763 13280 20904 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 20898 13268 20904 13280
rect 20956 13308 20962 13320
rect 21361 13311 21419 13317
rect 21361 13308 21373 13311
rect 20956 13280 21373 13308
rect 20956 13268 20962 13280
rect 21361 13277 21373 13280
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 21634 13308 21640 13320
rect 21591 13280 21640 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22649 13311 22707 13317
rect 22649 13308 22661 13311
rect 22244 13280 22661 13308
rect 22244 13268 22250 13280
rect 22649 13277 22661 13280
rect 22695 13277 22707 13311
rect 22649 13271 22707 13277
rect 22738 13268 22744 13320
rect 22796 13308 22802 13320
rect 23753 13311 23811 13317
rect 23753 13308 23765 13311
rect 22796 13280 23765 13308
rect 22796 13268 22802 13280
rect 23753 13277 23765 13280
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 18230 13240 18236 13252
rect 18191 13212 18236 13240
rect 18230 13200 18236 13212
rect 18288 13200 18294 13252
rect 17494 13172 17500 13184
rect 16448 13144 17500 13172
rect 16448 13132 16454 13144
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 25130 13172 25136 13184
rect 25091 13144 25136 13172
rect 25130 13132 25136 13144
rect 25188 13132 25194 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1302 12928 1308 12980
rect 1360 12968 1366 12980
rect 3418 12968 3424 12980
rect 1360 12940 3096 12968
rect 1360 12928 1366 12940
rect 1581 12903 1639 12909
rect 1581 12869 1593 12903
rect 1627 12900 1639 12903
rect 2222 12900 2228 12912
rect 1627 12872 2228 12900
rect 1627 12869 1639 12872
rect 1581 12863 1639 12869
rect 2222 12860 2228 12872
rect 2280 12860 2286 12912
rect 937 12835 995 12841
rect 937 12801 949 12835
rect 983 12832 995 12835
rect 2041 12835 2099 12841
rect 2041 12832 2053 12835
rect 983 12804 2053 12832
rect 983 12801 995 12804
rect 937 12795 995 12801
rect 2041 12801 2053 12804
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 2314 12832 2320 12844
rect 2179 12804 2320 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 2314 12792 2320 12804
rect 2372 12792 2378 12844
rect 1946 12724 1952 12776
rect 2004 12764 2010 12776
rect 2682 12764 2688 12776
rect 2004 12736 2688 12764
rect 2004 12724 2010 12736
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 3068 12764 3096 12940
rect 3160 12940 3424 12968
rect 3160 12912 3188 12940
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4571 12940 5181 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 5169 12937 5181 12940
rect 5215 12968 5227 12971
rect 5350 12968 5356 12980
rect 5215 12940 5356 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 5994 12968 6000 12980
rect 5859 12940 6000 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 7742 12968 7748 12980
rect 7703 12940 7748 12968
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 9122 12928 9128 12940
rect 9180 12968 9186 12980
rect 9398 12968 9404 12980
rect 9180 12940 9404 12968
rect 9180 12928 9186 12940
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 10284 12940 10701 12968
rect 10284 12928 10290 12940
rect 10689 12937 10701 12940
rect 10735 12968 10747 12971
rect 10962 12968 10968 12980
rect 10735 12940 10968 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12342 12968 12348 12980
rect 12299 12940 12348 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 13630 12968 13636 12980
rect 13543 12940 13636 12968
rect 13630 12928 13636 12940
rect 13688 12968 13694 12980
rect 14090 12968 14096 12980
rect 13688 12940 14096 12968
rect 13688 12928 13694 12940
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 16206 12928 16212 12980
rect 16264 12968 16270 12980
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 16264 12940 17141 12968
rect 16264 12928 16270 12940
rect 17129 12937 17141 12940
rect 17175 12968 17187 12971
rect 17405 12971 17463 12977
rect 17405 12968 17417 12971
rect 17175 12940 17417 12968
rect 17175 12937 17187 12940
rect 17129 12931 17187 12937
rect 17405 12937 17417 12940
rect 17451 12937 17463 12971
rect 17405 12931 17463 12937
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17681 12971 17739 12977
rect 17681 12968 17693 12971
rect 17552 12940 17693 12968
rect 17552 12928 17558 12940
rect 17681 12937 17693 12940
rect 17727 12937 17739 12971
rect 17681 12931 17739 12937
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19392 12940 19441 12968
rect 19392 12928 19398 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 19610 12928 19616 12980
rect 19668 12968 19674 12980
rect 19889 12971 19947 12977
rect 19889 12968 19901 12971
rect 19668 12940 19901 12968
rect 19668 12928 19674 12940
rect 19889 12937 19901 12940
rect 19935 12937 19947 12971
rect 19889 12931 19947 12937
rect 3142 12860 3148 12912
rect 3200 12860 3206 12912
rect 7285 12903 7343 12909
rect 7285 12869 7297 12903
rect 7331 12900 7343 12903
rect 7926 12900 7932 12912
rect 7331 12872 7932 12900
rect 7331 12869 7343 12872
rect 7285 12863 7343 12869
rect 7926 12860 7932 12872
rect 7984 12900 7990 12912
rect 13541 12903 13599 12909
rect 7984 12872 8340 12900
rect 7984 12860 7990 12872
rect 5534 12832 5540 12844
rect 5495 12804 5540 12832
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 8312 12841 8340 12872
rect 13541 12869 13553 12903
rect 13587 12900 13599 12903
rect 16577 12903 16635 12909
rect 13587 12872 15148 12900
rect 13587 12869 13599 12872
rect 13541 12863 13599 12869
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7576 12804 8217 12832
rect 7576 12776 7604 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9824 12804 9873 12832
rect 9824 12792 9830 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13219 12804 14197 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 14185 12801 14197 12804
rect 14231 12832 14243 12835
rect 14642 12832 14648 12844
rect 14231 12804 14648 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 15120 12841 15148 12872
rect 16577 12869 16589 12903
rect 16623 12900 16635 12903
rect 18506 12900 18512 12912
rect 16623 12872 18512 12900
rect 16623 12869 16635 12872
rect 16577 12863 16635 12869
rect 18506 12860 18512 12872
rect 18564 12900 18570 12912
rect 19904 12900 19932 12931
rect 22462 12928 22468 12980
rect 22520 12968 22526 12980
rect 22649 12971 22707 12977
rect 22649 12968 22661 12971
rect 22520 12940 22661 12968
rect 22520 12928 22526 12940
rect 22649 12937 22661 12940
rect 22695 12937 22707 12971
rect 23014 12968 23020 12980
rect 22975 12940 23020 12968
rect 22649 12931 22707 12937
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 23477 12971 23535 12977
rect 23477 12937 23489 12971
rect 23523 12968 23535 12971
rect 24118 12968 24124 12980
rect 23523 12940 24124 12968
rect 23523 12937 23535 12940
rect 23477 12931 23535 12937
rect 24118 12928 24124 12940
rect 24176 12928 24182 12980
rect 20070 12900 20076 12912
rect 18564 12872 18644 12900
rect 18564 12860 18570 12872
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 15151 12804 15332 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 3068 12736 3157 12764
rect 3145 12733 3157 12736
rect 3191 12764 3203 12767
rect 4706 12764 4712 12776
rect 3191 12736 4712 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 5258 12724 5264 12776
rect 5316 12764 5322 12776
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5316 12736 5641 12764
rect 5316 12724 5322 12736
rect 5629 12733 5641 12736
rect 5675 12764 5687 12767
rect 6181 12767 6239 12773
rect 6181 12764 6193 12767
rect 5675 12736 6193 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 6181 12733 6193 12736
rect 6227 12733 6239 12767
rect 7558 12764 7564 12776
rect 7519 12736 7564 12764
rect 6181 12727 6239 12733
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 8110 12764 8116 12776
rect 8071 12736 8116 12764
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 9582 12764 9588 12776
rect 9088 12736 9588 12764
rect 9088 12724 9094 12736
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 11054 12764 11060 12776
rect 11015 12736 11060 12764
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13504 12736 14013 12764
rect 13504 12724 13510 12736
rect 14001 12733 14013 12736
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 15197 12767 15255 12773
rect 15197 12733 15209 12767
rect 15243 12733 15255 12767
rect 15304 12764 15332 12804
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 17310 12832 17316 12844
rect 17184 12804 17316 12832
rect 17184 12792 17190 12804
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 18616 12841 18644 12872
rect 19904 12872 20076 12900
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12832 18659 12835
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18647 12804 19073 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19904 12832 19932 12872
rect 20070 12860 20076 12872
rect 20128 12860 20134 12912
rect 23750 12860 23756 12912
rect 23808 12900 23814 12912
rect 24946 12900 24952 12912
rect 23808 12872 24952 12900
rect 23808 12860 23814 12872
rect 24946 12860 24952 12872
rect 25004 12900 25010 12912
rect 25004 12872 25084 12900
rect 25004 12860 25010 12872
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 19904 12804 20361 12832
rect 19061 12795 19119 12801
rect 20349 12801 20361 12804
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 23474 12832 23480 12844
rect 22428 12804 23480 12832
rect 22428 12792 22434 12804
rect 23474 12792 23480 12804
rect 23532 12832 23538 12844
rect 25056 12841 25084 12872
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23532 12804 24225 12832
rect 23532 12792 23538 12804
rect 24213 12801 24225 12804
rect 24259 12832 24271 12835
rect 24857 12835 24915 12841
rect 24857 12832 24869 12835
rect 24259 12804 24869 12832
rect 24259 12801 24271 12804
rect 24213 12795 24271 12801
rect 24857 12801 24869 12804
rect 24903 12801 24915 12835
rect 24857 12795 24915 12801
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 25087 12804 25421 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 15470 12773 15476 12776
rect 15464 12764 15476 12773
rect 15304 12736 15476 12764
rect 15197 12727 15255 12733
rect 15464 12727 15476 12736
rect 2593 12699 2651 12705
rect 2593 12696 2605 12699
rect 1964 12668 2605 12696
rect 1964 12640 1992 12668
rect 2593 12665 2605 12668
rect 2639 12665 2651 12699
rect 3390 12699 3448 12705
rect 3390 12696 3402 12699
rect 2593 12659 2651 12665
rect 2976 12668 3402 12696
rect 2976 12640 3004 12668
rect 3390 12665 3402 12668
rect 3436 12665 3448 12699
rect 3390 12659 3448 12665
rect 7926 12656 7932 12708
rect 7984 12696 7990 12708
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 7984 12668 9689 12696
rect 7984 12656 7990 12668
rect 9677 12665 9689 12668
rect 9723 12696 9735 12699
rect 9858 12696 9864 12708
rect 9723 12668 9864 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 10042 12656 10048 12708
rect 10100 12696 10106 12708
rect 10413 12699 10471 12705
rect 10413 12696 10425 12699
rect 10100 12668 10425 12696
rect 10100 12656 10106 12668
rect 10413 12665 10425 12668
rect 10459 12696 10471 12699
rect 10870 12696 10876 12708
rect 10459 12668 10876 12696
rect 10459 12665 10471 12668
rect 10413 12659 10471 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 11333 12699 11391 12705
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 12066 12696 12072 12708
rect 11379 12668 12072 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 15212 12696 15240 12727
rect 15470 12724 15476 12727
rect 15528 12724 15534 12776
rect 17494 12764 17500 12776
rect 17455 12736 17500 12764
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 17770 12724 17776 12776
rect 17828 12764 17834 12776
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 17828 12736 17877 12764
rect 17828 12724 17834 12736
rect 17865 12733 17877 12736
rect 17911 12764 17923 12767
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 17911 12736 20085 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 19076 12708 19104 12736
rect 20073 12733 20085 12736
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 16390 12696 16396 12708
rect 15212 12668 16396 12696
rect 16390 12656 16396 12668
rect 16448 12656 16454 12708
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 18417 12699 18475 12705
rect 18417 12696 18429 12699
rect 17451 12668 18429 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 18417 12665 18429 12668
rect 18463 12665 18475 12699
rect 18417 12659 18475 12665
rect 19058 12656 19064 12708
rect 19116 12656 19122 12708
rect 20088 12696 20116 12727
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 20605 12767 20663 12773
rect 20605 12764 20617 12767
rect 20496 12736 20617 12764
rect 20496 12724 20502 12736
rect 20605 12733 20617 12736
rect 20651 12733 20663 12767
rect 20605 12727 20663 12733
rect 20714 12696 20720 12708
rect 20088 12668 20720 12696
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 21266 12656 21272 12708
rect 21324 12696 21330 12708
rect 23937 12699 23995 12705
rect 23937 12696 23949 12699
rect 21324 12668 23949 12696
rect 21324 12656 21330 12668
rect 23937 12665 23949 12668
rect 23983 12696 23995 12699
rect 24765 12699 24823 12705
rect 24765 12696 24777 12699
rect 23983 12668 24777 12696
rect 23983 12665 23995 12668
rect 23937 12659 23995 12665
rect 24765 12665 24777 12668
rect 24811 12696 24823 12699
rect 25774 12696 25780 12708
rect 24811 12668 25780 12696
rect 24811 12665 24823 12668
rect 24765 12659 24823 12665
rect 25774 12656 25780 12668
rect 25832 12656 25838 12708
rect 1946 12628 1952 12640
rect 1907 12600 1952 12628
rect 1946 12588 1952 12600
rect 2004 12588 2010 12640
rect 2958 12628 2964 12640
rect 2919 12600 2964 12628
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 6638 12628 6644 12640
rect 6599 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 9306 12628 9312 12640
rect 9267 12600 9312 12628
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9769 12631 9827 12637
rect 9769 12628 9781 12631
rect 9456 12600 9781 12628
rect 9456 12588 9462 12600
rect 9769 12597 9781 12600
rect 9815 12628 9827 12631
rect 10686 12628 10692 12640
rect 9815 12600 10692 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 12621 12631 12679 12637
rect 12621 12597 12633 12631
rect 12667 12628 12679 12631
rect 13722 12628 13728 12640
rect 12667 12600 13728 12628
rect 12667 12597 12679 12600
rect 12621 12591 12679 12597
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 14093 12631 14151 12637
rect 14093 12597 14105 12631
rect 14139 12628 14151 12631
rect 14366 12628 14372 12640
rect 14139 12600 14372 12628
rect 14139 12597 14151 12600
rect 14093 12591 14151 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 17034 12628 17040 12640
rect 16632 12600 17040 12628
rect 16632 12588 16638 12600
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 18046 12628 18052 12640
rect 18007 12600 18052 12628
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 18509 12631 18567 12637
rect 18509 12628 18521 12631
rect 18380 12600 18521 12628
rect 18380 12588 18386 12600
rect 18509 12597 18521 12600
rect 18555 12597 18567 12631
rect 18509 12591 18567 12597
rect 21634 12588 21640 12640
rect 21692 12628 21698 12640
rect 21729 12631 21787 12637
rect 21729 12628 21741 12631
rect 21692 12600 21741 12628
rect 21692 12588 21698 12600
rect 21729 12597 21741 12600
rect 21775 12628 21787 12631
rect 22281 12631 22339 12637
rect 22281 12628 22293 12631
rect 21775 12600 22293 12628
rect 21775 12597 21787 12600
rect 21729 12591 21787 12597
rect 22281 12597 22293 12600
rect 22327 12597 22339 12631
rect 22281 12591 22339 12597
rect 23014 12588 23020 12640
rect 23072 12628 23078 12640
rect 24118 12628 24124 12640
rect 23072 12600 24124 12628
rect 23072 12588 23078 12600
rect 24118 12588 24124 12600
rect 24176 12588 24182 12640
rect 24397 12631 24455 12637
rect 24397 12597 24409 12631
rect 24443 12628 24455 12631
rect 24670 12628 24676 12640
rect 24443 12600 24676 12628
rect 24443 12597 24455 12600
rect 24397 12591 24455 12597
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 25406 12588 25412 12640
rect 25464 12628 25470 12640
rect 25869 12631 25927 12637
rect 25869 12628 25881 12631
rect 25464 12600 25881 12628
rect 25464 12588 25470 12600
rect 25869 12597 25881 12600
rect 25915 12628 25927 12631
rect 26145 12631 26203 12637
rect 26145 12628 26157 12631
rect 25915 12600 26157 12628
rect 25915 12597 25927 12600
rect 25869 12591 25927 12597
rect 26145 12597 26157 12600
rect 26191 12597 26203 12631
rect 26145 12591 26203 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1210 12384 1216 12436
rect 1268 12424 1274 12436
rect 1673 12427 1731 12433
rect 1673 12424 1685 12427
rect 1268 12396 1685 12424
rect 1268 12384 1274 12396
rect 1673 12393 1685 12396
rect 1719 12393 1731 12427
rect 1673 12387 1731 12393
rect 1688 12356 1716 12387
rect 2130 12384 2136 12436
rect 2188 12424 2194 12436
rect 3510 12424 3516 12436
rect 2188 12396 2820 12424
rect 3471 12396 3516 12424
rect 2188 12384 2194 12396
rect 2792 12356 2820 12396
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 4246 12424 4252 12436
rect 4207 12396 4252 12424
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 4522 12424 4528 12436
rect 4479 12396 4528 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 5997 12427 6055 12433
rect 5997 12424 6009 12427
rect 4764 12396 6009 12424
rect 4764 12384 4770 12396
rect 5997 12393 6009 12396
rect 6043 12393 6055 12427
rect 5997 12387 6055 12393
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 8352 12396 8769 12424
rect 8352 12384 8358 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 8757 12387 8815 12393
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 11514 12424 11520 12436
rect 9916 12396 11520 12424
rect 9916 12384 9922 12396
rect 11514 12384 11520 12396
rect 11572 12384 11578 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 11664 12396 12265 12424
rect 11664 12384 11670 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 12253 12387 12311 12393
rect 13173 12427 13231 12433
rect 13173 12393 13185 12427
rect 13219 12424 13231 12427
rect 13630 12424 13636 12436
rect 13219 12396 13636 12424
rect 13219 12393 13231 12396
rect 13173 12387 13231 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 13998 12424 14004 12436
rect 13872 12396 14004 12424
rect 13872 12384 13878 12396
rect 13998 12384 14004 12396
rect 14056 12384 14062 12436
rect 15105 12427 15163 12433
rect 15105 12393 15117 12427
rect 15151 12424 15163 12427
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15151 12396 15301 12424
rect 15151 12393 15163 12396
rect 15105 12387 15163 12393
rect 15289 12393 15301 12396
rect 15335 12424 15347 12427
rect 15746 12424 15752 12436
rect 15335 12396 15752 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 17402 12424 17408 12436
rect 17363 12396 17408 12424
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 19337 12427 19395 12433
rect 19337 12393 19349 12427
rect 19383 12424 19395 12427
rect 19426 12424 19432 12436
rect 19383 12396 19432 12424
rect 19383 12393 19395 12396
rect 19337 12387 19395 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 20438 12424 20444 12436
rect 20399 12396 20444 12424
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 20898 12424 20904 12436
rect 20859 12396 20904 12424
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 21910 12424 21916 12436
rect 21871 12396 21916 12424
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 23934 12384 23940 12436
rect 23992 12424 23998 12436
rect 24118 12424 24124 12436
rect 23992 12396 24124 12424
rect 23992 12384 23998 12396
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 24854 12424 24860 12436
rect 24815 12396 24860 12424
rect 24854 12384 24860 12396
rect 24912 12384 24918 12436
rect 3418 12356 3424 12368
rect 1688 12328 2728 12356
rect 2792 12328 3424 12356
rect 1670 12248 1676 12300
rect 1728 12288 1734 12300
rect 2041 12291 2099 12297
rect 2041 12288 2053 12291
rect 1728 12260 2053 12288
rect 1728 12248 1734 12260
rect 2041 12257 2053 12260
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2590 12288 2596 12300
rect 2179 12260 2596 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 2700 12288 2728 12328
rect 3418 12316 3424 12328
rect 3476 12316 3482 12368
rect 4264 12356 4292 12384
rect 4893 12359 4951 12365
rect 4893 12356 4905 12359
rect 4264 12328 4905 12356
rect 4893 12325 4905 12328
rect 4939 12325 4951 12359
rect 8570 12356 8576 12368
rect 4893 12319 4951 12325
rect 6472 12328 8576 12356
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 2700 12260 3801 12288
rect 3789 12257 3801 12260
rect 3835 12257 3847 12291
rect 3789 12251 3847 12257
rect 4801 12291 4859 12297
rect 4801 12257 4813 12291
rect 4847 12288 4859 12291
rect 5350 12288 5356 12300
rect 4847 12260 5356 12288
rect 4847 12257 4859 12260
rect 4801 12251 4859 12257
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 6472 12297 6500 12328
rect 8570 12316 8576 12328
rect 8628 12356 8634 12368
rect 8628 12328 9536 12356
rect 8628 12316 8634 12328
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 6227 12260 6469 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 7092 12291 7150 12297
rect 7092 12257 7104 12291
rect 7138 12288 7150 12291
rect 7374 12288 7380 12300
rect 7138 12260 7380 12288
rect 7138 12257 7150 12260
rect 7092 12251 7150 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 9508 12297 9536 12328
rect 9582 12316 9588 12368
rect 9640 12356 9646 12368
rect 10410 12356 10416 12368
rect 9640 12328 10416 12356
rect 9640 12316 9646 12328
rect 10410 12316 10416 12328
rect 10468 12316 10474 12368
rect 10588 12359 10646 12365
rect 10588 12325 10600 12359
rect 10634 12356 10646 12359
rect 10686 12356 10692 12368
rect 10634 12328 10692 12356
rect 10634 12325 10646 12328
rect 10588 12319 10646 12325
rect 10686 12316 10692 12328
rect 10744 12316 10750 12368
rect 14737 12359 14795 12365
rect 14737 12356 14749 12359
rect 13648 12328 14749 12356
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 2314 12220 2320 12232
rect 2227 12192 2320 12220
rect 2314 12180 2320 12192
rect 2372 12220 2378 12232
rect 3145 12223 3203 12229
rect 3145 12220 3157 12223
rect 2372 12192 3157 12220
rect 2372 12180 2378 12192
rect 3145 12189 3157 12192
rect 3191 12220 3203 12223
rect 3234 12220 3240 12232
rect 3191 12192 3240 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3234 12180 3240 12192
rect 3292 12220 3298 12232
rect 4522 12220 4528 12232
rect 3292 12192 4528 12220
rect 3292 12180 3298 12192
rect 4522 12180 4528 12192
rect 4580 12220 4586 12232
rect 5077 12223 5135 12229
rect 5077 12220 5089 12223
rect 4580 12192 5089 12220
rect 4580 12180 4586 12192
rect 5077 12189 5089 12192
rect 5123 12220 5135 12223
rect 5442 12220 5448 12232
rect 5123 12192 5448 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 6822 12220 6828 12232
rect 6783 12192 6828 12220
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 1486 12112 1492 12164
rect 1544 12152 1550 12164
rect 2130 12152 2136 12164
rect 1544 12124 2136 12152
rect 1544 12112 1550 12124
rect 2130 12112 2136 12124
rect 2188 12112 2194 12164
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 4890 12152 4896 12164
rect 4764 12124 4896 12152
rect 4764 12112 4770 12124
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 5905 12155 5963 12161
rect 5905 12121 5917 12155
rect 5951 12152 5963 12155
rect 6270 12152 6276 12164
rect 5951 12124 6276 12152
rect 5951 12121 5963 12124
rect 5905 12115 5963 12121
rect 6270 12112 6276 12124
rect 6328 12112 6334 12164
rect 9214 12112 9220 12164
rect 9272 12152 9278 12164
rect 9309 12155 9367 12161
rect 9309 12152 9321 12155
rect 9272 12124 9321 12152
rect 9272 12112 9278 12124
rect 9309 12121 9321 12124
rect 9355 12152 9367 12155
rect 10336 12152 10364 12180
rect 13648 12161 13676 12328
rect 14737 12325 14749 12328
rect 14783 12356 14795 12359
rect 15194 12356 15200 12368
rect 14783 12328 15200 12356
rect 14783 12325 14795 12328
rect 14737 12319 14795 12325
rect 15194 12316 15200 12328
rect 15252 12316 15258 12368
rect 15838 12316 15844 12368
rect 15896 12316 15902 12368
rect 20070 12356 20076 12368
rect 17972 12328 20076 12356
rect 13722 12248 13728 12300
rect 13780 12288 13786 12300
rect 13998 12288 14004 12300
rect 13780 12260 14004 12288
rect 13780 12248 13786 12260
rect 13998 12248 14004 12260
rect 14056 12248 14062 12300
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15528 12260 15669 12288
rect 15528 12248 15534 12260
rect 15657 12257 15669 12260
rect 15703 12288 15715 12291
rect 15856 12288 15884 12316
rect 16850 12288 16856 12300
rect 15703 12260 15884 12288
rect 16811 12260 16856 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 17972 12297 18000 12328
rect 20070 12316 20076 12328
rect 20128 12356 20134 12368
rect 22738 12356 22744 12368
rect 20128 12328 22744 12356
rect 20128 12316 20134 12328
rect 22738 12316 22744 12328
rect 22796 12316 22802 12368
rect 24578 12356 24584 12368
rect 23308 12328 24584 12356
rect 17957 12291 18015 12297
rect 17957 12257 17969 12291
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 18224 12291 18282 12297
rect 18224 12257 18236 12291
rect 18270 12288 18282 12291
rect 18598 12288 18604 12300
rect 18270 12260 18604 12288
rect 18270 12257 18282 12260
rect 18224 12251 18282 12257
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19392 12260 19993 12288
rect 19392 12248 19398 12260
rect 19981 12257 19993 12260
rect 20027 12288 20039 12291
rect 21269 12291 21327 12297
rect 21269 12288 21281 12291
rect 20027 12260 21281 12288
rect 20027 12257 20039 12260
rect 19981 12251 20039 12257
rect 21269 12257 21281 12260
rect 21315 12257 21327 12291
rect 23198 12288 23204 12300
rect 23159 12260 23204 12288
rect 21269 12251 21327 12257
rect 23198 12248 23204 12260
rect 23256 12248 23262 12300
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14090 12220 14096 12232
rect 13964 12192 14096 12220
rect 13964 12180 13970 12192
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14642 12220 14648 12232
rect 14323 12192 14648 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 15746 12220 15752 12232
rect 15707 12192 15752 12220
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12220 15991 12223
rect 16022 12220 16028 12232
rect 15979 12192 16028 12220
rect 15979 12189 15991 12192
rect 15933 12183 15991 12189
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 21358 12220 21364 12232
rect 20772 12192 21364 12220
rect 20772 12180 20778 12192
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21508 12192 21553 12220
rect 21508 12180 21514 12192
rect 22830 12180 22836 12232
rect 22888 12220 22894 12232
rect 23308 12229 23336 12328
rect 24578 12316 24584 12328
rect 24636 12316 24642 12368
rect 23934 12248 23940 12300
rect 23992 12288 23998 12300
rect 24765 12291 24823 12297
rect 24765 12288 24777 12291
rect 23992 12260 24777 12288
rect 23992 12248 23998 12260
rect 24765 12257 24777 12260
rect 24811 12257 24823 12291
rect 24765 12251 24823 12257
rect 23293 12223 23351 12229
rect 23293 12220 23305 12223
rect 22888 12192 23305 12220
rect 22888 12180 22894 12192
rect 23293 12189 23305 12192
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 23382 12180 23388 12232
rect 23440 12220 23446 12232
rect 23477 12223 23535 12229
rect 23477 12220 23489 12223
rect 23440 12192 23489 12220
rect 23440 12180 23446 12192
rect 23477 12189 23489 12192
rect 23523 12220 23535 12223
rect 23750 12220 23756 12232
rect 23523 12192 23756 12220
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 23750 12180 23756 12192
rect 23808 12180 23814 12232
rect 24213 12223 24271 12229
rect 24213 12189 24225 12223
rect 24259 12220 24271 12223
rect 25041 12223 25099 12229
rect 25041 12220 25053 12223
rect 24259 12192 25053 12220
rect 24259 12189 24271 12192
rect 24213 12183 24271 12189
rect 25041 12189 25053 12192
rect 25087 12220 25099 12223
rect 25130 12220 25136 12232
rect 25087 12192 25136 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 25130 12180 25136 12192
rect 25188 12180 25194 12232
rect 9355 12124 10364 12152
rect 13633 12155 13691 12161
rect 9355 12121 9367 12124
rect 9309 12115 9367 12121
rect 13633 12121 13645 12155
rect 13679 12121 13691 12155
rect 22738 12152 22744 12164
rect 22651 12124 22744 12152
rect 13633 12115 13691 12121
rect 22738 12112 22744 12124
rect 22796 12152 22802 12164
rect 22922 12152 22928 12164
rect 22796 12124 22928 12152
rect 22796 12112 22802 12124
rect 22922 12112 22928 12124
rect 22980 12112 22986 12164
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 2590 12084 2596 12096
rect 2464 12056 2596 12084
rect 2464 12044 2470 12056
rect 2590 12044 2596 12056
rect 2648 12084 2654 12096
rect 2685 12087 2743 12093
rect 2685 12084 2697 12087
rect 2648 12056 2697 12084
rect 2648 12044 2654 12056
rect 2685 12053 2697 12056
rect 2731 12053 2743 12087
rect 2685 12047 2743 12053
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 5224 12056 5457 12084
rect 5224 12044 5230 12056
rect 5445 12053 5457 12056
rect 5491 12053 5503 12087
rect 8202 12084 8208 12096
rect 8163 12056 8208 12084
rect 5445 12047 5503 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 8904 12056 9137 12084
rect 8904 12044 8910 12056
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 9950 12084 9956 12096
rect 9911 12056 9956 12084
rect 9125 12047 9183 12053
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11112 12056 11713 12084
rect 11112 12044 11118 12056
rect 11701 12053 11713 12056
rect 11747 12053 11759 12087
rect 11701 12047 11759 12053
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 12713 12087 12771 12093
rect 12713 12084 12725 12087
rect 11848 12056 12725 12084
rect 11848 12044 11854 12056
rect 12713 12053 12725 12056
rect 12759 12084 12771 12087
rect 13446 12084 13452 12096
rect 12759 12056 13452 12084
rect 12759 12053 12771 12056
rect 12713 12047 12771 12053
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 13541 12087 13599 12093
rect 13541 12053 13553 12087
rect 13587 12084 13599 12087
rect 14366 12084 14372 12096
rect 13587 12056 14372 12084
rect 13587 12053 13599 12056
rect 13541 12047 13599 12053
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 16393 12087 16451 12093
rect 16393 12053 16405 12087
rect 16439 12084 16451 12087
rect 16482 12084 16488 12096
rect 16439 12056 16488 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 16761 12087 16819 12093
rect 16761 12053 16773 12087
rect 16807 12084 16819 12087
rect 16850 12084 16856 12096
rect 16807 12056 16856 12084
rect 16807 12053 16819 12056
rect 16761 12047 16819 12053
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17037 12087 17095 12093
rect 17037 12053 17049 12087
rect 17083 12084 17095 12087
rect 17310 12084 17316 12096
rect 17083 12056 17316 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 17770 12084 17776 12096
rect 17731 12056 17776 12084
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 18690 12084 18696 12096
rect 18012 12056 18696 12084
rect 18012 12044 18018 12056
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 22370 12084 22376 12096
rect 22331 12056 22376 12084
rect 22370 12044 22376 12056
rect 22428 12044 22434 12096
rect 22833 12087 22891 12093
rect 22833 12053 22845 12087
rect 22879 12084 22891 12087
rect 23106 12084 23112 12096
rect 22879 12056 23112 12084
rect 22879 12053 22891 12056
rect 22833 12047 22891 12053
rect 23106 12044 23112 12056
rect 23164 12044 23170 12096
rect 24397 12087 24455 12093
rect 24397 12053 24409 12087
rect 24443 12084 24455 12087
rect 24762 12084 24768 12096
rect 24443 12056 24768 12084
rect 24443 12053 24455 12056
rect 24397 12047 24455 12053
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 25406 12044 25412 12096
rect 25464 12084 25470 12096
rect 25501 12087 25559 12093
rect 25501 12084 25513 12087
rect 25464 12056 25513 12084
rect 25464 12044 25470 12056
rect 25501 12053 25513 12056
rect 25547 12084 25559 12087
rect 25866 12084 25872 12096
rect 25547 12056 25872 12084
rect 25547 12053 25559 12056
rect 25501 12047 25559 12053
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1489 11883 1547 11889
rect 1489 11849 1501 11883
rect 1535 11880 1547 11883
rect 1670 11880 1676 11892
rect 1535 11852 1676 11880
rect 1535 11849 1547 11852
rect 1489 11843 1547 11849
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2682 11880 2688 11892
rect 2464 11852 2688 11880
rect 2464 11840 2470 11852
rect 2682 11840 2688 11852
rect 2740 11880 2746 11892
rect 3697 11883 3755 11889
rect 3697 11880 3709 11883
rect 2740 11852 3709 11880
rect 2740 11840 2746 11852
rect 3697 11849 3709 11852
rect 3743 11849 3755 11883
rect 3697 11843 3755 11849
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 5534 11880 5540 11892
rect 4203 11852 5540 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7653 11883 7711 11889
rect 7653 11880 7665 11883
rect 7248 11852 7665 11880
rect 7248 11840 7254 11852
rect 7653 11849 7665 11852
rect 7699 11849 7711 11883
rect 10778 11880 10784 11892
rect 10739 11852 10784 11880
rect 7653 11843 7711 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14148 11852 14381 11880
rect 14148 11840 14154 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15804 11852 15853 11880
rect 15804 11840 15810 11852
rect 15841 11849 15853 11852
rect 15887 11849 15899 11883
rect 15841 11843 15899 11849
rect 16942 11840 16948 11892
rect 17000 11880 17006 11892
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 17000 11852 17049 11880
rect 17000 11840 17006 11852
rect 17037 11849 17049 11852
rect 17083 11849 17095 11883
rect 17037 11843 17095 11849
rect 17589 11883 17647 11889
rect 17589 11849 17601 11883
rect 17635 11880 17647 11883
rect 18598 11880 18604 11892
rect 17635 11852 18092 11880
rect 18559 11852 18604 11880
rect 17635 11849 17647 11852
rect 17589 11843 17647 11849
rect 1118 11772 1124 11824
rect 1176 11812 1182 11824
rect 1578 11812 1584 11824
rect 1176 11784 1584 11812
rect 1176 11772 1182 11784
rect 1578 11772 1584 11784
rect 1636 11772 1642 11824
rect 5905 11815 5963 11821
rect 5905 11812 5917 11815
rect 5368 11784 5917 11812
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1670 11744 1676 11756
rect 1360 11716 1676 11744
rect 1360 11704 1366 11716
rect 1670 11704 1676 11716
rect 1728 11744 1734 11756
rect 1765 11747 1823 11753
rect 1765 11744 1777 11747
rect 1728 11716 1777 11744
rect 1728 11704 1734 11716
rect 1765 11713 1777 11716
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 5074 11704 5080 11756
rect 5132 11744 5138 11756
rect 5368 11753 5396 11784
rect 5905 11781 5917 11784
rect 5951 11781 5963 11815
rect 5905 11775 5963 11781
rect 9125 11815 9183 11821
rect 9125 11781 9137 11815
rect 9171 11812 9183 11815
rect 9582 11812 9588 11824
rect 9171 11784 9588 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 10410 11772 10416 11824
rect 10468 11812 10474 11824
rect 11790 11812 11796 11824
rect 10468 11784 11796 11812
rect 10468 11772 10474 11784
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 12069 11815 12127 11821
rect 12069 11812 12081 11815
rect 11940 11784 12081 11812
rect 11940 11772 11946 11784
rect 12069 11781 12081 11784
rect 12115 11812 12127 11815
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 12115 11784 12173 11812
rect 12115 11781 12127 11784
rect 12069 11775 12127 11781
rect 12161 11781 12173 11784
rect 12207 11781 12219 11815
rect 12161 11775 12219 11781
rect 15286 11772 15292 11824
rect 15344 11812 15350 11824
rect 16025 11815 16083 11821
rect 16025 11812 16037 11815
rect 15344 11784 16037 11812
rect 15344 11772 15350 11784
rect 16025 11781 16037 11784
rect 16071 11812 16083 11815
rect 16666 11812 16672 11824
rect 16071 11784 16672 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 17678 11812 17684 11824
rect 17639 11784 17684 11812
rect 17678 11772 17684 11784
rect 17736 11772 17742 11824
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 17828 11784 17908 11812
rect 17828 11772 17834 11784
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 5132 11716 5365 11744
rect 5132 11704 5138 11716
rect 5353 11713 5365 11716
rect 5399 11713 5411 11747
rect 5534 11744 5540 11756
rect 5495 11716 5540 11744
rect 5353 11707 5411 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7064 11716 7573 11744
rect 7064 11704 7070 11716
rect 7561 11713 7573 11716
rect 7607 11744 7619 11747
rect 8202 11744 8208 11756
rect 7607 11716 8208 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9766 11744 9772 11756
rect 8904 11716 9772 11744
rect 8904 11704 8910 11716
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 11422 11744 11428 11756
rect 11383 11716 11428 11744
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 16577 11747 16635 11753
rect 16577 11744 16589 11747
rect 16540 11716 16589 11744
rect 16540 11704 16546 11716
rect 16577 11713 16589 11716
rect 16623 11713 16635 11747
rect 16577 11707 16635 11713
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 2021 11679 2079 11685
rect 2021 11676 2033 11679
rect 1636 11648 2033 11676
rect 1636 11636 1642 11648
rect 2021 11645 2033 11648
rect 2067 11676 2079 11679
rect 2590 11676 2596 11688
rect 2067 11648 2596 11676
rect 2067 11645 2079 11648
rect 2021 11639 2079 11645
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8294 11676 8300 11688
rect 8159 11648 8300 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8294 11636 8300 11648
rect 8352 11676 8358 11688
rect 9306 11676 9312 11688
rect 8352 11648 9312 11676
rect 8352 11636 8358 11648
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 9582 11636 9588 11688
rect 9640 11676 9646 11688
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9640 11648 9689 11676
rect 9640 11636 9646 11648
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 9677 11639 9735 11645
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 10376 11648 12449 11676
rect 10376 11636 10382 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 1489 11611 1547 11617
rect 1489 11577 1501 11611
rect 1535 11608 1547 11611
rect 1673 11611 1731 11617
rect 1673 11608 1685 11611
rect 1535 11580 1685 11608
rect 1535 11577 1547 11580
rect 1489 11571 1547 11577
rect 1673 11577 1685 11580
rect 1719 11608 1731 11611
rect 2406 11608 2412 11620
rect 1719 11580 2412 11608
rect 1719 11577 1731 11580
rect 1673 11571 1731 11577
rect 2406 11568 2412 11580
rect 2464 11568 2470 11620
rect 2958 11568 2964 11620
rect 3016 11568 3022 11620
rect 4525 11611 4583 11617
rect 4525 11577 4537 11611
rect 4571 11608 4583 11611
rect 5350 11608 5356 11620
rect 4571 11580 5356 11608
rect 4571 11577 4583 11580
rect 4525 11571 4583 11577
rect 5350 11568 5356 11580
rect 5408 11608 5414 11620
rect 6178 11608 6184 11620
rect 5408 11580 6184 11608
rect 5408 11568 5414 11580
rect 6178 11568 6184 11580
rect 6236 11568 6242 11620
rect 6641 11611 6699 11617
rect 6641 11577 6653 11611
rect 6687 11608 6699 11611
rect 8021 11611 8079 11617
rect 8021 11608 8033 11611
rect 6687 11580 8033 11608
rect 6687 11577 6699 11580
rect 6641 11571 6699 11577
rect 8021 11577 8033 11580
rect 8067 11608 8079 11611
rect 8067 11580 9260 11608
rect 8067 11577 8079 11580
rect 8021 11571 8079 11577
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2976 11540 3004 11568
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 2188 11512 3157 11540
rect 2188 11500 2194 11512
rect 3145 11509 3157 11512
rect 3191 11509 3203 11543
rect 4890 11540 4896 11552
rect 4851 11512 4896 11540
rect 3145 11503 3203 11509
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5261 11543 5319 11549
rect 5261 11540 5273 11543
rect 5224 11512 5273 11540
rect 5224 11500 5230 11512
rect 5261 11509 5273 11512
rect 5307 11509 5319 11543
rect 5261 11503 5319 11509
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7374 11540 7380 11552
rect 7147 11512 7380 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 7374 11500 7380 11512
rect 7432 11540 7438 11552
rect 8665 11543 8723 11549
rect 8665 11540 8677 11543
rect 7432 11512 8677 11540
rect 7432 11500 7438 11512
rect 8665 11509 8677 11512
rect 8711 11540 8723 11543
rect 8846 11540 8852 11552
rect 8711 11512 8852 11540
rect 8711 11509 8723 11512
rect 8665 11503 8723 11509
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9232 11549 9260 11580
rect 9766 11568 9772 11620
rect 9824 11608 9830 11620
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 9824 11580 10609 11608
rect 9824 11568 9830 11580
rect 10597 11577 10609 11580
rect 10643 11608 10655 11611
rect 11241 11611 11299 11617
rect 11241 11608 11253 11611
rect 10643 11580 11253 11608
rect 10643 11577 10655 11580
rect 10597 11571 10655 11577
rect 11241 11577 11253 11580
rect 11287 11577 11299 11611
rect 12452 11608 12480 11639
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 12693 11679 12751 11685
rect 12693 11676 12705 11679
rect 12584 11648 12705 11676
rect 12584 11636 12590 11648
rect 12693 11645 12705 11648
rect 12739 11645 12751 11679
rect 14918 11676 14924 11688
rect 14879 11648 14924 11676
rect 12693 11639 12751 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11676 16451 11679
rect 17770 11676 17776 11688
rect 16439 11648 17776 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 17880 11685 17908 11784
rect 18064 11688 18092 11852
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19245 11883 19303 11889
rect 19245 11849 19257 11883
rect 19291 11880 19303 11883
rect 19334 11880 19340 11892
rect 19291 11852 19340 11880
rect 19291 11849 19303 11852
rect 19245 11843 19303 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 20717 11883 20775 11889
rect 20717 11880 20729 11883
rect 20496 11852 20729 11880
rect 20496 11840 20502 11852
rect 20717 11849 20729 11852
rect 20763 11880 20775 11883
rect 21269 11883 21327 11889
rect 21269 11880 21281 11883
rect 20763 11852 21281 11880
rect 20763 11849 20775 11852
rect 20717 11843 20775 11849
rect 21269 11849 21281 11852
rect 21315 11880 21327 11883
rect 21450 11880 21456 11892
rect 21315 11852 21456 11880
rect 21315 11849 21327 11852
rect 21269 11843 21327 11849
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 22462 11840 22468 11892
rect 22520 11880 22526 11892
rect 23198 11880 23204 11892
rect 22520 11852 23204 11880
rect 22520 11840 22526 11852
rect 23198 11840 23204 11852
rect 23256 11880 23262 11892
rect 23293 11883 23351 11889
rect 23293 11880 23305 11883
rect 23256 11852 23305 11880
rect 23256 11840 23262 11852
rect 23293 11849 23305 11852
rect 23339 11849 23351 11883
rect 23934 11880 23940 11892
rect 23895 11852 23940 11880
rect 23293 11843 23351 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 20622 11772 20628 11824
rect 20680 11812 20686 11824
rect 21729 11815 21787 11821
rect 21729 11812 21741 11815
rect 20680 11784 21741 11812
rect 20680 11772 20686 11784
rect 21729 11781 21741 11784
rect 21775 11781 21787 11815
rect 21729 11775 21787 11781
rect 17865 11679 17923 11685
rect 17865 11645 17877 11679
rect 17911 11645 17923 11679
rect 18046 11676 18052 11688
rect 18007 11648 18052 11676
rect 17865 11639 17923 11645
rect 14550 11608 14556 11620
rect 12452 11580 14556 11608
rect 11241 11571 11299 11577
rect 14550 11568 14556 11580
rect 14608 11568 14614 11620
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 14829 11611 14887 11617
rect 14829 11608 14841 11611
rect 14700 11580 14841 11608
rect 14700 11568 14706 11580
rect 14829 11577 14841 11580
rect 14875 11608 14887 11611
rect 16022 11608 16028 11620
rect 14875 11580 16028 11608
rect 14875 11577 14887 11580
rect 14829 11571 14887 11577
rect 16022 11568 16028 11580
rect 16080 11568 16086 11620
rect 17880 11608 17908 11639
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 19337 11679 19395 11685
rect 19337 11645 19349 11679
rect 19383 11645 19395 11679
rect 19337 11639 19395 11645
rect 17788 11580 17908 11608
rect 19352 11608 19380 11639
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 19593 11679 19651 11685
rect 19593 11676 19605 11679
rect 19484 11648 19605 11676
rect 19484 11636 19490 11648
rect 19593 11645 19605 11648
rect 19639 11645 19651 11679
rect 21744 11676 21772 11775
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22465 11747 22523 11753
rect 22465 11744 22477 11747
rect 22060 11716 22477 11744
rect 22060 11704 22066 11716
rect 22465 11713 22477 11716
rect 22511 11713 22523 11747
rect 22465 11707 22523 11713
rect 22278 11676 22284 11688
rect 21744 11648 22284 11676
rect 19593 11639 19651 11645
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 22922 11636 22928 11688
rect 22980 11676 22986 11688
rect 24121 11679 24179 11685
rect 24121 11676 24133 11679
rect 22980 11648 24133 11676
rect 22980 11636 22986 11648
rect 24121 11645 24133 11648
rect 24167 11676 24179 11679
rect 25406 11676 25412 11688
rect 24167 11648 25412 11676
rect 24167 11645 24179 11648
rect 24121 11639 24179 11645
rect 25406 11636 25412 11648
rect 25464 11636 25470 11688
rect 20070 11608 20076 11620
rect 19352 11580 20076 11608
rect 17788 11552 17816 11580
rect 20070 11568 20076 11580
rect 20128 11568 20134 11620
rect 24388 11611 24446 11617
rect 24388 11577 24400 11611
rect 24434 11608 24446 11611
rect 25038 11608 25044 11620
rect 24434 11580 25044 11608
rect 24434 11577 24446 11580
rect 24388 11571 24446 11577
rect 25038 11568 25044 11580
rect 25096 11568 25102 11620
rect 9217 11543 9275 11549
rect 9217 11509 9229 11543
rect 9263 11509 9275 11543
rect 9582 11540 9588 11552
rect 9543 11512 9588 11540
rect 9217 11503 9275 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10229 11543 10287 11549
rect 10229 11540 10241 11543
rect 9916 11512 10241 11540
rect 9916 11500 9922 11512
rect 10229 11509 10241 11512
rect 10275 11540 10287 11543
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 10275 11512 11161 11540
rect 10275 11509 10287 11512
rect 10229 11503 10287 11509
rect 11149 11509 11161 11512
rect 11195 11509 11207 11543
rect 11149 11503 11207 11509
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11664 11512 11805 11540
rect 11664 11500 11670 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12069 11543 12127 11549
rect 12069 11509 12081 11543
rect 12115 11540 12127 11543
rect 12526 11540 12532 11552
rect 12115 11512 12532 11540
rect 12115 11509 12127 11512
rect 12069 11503 12127 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 15102 11540 15108 11552
rect 15063 11512 15108 11540
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 16485 11543 16543 11549
rect 16485 11509 16497 11543
rect 16531 11540 16543 11543
rect 16850 11540 16856 11552
rect 16531 11512 16856 11540
rect 16531 11509 16543 11512
rect 16485 11503 16543 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17770 11500 17776 11552
rect 17828 11500 17834 11552
rect 18233 11543 18291 11549
rect 18233 11509 18245 11543
rect 18279 11540 18291 11543
rect 18966 11540 18972 11552
rect 18279 11512 18972 11540
rect 18279 11509 18291 11512
rect 18233 11503 18291 11509
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 21910 11540 21916 11552
rect 21871 11512 21916 11540
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 22373 11543 22431 11549
rect 22373 11509 22385 11543
rect 22419 11540 22431 11543
rect 22646 11540 22652 11552
rect 22419 11512 22652 11540
rect 22419 11509 22431 11512
rect 22373 11503 22431 11509
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 22738 11500 22744 11552
rect 22796 11540 22802 11552
rect 22925 11543 22983 11549
rect 22925 11540 22937 11543
rect 22796 11512 22937 11540
rect 22796 11500 22802 11512
rect 22925 11509 22937 11512
rect 22971 11509 22983 11543
rect 22925 11503 22983 11509
rect 25130 11500 25136 11552
rect 25188 11540 25194 11552
rect 25501 11543 25559 11549
rect 25501 11540 25513 11543
rect 25188 11512 25513 11540
rect 25188 11500 25194 11512
rect 25501 11509 25513 11512
rect 25547 11509 25559 11543
rect 25501 11503 25559 11509
rect 25866 11500 25872 11552
rect 25924 11540 25930 11552
rect 26053 11543 26111 11549
rect 26053 11540 26065 11543
rect 25924 11512 26065 11540
rect 25924 11500 25930 11512
rect 26053 11509 26065 11512
rect 26099 11509 26111 11543
rect 26053 11503 26111 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1581 11339 1639 11345
rect 1581 11336 1593 11339
rect 1452 11308 1593 11336
rect 1452 11296 1458 11308
rect 1581 11305 1593 11308
rect 1627 11305 1639 11339
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 1581 11299 1639 11305
rect 2038 11296 2044 11308
rect 2096 11336 2102 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 2096 11308 3341 11336
rect 2096 11296 2102 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 4522 11336 4528 11348
rect 4483 11308 4528 11336
rect 3329 11299 3387 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 5626 11336 5632 11348
rect 5500 11308 5632 11336
rect 5500 11296 5506 11308
rect 5626 11296 5632 11308
rect 5684 11336 5690 11348
rect 6089 11339 6147 11345
rect 6089 11336 6101 11339
rect 5684 11308 6101 11336
rect 5684 11296 5690 11308
rect 6089 11305 6101 11308
rect 6135 11305 6147 11339
rect 8294 11336 8300 11348
rect 8255 11308 8300 11336
rect 6089 11299 6147 11305
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11336 8634 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 8628 11308 8769 11336
rect 8628 11296 8634 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 9858 11296 9864 11348
rect 9916 11296 9922 11348
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 14056 11308 14197 11336
rect 14056 11296 14062 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14550 11336 14556 11348
rect 14511 11308 14556 11336
rect 14185 11299 14243 11305
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 16114 11336 16120 11348
rect 15519 11308 16120 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16393 11339 16451 11345
rect 16393 11336 16405 11339
rect 16356 11308 16405 11336
rect 16356 11296 16362 11308
rect 16393 11305 16405 11308
rect 16439 11305 16451 11339
rect 16393 11299 16451 11305
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16724 11308 16773 11336
rect 16724 11296 16730 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 19058 11336 19064 11348
rect 19019 11308 19064 11336
rect 16761 11299 16819 11305
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 20714 11336 20720 11348
rect 20675 11308 20720 11336
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 21266 11336 21272 11348
rect 21227 11308 21272 11336
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 22002 11336 22008 11348
rect 21915 11308 22008 11336
rect 22002 11296 22008 11308
rect 22060 11336 22066 11348
rect 24305 11339 24363 11345
rect 24305 11336 24317 11339
rect 22060 11308 24317 11336
rect 22060 11296 22066 11308
rect 24305 11305 24317 11308
rect 24351 11305 24363 11339
rect 24854 11336 24860 11348
rect 24815 11308 24860 11336
rect 24305 11299 24363 11305
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25038 11296 25044 11348
rect 25096 11336 25102 11348
rect 25225 11339 25283 11345
rect 25225 11336 25237 11339
rect 25096 11308 25237 11336
rect 25096 11296 25102 11308
rect 25225 11305 25237 11308
rect 25271 11305 25283 11339
rect 25225 11299 25283 11305
rect 2685 11271 2743 11277
rect 2685 11237 2697 11271
rect 2731 11268 2743 11271
rect 2866 11268 2872 11280
rect 2731 11240 2872 11268
rect 2731 11237 2743 11240
rect 2685 11231 2743 11237
rect 2866 11228 2872 11240
rect 2924 11228 2930 11280
rect 4798 11228 4804 11280
rect 4856 11268 4862 11280
rect 4954 11271 5012 11277
rect 4954 11268 4966 11271
rect 4856 11240 4966 11268
rect 4856 11228 4862 11240
rect 4954 11237 4966 11240
rect 5000 11268 5012 11271
rect 5534 11268 5540 11280
rect 5000 11240 5540 11268
rect 5000 11237 5012 11240
rect 4954 11231 5012 11237
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 7561 11271 7619 11277
rect 7561 11237 7573 11271
rect 7607 11268 7619 11271
rect 7834 11268 7840 11280
rect 7607 11240 7840 11268
rect 7607 11237 7619 11240
rect 7561 11231 7619 11237
rect 7834 11228 7840 11240
rect 7892 11268 7898 11280
rect 9122 11268 9128 11280
rect 7892 11240 9128 11268
rect 7892 11228 7898 11240
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 9309 11271 9367 11277
rect 9309 11237 9321 11271
rect 9355 11268 9367 11271
rect 9582 11268 9588 11280
rect 9355 11240 9588 11268
rect 9355 11237 9367 11240
rect 9309 11231 9367 11237
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 1949 11203 2007 11209
rect 1949 11200 1961 11203
rect 1452 11172 1961 11200
rect 1452 11160 1458 11172
rect 1949 11169 1961 11172
rect 1995 11200 2007 11203
rect 3697 11203 3755 11209
rect 3697 11200 3709 11203
rect 1995 11172 3709 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 3697 11169 3709 11172
rect 3743 11169 3755 11203
rect 3697 11163 3755 11169
rect 6270 11160 6276 11212
rect 6328 11200 6334 11212
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 6328 11172 6745 11200
rect 6328 11160 6334 11172
rect 6733 11169 6745 11172
rect 6779 11200 6791 11203
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6779 11172 7113 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 7101 11169 7113 11172
rect 7147 11200 7159 11203
rect 8202 11200 8208 11212
rect 7147 11172 8208 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8938 11200 8944 11212
rect 8899 11172 8944 11200
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9876 11144 9904 11296
rect 10137 11271 10195 11277
rect 10137 11237 10149 11271
rect 10183 11268 10195 11271
rect 11422 11268 11428 11280
rect 10183 11240 11428 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 11422 11228 11428 11240
rect 11480 11228 11486 11280
rect 13354 11228 13360 11280
rect 13412 11268 13418 11280
rect 13541 11271 13599 11277
rect 13541 11268 13553 11271
rect 13412 11240 13553 11268
rect 13412 11228 13418 11240
rect 13541 11237 13553 11240
rect 13587 11268 13599 11271
rect 13722 11268 13728 11280
rect 13587 11240 13728 11268
rect 13587 11237 13599 11240
rect 13541 11231 13599 11237
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 16209 11271 16267 11277
rect 16209 11237 16221 11271
rect 16255 11268 16267 11271
rect 17497 11271 17555 11277
rect 16255 11240 16988 11268
rect 16255 11237 16267 11240
rect 16209 11231 16267 11237
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 10485 11203 10543 11209
rect 10485 11200 10497 11203
rect 10376 11172 10497 11200
rect 10376 11160 10382 11172
rect 10485 11169 10497 11172
rect 10531 11169 10543 11203
rect 10485 11163 10543 11169
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15378 11200 15384 11212
rect 15335 11172 15384 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15378 11160 15384 11172
rect 15436 11200 15442 11212
rect 15746 11200 15752 11212
rect 15436 11172 15752 11200
rect 15436 11160 15442 11172
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 2130 11132 2136 11144
rect 2091 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 2792 11104 4721 11132
rect 2038 11024 2044 11076
rect 2096 11064 2102 11076
rect 2406 11064 2412 11076
rect 2096 11036 2412 11064
rect 2096 11024 2102 11036
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 937 10999 995 11005
rect 937 10965 949 10999
rect 983 10996 995 10999
rect 1486 10996 1492 11008
rect 983 10968 1492 10996
rect 983 10965 995 10968
rect 937 10959 995 10965
rect 1486 10956 1492 10968
rect 1544 10956 1550 11008
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 2792 10996 2820 11104
rect 4709 11101 4721 11104
rect 4755 11101 4767 11135
rect 7653 11135 7711 11141
rect 7653 11132 7665 11135
rect 4709 11095 4767 11101
rect 6932 11104 7665 11132
rect 4724 11008 4752 11095
rect 6932 11064 6960 11104
rect 7653 11101 7665 11104
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 8018 11132 8024 11144
rect 7883 11104 8024 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 10192 11104 10241 11132
rect 10192 11092 10198 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 10229 11095 10287 11101
rect 12176 11104 12541 11132
rect 7190 11064 7196 11076
rect 6840 11036 6960 11064
rect 7151 11036 7196 11064
rect 2958 10996 2964 11008
rect 1728 10968 2820 10996
rect 2919 10968 2964 10996
rect 1728 10956 1734 10968
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 4706 10956 4712 11008
rect 4764 10956 4770 11008
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 6840 10996 6868 11036
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 11514 11024 11520 11076
rect 11572 11064 11578 11076
rect 12176 11073 12204 11104
rect 12529 11101 12541 11104
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13633 11135 13691 11141
rect 13633 11132 13645 11135
rect 13412 11104 13645 11132
rect 13412 11092 13418 11104
rect 13633 11101 13645 11104
rect 13679 11101 13691 11135
rect 13633 11095 13691 11101
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 13814 11132 13820 11144
rect 13771 11104 13820 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 12161 11067 12219 11073
rect 12161 11064 12173 11067
rect 11572 11036 12173 11064
rect 11572 11024 11578 11036
rect 12161 11033 12173 11036
rect 12207 11033 12219 11067
rect 13078 11064 13084 11076
rect 13039 11036 13084 11064
rect 12161 11027 12219 11033
rect 13078 11024 13084 11036
rect 13136 11064 13142 11076
rect 13740 11064 13768 11095
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16022 11132 16028 11144
rect 15979 11104 16028 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16960 11141 16988 11240
rect 17497 11237 17509 11271
rect 17543 11268 17555 11271
rect 17862 11268 17868 11280
rect 17543 11240 17868 11268
rect 17543 11237 17555 11240
rect 17497 11231 17555 11237
rect 17862 11228 17868 11240
rect 17920 11228 17926 11280
rect 19429 11271 19487 11277
rect 19429 11237 19441 11271
rect 19475 11268 19487 11271
rect 20254 11268 20260 11280
rect 19475 11240 20260 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 20254 11228 20260 11240
rect 20312 11228 20318 11280
rect 21910 11228 21916 11280
rect 21968 11268 21974 11280
rect 22833 11271 22891 11277
rect 22833 11268 22845 11271
rect 21968 11240 22845 11268
rect 21968 11228 21974 11240
rect 22833 11237 22845 11240
rect 22879 11268 22891 11271
rect 23382 11268 23388 11280
rect 22879 11240 23388 11268
rect 22879 11237 22891 11240
rect 22833 11231 22891 11237
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 18012 11172 18337 11200
rect 18012 11160 18018 11172
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 18325 11163 18383 11169
rect 19521 11203 19579 11209
rect 19521 11169 19533 11203
rect 19567 11169 19579 11203
rect 22922 11200 22928 11212
rect 22883 11172 22928 11200
rect 19521 11163 19579 11169
rect 16853 11135 16911 11141
rect 16853 11101 16865 11135
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11132 17003 11135
rect 17678 11132 17684 11144
rect 16991 11104 17684 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 14918 11064 14924 11076
rect 13136 11036 13768 11064
rect 14879 11036 14924 11064
rect 13136 11024 13142 11036
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 16868 11064 16896 11095
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 18417 11135 18475 11141
rect 18417 11132 18429 11135
rect 18104 11104 18429 11132
rect 18104 11092 18110 11104
rect 18417 11101 18429 11104
rect 18463 11101 18475 11135
rect 18417 11095 18475 11101
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 19536 11132 19564 11163
rect 22922 11160 22928 11172
rect 22980 11160 22986 11212
rect 23198 11209 23204 11212
rect 23192 11200 23204 11209
rect 23159 11172 23204 11200
rect 23192 11163 23204 11172
rect 23198 11160 23204 11163
rect 23256 11160 23262 11212
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 18647 11104 18736 11132
rect 19536 11104 20177 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 17862 11064 17868 11076
rect 16868 11036 17868 11064
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 17957 11067 18015 11073
rect 17957 11033 17969 11067
rect 18003 11064 18015 11067
rect 18322 11064 18328 11076
rect 18003 11036 18328 11064
rect 18003 11033 18015 11036
rect 17957 11027 18015 11033
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 11606 10996 11612 11008
rect 6512 10968 6868 10996
rect 11567 10968 11612 10996
rect 6512 10956 6518 10968
rect 11606 10956 11612 10968
rect 11664 10956 11670 11008
rect 13170 10996 13176 11008
rect 13131 10968 13176 10996
rect 13170 10956 13176 10968
rect 13228 10956 13234 11008
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 16206 10996 16212 11008
rect 14884 10968 16212 10996
rect 14884 10956 14890 10968
rect 16206 10956 16212 10968
rect 16264 10996 16270 11008
rect 18138 10996 18144 11008
rect 16264 10968 18144 10996
rect 16264 10956 16270 10968
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 18598 10956 18604 11008
rect 18656 10996 18662 11008
rect 18708 10996 18736 11104
rect 20165 11101 20177 11104
rect 20211 11132 20223 11135
rect 20346 11132 20352 11144
rect 20211 11104 20352 11132
rect 20211 11101 20223 11104
rect 20165 11095 20223 11101
rect 20346 11092 20352 11104
rect 20404 11092 20410 11144
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20864 11104 21373 11132
rect 20864 11092 20870 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 21453 11135 21511 11141
rect 21453 11101 21465 11135
rect 21499 11101 21511 11135
rect 25406 11132 25412 11144
rect 25367 11104 25412 11132
rect 21453 11095 21511 11101
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20530 11064 20536 11076
rect 19751 11036 20536 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 20898 11064 20904 11076
rect 20859 11036 20904 11064
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 21468 11064 21496 11095
rect 25406 11092 25412 11104
rect 25464 11092 25470 11144
rect 21008 11036 21496 11064
rect 20070 10996 20076 11008
rect 18656 10968 20076 10996
rect 18656 10956 18662 10968
rect 20070 10956 20076 10968
rect 20128 10996 20134 11008
rect 21008 10996 21036 11036
rect 22462 11024 22468 11076
rect 22520 11064 22526 11076
rect 22922 11064 22928 11076
rect 22520 11036 22928 11064
rect 22520 11024 22526 11036
rect 22922 11024 22928 11036
rect 22980 11024 22986 11076
rect 20128 10968 21036 10996
rect 22373 10999 22431 11005
rect 20128 10956 20134 10968
rect 22373 10965 22385 10999
rect 22419 10996 22431 10999
rect 22646 10996 22652 11008
rect 22419 10968 22652 10996
rect 22419 10965 22431 10968
rect 22373 10959 22431 10965
rect 22646 10956 22652 10968
rect 22704 10956 22710 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4433 10795 4491 10801
rect 4433 10792 4445 10795
rect 4212 10764 4445 10792
rect 4212 10752 4218 10764
rect 4433 10761 4445 10764
rect 4479 10761 4491 10795
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 4433 10755 4491 10761
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6512 10764 6561 10792
rect 6512 10752 6518 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 7098 10792 7104 10804
rect 6549 10755 6607 10761
rect 6840 10764 7104 10792
rect 4706 10684 4712 10736
rect 4764 10724 4770 10736
rect 6840 10724 6868 10764
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 11330 10792 11336 10804
rect 9824 10764 11336 10792
rect 9824 10752 9830 10764
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 11514 10792 11520 10804
rect 11475 10764 11520 10792
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 14921 10795 14979 10801
rect 14921 10792 14933 10795
rect 13780 10764 14933 10792
rect 13780 10752 13786 10764
rect 14921 10761 14933 10764
rect 14967 10761 14979 10795
rect 14921 10755 14979 10761
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15654 10792 15660 10804
rect 15436 10764 15660 10792
rect 15436 10752 15442 10764
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 16853 10795 16911 10801
rect 16853 10792 16865 10795
rect 16632 10764 16865 10792
rect 16632 10752 16638 10764
rect 16853 10761 16865 10764
rect 16899 10761 16911 10795
rect 20070 10792 20076 10804
rect 20031 10764 20076 10792
rect 16853 10755 16911 10761
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 20441 10795 20499 10801
rect 20441 10761 20453 10795
rect 20487 10792 20499 10795
rect 21266 10792 21272 10804
rect 20487 10764 21272 10792
rect 20487 10761 20499 10764
rect 20441 10755 20499 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 22278 10792 22284 10804
rect 21744 10764 22284 10792
rect 4764 10696 6868 10724
rect 4764 10684 4770 10696
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4890 10656 4896 10668
rect 4019 10628 4896 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 6840 10665 6868 10696
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10137 10727 10195 10733
rect 10137 10724 10149 10727
rect 9732 10696 10149 10724
rect 9732 10684 9738 10696
rect 10137 10693 10149 10696
rect 10183 10693 10195 10727
rect 17402 10724 17408 10736
rect 17363 10696 17408 10724
rect 10137 10687 10195 10693
rect 17402 10684 17408 10696
rect 17460 10724 17466 10736
rect 17954 10724 17960 10736
rect 17460 10696 17960 10724
rect 17460 10684 17466 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10686 10656 10692 10668
rect 10091 10628 10692 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 1940 10591 1998 10597
rect 1940 10557 1952 10591
rect 1986 10588 1998 10591
rect 2958 10588 2964 10600
rect 1986 10560 2964 10588
rect 1986 10557 1998 10560
rect 1940 10551 1998 10557
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 5000 10588 5028 10619
rect 10686 10616 10692 10628
rect 10744 10656 10750 10668
rect 11606 10656 11612 10668
rect 10744 10628 11612 10656
rect 10744 10616 10750 10628
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 21744 10665 21772 10764
rect 22278 10752 22284 10764
rect 22336 10792 22342 10804
rect 22830 10792 22836 10804
rect 22336 10764 22836 10792
rect 22336 10752 22342 10764
rect 22830 10752 22836 10764
rect 22888 10752 22894 10804
rect 24026 10752 24032 10804
rect 24084 10792 24090 10804
rect 24213 10795 24271 10801
rect 24213 10792 24225 10795
rect 24084 10764 24225 10792
rect 24084 10752 24090 10764
rect 24213 10761 24225 10764
rect 24259 10761 24271 10795
rect 25866 10792 25872 10804
rect 25827 10764 25872 10792
rect 24213 10755 24271 10761
rect 21729 10659 21787 10665
rect 21729 10625 21741 10659
rect 21775 10625 21787 10659
rect 21910 10656 21916 10668
rect 21871 10628 21916 10656
rect 21729 10619 21787 10625
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 6270 10588 6276 10600
rect 4387 10560 6276 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 10134 10588 10140 10600
rect 9355 10560 10140 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 10134 10548 10140 10560
rect 10192 10588 10198 10600
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10192 10560 10609 10588
rect 10192 10548 10198 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 13035 10560 15485 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 15473 10557 15485 10560
rect 15519 10588 15531 10591
rect 16298 10588 16304 10600
rect 15519 10560 16304 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 1118 10480 1124 10532
rect 1176 10520 1182 10532
rect 1670 10520 1676 10532
rect 1176 10492 1676 10520
rect 1176 10480 1182 10492
rect 1670 10480 1676 10492
rect 1728 10480 1734 10532
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 4801 10523 4859 10529
rect 4801 10520 4813 10523
rect 4672 10492 4813 10520
rect 4672 10480 4678 10492
rect 4801 10489 4813 10492
rect 4847 10520 4859 10523
rect 5813 10523 5871 10529
rect 5813 10520 5825 10523
rect 4847 10492 5825 10520
rect 4847 10489 4859 10492
rect 4801 10483 4859 10489
rect 5813 10489 5825 10492
rect 5859 10489 5871 10523
rect 6288 10520 6316 10548
rect 7070 10523 7128 10529
rect 7070 10520 7082 10523
rect 6288 10492 7082 10520
rect 5813 10483 5871 10489
rect 7070 10489 7082 10492
rect 7116 10489 7128 10523
rect 7070 10483 7128 10489
rect 9677 10523 9735 10529
rect 9677 10489 9689 10523
rect 9723 10520 9735 10523
rect 10318 10520 10324 10532
rect 9723 10492 10324 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10505 10523 10563 10529
rect 10505 10489 10517 10523
rect 10551 10520 10563 10523
rect 10686 10520 10692 10532
rect 10551 10492 10692 10520
rect 10551 10489 10563 10492
rect 10505 10483 10563 10489
rect 10686 10480 10692 10492
rect 10744 10520 10750 10532
rect 11149 10523 11207 10529
rect 11149 10520 11161 10523
rect 10744 10492 11161 10520
rect 10744 10480 10750 10492
rect 11149 10489 11161 10492
rect 11195 10489 11207 10523
rect 11149 10483 11207 10489
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 13078 10520 13084 10532
rect 12299 10492 13084 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 13078 10480 13084 10492
rect 13136 10520 13142 10532
rect 13256 10523 13314 10529
rect 13256 10520 13268 10523
rect 13136 10492 13268 10520
rect 13136 10480 13142 10492
rect 13256 10489 13268 10492
rect 13302 10520 13314 10523
rect 13722 10520 13728 10532
rect 13302 10492 13728 10520
rect 13302 10489 13314 10492
rect 13256 10483 13314 10489
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 15381 10523 15439 10529
rect 15381 10489 15393 10523
rect 15427 10520 15439 10523
rect 15740 10523 15798 10529
rect 15740 10520 15752 10523
rect 15427 10492 15752 10520
rect 15427 10489 15439 10492
rect 15381 10483 15439 10489
rect 15740 10489 15752 10492
rect 15786 10520 15798 10523
rect 15838 10520 15844 10532
rect 15786 10492 15844 10520
rect 15786 10489 15798 10492
rect 15740 10483 15798 10489
rect 15838 10480 15844 10492
rect 15896 10480 15902 10532
rect 17678 10480 17684 10532
rect 17736 10520 17742 10532
rect 18294 10523 18352 10529
rect 18294 10520 18306 10523
rect 17736 10492 18306 10520
rect 17736 10480 17742 10492
rect 18294 10489 18306 10492
rect 18340 10489 18352 10523
rect 21082 10520 21088 10532
rect 21043 10492 21088 10520
rect 18294 10483 18352 10489
rect 21082 10480 21088 10492
rect 21140 10520 21146 10532
rect 21637 10523 21695 10529
rect 21637 10520 21649 10523
rect 21140 10492 21649 10520
rect 21140 10480 21146 10492
rect 21637 10489 21649 10492
rect 21683 10489 21695 10523
rect 24228 10520 24256 10755
rect 25866 10752 25872 10764
rect 25924 10752 25930 10804
rect 25409 10727 25467 10733
rect 25409 10724 25421 10727
rect 24872 10696 25421 10724
rect 24762 10616 24768 10668
rect 24820 10656 24826 10668
rect 24872 10665 24900 10696
rect 25409 10693 25421 10696
rect 25455 10693 25467 10727
rect 25409 10687 25467 10693
rect 24857 10659 24915 10665
rect 24857 10656 24869 10659
rect 24820 10628 24869 10656
rect 24820 10616 24826 10628
rect 24857 10625 24869 10628
rect 24903 10625 24915 10659
rect 24857 10619 24915 10625
rect 25041 10659 25099 10665
rect 25041 10625 25053 10659
rect 25087 10656 25099 10659
rect 25130 10656 25136 10668
rect 25087 10628 25136 10656
rect 25087 10625 25099 10628
rect 25041 10619 25099 10625
rect 24302 10548 24308 10600
rect 24360 10588 24366 10600
rect 25056 10588 25084 10619
rect 25130 10616 25136 10628
rect 25188 10616 25194 10668
rect 24360 10560 25084 10588
rect 24360 10548 24366 10560
rect 24765 10523 24823 10529
rect 24765 10520 24777 10523
rect 24228 10492 24777 10520
rect 21637 10483 21695 10489
rect 24765 10489 24777 10492
rect 24811 10489 24823 10523
rect 24765 10483 24823 10489
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 1636 10424 3065 10452
rect 1636 10412 1642 10424
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3053 10415 3111 10421
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6181 10455 6239 10461
rect 6181 10452 6193 10455
rect 6052 10424 6193 10452
rect 6052 10412 6058 10424
rect 6181 10421 6193 10424
rect 6227 10421 6239 10455
rect 6181 10415 6239 10421
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 8018 10452 8024 10464
rect 7340 10424 8024 10452
rect 7340 10412 7346 10424
rect 8018 10412 8024 10424
rect 8076 10452 8082 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 8076 10424 8217 10452
rect 8076 10412 8082 10424
rect 8205 10421 8217 10424
rect 8251 10452 8263 10455
rect 8757 10455 8815 10461
rect 8757 10452 8769 10455
rect 8251 10424 8769 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 8757 10421 8769 10424
rect 8803 10421 8815 10455
rect 10336 10452 10364 10480
rect 10778 10452 10784 10464
rect 10336 10424 10784 10452
rect 8757 10415 8815 10421
rect 10778 10412 10784 10424
rect 10836 10452 10842 10464
rect 11422 10452 11428 10464
rect 10836 10424 11428 10452
rect 10836 10412 10842 10424
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13354 10452 13360 10464
rect 12943 10424 13360 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 13688 10424 14381 10452
rect 13688 10412 13694 10424
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 14369 10415 14427 10421
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 17460 10424 17785 10452
rect 17460 10412 17466 10424
rect 17773 10421 17785 10424
rect 17819 10452 17831 10455
rect 18046 10452 18052 10464
rect 17819 10424 18052 10452
rect 17819 10421 17831 10424
rect 17773 10415 17831 10421
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19429 10455 19487 10461
rect 19429 10452 19441 10455
rect 19392 10424 19441 10452
rect 19392 10412 19398 10424
rect 19429 10421 19441 10424
rect 19475 10421 19487 10455
rect 20806 10452 20812 10464
rect 20767 10424 20812 10452
rect 19429 10415 19487 10421
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 21269 10455 21327 10461
rect 21269 10421 21281 10455
rect 21315 10452 21327 10455
rect 21818 10452 21824 10464
rect 21315 10424 21824 10452
rect 21315 10421 21327 10424
rect 21269 10415 21327 10421
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 23017 10455 23075 10461
rect 23017 10421 23029 10455
rect 23063 10452 23075 10455
rect 23198 10452 23204 10464
rect 23063 10424 23204 10452
rect 23063 10421 23075 10424
rect 23017 10415 23075 10421
rect 23198 10412 23204 10424
rect 23256 10412 23262 10464
rect 23385 10455 23443 10461
rect 23385 10421 23397 10455
rect 23431 10452 23443 10455
rect 23658 10452 23664 10464
rect 23431 10424 23664 10452
rect 23431 10421 23443 10424
rect 23385 10415 23443 10421
rect 23658 10412 23664 10424
rect 23716 10412 23722 10464
rect 23937 10455 23995 10461
rect 23937 10421 23949 10455
rect 23983 10452 23995 10455
rect 24302 10452 24308 10464
rect 23983 10424 24308 10452
rect 23983 10421 23995 10424
rect 23937 10415 23995 10421
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 24397 10455 24455 10461
rect 24397 10421 24409 10455
rect 24443 10452 24455 10455
rect 24670 10452 24676 10464
rect 24443 10424 24676 10452
rect 24443 10421 24455 10424
rect 24397 10415 24455 10421
rect 24670 10412 24676 10424
rect 24728 10412 24734 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1397 10251 1455 10257
rect 1397 10217 1409 10251
rect 1443 10248 1455 10251
rect 1946 10248 1952 10260
rect 1443 10220 1952 10248
rect 1443 10217 1455 10220
rect 1397 10211 1455 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2866 10248 2872 10260
rect 2823 10220 2872 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3292 10220 3433 10248
rect 3292 10208 3298 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 6270 10248 6276 10260
rect 6231 10220 6276 10248
rect 3421 10211 3479 10217
rect 6270 10208 6276 10220
rect 6328 10248 6334 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6328 10220 6837 10248
rect 6328 10208 6334 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 6825 10211 6883 10217
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7834 10248 7840 10260
rect 7331 10220 7840 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 9582 10248 9588 10260
rect 8435 10220 9588 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10180 2375 10183
rect 3602 10180 3608 10192
rect 2363 10152 3608 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2130 10112 2136 10124
rect 1995 10084 2136 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 3068 10056 3096 10152
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 4246 10180 4252 10192
rect 4207 10152 4252 10180
rect 4246 10140 4252 10152
rect 4304 10140 4310 10192
rect 5160 10183 5218 10189
rect 5160 10149 5172 10183
rect 5206 10180 5218 10183
rect 5442 10180 5448 10192
rect 5206 10152 5448 10180
rect 5206 10149 5218 10152
rect 5160 10143 5218 10149
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 7742 10140 7748 10192
rect 7800 10180 7806 10192
rect 8404 10180 8432 10211
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 11422 10248 11428 10260
rect 11383 10220 11428 10248
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11977 10251 12035 10257
rect 11977 10248 11989 10251
rect 11572 10220 11989 10248
rect 11572 10208 11578 10220
rect 11977 10217 11989 10220
rect 12023 10248 12035 10251
rect 12526 10248 12532 10260
rect 12023 10220 12532 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 12621 10251 12679 10257
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 13170 10248 13176 10260
rect 12667 10220 13176 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 13170 10208 13176 10220
rect 13228 10248 13234 10260
rect 13449 10251 13507 10257
rect 13449 10248 13461 10251
rect 13228 10220 13461 10248
rect 13228 10208 13234 10220
rect 13449 10217 13461 10220
rect 13495 10217 13507 10251
rect 13449 10211 13507 10217
rect 13538 10208 13544 10260
rect 13596 10248 13602 10260
rect 14461 10251 14519 10257
rect 14461 10248 14473 10251
rect 13596 10220 14473 10248
rect 13596 10208 13602 10220
rect 14461 10217 14473 10220
rect 14507 10217 14519 10251
rect 15102 10248 15108 10260
rect 15063 10220 15108 10248
rect 14461 10211 14519 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15286 10248 15292 10260
rect 15247 10220 15292 10248
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 17678 10208 17684 10220
rect 17736 10248 17742 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 17736 10220 18245 10248
rect 17736 10208 17742 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18233 10211 18291 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19576 10220 19717 10248
rect 19576 10208 19582 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 21910 10248 21916 10260
rect 21871 10220 21916 10248
rect 19705 10211 19763 10217
rect 21910 10208 21916 10220
rect 21968 10208 21974 10260
rect 22646 10248 22652 10260
rect 22607 10220 22652 10248
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 23014 10208 23020 10260
rect 23072 10248 23078 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 23072 10220 23121 10248
rect 23072 10208 23078 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 23109 10211 23167 10217
rect 24213 10251 24271 10257
rect 24213 10217 24225 10251
rect 24259 10248 24271 10251
rect 24302 10248 24308 10260
rect 24259 10220 24308 10248
rect 24259 10217 24271 10220
rect 24213 10211 24271 10217
rect 24302 10208 24308 10220
rect 24360 10208 24366 10260
rect 7800 10152 8432 10180
rect 7800 10140 7806 10152
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 8536 10152 8581 10180
rect 8536 10140 8542 10152
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 16574 10189 16580 10192
rect 10290 10183 10348 10189
rect 10290 10180 10302 10183
rect 10100 10152 10302 10180
rect 10100 10140 10106 10152
rect 10290 10149 10302 10152
rect 10336 10149 10348 10183
rect 16568 10180 16580 10189
rect 16535 10152 16580 10180
rect 10290 10143 10348 10149
rect 16568 10143 16580 10152
rect 16574 10140 16580 10143
rect 16632 10140 16638 10192
rect 19426 10140 19432 10192
rect 19484 10180 19490 10192
rect 19613 10183 19671 10189
rect 19613 10180 19625 10183
rect 19484 10152 19625 10180
rect 19484 10140 19490 10152
rect 19613 10149 19625 10152
rect 19659 10149 19671 10183
rect 19613 10143 19671 10149
rect 21361 10183 21419 10189
rect 21361 10149 21373 10183
rect 21407 10180 21419 10183
rect 21542 10180 21548 10192
rect 21407 10152 21548 10180
rect 21407 10149 21419 10152
rect 21361 10143 21419 10149
rect 21542 10140 21548 10152
rect 21600 10140 21606 10192
rect 22370 10140 22376 10192
rect 22428 10180 22434 10192
rect 25409 10183 25467 10189
rect 25409 10180 25421 10183
rect 22428 10152 25421 10180
rect 22428 10140 22434 10152
rect 25409 10149 25421 10152
rect 25455 10149 25467 10183
rect 25409 10143 25467 10149
rect 4706 10072 4712 10124
rect 4764 10112 4770 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4764 10084 4905 10112
rect 4764 10072 4770 10084
rect 4893 10081 4905 10084
rect 4939 10081 4951 10115
rect 8386 10112 8392 10124
rect 4893 10075 4951 10081
rect 5000 10084 8392 10112
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 3050 10044 3056 10056
rect 2963 10016 3056 10044
rect 2869 10007 2927 10013
rect 2406 9976 2412 9988
rect 2367 9948 2412 9976
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 2884 9976 2912 10007
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 5000 10044 5028 10084
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 12584 10084 14105 10112
rect 12584 10072 12590 10084
rect 14093 10081 14105 10084
rect 14139 10112 14151 10115
rect 15746 10112 15752 10124
rect 14139 10084 15752 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 16298 10112 16304 10124
rect 16259 10084 16304 10112
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10112 21327 10115
rect 22002 10112 22008 10124
rect 21315 10084 22008 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 23017 10115 23075 10121
rect 23017 10081 23029 10115
rect 23063 10112 23075 10115
rect 23474 10112 23480 10124
rect 23063 10084 23480 10112
rect 23063 10081 23075 10084
rect 23017 10075 23075 10081
rect 23474 10072 23480 10084
rect 23532 10072 23538 10124
rect 24765 10115 24823 10121
rect 24765 10081 24777 10115
rect 24811 10112 24823 10115
rect 25038 10112 25044 10124
rect 24811 10084 25044 10112
rect 24811 10081 24823 10084
rect 24765 10075 24823 10081
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 8662 10044 8668 10056
rect 4120 10016 5028 10044
rect 8623 10016 8668 10044
rect 4120 10004 4126 10016
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 10008 10016 10057 10044
rect 10008 10004 10014 10016
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10044 13047 10047
rect 13538 10044 13544 10056
rect 13035 10016 13544 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 13630 10004 13636 10056
rect 13688 10044 13694 10056
rect 19334 10044 19340 10056
rect 13688 10016 13733 10044
rect 19076 10016 19340 10044
rect 13688 10004 13694 10016
rect 3510 9976 3516 9988
rect 2884 9948 3516 9976
rect 3510 9936 3516 9948
rect 3568 9936 3574 9988
rect 8938 9936 8944 9988
rect 8996 9976 9002 9988
rect 9125 9979 9183 9985
rect 9125 9976 9137 9979
rect 8996 9948 9137 9976
rect 8996 9936 9002 9948
rect 9125 9945 9137 9948
rect 9171 9976 9183 9979
rect 9490 9976 9496 9988
rect 9171 9948 9496 9976
rect 9171 9945 9183 9948
rect 9125 9939 9183 9945
rect 9490 9936 9496 9948
rect 9548 9936 9554 9988
rect 16114 9976 16120 9988
rect 16075 9948 16120 9976
rect 16114 9936 16120 9948
rect 16172 9936 16178 9988
rect 3881 9911 3939 9917
rect 3881 9877 3893 9911
rect 3927 9908 3939 9911
rect 3970 9908 3976 9920
rect 3927 9880 3976 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 3970 9868 3976 9880
rect 4028 9868 4034 9920
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 5074 9908 5080 9920
rect 4755 9880 5080 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 8260 9880 9413 9908
rect 8260 9868 8266 9880
rect 9401 9877 9413 9880
rect 9447 9908 9459 9911
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9447 9880 9965 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9953 9877 9965 9880
rect 9999 9908 10011 9911
rect 10962 9908 10968 9920
rect 9999 9880 10968 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13446 9908 13452 9920
rect 13127 9880 13452 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 17678 9908 17684 9920
rect 17276 9880 17684 9908
rect 17276 9868 17282 9880
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 18414 9868 18420 9920
rect 18472 9908 18478 9920
rect 18874 9908 18880 9920
rect 18472 9880 18880 9908
rect 18472 9868 18478 9880
rect 18874 9868 18880 9880
rect 18932 9908 18938 9920
rect 19076 9917 19104 10016
rect 19334 10004 19340 10016
rect 19392 10044 19398 10056
rect 19797 10047 19855 10053
rect 19797 10044 19809 10047
rect 19392 10016 19809 10044
rect 19392 10004 19398 10016
rect 19797 10013 19809 10016
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 20254 10004 20260 10056
rect 20312 10044 20318 10056
rect 20349 10047 20407 10053
rect 20349 10044 20361 10047
rect 20312 10016 20361 10044
rect 20312 10004 20318 10016
rect 20349 10013 20361 10016
rect 20395 10044 20407 10047
rect 20625 10047 20683 10053
rect 20625 10044 20637 10047
rect 20395 10016 20637 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 20625 10013 20637 10016
rect 20671 10044 20683 10047
rect 20990 10044 20996 10056
rect 20671 10016 20996 10044
rect 20671 10013 20683 10016
rect 20625 10007 20683 10013
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21910 10044 21916 10056
rect 21591 10016 21916 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 20714 9936 20720 9988
rect 20772 9976 20778 9988
rect 21560 9976 21588 10007
rect 21910 10004 21916 10016
rect 21968 10004 21974 10056
rect 23198 10004 23204 10056
rect 23256 10044 23262 10056
rect 24854 10044 24860 10056
rect 23256 10016 23301 10044
rect 24815 10016 24860 10044
rect 23256 10004 23262 10016
rect 24854 10004 24860 10016
rect 24912 10004 24918 10056
rect 24946 10004 24952 10056
rect 25004 10044 25010 10056
rect 25004 10016 25049 10044
rect 25004 10004 25010 10016
rect 20772 9948 21588 9976
rect 20772 9936 20778 9948
rect 24026 9936 24032 9988
rect 24084 9976 24090 9988
rect 24578 9976 24584 9988
rect 24084 9948 24584 9976
rect 24084 9936 24090 9948
rect 24578 9936 24584 9948
rect 24636 9936 24642 9988
rect 19061 9911 19119 9917
rect 19061 9908 19073 9911
rect 18932 9880 19073 9908
rect 18932 9868 18938 9880
rect 19061 9877 19073 9880
rect 19107 9877 19119 9911
rect 19242 9908 19248 9920
rect 19203 9880 19248 9908
rect 19061 9871 19119 9877
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 20901 9911 20959 9917
rect 20901 9877 20913 9911
rect 20947 9908 20959 9911
rect 21726 9908 21732 9920
rect 20947 9880 21732 9908
rect 20947 9877 20959 9880
rect 20901 9871 20959 9877
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 22278 9868 22284 9920
rect 22336 9908 22342 9920
rect 22373 9911 22431 9917
rect 22373 9908 22385 9911
rect 22336 9880 22385 9908
rect 22336 9868 22342 9880
rect 22373 9877 22385 9880
rect 22419 9908 22431 9911
rect 23658 9908 23664 9920
rect 22419 9880 23664 9908
rect 22419 9877 22431 9880
rect 22373 9871 22431 9877
rect 23658 9868 23664 9880
rect 23716 9908 23722 9920
rect 23753 9911 23811 9917
rect 23753 9908 23765 9911
rect 23716 9880 23765 9908
rect 23716 9868 23722 9880
rect 23753 9877 23765 9880
rect 23799 9877 23811 9911
rect 23753 9871 23811 9877
rect 24397 9911 24455 9917
rect 24397 9877 24409 9911
rect 24443 9908 24455 9911
rect 24670 9908 24676 9920
rect 24443 9880 24676 9908
rect 24443 9877 24455 9880
rect 24397 9871 24455 9877
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 24854 9868 24860 9920
rect 24912 9908 24918 9920
rect 26050 9908 26056 9920
rect 24912 9880 26056 9908
rect 24912 9868 24918 9880
rect 26050 9868 26056 9880
rect 26108 9868 26114 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 3510 9704 3516 9716
rect 2976 9676 3516 9704
rect 1394 9636 1400 9648
rect 1355 9608 1400 9636
rect 1394 9596 1400 9608
rect 1452 9596 1458 9648
rect 2501 9639 2559 9645
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 2976 9636 3004 9676
rect 3510 9664 3516 9676
rect 3568 9704 3574 9716
rect 4246 9704 4252 9716
rect 3568 9676 4252 9704
rect 3568 9664 3574 9676
rect 4246 9664 4252 9676
rect 4304 9664 4310 9716
rect 4614 9704 4620 9716
rect 4575 9676 4620 9704
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 9677 9707 9735 9713
rect 9677 9704 9689 9707
rect 8720 9676 9689 9704
rect 8720 9664 8726 9676
rect 9677 9673 9689 9676
rect 9723 9704 9735 9707
rect 10042 9704 10048 9716
rect 9723 9676 10048 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 10229 9707 10287 9713
rect 10229 9673 10241 9707
rect 10275 9704 10287 9707
rect 10686 9704 10692 9716
rect 10275 9676 10692 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 11514 9704 11520 9716
rect 11112 9676 11520 9704
rect 11112 9664 11118 9676
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 12308 9676 12664 9704
rect 12308 9664 12314 9676
rect 2547 9608 3004 9636
rect 3053 9639 3111 9645
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3878 9636 3884 9648
rect 3099 9608 3884 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 5442 9636 5448 9648
rect 4571 9608 5448 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 1578 9528 1584 9580
rect 1636 9568 1642 9580
rect 1946 9568 1952 9580
rect 1636 9540 1952 9568
rect 1636 9528 1642 9540
rect 1946 9528 1952 9540
rect 2004 9528 2010 9580
rect 5184 9577 5212 9608
rect 5442 9596 5448 9608
rect 5500 9636 5506 9648
rect 5629 9639 5687 9645
rect 5629 9636 5641 9639
rect 5500 9608 5641 9636
rect 5500 9596 5506 9608
rect 5629 9605 5641 9608
rect 5675 9605 5687 9639
rect 5629 9599 5687 9605
rect 7285 9639 7343 9645
rect 7285 9605 7297 9639
rect 7331 9636 7343 9639
rect 7742 9636 7748 9648
rect 7331 9608 7748 9636
rect 7331 9605 7343 9608
rect 7285 9599 7343 9605
rect 7742 9596 7748 9608
rect 7800 9596 7806 9648
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 9125 9639 9183 9645
rect 9125 9636 9137 9639
rect 8904 9608 9137 9636
rect 8904 9596 8910 9608
rect 9125 9605 9137 9608
rect 9171 9605 9183 9639
rect 10060 9636 10088 9664
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 10060 9608 11989 9636
rect 9125 9599 9183 9605
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5215 9540 5249 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 2314 9500 2320 9512
rect 1903 9472 2320 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3476 9472 3525 9500
rect 3476 9460 3482 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3712 9500 3740 9531
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 10778 9568 10784 9580
rect 10739 9540 10784 9568
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 11992 9568 12020 9599
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12636 9636 12664 9676
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16853 9707 16911 9713
rect 16853 9704 16865 9707
rect 16632 9676 16865 9704
rect 16632 9664 16638 9676
rect 16853 9673 16865 9676
rect 16899 9704 16911 9707
rect 17773 9707 17831 9713
rect 17773 9704 17785 9707
rect 16899 9676 17785 9704
rect 16899 9673 16911 9676
rect 16853 9667 16911 9673
rect 17773 9673 17785 9676
rect 17819 9704 17831 9707
rect 19337 9707 19395 9713
rect 17819 9676 18184 9704
rect 17819 9673 17831 9676
rect 17773 9667 17831 9673
rect 12492 9608 12664 9636
rect 12492 9596 12498 9608
rect 12894 9596 12900 9648
rect 12952 9636 12958 9648
rect 12989 9639 13047 9645
rect 12989 9636 13001 9639
rect 12952 9608 13001 9636
rect 12952 9596 12958 9608
rect 12989 9605 13001 9608
rect 13035 9605 13047 9639
rect 12989 9599 13047 9605
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 15930 9636 15936 9648
rect 15887 9608 15936 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 12526 9568 12532 9580
rect 11992 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3712 9472 4169 9500
rect 3513 9463 3571 9469
rect 4157 9469 4169 9472
rect 4203 9500 4215 9503
rect 7392 9500 7420 9528
rect 4203 9472 7420 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7708 9472 7757 9500
rect 7708 9460 7714 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 7745 9463 7803 9469
rect 10594 9460 10600 9472
rect 10652 9500 10658 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 10652 9472 11621 9500
rect 10652 9460 10658 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 13004 9500 13032 9599
rect 15930 9596 15936 9608
rect 15988 9596 15994 9648
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 18012 9608 18061 9636
rect 18012 9596 18018 9608
rect 18049 9605 18061 9608
rect 18095 9605 18107 9639
rect 18156 9636 18184 9676
rect 19337 9673 19349 9707
rect 19383 9704 19395 9707
rect 19518 9704 19524 9716
rect 19383 9676 19524 9704
rect 19383 9673 19395 9676
rect 19337 9667 19395 9673
rect 19518 9664 19524 9676
rect 19576 9664 19582 9716
rect 22373 9707 22431 9713
rect 22373 9673 22385 9707
rect 22419 9704 22431 9707
rect 23014 9704 23020 9716
rect 22419 9676 23020 9704
rect 22419 9673 22431 9676
rect 22373 9667 22431 9673
rect 23014 9664 23020 9676
rect 23072 9704 23078 9716
rect 23934 9704 23940 9716
rect 23072 9676 23940 9704
rect 23072 9664 23078 9676
rect 23934 9664 23940 9676
rect 23992 9664 23998 9716
rect 24029 9707 24087 9713
rect 24029 9673 24041 9707
rect 24075 9704 24087 9707
rect 24854 9704 24860 9716
rect 24075 9676 24860 9704
rect 24075 9673 24087 9676
rect 24029 9667 24087 9673
rect 22649 9639 22707 9645
rect 18156 9608 18644 9636
rect 18049 9599 18107 9605
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 16393 9571 16451 9577
rect 16393 9568 16405 9571
rect 15712 9540 16405 9568
rect 15712 9528 15718 9540
rect 16393 9537 16405 9540
rect 16439 9537 16451 9571
rect 16393 9531 16451 9537
rect 17497 9571 17555 9577
rect 17497 9537 17509 9571
rect 17543 9568 17555 9571
rect 18506 9568 18512 9580
rect 17543 9540 18512 9568
rect 17543 9537 17555 9540
rect 17497 9531 17555 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18616 9577 18644 9608
rect 22649 9605 22661 9639
rect 22695 9636 22707 9639
rect 23290 9636 23296 9648
rect 22695 9608 23296 9636
rect 22695 9605 22707 9608
rect 22649 9599 22707 9605
rect 23290 9596 23296 9608
rect 23348 9596 23354 9648
rect 23382 9596 23388 9648
rect 23440 9636 23446 9648
rect 24044 9636 24072 9667
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 23440 9608 24072 9636
rect 23440 9596 23446 9608
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 23658 9528 23664 9580
rect 23716 9568 23722 9580
rect 24121 9571 24179 9577
rect 24121 9568 24133 9571
rect 23716 9540 24133 9568
rect 23716 9528 23722 9540
rect 24121 9537 24133 9540
rect 24167 9537 24179 9571
rect 24121 9531 24179 9537
rect 13173 9503 13231 9509
rect 13173 9500 13185 9503
rect 13004 9472 13185 9500
rect 11609 9463 11667 9469
rect 13173 9469 13185 9472
rect 13219 9469 13231 9503
rect 13173 9463 13231 9469
rect 16114 9460 16120 9512
rect 16172 9500 16178 9512
rect 16209 9503 16267 9509
rect 16209 9500 16221 9503
rect 16172 9472 16221 9500
rect 16172 9460 16178 9472
rect 16209 9469 16221 9472
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 17402 9500 17408 9512
rect 17184 9472 17408 9500
rect 17184 9460 17190 9472
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 18322 9460 18328 9512
rect 18380 9500 18386 9512
rect 18417 9503 18475 9509
rect 18417 9500 18429 9503
rect 18380 9472 18429 9500
rect 18380 9460 18386 9472
rect 18417 9469 18429 9472
rect 18463 9469 18475 9503
rect 18417 9463 18475 9469
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 18932 9472 19625 9500
rect 18932 9460 18938 9472
rect 19613 9469 19625 9472
rect 19659 9500 19671 9503
rect 21450 9500 21456 9512
rect 19659 9472 21456 9500
rect 19659 9469 19671 9472
rect 19613 9463 19671 9469
rect 21450 9460 21456 9472
rect 21508 9500 21514 9512
rect 22278 9500 22284 9512
rect 21508 9472 22284 9500
rect 21508 9460 21514 9472
rect 22278 9460 22284 9472
rect 22336 9460 22342 9512
rect 22462 9500 22468 9512
rect 22423 9472 22468 9500
rect 22462 9460 22468 9472
rect 22520 9500 22526 9512
rect 23017 9503 23075 9509
rect 23017 9500 23029 9503
rect 22520 9472 23029 9500
rect 22520 9460 22526 9472
rect 23017 9469 23029 9472
rect 23063 9469 23075 9503
rect 23017 9463 23075 9469
rect 24210 9460 24216 9512
rect 24268 9500 24274 9512
rect 24377 9503 24435 9509
rect 24377 9500 24389 9503
rect 24268 9472 24389 9500
rect 24268 9460 24274 9472
rect 24377 9469 24389 9472
rect 24423 9469 24435 9503
rect 24377 9463 24435 9469
rect 24946 9460 24952 9512
rect 25004 9500 25010 9512
rect 26053 9503 26111 9509
rect 26053 9500 26065 9503
rect 25004 9472 26065 9500
rect 25004 9460 25010 9472
rect 26053 9469 26065 9472
rect 26099 9469 26111 9503
rect 26053 9463 26111 9469
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 2222 9432 2228 9444
rect 1811 9404 2228 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 2222 9392 2228 9404
rect 2280 9392 2286 9444
rect 4985 9435 5043 9441
rect 4985 9401 4997 9435
rect 5031 9432 5043 9435
rect 5350 9432 5356 9444
rect 5031 9404 5356 9432
rect 5031 9401 5043 9404
rect 4985 9395 5043 9401
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 7006 9392 7012 9444
rect 7064 9432 7070 9444
rect 7834 9432 7840 9444
rect 7064 9404 7840 9432
rect 7064 9392 7070 9404
rect 7834 9392 7840 9404
rect 7892 9432 7898 9444
rect 7990 9435 8048 9441
rect 7990 9432 8002 9435
rect 7892 9404 8002 9432
rect 7892 9392 7898 9404
rect 7990 9401 8002 9404
rect 8036 9401 8048 9435
rect 7990 9395 8048 9401
rect 12713 9435 12771 9441
rect 12713 9401 12725 9435
rect 12759 9432 12771 9435
rect 13630 9432 13636 9444
rect 12759 9404 13636 9432
rect 12759 9401 12771 9404
rect 12713 9395 12771 9401
rect 13630 9392 13636 9404
rect 13688 9392 13694 9444
rect 14918 9432 14924 9444
rect 14879 9404 14924 9432
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 16301 9435 16359 9441
rect 16301 9432 16313 9435
rect 15304 9404 16313 9432
rect 15304 9376 15332 9404
rect 16301 9401 16313 9404
rect 16347 9401 16359 9435
rect 16301 9395 16359 9401
rect 19880 9435 19938 9441
rect 19880 9401 19892 9435
rect 19926 9432 19938 9435
rect 20254 9432 20260 9444
rect 19926 9404 20260 9432
rect 19926 9401 19938 9404
rect 19880 9395 19938 9401
rect 20254 9392 20260 9404
rect 20312 9392 20318 9444
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 3292 9336 3433 9364
rect 3292 9324 3298 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 5074 9364 5080 9376
rect 5035 9336 5080 9364
rect 3421 9327 3479 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6549 9367 6607 9373
rect 6549 9333 6561 9367
rect 6595 9364 6607 9367
rect 6730 9364 6736 9376
rect 6595 9336 6736 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 10744 9336 11253 9364
rect 10744 9324 10750 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 15286 9364 15292 9376
rect 15247 9336 15292 9364
rect 11241 9327 11299 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 15654 9364 15660 9376
rect 15615 9336 15660 9364
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 18046 9364 18052 9376
rect 17092 9336 18052 9364
rect 17092 9324 17098 9336
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 20990 9364 20996 9376
rect 20951 9336 20996 9364
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 21542 9364 21548 9376
rect 21503 9336 21548 9364
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 21910 9364 21916 9376
rect 21871 9336 21916 9364
rect 21910 9324 21916 9336
rect 21968 9324 21974 9376
rect 23474 9364 23480 9376
rect 23435 9336 23480 9364
rect 23474 9324 23480 9336
rect 23532 9324 23538 9376
rect 25498 9364 25504 9376
rect 25459 9336 25504 9364
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1397 9163 1455 9169
rect 1397 9129 1409 9163
rect 1443 9160 1455 9163
rect 1854 9160 1860 9172
rect 1443 9132 1860 9160
rect 1443 9129 1455 9132
rect 1397 9123 1455 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2409 9163 2467 9169
rect 2004 9132 2049 9160
rect 2004 9120 2010 9132
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2590 9160 2596 9172
rect 2455 9132 2596 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 5537 9163 5595 9169
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 6086 9160 6092 9172
rect 5583 9132 6092 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 7834 9120 7840 9172
rect 7892 9160 7898 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 7892 9132 8493 9160
rect 7892 9120 7898 9132
rect 8481 9129 8493 9132
rect 8527 9129 8539 9163
rect 8481 9123 8539 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 10192 9132 10425 9160
rect 10192 9120 10198 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 10413 9123 10471 9129
rect 10778 9120 10784 9172
rect 10836 9120 10842 9172
rect 12342 9120 12348 9172
rect 12400 9120 12406 9172
rect 14642 9120 14648 9172
rect 14700 9160 14706 9172
rect 15378 9160 15384 9172
rect 14700 9132 15384 9160
rect 14700 9120 14706 9132
rect 15378 9120 15384 9132
rect 15436 9120 15442 9172
rect 16758 9120 16764 9172
rect 16816 9160 16822 9172
rect 17129 9163 17187 9169
rect 17129 9160 17141 9163
rect 16816 9132 17141 9160
rect 16816 9120 16822 9132
rect 17129 9129 17141 9132
rect 17175 9129 17187 9163
rect 17129 9123 17187 9129
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 18322 9160 18328 9172
rect 17635 9132 18328 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 18322 9120 18328 9132
rect 18380 9120 18386 9172
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 18472 9132 18705 9160
rect 18472 9120 18478 9132
rect 18693 9129 18705 9132
rect 18739 9129 18751 9163
rect 18693 9123 18751 9129
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 19245 9163 19303 9169
rect 19245 9160 19257 9163
rect 18840 9132 19257 9160
rect 18840 9120 18846 9132
rect 19245 9129 19257 9132
rect 19291 9129 19303 9163
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 19245 9123 19303 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 21266 9160 21272 9172
rect 21227 9132 21272 9160
rect 21266 9120 21272 9132
rect 21324 9160 21330 9172
rect 22094 9160 22100 9172
rect 21324 9132 22100 9160
rect 21324 9120 21330 9132
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22741 9163 22799 9169
rect 22741 9129 22753 9163
rect 22787 9160 22799 9163
rect 23198 9160 23204 9172
rect 22787 9132 23204 9160
rect 22787 9129 22799 9132
rect 22741 9123 22799 9129
rect 23198 9120 23204 9132
rect 23256 9160 23262 9172
rect 24489 9163 24547 9169
rect 24489 9160 24501 9163
rect 23256 9132 24501 9160
rect 23256 9120 23262 9132
rect 24489 9129 24501 9132
rect 24535 9129 24547 9163
rect 24489 9123 24547 9129
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 3786 9092 3792 9104
rect 2832 9064 3792 9092
rect 2832 9052 2838 9064
rect 3786 9052 3792 9064
rect 3844 9052 3850 9104
rect 5994 9092 6000 9104
rect 5955 9064 6000 9092
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 7368 9095 7426 9101
rect 7368 9061 7380 9095
rect 7414 9092 7426 9095
rect 8018 9092 8024 9104
rect 7414 9064 8024 9092
rect 7414 9061 7426 9064
rect 7368 9055 7426 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 10321 9095 10379 9101
rect 10321 9061 10333 9095
rect 10367 9092 10379 9095
rect 10796 9092 10824 9120
rect 10367 9064 11008 9092
rect 10367 9061 10379 9064
rect 10321 9055 10379 9061
rect 2130 8984 2136 9036
rect 2188 9024 2194 9036
rect 2317 9027 2375 9033
rect 2317 9024 2329 9027
rect 2188 8996 2329 9024
rect 2188 8984 2194 8996
rect 2317 8993 2329 8996
rect 2363 9024 2375 9027
rect 5905 9027 5963 9033
rect 2363 8996 3004 9024
rect 2363 8993 2375 8996
rect 2317 8987 2375 8993
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 2976 8956 3004 8996
rect 5905 8993 5917 9027
rect 5951 9024 5963 9027
rect 6454 9024 6460 9036
rect 5951 8996 6460 9024
rect 5951 8993 5963 8996
rect 5905 8987 5963 8993
rect 6454 8984 6460 8996
rect 6512 9024 6518 9036
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 6512 8996 9045 9024
rect 6512 8984 6518 8996
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 9033 8987 9091 8993
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10778 9024 10784 9036
rect 9999 8996 10784 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10980 8968 11008 9064
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12360 9033 12388 9120
rect 12437 9095 12495 9101
rect 12437 9061 12449 9095
rect 12483 9092 12495 9095
rect 15838 9092 15844 9104
rect 12483 9064 15844 9092
rect 12483 9061 12495 9064
rect 12437 9055 12495 9061
rect 12345 9027 12403 9033
rect 12345 9024 12357 9027
rect 12032 8996 12357 9024
rect 12032 8984 12038 8996
rect 12345 8993 12357 8996
rect 12391 8993 12403 9027
rect 12345 8987 12403 8993
rect 3050 8956 3056 8968
rect 2963 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8956 3114 8968
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 3108 8928 4353 8956
rect 3108 8916 3114 8928
rect 4341 8925 4353 8928
rect 4387 8925 4399 8959
rect 4522 8956 4528 8968
rect 4483 8928 4528 8956
rect 4341 8919 4399 8925
rect 2590 8848 2596 8900
rect 2648 8888 2654 8900
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 2648 8860 3801 8888
rect 2648 8848 2654 8860
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 4356 8888 4384 8919
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 6086 8956 6092 8968
rect 6047 8928 6092 8956
rect 6086 8916 6092 8928
rect 6144 8956 6150 8968
rect 7006 8956 7012 8968
rect 6144 8928 7012 8956
rect 6144 8916 6150 8928
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 10870 8956 10876 8968
rect 7156 8928 7201 8956
rect 10831 8928 10876 8956
rect 7156 8916 7162 8928
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 12526 8956 12532 8968
rect 11020 8928 11113 8956
rect 12487 8928 12532 8956
rect 11020 8916 11026 8928
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 4890 8888 4896 8900
rect 4356 8860 4896 8888
rect 3789 8851 3847 8857
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 10888 8888 10916 8916
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 10888 8860 11989 8888
rect 11977 8857 11989 8860
rect 12023 8857 12035 8891
rect 11977 8851 12035 8857
rect 3418 8820 3424 8832
rect 3379 8792 3424 8820
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 4062 8820 4068 8832
rect 3568 8792 4068 8820
rect 3568 8780 3574 8792
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4982 8820 4988 8832
rect 4943 8792 4988 8820
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5350 8820 5356 8832
rect 5311 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 7098 8820 7104 8832
rect 6963 8792 7104 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9401 8823 9459 8829
rect 9401 8820 9413 8823
rect 9180 8792 9413 8820
rect 9180 8780 9186 8792
rect 9401 8789 9413 8792
rect 9447 8789 9459 8823
rect 9401 8783 9459 8789
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11514 8820 11520 8832
rect 11204 8792 11520 8820
rect 11204 8780 11210 8792
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11756 8792 11897 8820
rect 11756 8780 11762 8792
rect 11885 8789 11897 8792
rect 11931 8820 11943 8823
rect 12636 8820 12664 9064
rect 15838 9052 15844 9064
rect 15896 9052 15902 9104
rect 18046 9092 18052 9104
rect 18007 9064 18052 9092
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 18138 9052 18144 9104
rect 18196 9092 18202 9104
rect 19058 9092 19064 9104
rect 18196 9064 18241 9092
rect 19019 9064 19064 9092
rect 18196 9052 18202 9064
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 23658 9092 23664 9104
rect 23124 9064 23664 9092
rect 13630 9033 13636 9036
rect 13624 9024 13636 9033
rect 13543 8996 13636 9024
rect 13624 8987 13636 8996
rect 13688 9024 13694 9036
rect 15378 9024 15384 9036
rect 13688 8996 15384 9024
rect 13630 8984 13636 8987
rect 13688 8984 13694 8996
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 16482 9024 16488 9036
rect 16443 8996 16488 9024
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19613 9027 19671 9033
rect 19613 9024 19625 9027
rect 19392 8996 19625 9024
rect 19392 8984 19398 8996
rect 19613 8993 19625 8996
rect 19659 9024 19671 9027
rect 19659 8996 19840 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13228 8928 13369 8956
rect 13228 8916 13234 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 16022 8916 16028 8968
rect 16080 8956 16086 8968
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16080 8928 16589 8956
rect 16080 8916 16086 8928
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 16577 8919 16635 8925
rect 16669 8959 16727 8965
rect 16669 8925 16681 8959
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8956 18383 8959
rect 18598 8956 18604 8968
rect 18371 8928 18604 8956
rect 18371 8925 18383 8928
rect 18325 8919 18383 8925
rect 16684 8888 16712 8919
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19576 8928 19717 8956
rect 19576 8916 19582 8928
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 15948 8860 16712 8888
rect 15948 8832 15976 8860
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 17681 8891 17739 8897
rect 17681 8888 17693 8891
rect 16908 8860 17693 8888
rect 16908 8848 16914 8860
rect 17681 8857 17693 8860
rect 17727 8857 17739 8891
rect 19812 8888 19840 8996
rect 20254 8984 20260 9036
rect 20312 9024 20318 9036
rect 21082 9024 21088 9036
rect 20312 8996 21088 9024
rect 20312 8984 20318 8996
rect 21082 8984 21088 8996
rect 21140 9024 21146 9036
rect 23124 9033 23152 9064
rect 23658 9052 23664 9064
rect 23716 9092 23722 9104
rect 25409 9095 25467 9101
rect 25409 9092 25421 9095
rect 23716 9064 25421 9092
rect 23716 9052 23722 9064
rect 25409 9061 25421 9064
rect 25455 9092 25467 9095
rect 25590 9092 25596 9104
rect 25455 9064 25596 9092
rect 25455 9061 25467 9064
rect 25409 9055 25467 9061
rect 25590 9052 25596 9064
rect 25648 9052 25654 9104
rect 23382 9033 23388 9036
rect 23109 9027 23167 9033
rect 21140 8996 21496 9024
rect 21140 8984 21146 8996
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20162 8956 20168 8968
rect 19935 8928 20168 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20162 8916 20168 8928
rect 20220 8956 20226 8968
rect 20990 8956 20996 8968
rect 20220 8928 20996 8956
rect 20220 8916 20226 8928
rect 20990 8916 20996 8928
rect 21048 8916 21054 8968
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 21468 8965 21496 8996
rect 23109 8993 23121 9027
rect 23155 8993 23167 9027
rect 23376 9024 23388 9033
rect 23343 8996 23388 9024
rect 23109 8987 23167 8993
rect 23376 8987 23388 8996
rect 23382 8984 23388 8987
rect 23440 8984 23446 9036
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 20901 8891 20959 8897
rect 20901 8888 20913 8891
rect 19812 8860 20913 8888
rect 17681 8851 17739 8857
rect 20901 8857 20913 8860
rect 20947 8857 20959 8891
rect 21376 8888 21404 8916
rect 22281 8891 22339 8897
rect 22281 8888 22293 8891
rect 21376 8860 22293 8888
rect 20901 8851 20959 8857
rect 22281 8857 22293 8860
rect 22327 8857 22339 8891
rect 22281 8851 22339 8857
rect 25774 8848 25780 8900
rect 25832 8888 25838 8900
rect 25958 8888 25964 8900
rect 25832 8860 25964 8888
rect 25832 8848 25838 8860
rect 25958 8848 25964 8860
rect 26016 8848 26022 8900
rect 11931 8792 12664 8820
rect 13265 8823 13323 8829
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 13265 8789 13277 8823
rect 13311 8820 13323 8823
rect 13998 8820 14004 8832
rect 13311 8792 14004 8820
rect 13311 8789 13323 8792
rect 13265 8783 13323 8789
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 14826 8820 14832 8832
rect 14783 8792 14832 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 14826 8780 14832 8792
rect 14884 8820 14890 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 14884 8792 15485 8820
rect 14884 8780 14890 8792
rect 15473 8789 15485 8792
rect 15519 8789 15531 8823
rect 15930 8820 15936 8832
rect 15891 8792 15936 8820
rect 15473 8783 15531 8789
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 16114 8820 16120 8832
rect 16075 8792 16120 8820
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 20714 8820 20720 8832
rect 20675 8792 20720 8820
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 21266 8780 21272 8832
rect 21324 8820 21330 8832
rect 21913 8823 21971 8829
rect 21913 8820 21925 8823
rect 21324 8792 21925 8820
rect 21324 8780 21330 8792
rect 21913 8789 21925 8792
rect 21959 8789 21971 8823
rect 25038 8820 25044 8832
rect 24999 8792 25044 8820
rect 21913 8783 21971 8789
rect 25038 8780 25044 8792
rect 25096 8780 25102 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2866 8616 2872 8628
rect 1811 8588 2872 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2866 8576 2872 8588
rect 2924 8616 2930 8628
rect 3602 8616 3608 8628
rect 2924 8588 3608 8616
rect 2924 8576 2930 8588
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 3786 8616 3792 8628
rect 3747 8588 3792 8616
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 6086 8616 6092 8628
rect 5675 8588 6092 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6362 8616 6368 8628
rect 6236 8588 6368 8616
rect 6236 8576 6242 8588
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 8202 8616 8208 8628
rect 7024 8588 8208 8616
rect 3237 8551 3295 8557
rect 3237 8517 3249 8551
rect 3283 8548 3295 8551
rect 3326 8548 3332 8560
rect 3283 8520 3332 8548
rect 3283 8517 3295 8520
rect 3237 8511 3295 8517
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 4338 8548 4344 8560
rect 4299 8520 4344 8548
rect 4338 8508 4344 8520
rect 4396 8508 4402 8560
rect 7024 8492 7052 8588
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 9582 8616 9588 8628
rect 9263 8588 9588 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10042 8616 10048 8628
rect 9999 8588 10048 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10042 8576 10048 8588
rect 10100 8576 10106 8628
rect 10413 8619 10471 8625
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10686 8616 10692 8628
rect 10459 8588 10692 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13538 8616 13544 8628
rect 12492 8588 12537 8616
rect 13499 8588 13544 8616
rect 12492 8576 12498 8588
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 15378 8616 15384 8628
rect 15339 8588 15384 8616
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15841 8619 15899 8625
rect 15841 8585 15853 8619
rect 15887 8616 15899 8619
rect 16850 8616 16856 8628
rect 15887 8588 16856 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 17773 8619 17831 8625
rect 17773 8585 17785 8619
rect 17819 8616 17831 8619
rect 18046 8616 18052 8628
rect 17819 8588 18052 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 18233 8619 18291 8625
rect 18233 8616 18245 8619
rect 18196 8588 18245 8616
rect 18196 8576 18202 8588
rect 18233 8585 18245 8588
rect 18279 8585 18291 8619
rect 18598 8616 18604 8628
rect 18559 8588 18604 8616
rect 18233 8579 18291 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 20349 8619 20407 8625
rect 20349 8616 20361 8619
rect 20312 8588 20361 8616
rect 20312 8576 20318 8588
rect 20349 8585 20361 8588
rect 20395 8585 20407 8619
rect 20349 8579 20407 8585
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 21910 8616 21916 8628
rect 21416 8588 21916 8616
rect 21416 8576 21422 8588
rect 21910 8576 21916 8588
rect 21968 8576 21974 8628
rect 25590 8616 25596 8628
rect 25551 8588 25596 8616
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 8018 8508 8024 8560
rect 8076 8548 8082 8560
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 8076 8520 8401 8548
rect 8076 8508 8082 8520
rect 8389 8517 8401 8520
rect 8435 8517 8447 8551
rect 10060 8548 10088 8576
rect 10060 8520 11008 8548
rect 8389 8511 8447 8517
rect 4890 8480 4896 8492
rect 4851 8452 4896 8480
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 7006 8480 7012 8492
rect 6919 8452 7012 8480
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 10870 8480 10876 8492
rect 9631 8452 10876 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 10980 8489 11008 8520
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 14369 8551 14427 8557
rect 14369 8548 14381 8551
rect 13872 8520 14381 8548
rect 13872 8508 13878 8520
rect 14369 8517 14381 8520
rect 14415 8517 14427 8551
rect 14369 8511 14427 8517
rect 14550 8508 14556 8560
rect 14608 8548 14614 8560
rect 14826 8548 14832 8560
rect 14608 8520 14832 8548
rect 14608 8508 14614 8520
rect 14826 8508 14832 8520
rect 14884 8548 14890 8560
rect 14884 8520 14964 8548
rect 14884 8508 14890 8520
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12584 8452 13001 8480
rect 12584 8440 12590 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14936 8489 14964 8520
rect 20622 8508 20628 8560
rect 20680 8548 20686 8560
rect 21453 8551 21511 8557
rect 21453 8548 21465 8551
rect 20680 8520 21465 8548
rect 20680 8508 20686 8520
rect 21453 8517 21465 8520
rect 21499 8517 21511 8551
rect 21453 8511 21511 8517
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13780 8452 14105 8480
rect 13780 8440 13786 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8449 14979 8483
rect 16942 8480 16948 8492
rect 16903 8452 16948 8480
rect 14921 8443 14979 8449
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 18969 8483 19027 8489
rect 18969 8480 18981 8483
rect 18932 8452 18981 8480
rect 18932 8440 18938 8452
rect 18969 8449 18981 8452
rect 19015 8449 19027 8483
rect 18969 8443 19027 8449
rect 21266 8440 21272 8492
rect 21324 8480 21330 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21324 8452 22017 8480
rect 21324 8440 21330 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 23658 8480 23664 8492
rect 23619 8452 23664 8480
rect 22005 8443 22063 8449
rect 23658 8440 23664 8452
rect 23716 8440 23722 8492
rect 2130 8421 2136 8424
rect 1857 8415 1915 8421
rect 1857 8381 1869 8415
rect 1903 8381 1915 8415
rect 2124 8412 2136 8421
rect 2091 8384 2136 8412
rect 1857 8375 1915 8381
rect 2124 8375 2136 8384
rect 1872 8344 1900 8375
rect 2130 8372 2136 8375
rect 2188 8372 2194 8424
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4706 8412 4712 8424
rect 4295 8384 4712 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 6638 8412 6644 8424
rect 6551 8384 6644 8412
rect 6638 8372 6644 8384
rect 6696 8412 6702 8424
rect 7282 8421 7288 8424
rect 7276 8412 7288 8421
rect 6696 8384 7288 8412
rect 6696 8372 6702 8384
rect 7276 8375 7288 8384
rect 7282 8372 7288 8375
rect 7340 8372 7346 8424
rect 9766 8412 9772 8424
rect 9679 8384 9772 8412
rect 2314 8344 2320 8356
rect 1872 8316 2320 8344
rect 2314 8304 2320 8316
rect 2372 8304 2378 8356
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 4801 8347 4859 8353
rect 4801 8344 4813 8347
rect 4212 8316 4813 8344
rect 4212 8304 4218 8316
rect 4801 8313 4813 8316
rect 4847 8344 4859 8347
rect 5442 8344 5448 8356
rect 4847 8316 5448 8344
rect 4847 8313 4859 8316
rect 4801 8307 4859 8313
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 9692 8344 9720 8384
rect 9766 8372 9772 8384
rect 9824 8412 9830 8424
rect 10229 8415 10287 8421
rect 10229 8412 10241 8415
rect 9824 8384 10241 8412
rect 9824 8372 9830 8384
rect 10229 8381 10241 8384
rect 10275 8412 10287 8415
rect 13998 8412 14004 8424
rect 10275 8384 10916 8412
rect 13959 8384 14004 8412
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 9600 8316 9720 8344
rect 6273 8279 6331 8285
rect 6273 8245 6285 8279
rect 6319 8276 6331 8279
rect 6362 8276 6368 8288
rect 6319 8248 6368 8276
rect 6319 8245 6331 8248
rect 6273 8239 6331 8245
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 8478 8236 8484 8288
rect 8536 8276 8542 8288
rect 9600 8276 9628 8316
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10778 8344 10784 8356
rect 10192 8316 10784 8344
rect 10192 8304 10198 8316
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 10888 8353 10916 8384
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8412 14795 8415
rect 14826 8412 14832 8424
rect 14783 8384 14832 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 14826 8372 14832 8384
rect 14884 8372 14890 8424
rect 16758 8412 16764 8424
rect 16719 8384 16764 8412
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 16908 8384 16953 8412
rect 16908 8372 16914 8384
rect 18414 8372 18420 8424
rect 18472 8412 18478 8424
rect 19225 8415 19283 8421
rect 19225 8412 19237 8415
rect 18472 8384 19237 8412
rect 18472 8372 18478 8384
rect 19225 8381 19237 8384
rect 19271 8412 19283 8415
rect 20993 8415 21051 8421
rect 19271 8381 19288 8412
rect 19225 8375 19288 8381
rect 20993 8381 21005 8415
rect 21039 8412 21051 8415
rect 21821 8415 21879 8421
rect 21821 8412 21833 8415
rect 21039 8384 21833 8412
rect 21039 8381 21051 8384
rect 20993 8375 21051 8381
rect 21821 8381 21833 8384
rect 21867 8412 21879 8415
rect 22278 8412 22284 8424
rect 21867 8384 22284 8412
rect 21867 8381 21879 8384
rect 21821 8375 21879 8381
rect 10873 8347 10931 8353
rect 10873 8313 10885 8347
rect 10919 8313 10931 8347
rect 10873 8307 10931 8313
rect 11701 8347 11759 8353
rect 11701 8313 11713 8347
rect 11747 8344 11759 8347
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 11747 8316 12909 8344
rect 11747 8313 11759 8316
rect 11701 8307 11759 8313
rect 12897 8313 12909 8316
rect 12943 8344 12955 8347
rect 13354 8344 13360 8356
rect 12943 8316 13360 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 13906 8344 13912 8356
rect 13867 8316 13912 8344
rect 13906 8304 13912 8316
rect 13964 8304 13970 8356
rect 15654 8304 15660 8356
rect 15712 8344 15718 8356
rect 16117 8347 16175 8353
rect 16117 8344 16129 8347
rect 15712 8316 16129 8344
rect 15712 8304 15718 8316
rect 16117 8313 16129 8316
rect 16163 8344 16175 8347
rect 16482 8344 16488 8356
rect 16163 8316 16488 8344
rect 16163 8313 16175 8316
rect 16117 8307 16175 8313
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 19260 8344 19288 8375
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 22738 8412 22744 8424
rect 22664 8384 22744 8412
rect 19334 8344 19340 8356
rect 19260 8316 19340 8344
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 21361 8347 21419 8353
rect 21361 8313 21373 8347
rect 21407 8344 21419 8347
rect 21913 8347 21971 8353
rect 21913 8344 21925 8347
rect 21407 8316 21925 8344
rect 21407 8313 21419 8316
rect 21361 8307 21419 8313
rect 21913 8313 21925 8316
rect 21959 8344 21971 8347
rect 22664 8344 22692 8384
rect 22738 8372 22744 8384
rect 22796 8412 22802 8424
rect 26234 8412 26240 8424
rect 22796 8384 26240 8412
rect 22796 8372 22802 8384
rect 26234 8372 26240 8384
rect 26292 8372 26298 8424
rect 23906 8347 23964 8353
rect 23906 8344 23918 8347
rect 21959 8316 22692 8344
rect 22756 8316 23918 8344
rect 21959 8313 21971 8316
rect 21913 8307 21971 8313
rect 11974 8276 11980 8288
rect 8536 8248 9628 8276
rect 11935 8248 11980 8276
rect 8536 8236 8542 8248
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 12805 8279 12863 8285
rect 12805 8276 12817 8279
rect 12768 8248 12817 8276
rect 12768 8236 12774 8248
rect 12805 8245 12817 8248
rect 12851 8245 12863 8279
rect 12805 8239 12863 8245
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 14829 8279 14887 8285
rect 14829 8276 14841 8279
rect 14516 8248 14841 8276
rect 14516 8236 14522 8248
rect 14829 8245 14841 8248
rect 14875 8245 14887 8279
rect 14829 8239 14887 8245
rect 16393 8279 16451 8285
rect 16393 8245 16405 8279
rect 16439 8276 16451 8279
rect 16758 8276 16764 8288
rect 16439 8248 16764 8276
rect 16439 8245 16451 8248
rect 16393 8239 16451 8245
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 22646 8236 22652 8288
rect 22704 8276 22710 8288
rect 22756 8285 22784 8316
rect 23906 8313 23918 8316
rect 23952 8313 23964 8347
rect 23906 8307 23964 8313
rect 22741 8279 22799 8285
rect 22741 8276 22753 8279
rect 22704 8248 22753 8276
rect 22704 8236 22710 8248
rect 22741 8245 22753 8248
rect 22787 8245 22799 8279
rect 22741 8239 22799 8245
rect 23201 8279 23259 8285
rect 23201 8245 23213 8279
rect 23247 8276 23259 8279
rect 23382 8276 23388 8288
rect 23247 8248 23388 8276
rect 23247 8245 23259 8248
rect 23201 8239 23259 8245
rect 23382 8236 23388 8248
rect 23440 8276 23446 8288
rect 23658 8276 23664 8288
rect 23440 8248 23664 8276
rect 23440 8236 23446 8248
rect 23658 8236 23664 8248
rect 23716 8276 23722 8288
rect 25041 8279 25099 8285
rect 25041 8276 25053 8279
rect 23716 8248 25053 8276
rect 23716 8236 23722 8248
rect 25041 8245 25053 8248
rect 25087 8245 25099 8279
rect 25041 8239 25099 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2130 8072 2136 8084
rect 1995 8044 2136 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2130 8032 2136 8044
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2406 8072 2412 8084
rect 2367 8044 2412 8072
rect 2225 8035 2283 8041
rect 2240 8004 2268 8035
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4522 8072 4528 8084
rect 3927 8044 4528 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4522 8032 4528 8044
rect 4580 8072 4586 8084
rect 4893 8075 4951 8081
rect 4893 8072 4905 8075
rect 4580 8044 4905 8072
rect 4580 8032 4586 8044
rect 4893 8041 4905 8044
rect 4939 8041 4951 8075
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 4893 8035 4951 8041
rect 5534 8032 5540 8044
rect 5592 8072 5598 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5592 8044 5917 8072
rect 5592 8032 5598 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 5905 8035 5963 8041
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6328 8044 6837 8072
rect 6328 8032 6334 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7248 8044 7849 8072
rect 7248 8032 7254 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 10413 8075 10471 8081
rect 10413 8072 10425 8075
rect 10192 8044 10425 8072
rect 10192 8032 10198 8044
rect 10413 8041 10425 8044
rect 10459 8041 10471 8075
rect 10413 8035 10471 8041
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 10962 8072 10968 8084
rect 10919 8044 10968 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 12345 8075 12403 8081
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12526 8072 12532 8084
rect 12391 8044 12532 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13357 8075 13415 8081
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13906 8072 13912 8084
rect 13403 8044 13912 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 2240 7976 3096 8004
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 2958 7936 2964 7948
rect 2823 7908 2964 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 2866 7868 2872 7880
rect 2827 7840 2872 7868
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3068 7877 3096 7976
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4341 8007 4399 8013
rect 4341 8004 4353 8007
rect 4212 7976 4353 8004
rect 4212 7964 4218 7976
rect 4341 7973 4353 7976
rect 4387 7973 4399 8007
rect 4341 7967 4399 7973
rect 7561 8007 7619 8013
rect 7561 7973 7573 8007
rect 7607 8004 7619 8007
rect 8018 8004 8024 8016
rect 7607 7976 8024 8004
rect 7607 7973 7619 7976
rect 7561 7967 7619 7973
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 3878 7936 3884 7948
rect 3559 7908 3884 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3878 7896 3884 7908
rect 3936 7896 3942 7948
rect 5258 7936 5264 7948
rect 5000 7908 5264 7936
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3234 7868 3240 7880
rect 3099 7840 3240 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 5000 7877 5028 7908
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 4985 7871 5043 7877
rect 4985 7868 4997 7871
rect 4488 7840 4997 7868
rect 4488 7828 4494 7840
rect 4985 7837 4997 7840
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5534 7868 5540 7880
rect 5215 7840 5540 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6788 7840 6929 7868
rect 6788 7828 6794 7840
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7868 7159 7871
rect 7374 7868 7380 7880
rect 7147 7840 7380 7868
rect 7147 7837 7159 7840
rect 7101 7831 7159 7837
rect 7374 7828 7380 7840
rect 7432 7868 7438 7880
rect 7576 7868 7604 7967
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 11146 7964 11152 8016
rect 11204 8013 11210 8016
rect 11204 8007 11268 8013
rect 11204 7973 11222 8007
rect 11256 7973 11268 8007
rect 11204 7967 11268 7973
rect 11204 7964 11210 7967
rect 11422 7964 11428 8016
rect 11480 8004 11486 8016
rect 13372 8004 13400 8035
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 14458 8072 14464 8084
rect 14419 8044 14464 8072
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 14792 8044 15301 8072
rect 14792 8032 14798 8044
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 15289 8035 15347 8041
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 16080 8044 16129 8072
rect 16080 8032 16086 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 17552 8044 17693 8072
rect 17552 8032 17558 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 19058 8072 19064 8084
rect 19019 8044 19064 8072
rect 17681 8035 17739 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19150 8032 19156 8084
rect 19208 8072 19214 8084
rect 19429 8075 19487 8081
rect 19429 8072 19441 8075
rect 19208 8044 19441 8072
rect 19208 8032 19214 8044
rect 19429 8041 19441 8044
rect 19475 8072 19487 8075
rect 19978 8072 19984 8084
rect 19475 8044 19984 8072
rect 19475 8041 19487 8044
rect 19429 8035 19487 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20162 8072 20168 8084
rect 20123 8044 20168 8072
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20533 8075 20591 8081
rect 20533 8041 20545 8075
rect 20579 8072 20591 8075
rect 20622 8072 20628 8084
rect 20579 8044 20628 8072
rect 20579 8041 20591 8044
rect 20533 8035 20591 8041
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 21082 8072 21088 8084
rect 21043 8044 21088 8072
rect 21082 8032 21088 8044
rect 21140 8032 21146 8084
rect 21174 8032 21180 8084
rect 21232 8072 21238 8084
rect 21634 8072 21640 8084
rect 21232 8044 21640 8072
rect 21232 8032 21238 8044
rect 21634 8032 21640 8044
rect 21692 8072 21698 8084
rect 21913 8075 21971 8081
rect 21913 8072 21925 8075
rect 21692 8044 21925 8072
rect 21692 8032 21698 8044
rect 21913 8041 21925 8044
rect 21959 8041 21971 8075
rect 21913 8035 21971 8041
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22152 8044 22937 8072
rect 22152 8032 22158 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 23109 8075 23167 8081
rect 23109 8041 23121 8075
rect 23155 8041 23167 8075
rect 23109 8035 23167 8041
rect 14826 8004 14832 8016
rect 11480 7976 13400 8004
rect 14787 7976 14832 8004
rect 11480 7964 11486 7976
rect 14826 7964 14832 7976
rect 14884 7964 14890 8016
rect 18325 8007 18383 8013
rect 18325 7973 18337 8007
rect 18371 8004 18383 8007
rect 19518 8004 19524 8016
rect 18371 7976 19524 8004
rect 18371 7973 18383 7976
rect 18325 7967 18383 7973
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 20714 7964 20720 8016
rect 20772 8004 20778 8016
rect 20772 7976 22048 8004
rect 20772 7964 20778 7976
rect 8386 7936 8392 7948
rect 8347 7908 8392 7936
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10962 7936 10968 7948
rect 9824 7908 10968 7936
rect 9824 7896 9830 7908
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 13814 7936 13820 7948
rect 13775 7908 13820 7936
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 13964 7908 14009 7936
rect 13964 7896 13970 7908
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 16557 7939 16615 7945
rect 16557 7936 16569 7939
rect 15988 7908 16569 7936
rect 15988 7896 15994 7908
rect 16557 7905 16569 7908
rect 16603 7936 16615 7939
rect 16942 7936 16948 7948
rect 16603 7908 16948 7936
rect 16603 7905 16615 7908
rect 16557 7899 16615 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18969 7939 19027 7945
rect 18969 7936 18981 7939
rect 18012 7908 18981 7936
rect 18012 7896 18018 7908
rect 18969 7905 18981 7908
rect 19015 7936 19027 7939
rect 19058 7936 19064 7948
rect 19015 7908 19064 7936
rect 19015 7905 19027 7908
rect 18969 7899 19027 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 22020 7936 22048 7976
rect 22554 7964 22560 8016
rect 22612 8004 22618 8016
rect 23124 8004 23152 8035
rect 23474 8032 23480 8084
rect 23532 8072 23538 8084
rect 25041 8075 25099 8081
rect 23532 8044 23888 8072
rect 23532 8032 23538 8044
rect 22612 7976 23152 8004
rect 22612 7964 22618 7976
rect 23290 7964 23296 8016
rect 23348 8004 23354 8016
rect 23750 8004 23756 8016
rect 23348 7976 23756 8004
rect 23348 7964 23354 7976
rect 23750 7964 23756 7976
rect 23808 7964 23814 8016
rect 23860 8004 23888 8044
rect 25041 8041 25053 8075
rect 25087 8072 25099 8075
rect 25406 8072 25412 8084
rect 25087 8044 25412 8072
rect 25087 8041 25099 8044
rect 25041 8035 25099 8041
rect 25406 8032 25412 8044
rect 25464 8032 25470 8084
rect 27246 8004 27252 8016
rect 23860 7976 27252 8004
rect 27246 7964 27252 7976
rect 27304 7964 27310 8016
rect 22646 7936 22652 7948
rect 19392 7908 19656 7936
rect 22020 7908 22140 7936
rect 22607 7908 22652 7936
rect 19392 7896 19398 7908
rect 7432 7840 7604 7868
rect 7432 7828 7438 7840
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8478 7868 8484 7880
rect 8076 7840 8484 7868
rect 8076 7828 8082 7840
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 8662 7868 8668 7880
rect 8623 7840 8668 7868
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 9950 7868 9956 7880
rect 9911 7840 9956 7868
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 13998 7868 14004 7880
rect 13959 7840 14004 7868
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 19628 7877 19656 7908
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 20438 7868 20444 7880
rect 19659 7840 20444 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 4525 7803 4583 7809
rect 4525 7769 4537 7803
rect 4571 7800 4583 7803
rect 5350 7800 5356 7812
rect 4571 7772 5356 7800
rect 4571 7769 4583 7772
rect 4525 7763 4583 7769
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 6454 7800 6460 7812
rect 6415 7772 6460 7800
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 18598 7800 18604 7812
rect 18559 7772 18604 7800
rect 18598 7760 18604 7772
rect 18656 7760 18662 7812
rect 19426 7760 19432 7812
rect 19484 7800 19490 7812
rect 19536 7800 19564 7831
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 21174 7828 21180 7880
rect 21232 7868 21238 7880
rect 22112 7877 22140 7908
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 23474 7936 23480 7948
rect 23435 7908 23480 7936
rect 23474 7896 23480 7908
rect 23532 7936 23538 7948
rect 24121 7939 24179 7945
rect 24121 7936 24133 7939
rect 23532 7908 24133 7936
rect 23532 7896 23538 7908
rect 24121 7905 24133 7908
rect 24167 7905 24179 7939
rect 24121 7899 24179 7905
rect 22005 7871 22063 7877
rect 22005 7868 22017 7871
rect 21232 7840 22017 7868
rect 21232 7828 21238 7840
rect 22005 7837 22017 7840
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 23569 7871 23627 7877
rect 23569 7837 23581 7871
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 19484 7772 19564 7800
rect 19484 7760 19490 7772
rect 23474 7760 23480 7812
rect 23532 7800 23538 7812
rect 23584 7800 23612 7831
rect 23658 7828 23664 7880
rect 23716 7868 23722 7880
rect 25130 7868 25136 7880
rect 23716 7840 23761 7868
rect 25091 7840 25136 7868
rect 23716 7828 23722 7840
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 25317 7871 25375 7877
rect 25317 7837 25329 7871
rect 25363 7868 25375 7871
rect 25682 7868 25688 7880
rect 25363 7840 25688 7868
rect 25363 7837 25375 7840
rect 25317 7831 25375 7837
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 23532 7772 23612 7800
rect 23532 7760 23538 7772
rect 23750 7760 23756 7812
rect 23808 7800 23814 7812
rect 24673 7803 24731 7809
rect 24673 7800 24685 7803
rect 23808 7772 24685 7800
rect 23808 7760 23814 7772
rect 24673 7769 24685 7772
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 6270 7732 6276 7744
rect 6231 7704 6276 7732
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8110 7732 8116 7744
rect 8067 7704 8116 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 9033 7735 9091 7741
rect 9033 7732 9045 7735
rect 8996 7704 9045 7732
rect 8996 7692 9002 7704
rect 9033 7701 9045 7704
rect 9079 7701 9091 7735
rect 9490 7732 9496 7744
rect 9451 7704 9496 7732
rect 9033 7695 9091 7701
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12768 7704 12909 7732
rect 12768 7692 12774 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 12897 7695 12955 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 15930 7732 15936 7744
rect 15887 7704 15936 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 18782 7732 18788 7744
rect 18743 7704 18788 7732
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 21545 7735 21603 7741
rect 21545 7701 21557 7735
rect 21591 7732 21603 7735
rect 22094 7732 22100 7744
rect 21591 7704 22100 7732
rect 21591 7701 21603 7704
rect 21545 7695 21603 7701
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 24210 7692 24216 7744
rect 24268 7732 24274 7744
rect 24489 7735 24547 7741
rect 24489 7732 24501 7735
rect 24268 7704 24501 7732
rect 24268 7692 24274 7704
rect 24489 7701 24501 7704
rect 24535 7701 24547 7735
rect 24489 7695 24547 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 2498 7528 2504 7540
rect 1627 7500 2504 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 3602 7528 3608 7540
rect 3563 7500 3608 7528
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6052 7500 6837 7528
rect 6052 7488 6058 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 8662 7488 8668 7540
rect 8720 7528 8726 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 8720 7500 9597 7528
rect 8720 7488 8726 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 9585 7491 9643 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12526 7528 12532 7540
rect 12299 7500 12532 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13722 7528 13728 7540
rect 13311 7500 13728 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 15565 7531 15623 7537
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 16114 7528 16120 7540
rect 15611 7500 16120 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 16114 7488 16120 7500
rect 16172 7488 16178 7540
rect 19150 7528 19156 7540
rect 19111 7500 19156 7528
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 19797 7531 19855 7537
rect 19797 7528 19809 7531
rect 19576 7500 19809 7528
rect 19576 7488 19582 7500
rect 19797 7497 19809 7500
rect 19843 7497 19855 7531
rect 19797 7491 19855 7497
rect 20438 7488 20444 7540
rect 20496 7528 20502 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 20496 7500 20821 7528
rect 20496 7488 20502 7500
rect 20809 7497 20821 7500
rect 20855 7528 20867 7531
rect 21266 7528 21272 7540
rect 20855 7500 21272 7528
rect 20855 7497 20867 7500
rect 20809 7491 20867 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 21361 7531 21419 7537
rect 21361 7497 21373 7531
rect 21407 7528 21419 7531
rect 21450 7528 21456 7540
rect 21407 7500 21456 7528
rect 21407 7497 21419 7500
rect 21361 7491 21419 7497
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 21634 7488 21640 7540
rect 21692 7528 21698 7540
rect 21821 7531 21879 7537
rect 21821 7528 21833 7531
rect 21692 7500 21833 7528
rect 21692 7488 21698 7500
rect 21821 7497 21833 7500
rect 21867 7497 21879 7531
rect 22002 7528 22008 7540
rect 21963 7500 22008 7528
rect 21821 7491 21879 7497
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 23201 7531 23259 7537
rect 23201 7497 23213 7531
rect 23247 7528 23259 7531
rect 23658 7528 23664 7540
rect 23247 7500 23664 7528
rect 23247 7497 23259 7500
rect 23201 7491 23259 7497
rect 23658 7488 23664 7500
rect 23716 7488 23722 7540
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 24029 7531 24087 7537
rect 24029 7528 24041 7531
rect 23992 7500 24041 7528
rect 23992 7488 23998 7500
rect 24029 7497 24041 7500
rect 24075 7497 24087 7531
rect 24029 7491 24087 7497
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 5316 7432 6040 7460
rect 5316 7420 5322 7432
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2130 7352 2136 7404
rect 2188 7392 2194 7404
rect 2188 7364 2233 7392
rect 2188 7352 2194 7364
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 3936 7364 4169 7392
rect 3936 7352 3942 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5592 7364 5733 7392
rect 5592 7352 5598 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 6012 7392 6040 7432
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 6641 7463 6699 7469
rect 6641 7460 6653 7463
rect 6420 7432 6653 7460
rect 6420 7420 6426 7432
rect 6641 7429 6653 7432
rect 6687 7460 6699 7463
rect 8573 7463 8631 7469
rect 6687 7432 7420 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 7392 7404 7420 7432
rect 8573 7429 8585 7463
rect 8619 7460 8631 7463
rect 9490 7460 9496 7472
rect 8619 7432 9496 7460
rect 8619 7429 8631 7432
rect 8573 7423 8631 7429
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 6012 7364 6960 7392
rect 5721 7355 5779 7361
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7324 2743 7327
rect 2866 7324 2872 7336
rect 2731 7296 2872 7324
rect 2731 7293 2743 7296
rect 2685 7287 2743 7293
rect 2866 7284 2872 7296
rect 2924 7324 2930 7336
rect 3602 7324 3608 7336
rect 2924 7296 3608 7324
rect 2924 7284 2930 7296
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 4755 7296 5641 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 5629 7293 5641 7296
rect 5675 7324 5687 7327
rect 6822 7324 6828 7336
rect 5675 7296 6828 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6932 7324 6960 7364
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7248 7364 7297 7392
rect 7248 7352 7254 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7285 7355 7343 7361
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 9214 7392 9220 7404
rect 7432 7364 7477 7392
rect 9175 7364 9220 7392
rect 7432 7352 7438 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 10870 7392 10876 7404
rect 10827 7364 10876 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 16132 7392 16160 7488
rect 16301 7463 16359 7469
rect 16301 7429 16313 7463
rect 16347 7460 16359 7463
rect 21174 7460 21180 7472
rect 16347 7432 17080 7460
rect 21135 7432 21180 7460
rect 16347 7429 16359 7432
rect 16301 7423 16359 7429
rect 17052 7401 17080 7432
rect 21174 7420 21180 7432
rect 21232 7420 21238 7472
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16132 7364 16865 7392
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17494 7392 17500 7404
rect 17083 7364 17500 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 17770 7352 17776 7404
rect 17828 7392 17834 7404
rect 18509 7395 18567 7401
rect 18509 7392 18521 7395
rect 17828 7364 18521 7392
rect 17828 7352 17834 7364
rect 18509 7361 18521 7364
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 18601 7395 18659 7401
rect 18601 7361 18613 7395
rect 18647 7361 18659 7395
rect 20438 7392 20444 7404
rect 20351 7364 20444 7392
rect 18601 7355 18659 7361
rect 8386 7324 8392 7336
rect 6932 7296 8392 7324
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 10505 7327 10563 7333
rect 10505 7324 10517 7327
rect 9548 7296 10517 7324
rect 9548 7284 9554 7296
rect 10505 7293 10517 7296
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 13630 7333 13636 7336
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 13228 7296 13369 7324
rect 13228 7284 13234 7296
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 13624 7324 13636 7333
rect 13543 7296 13636 7324
rect 13357 7287 13415 7293
rect 13624 7287 13636 7296
rect 13688 7324 13694 7336
rect 14550 7324 14556 7336
rect 13688 7296 14556 7324
rect 3513 7259 3571 7265
rect 3513 7225 3525 7259
rect 3559 7256 3571 7259
rect 3878 7256 3884 7268
rect 3559 7228 3884 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3878 7216 3884 7228
rect 3936 7256 3942 7268
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 3936 7228 4077 7256
rect 3936 7216 3942 7228
rect 4065 7225 4077 7228
rect 4111 7225 4123 7259
rect 4065 7219 4123 7225
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 5123 7228 5549 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5537 7225 5549 7228
rect 5583 7256 5595 7259
rect 6454 7256 6460 7268
rect 5583 7228 6460 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 13372 7256 13400 7287
rect 13630 7284 13636 7287
rect 13688 7284 13694 7296
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 16758 7324 16764 7336
rect 16632 7296 16764 7324
rect 16632 7284 16638 7296
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18104 7296 18429 7324
rect 18104 7284 18110 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18616 7324 18644 7355
rect 20438 7352 20444 7364
rect 20496 7392 20502 7404
rect 21082 7392 21088 7404
rect 20496 7364 21088 7392
rect 20496 7352 20502 7364
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 22646 7392 22652 7404
rect 22607 7364 22652 7392
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 18417 7287 18475 7293
rect 18524 7296 18644 7324
rect 20257 7327 20315 7333
rect 13722 7256 13728 7268
rect 13372 7228 13728 7256
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 17405 7259 17463 7265
rect 17405 7256 17417 7259
rect 14332 7228 17417 7256
rect 14332 7216 14338 7228
rect 17405 7225 17417 7228
rect 17451 7256 17463 7259
rect 17678 7256 17684 7268
rect 17451 7228 17684 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 17678 7216 17684 7228
rect 17736 7256 17742 7268
rect 18524 7256 18552 7296
rect 20257 7293 20269 7327
rect 20303 7324 20315 7327
rect 20622 7324 20628 7336
rect 20303 7296 20628 7324
rect 20303 7293 20315 7296
rect 20257 7287 20315 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 21542 7324 21548 7336
rect 21503 7296 21548 7324
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 24044 7324 24072 7491
rect 25130 7488 25136 7540
rect 25188 7488 25194 7540
rect 25406 7488 25412 7540
rect 25464 7528 25470 7540
rect 25593 7531 25651 7537
rect 25593 7528 25605 7531
rect 25464 7500 25605 7528
rect 25464 7488 25470 7500
rect 25593 7497 25605 7500
rect 25639 7497 25651 7531
rect 25593 7491 25651 7497
rect 25682 7488 25688 7540
rect 25740 7528 25746 7540
rect 25961 7531 26019 7537
rect 25961 7528 25973 7531
rect 25740 7500 25973 7528
rect 25740 7488 25746 7500
rect 25961 7497 25973 7500
rect 26007 7497 26019 7531
rect 25961 7491 26019 7497
rect 25148 7460 25176 7488
rect 26329 7463 26387 7469
rect 26329 7460 26341 7463
rect 25148 7432 26341 7460
rect 26329 7429 26341 7432
rect 26375 7429 26387 7463
rect 26329 7423 26387 7429
rect 24946 7352 24952 7404
rect 25004 7392 25010 7404
rect 25133 7395 25191 7401
rect 25133 7392 25145 7395
rect 25004 7364 25145 7392
rect 25004 7352 25010 7364
rect 25133 7361 25145 7364
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 25041 7327 25099 7333
rect 25041 7324 25053 7327
rect 21652 7296 22508 7324
rect 24044 7296 25053 7324
rect 17736 7228 18552 7256
rect 17736 7216 17742 7228
rect 18598 7216 18604 7268
rect 18656 7256 18662 7268
rect 20165 7259 20223 7265
rect 20165 7256 20177 7259
rect 18656 7228 20177 7256
rect 18656 7216 18662 7228
rect 20165 7225 20177 7228
rect 20211 7225 20223 7259
rect 20165 7219 20223 7225
rect 20806 7216 20812 7268
rect 20864 7256 20870 7268
rect 21652 7256 21680 7296
rect 22370 7256 22376 7268
rect 20864 7228 21680 7256
rect 22331 7228 22376 7256
rect 20864 7216 20870 7228
rect 22370 7216 22376 7228
rect 22428 7216 22434 7268
rect 22480 7256 22508 7296
rect 25041 7293 25053 7296
rect 25087 7293 25099 7327
rect 25041 7287 25099 7293
rect 24489 7259 24547 7265
rect 24489 7256 24501 7259
rect 22480 7228 24501 7256
rect 24489 7225 24501 7228
rect 24535 7256 24547 7259
rect 24535 7228 24992 7256
rect 24535 7225 24547 7228
rect 24489 7219 24547 7225
rect 1578 7148 1584 7200
rect 1636 7188 1642 7200
rect 1949 7191 2007 7197
rect 1949 7188 1961 7191
rect 1636 7160 1961 7188
rect 1636 7148 1642 7160
rect 1949 7157 1961 7160
rect 1995 7157 2007 7191
rect 1949 7151 2007 7157
rect 2590 7148 2596 7200
rect 2648 7188 2654 7200
rect 2958 7188 2964 7200
rect 2648 7160 2964 7188
rect 2648 7148 2654 7160
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 3973 7191 4031 7197
rect 3973 7188 3985 7191
rect 3844 7160 3985 7188
rect 3844 7148 3850 7160
rect 3973 7157 3985 7160
rect 4019 7157 4031 7191
rect 3973 7151 4031 7157
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 4488 7160 6193 7188
rect 4488 7148 4494 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 6181 7151 6239 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8018 7188 8024 7200
rect 7800 7160 8024 7188
rect 7800 7148 7806 7160
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 8938 7188 8944 7200
rect 8899 7160 8944 7188
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 10042 7188 10048 7200
rect 9088 7160 9133 7188
rect 10003 7160 10048 7188
rect 9088 7148 9094 7160
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10597 7191 10655 7197
rect 10192 7160 10237 7188
rect 10192 7148 10198 7160
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 10778 7188 10784 7200
rect 10643 7160 10784 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11146 7188 11152 7200
rect 11107 7160 11152 7188
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14737 7191 14795 7197
rect 14737 7188 14749 7191
rect 14056 7160 14749 7188
rect 14056 7148 14062 7160
rect 14737 7157 14749 7160
rect 14783 7157 14795 7191
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 14737 7151 14795 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16393 7191 16451 7197
rect 16393 7157 16405 7191
rect 16439 7188 16451 7191
rect 16482 7188 16488 7200
rect 16439 7160 16488 7188
rect 16439 7157 16451 7160
rect 16393 7151 16451 7157
rect 16482 7148 16488 7160
rect 16540 7148 16546 7200
rect 17770 7188 17776 7200
rect 17731 7160 17776 7188
rect 17770 7148 17776 7160
rect 17828 7148 17834 7200
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 18012 7160 18061 7188
rect 18012 7148 18018 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 19426 7188 19432 7200
rect 19387 7160 19432 7188
rect 18049 7151 18107 7157
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 22462 7188 22468 7200
rect 22423 7160 22468 7188
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 24581 7191 24639 7197
rect 24581 7157 24593 7191
rect 24627 7188 24639 7191
rect 24762 7188 24768 7200
rect 24627 7160 24768 7188
rect 24627 7157 24639 7160
rect 24581 7151 24639 7157
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 24964 7197 24992 7228
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25222 7188 25228 7200
rect 24995 7160 25228 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25222 7148 25228 7160
rect 25280 7148 25286 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2608 6956 2912 6984
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 2608 6848 2636 6956
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 2777 6919 2835 6925
rect 2777 6916 2789 6919
rect 2740 6888 2789 6916
rect 2740 6876 2746 6888
rect 2777 6885 2789 6888
rect 2823 6885 2835 6919
rect 2777 6879 2835 6885
rect 2363 6820 2636 6848
rect 2884 6848 2912 6956
rect 4522 6944 4528 6996
rect 4580 6984 4586 6996
rect 4617 6987 4675 6993
rect 4617 6984 4629 6987
rect 4580 6956 4629 6984
rect 4580 6944 4586 6956
rect 4617 6953 4629 6956
rect 4663 6984 4675 6987
rect 4798 6984 4804 6996
rect 4663 6956 4804 6984
rect 4663 6953 4675 6956
rect 4617 6947 4675 6953
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5629 6987 5687 6993
rect 5629 6984 5641 6987
rect 5592 6956 5641 6984
rect 5592 6944 5598 6956
rect 5629 6953 5641 6956
rect 5675 6953 5687 6987
rect 5629 6947 5687 6953
rect 5813 6987 5871 6993
rect 5813 6953 5825 6987
rect 5859 6984 5871 6987
rect 6178 6984 6184 6996
rect 5859 6956 6184 6984
rect 5859 6953 5871 6956
rect 5813 6947 5871 6953
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7745 6987 7803 6993
rect 7745 6984 7757 6987
rect 7340 6956 7757 6984
rect 7340 6944 7346 6956
rect 7745 6953 7757 6956
rect 7791 6984 7803 6987
rect 7926 6984 7932 6996
rect 7791 6956 7932 6984
rect 7791 6953 7803 6956
rect 7745 6947 7803 6953
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9272 6956 9413 6984
rect 9272 6944 9278 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9401 6947 9459 6953
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 11977 6987 12035 6993
rect 11977 6984 11989 6987
rect 11204 6956 11989 6984
rect 11204 6944 11210 6956
rect 11977 6953 11989 6956
rect 12023 6953 12035 6987
rect 12618 6984 12624 6996
rect 12579 6956 12624 6984
rect 11977 6947 12035 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 13998 6984 14004 6996
rect 12952 6956 14004 6984
rect 12952 6944 12958 6956
rect 13998 6944 14004 6956
rect 14056 6984 14062 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 14056 6956 14105 6984
rect 14056 6944 14062 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 15988 6956 17509 6984
rect 15988 6944 15994 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 20257 6987 20315 6993
rect 20257 6953 20269 6987
rect 20303 6984 20315 6987
rect 20438 6984 20444 6996
rect 20303 6956 20444 6984
rect 20303 6953 20315 6956
rect 20257 6947 20315 6953
rect 20438 6944 20444 6956
rect 20496 6944 20502 6996
rect 20714 6984 20720 6996
rect 20675 6956 20720 6984
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 21450 6984 21456 6996
rect 20916 6956 21456 6984
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 8573 6919 8631 6925
rect 8573 6916 8585 6919
rect 4120 6888 8585 6916
rect 4120 6876 4126 6888
rect 8573 6885 8585 6888
rect 8619 6916 8631 6919
rect 9030 6916 9036 6928
rect 8619 6888 9036 6916
rect 8619 6885 8631 6888
rect 8573 6879 8631 6885
rect 9030 6876 9036 6888
rect 9088 6876 9094 6928
rect 9950 6876 9956 6928
rect 10008 6916 10014 6928
rect 12636 6916 12664 6944
rect 10008 6888 12664 6916
rect 12989 6919 13047 6925
rect 10008 6876 10014 6888
rect 12989 6885 13001 6919
rect 13035 6916 13047 6919
rect 13630 6916 13636 6928
rect 13035 6888 13636 6916
rect 13035 6885 13047 6888
rect 12989 6879 13047 6885
rect 13630 6876 13636 6888
rect 13688 6876 13694 6928
rect 16574 6916 16580 6928
rect 16224 6888 16580 6916
rect 2884 6820 3096 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 3068 6792 3096 6820
rect 4706 6808 4712 6860
rect 4764 6848 4770 6860
rect 6178 6848 6184 6860
rect 4764 6820 4809 6848
rect 6139 6820 6184 6848
rect 4764 6808 4770 6820
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 9122 6848 9128 6860
rect 9083 6820 9128 6848
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 10042 6808 10048 6860
rect 10100 6848 10106 6860
rect 10870 6857 10876 6860
rect 10505 6851 10563 6857
rect 10505 6848 10517 6851
rect 10100 6820 10517 6848
rect 10100 6808 10106 6820
rect 10505 6817 10517 6820
rect 10551 6848 10563 6851
rect 10853 6851 10876 6857
rect 10853 6848 10865 6851
rect 10551 6820 10865 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 10853 6817 10865 6820
rect 10853 6811 10876 6817
rect 10870 6808 10876 6811
rect 10928 6808 10934 6860
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13136 6820 13461 6848
rect 13136 6808 13142 6820
rect 13449 6817 13461 6820
rect 13495 6848 13507 6851
rect 14274 6848 14280 6860
rect 13495 6820 14280 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 14274 6808 14280 6820
rect 14332 6848 14338 6860
rect 14550 6848 14556 6860
rect 14332 6820 14556 6848
rect 14332 6808 14338 6820
rect 14550 6808 14556 6820
rect 14608 6808 14614 6860
rect 14826 6848 14832 6860
rect 14787 6820 14832 6848
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 15746 6848 15752 6860
rect 15611 6820 15752 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16224 6848 16252 6888
rect 16574 6876 16580 6888
rect 16632 6876 16638 6928
rect 19521 6919 19579 6925
rect 19521 6916 19533 6919
rect 19260 6888 19533 6916
rect 19260 6860 19288 6888
rect 19521 6885 19533 6888
rect 19567 6885 19579 6919
rect 19521 6879 19579 6885
rect 20162 6876 20168 6928
rect 20220 6916 20226 6928
rect 20220 6888 20668 6916
rect 20220 6876 20226 6888
rect 16390 6857 16396 6860
rect 16384 6848 16396 6857
rect 16071 6820 16252 6848
rect 16351 6820 16396 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16384 6811 16396 6820
rect 16390 6808 16396 6811
rect 16448 6808 16454 6860
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18782 6848 18788 6860
rect 17920 6820 18788 6848
rect 17920 6808 17926 6820
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 19242 6808 19248 6860
rect 19300 6808 19306 6860
rect 20640 6848 20668 6888
rect 20916 6860 20944 6956
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 22370 6944 22376 6996
rect 22428 6984 22434 6996
rect 22925 6987 22983 6993
rect 22925 6984 22937 6987
rect 22428 6956 22937 6984
rect 22428 6944 22434 6956
rect 22925 6953 22937 6956
rect 22971 6984 22983 6987
rect 23750 6984 23756 6996
rect 22971 6956 23756 6984
rect 22971 6953 22983 6956
rect 22925 6947 22983 6953
rect 23750 6944 23756 6956
rect 23808 6944 23814 6996
rect 25590 6944 25596 6996
rect 25648 6984 25654 6996
rect 25777 6987 25835 6993
rect 25777 6984 25789 6987
rect 25648 6956 25789 6984
rect 25648 6944 25654 6956
rect 25777 6953 25789 6956
rect 25823 6953 25835 6987
rect 25777 6947 25835 6953
rect 22646 6876 22652 6928
rect 22704 6916 22710 6928
rect 25682 6916 25688 6928
rect 22704 6888 23796 6916
rect 22704 6876 22710 6888
rect 20898 6848 20904 6860
rect 20640 6820 20760 6848
rect 20811 6820 20904 6848
rect 1946 6740 1952 6792
rect 2004 6780 2010 6792
rect 2774 6780 2780 6792
rect 2004 6752 2780 6780
rect 2004 6740 2010 6752
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 2869 6783 2927 6789
rect 2869 6780 2881 6783
rect 2832 6752 2881 6780
rect 2832 6740 2838 6752
rect 2869 6749 2881 6752
rect 2915 6749 2927 6783
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 2869 6743 2927 6749
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 4798 6780 4804 6792
rect 4759 6752 4804 6780
rect 4798 6740 4804 6752
rect 4856 6740 4862 6792
rect 6270 6780 6276 6792
rect 6231 6752 6276 6780
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6454 6780 6460 6792
rect 6367 6752 6460 6780
rect 6454 6740 6460 6752
rect 6512 6780 6518 6792
rect 6638 6780 6644 6792
rect 6512 6752 6644 6780
rect 6512 6740 6518 6752
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8202 6780 8208 6792
rect 8067 6752 8208 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 9824 6752 10609 6780
rect 9824 6740 9830 6752
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13228 6752 13553 6780
rect 13228 6740 13234 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 5350 6712 5356 6724
rect 5311 6684 5356 6712
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 10137 6715 10195 6721
rect 10137 6681 10149 6715
rect 10183 6712 10195 6715
rect 13081 6715 13139 6721
rect 13081 6712 13093 6715
rect 10183 6684 10640 6712
rect 10183 6681 10195 6684
rect 10137 6675 10195 6681
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2038 6644 2044 6656
rect 1995 6616 2044 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2682 6644 2688 6656
rect 2455 6616 2688 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3016 6616 3617 6644
rect 3016 6604 3022 6616
rect 3605 6613 3617 6616
rect 3651 6644 3663 6647
rect 3786 6644 3792 6656
rect 3651 6616 3792 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4249 6647 4307 6653
rect 4249 6613 4261 6647
rect 4295 6644 4307 6647
rect 5442 6644 5448 6656
rect 4295 6616 5448 6644
rect 4295 6613 4307 6616
rect 4249 6607 4307 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6822 6644 6828 6656
rect 6696 6616 6828 6644
rect 6696 6604 6702 6616
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7006 6644 7012 6656
rect 6967 6616 7012 6644
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 8938 6644 8944 6656
rect 8899 6616 8944 6644
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 10612 6644 10640 6684
rect 11532 6684 13093 6712
rect 10778 6644 10784 6656
rect 10612 6616 10784 6644
rect 10778 6604 10784 6616
rect 10836 6644 10842 6656
rect 11532 6644 11560 6684
rect 13081 6681 13093 6684
rect 13127 6681 13139 6715
rect 13556 6712 13584 6743
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 16114 6780 16120 6792
rect 13688 6752 13733 6780
rect 16075 6752 16120 6780
rect 13688 6740 13694 6752
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 19150 6780 19156 6792
rect 18555 6752 19156 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6749 19855 6783
rect 20732 6780 20760 6820
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21157 6851 21215 6857
rect 21157 6848 21169 6851
rect 21048 6820 21169 6848
rect 21048 6808 21054 6820
rect 21157 6817 21169 6820
rect 21203 6817 21215 6851
rect 21157 6811 21215 6817
rect 23293 6851 23351 6857
rect 23293 6817 23305 6851
rect 23339 6848 23351 6851
rect 23474 6848 23480 6860
rect 23339 6820 23480 6848
rect 23339 6817 23351 6820
rect 23293 6811 23351 6817
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 23658 6857 23664 6860
rect 23652 6848 23664 6857
rect 23619 6820 23664 6848
rect 23652 6811 23664 6820
rect 23658 6808 23664 6811
rect 23716 6808 23722 6860
rect 23768 6848 23796 6888
rect 24872 6888 25688 6916
rect 24210 6848 24216 6860
rect 23768 6820 24216 6848
rect 24210 6808 24216 6820
rect 24268 6848 24274 6860
rect 24268 6820 24808 6848
rect 24268 6808 24274 6820
rect 21008 6780 21036 6808
rect 20732 6752 21036 6780
rect 19797 6743 19855 6749
rect 19628 6712 19656 6743
rect 13556 6684 16160 6712
rect 13081 6675 13139 6681
rect 10836 6616 11560 6644
rect 10836 6604 10842 6616
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13906 6644 13912 6656
rect 13228 6616 13912 6644
rect 13228 6604 13234 6616
rect 13906 6604 13912 6616
rect 13964 6644 13970 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 13964 6616 14473 6644
rect 13964 6604 13970 6616
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 16132 6644 16160 6684
rect 18524 6684 19656 6712
rect 19812 6712 19840 6743
rect 23382 6740 23388 6792
rect 23440 6780 23446 6792
rect 23440 6752 23485 6780
rect 23440 6740 23446 6752
rect 20714 6712 20720 6724
rect 19812 6684 20720 6712
rect 18524 6656 18552 6684
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 24780 6721 24808 6820
rect 24765 6715 24823 6721
rect 24765 6681 24777 6715
rect 24811 6681 24823 6715
rect 24765 6675 24823 6681
rect 17770 6644 17776 6656
rect 16132 6616 17776 6644
rect 14461 6607 14519 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18046 6644 18052 6656
rect 18007 6616 18052 6644
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 18506 6604 18512 6656
rect 18564 6604 18570 6656
rect 18598 6604 18604 6656
rect 18656 6644 18662 6656
rect 19153 6647 19211 6653
rect 18656 6616 18701 6644
rect 18656 6604 18662 6616
rect 19153 6613 19165 6647
rect 19199 6644 19211 6647
rect 19334 6644 19340 6656
rect 19199 6616 19340 6644
rect 19199 6613 19211 6616
rect 19153 6607 19211 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 22278 6644 22284 6656
rect 22239 6616 22284 6644
rect 22278 6604 22284 6616
rect 22336 6604 22342 6656
rect 23658 6604 23664 6656
rect 23716 6644 23722 6656
rect 24872 6644 24900 6888
rect 25682 6876 25688 6888
rect 25740 6876 25746 6928
rect 23716 6616 24900 6644
rect 23716 6604 23722 6616
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 25004 6616 25329 6644
rect 25004 6604 25010 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 25317 6607 25375 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1946 6440 1952 6452
rect 1907 6412 1952 6440
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 3786 6440 3792 6452
rect 2096 6412 3792 6440
rect 2096 6400 2102 6412
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4522 6440 4528 6452
rect 4479 6412 4528 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5074 6440 5080 6452
rect 5035 6412 5080 6440
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 7926 6440 7932 6452
rect 7887 6412 7932 6440
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9272 6412 9720 6440
rect 9272 6400 9278 6412
rect 4246 6332 4252 6384
rect 4304 6372 4310 6384
rect 4614 6372 4620 6384
rect 4304 6344 4620 6372
rect 4304 6332 4310 6344
rect 4614 6332 4620 6344
rect 4672 6332 4678 6384
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 6641 6375 6699 6381
rect 6641 6372 6653 6375
rect 6604 6344 6653 6372
rect 6604 6332 6610 6344
rect 6641 6341 6653 6344
rect 6687 6372 6699 6375
rect 7834 6372 7840 6384
rect 6687 6344 7840 6372
rect 6687 6341 6699 6344
rect 6641 6335 6699 6341
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 2314 6304 2320 6316
rect 1544 6276 2320 6304
rect 1544 6264 1550 6276
rect 2314 6264 2320 6276
rect 2372 6304 2378 6316
rect 2409 6307 2467 6313
rect 2409 6304 2421 6307
rect 2372 6276 2421 6304
rect 2372 6264 2378 6276
rect 2409 6273 2421 6276
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 2424 6236 2452 6267
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5408 6276 5549 6304
rect 5408 6264 5414 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5684 6276 5729 6304
rect 5684 6264 5690 6276
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7064 6276 7573 6304
rect 7064 6264 7070 6276
rect 7561 6273 7573 6276
rect 7607 6304 7619 6307
rect 8478 6304 8484 6316
rect 7607 6276 8484 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9692 6313 9720 6412
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 12986 6440 12992 6452
rect 12216 6412 12992 6440
rect 12216 6400 12222 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 14274 6440 14280 6452
rect 13955 6412 14280 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 18601 6443 18659 6449
rect 18601 6409 18613 6443
rect 18647 6440 18659 6443
rect 19242 6440 19248 6452
rect 18647 6412 19248 6440
rect 18647 6409 18659 6412
rect 18601 6403 18659 6409
rect 11330 6332 11336 6384
rect 11388 6372 11394 6384
rect 11885 6375 11943 6381
rect 11885 6372 11897 6375
rect 11388 6344 11897 6372
rect 11388 6332 11394 6344
rect 11885 6341 11897 6344
rect 11931 6372 11943 6375
rect 11931 6344 13124 6372
rect 11931 6341 11943 6344
rect 11885 6335 11943 6341
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 9723 6276 9996 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 4246 6236 4252 6248
rect 2424 6208 4252 6236
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6236 8631 6239
rect 8619 6208 9444 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 1302 6128 1308 6180
rect 1360 6168 1366 6180
rect 2225 6171 2283 6177
rect 2225 6168 2237 6171
rect 1360 6140 2237 6168
rect 1360 6128 1366 6140
rect 2225 6137 2237 6140
rect 2271 6137 2283 6171
rect 2225 6131 2283 6137
rect 1394 6100 1400 6112
rect 1355 6072 1400 6100
rect 1394 6060 1400 6072
rect 1452 6060 1458 6112
rect 2240 6100 2268 6131
rect 2406 6128 2412 6180
rect 2464 6168 2470 6180
rect 2676 6171 2734 6177
rect 2676 6168 2688 6171
rect 2464 6140 2688 6168
rect 2464 6128 2470 6140
rect 2676 6137 2688 6140
rect 2722 6137 2734 6171
rect 8846 6168 8852 6180
rect 8807 6140 8852 6168
rect 2676 6131 2734 6137
rect 8846 6128 8852 6140
rect 8904 6128 8910 6180
rect 9416 6112 9444 6208
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9824 6208 9873 6236
rect 9824 6196 9830 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9968 6236 9996 6276
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 13096 6313 13124 6344
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12676 6276 12909 6304
rect 12676 6264 12682 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6304 13139 6307
rect 13630 6304 13636 6316
rect 13127 6276 13636 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18616 6304 18644 6403
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 21545 6443 21603 6449
rect 21545 6409 21557 6443
rect 21591 6440 21603 6443
rect 22002 6440 22008 6452
rect 21591 6412 22008 6440
rect 21591 6409 21603 6412
rect 21545 6403 21603 6409
rect 22002 6400 22008 6412
rect 22060 6400 22066 6452
rect 22094 6400 22100 6452
rect 22152 6440 22158 6452
rect 22557 6443 22615 6449
rect 22557 6440 22569 6443
rect 22152 6412 22569 6440
rect 22152 6400 22158 6412
rect 22557 6409 22569 6412
rect 22603 6409 22615 6443
rect 22557 6403 22615 6409
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 23661 6443 23719 6449
rect 23661 6440 23673 6443
rect 23532 6412 23673 6440
rect 23532 6400 23538 6412
rect 23661 6409 23673 6412
rect 23707 6409 23719 6443
rect 23661 6403 23719 6409
rect 25590 6400 25596 6452
rect 25648 6440 25654 6452
rect 25958 6440 25964 6452
rect 25648 6412 25964 6440
rect 25648 6400 25654 6412
rect 25958 6400 25964 6412
rect 26016 6440 26022 6452
rect 26329 6443 26387 6449
rect 26329 6440 26341 6443
rect 26016 6412 26341 6440
rect 26016 6400 26022 6412
rect 26329 6409 26341 6412
rect 26375 6409 26387 6443
rect 26329 6403 26387 6409
rect 18690 6332 18696 6384
rect 18748 6372 18754 6384
rect 19061 6375 19119 6381
rect 19061 6372 19073 6375
rect 18748 6344 19073 6372
rect 18748 6332 18754 6344
rect 19061 6341 19073 6344
rect 19107 6341 19119 6375
rect 19061 6335 19119 6341
rect 20806 6332 20812 6384
rect 20864 6372 20870 6384
rect 22646 6372 22652 6384
rect 20864 6344 22652 6372
rect 20864 6332 20870 6344
rect 22646 6332 22652 6344
rect 22704 6332 22710 6384
rect 24118 6332 24124 6384
rect 24176 6372 24182 6384
rect 24302 6372 24308 6384
rect 24176 6344 24308 6372
rect 24176 6332 24182 6344
rect 24302 6332 24308 6344
rect 24360 6332 24366 6384
rect 24486 6332 24492 6384
rect 24544 6372 24550 6384
rect 25038 6372 25044 6384
rect 24544 6344 25044 6372
rect 24544 6332 24550 6344
rect 25038 6332 25044 6344
rect 25096 6332 25102 6384
rect 18095 6276 18644 6304
rect 19705 6307 19763 6313
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 19705 6273 19717 6307
rect 19751 6304 19763 6307
rect 20070 6304 20076 6316
rect 19751 6276 20076 6304
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21876 6276 22017 6304
rect 21876 6264 21882 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6304 22247 6307
rect 23477 6307 23535 6313
rect 23477 6304 23489 6307
rect 22235 6276 23489 6304
rect 22235 6273 22247 6276
rect 22189 6267 22247 6273
rect 23477 6273 23489 6276
rect 23523 6304 23535 6307
rect 23658 6304 23664 6316
rect 23523 6276 23664 6304
rect 23523 6273 23535 6276
rect 23477 6267 23535 6273
rect 10128 6239 10186 6245
rect 10128 6236 10140 6239
rect 9968 6208 10140 6236
rect 9861 6199 9919 6205
rect 10128 6205 10140 6208
rect 10174 6236 10186 6239
rect 11330 6236 11336 6248
rect 10174 6208 11336 6236
rect 10174 6205 10186 6208
rect 10128 6199 10186 6205
rect 11330 6196 11336 6208
rect 11388 6196 11394 6248
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11848 6208 12173 6236
rect 11848 6196 11854 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12176 6168 12204 6199
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 13872 6208 14105 6236
rect 13872 6196 13878 6208
rect 14093 6205 14105 6208
rect 14139 6236 14151 6239
rect 15194 6236 15200 6248
rect 14139 6208 15200 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 15194 6196 15200 6208
rect 15252 6236 15258 6248
rect 16114 6236 16120 6248
rect 15252 6208 16120 6236
rect 15252 6196 15258 6208
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16574 6236 16580 6248
rect 16535 6208 16580 6236
rect 16574 6196 16580 6208
rect 16632 6236 16638 6248
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 16632 6208 17325 6236
rect 16632 6196 16638 6208
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18877 6239 18935 6245
rect 18877 6236 18889 6239
rect 18564 6208 18889 6236
rect 18564 6196 18570 6208
rect 18877 6205 18889 6208
rect 18923 6205 18935 6239
rect 18877 6199 18935 6205
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 21913 6239 21971 6245
rect 21913 6236 21925 6239
rect 21784 6208 21925 6236
rect 21784 6196 21790 6208
rect 21913 6205 21925 6208
rect 21959 6236 21971 6239
rect 22094 6236 22100 6248
rect 21959 6208 22100 6236
rect 21959 6205 21971 6208
rect 21913 6199 21971 6205
rect 22094 6196 22100 6208
rect 22152 6196 22158 6248
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12176 6140 12817 6168
rect 12805 6137 12817 6140
rect 12851 6168 12863 6171
rect 12894 6168 12900 6180
rect 12851 6140 12900 6168
rect 12851 6137 12863 6140
rect 12805 6131 12863 6137
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 14338 6171 14396 6177
rect 14338 6168 14350 6171
rect 14056 6140 14350 6168
rect 14056 6128 14062 6140
rect 14338 6137 14350 6140
rect 14384 6137 14396 6171
rect 16850 6168 16856 6180
rect 16811 6140 16856 6168
rect 14338 6131 14396 6137
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 17865 6171 17923 6177
rect 17865 6137 17877 6171
rect 17911 6168 17923 6171
rect 19518 6168 19524 6180
rect 17911 6140 19524 6168
rect 17911 6137 17923 6140
rect 17865 6131 17923 6137
rect 19518 6128 19524 6140
rect 19576 6128 19582 6180
rect 21453 6171 21511 6177
rect 21453 6137 21465 6171
rect 21499 6168 21511 6171
rect 22204 6168 22232 6267
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 24210 6304 24216 6316
rect 24171 6276 24216 6304
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 25406 6304 25412 6316
rect 25367 6276 25412 6304
rect 25406 6264 25412 6276
rect 25464 6264 25470 6316
rect 23109 6239 23167 6245
rect 23109 6205 23121 6239
rect 23155 6236 23167 6239
rect 24118 6236 24124 6248
rect 23155 6208 24124 6236
rect 23155 6205 23167 6208
rect 23109 6199 23167 6205
rect 24118 6196 24124 6208
rect 24176 6196 24182 6248
rect 24854 6196 24860 6248
rect 24912 6236 24918 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 24912 6208 25237 6236
rect 24912 6196 24918 6208
rect 25225 6205 25237 6208
rect 25271 6236 25283 6239
rect 25961 6239 26019 6245
rect 25961 6236 25973 6239
rect 25271 6208 25973 6236
rect 25271 6205 25283 6208
rect 25225 6199 25283 6205
rect 25961 6205 25973 6208
rect 26007 6205 26019 6239
rect 25961 6199 26019 6205
rect 21499 6140 22232 6168
rect 21499 6137 21511 6140
rect 21453 6131 21511 6137
rect 23934 6128 23940 6180
rect 23992 6168 23998 6180
rect 24029 6171 24087 6177
rect 24029 6168 24041 6171
rect 23992 6140 24041 6168
rect 23992 6128 23998 6140
rect 24029 6137 24041 6140
rect 24075 6168 24087 6171
rect 24673 6171 24731 6177
rect 24673 6168 24685 6171
rect 24075 6140 24685 6168
rect 24075 6137 24087 6140
rect 24029 6131 24087 6137
rect 24673 6137 24685 6140
rect 24719 6137 24731 6171
rect 24673 6131 24731 6137
rect 2590 6100 2596 6112
rect 2240 6072 2596 6100
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 3660 6072 5457 6100
rect 3660 6060 3666 6072
rect 5445 6069 5457 6072
rect 5491 6100 5503 6103
rect 5994 6100 6000 6112
rect 5491 6072 6000 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5994 6060 6000 6072
rect 6052 6100 6058 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 6052 6072 6101 6100
rect 6052 6060 6058 6072
rect 6089 6069 6101 6072
rect 6135 6069 6147 6103
rect 6914 6100 6920 6112
rect 6875 6072 6920 6100
rect 6089 6063 6147 6069
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 7282 6100 7288 6112
rect 7243 6072 7288 6100
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 7432 6072 7477 6100
rect 7432 6060 7438 6072
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 8260 6072 8401 6100
rect 8260 6060 8266 6072
rect 8389 6069 8401 6072
rect 8435 6100 8447 6103
rect 8570 6100 8576 6112
rect 8435 6072 8576 6100
rect 8435 6069 8447 6072
rect 8389 6063 8447 6069
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 9398 6100 9404 6112
rect 9359 6072 9404 6100
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 11241 6103 11299 6109
rect 11241 6100 11253 6103
rect 10928 6072 11253 6100
rect 10928 6060 10934 6072
rect 11241 6069 11253 6072
rect 11287 6069 11299 6103
rect 11241 6063 11299 6069
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12492 6072 12537 6100
rect 12492 6060 12498 6072
rect 13078 6060 13084 6112
rect 13136 6100 13142 6112
rect 13446 6100 13452 6112
rect 13136 6072 13452 6100
rect 13136 6060 13142 6072
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 15470 6100 15476 6112
rect 15431 6072 15476 6100
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 16114 6100 16120 6112
rect 16075 6072 16120 6100
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19429 6103 19487 6109
rect 19429 6100 19441 6103
rect 19392 6072 19441 6100
rect 19392 6060 19398 6072
rect 19429 6069 19441 6072
rect 19475 6069 19487 6103
rect 20070 6100 20076 6112
rect 20031 6072 20076 6100
rect 19429 6063 19487 6069
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 20533 6103 20591 6109
rect 20533 6069 20545 6103
rect 20579 6100 20591 6103
rect 20714 6100 20720 6112
rect 20579 6072 20720 6100
rect 20579 6069 20591 6072
rect 20533 6063 20591 6069
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 22370 6100 22376 6112
rect 22060 6072 22376 6100
rect 22060 6060 22066 6072
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 25038 6100 25044 6112
rect 24999 6072 25044 6100
rect 25038 6060 25044 6072
rect 25096 6060 25102 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 2130 5896 2136 5908
rect 1820 5868 2136 5896
rect 1820 5856 1826 5868
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4798 5896 4804 5908
rect 3927 5868 4804 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4798 5856 4804 5868
rect 4856 5896 4862 5908
rect 5534 5896 5540 5908
rect 4856 5868 5540 5896
rect 4856 5856 4862 5868
rect 5534 5856 5540 5868
rect 5592 5896 5598 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 5592 5868 5733 5896
rect 5592 5856 5598 5868
rect 5721 5865 5733 5868
rect 5767 5865 5779 5899
rect 5721 5859 5779 5865
rect 6178 5856 6184 5908
rect 6236 5896 6242 5908
rect 6641 5899 6699 5905
rect 6641 5896 6653 5899
rect 6236 5868 6653 5896
rect 6236 5856 6242 5868
rect 6641 5865 6653 5868
rect 6687 5896 6699 5899
rect 6822 5896 6828 5908
rect 6687 5868 6828 5896
rect 6687 5865 6699 5868
rect 6641 5859 6699 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 7340 5868 9045 5896
rect 7340 5856 7346 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 9398 5856 9404 5908
rect 9456 5896 9462 5908
rect 10505 5899 10563 5905
rect 10505 5896 10517 5899
rect 9456 5868 10517 5896
rect 9456 5856 9462 5868
rect 10505 5865 10517 5868
rect 10551 5865 10563 5899
rect 13170 5896 13176 5908
rect 13131 5868 13176 5896
rect 10505 5859 10563 5865
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 13630 5856 13636 5908
rect 13688 5856 13694 5908
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 16390 5896 16396 5908
rect 16172 5868 16396 5896
rect 16172 5856 16178 5868
rect 16390 5856 16396 5868
rect 16448 5896 16454 5908
rect 16761 5899 16819 5905
rect 16761 5896 16773 5899
rect 16448 5868 16773 5896
rect 16448 5856 16454 5868
rect 16761 5865 16773 5868
rect 16807 5865 16819 5899
rect 17862 5896 17868 5908
rect 17823 5868 17868 5896
rect 16761 5859 16819 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18233 5899 18291 5905
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 19334 5896 19340 5908
rect 18279 5868 19340 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 19576 5868 20913 5896
rect 19576 5856 19582 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 21818 5856 21824 5908
rect 21876 5896 21882 5908
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 21876 5868 21925 5896
rect 21876 5856 21882 5868
rect 21913 5865 21925 5868
rect 21959 5865 21971 5899
rect 22370 5896 22376 5908
rect 22331 5868 22376 5896
rect 21913 5859 21971 5865
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 23934 5896 23940 5908
rect 23895 5868 23940 5896
rect 23934 5856 23940 5868
rect 23992 5856 23998 5908
rect 24305 5899 24363 5905
rect 24305 5865 24317 5899
rect 24351 5896 24363 5899
rect 24670 5896 24676 5908
rect 24351 5868 24676 5896
rect 24351 5865 24363 5868
rect 24305 5859 24363 5865
rect 24670 5856 24676 5868
rect 24728 5896 24734 5908
rect 24949 5899 25007 5905
rect 24949 5896 24961 5899
rect 24728 5868 24961 5896
rect 24728 5856 24734 5868
rect 24949 5865 24961 5868
rect 24995 5865 25007 5899
rect 24949 5859 25007 5865
rect 25038 5856 25044 5908
rect 25096 5896 25102 5908
rect 25317 5899 25375 5905
rect 25317 5896 25329 5899
rect 25096 5868 25329 5896
rect 25096 5856 25102 5868
rect 25317 5865 25329 5868
rect 25363 5896 25375 5899
rect 25685 5899 25743 5905
rect 25685 5896 25697 5899
rect 25363 5868 25697 5896
rect 25363 5865 25375 5868
rect 25317 5859 25375 5865
rect 25685 5865 25697 5868
rect 25731 5865 25743 5899
rect 25685 5859 25743 5865
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 4338 5828 4344 5840
rect 3844 5800 4344 5828
rect 3844 5788 3850 5800
rect 4338 5788 4344 5800
rect 4396 5828 4402 5840
rect 4586 5831 4644 5837
rect 4586 5828 4598 5831
rect 4396 5800 4598 5828
rect 4396 5788 4402 5800
rect 4586 5797 4598 5800
rect 4632 5797 4644 5831
rect 6270 5828 6276 5840
rect 6231 5800 6276 5828
rect 4586 5791 4644 5797
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 8938 5828 8944 5840
rect 7024 5800 8944 5828
rect 1486 5760 1492 5772
rect 1447 5732 1492 5760
rect 1486 5720 1492 5732
rect 1544 5720 1550 5772
rect 1762 5769 1768 5772
rect 1756 5760 1768 5769
rect 1723 5732 1768 5760
rect 1756 5723 1768 5732
rect 1762 5720 1768 5723
rect 1820 5720 1826 5772
rect 7024 5769 7052 5800
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 10413 5831 10471 5837
rect 10413 5797 10425 5831
rect 10459 5828 10471 5831
rect 10778 5828 10784 5840
rect 10459 5800 10784 5828
rect 10459 5797 10471 5800
rect 10413 5791 10471 5797
rect 10778 5788 10784 5800
rect 10836 5788 10842 5840
rect 13081 5831 13139 5837
rect 13081 5797 13093 5831
rect 13127 5828 13139 5831
rect 13648 5828 13676 5856
rect 13127 5800 13676 5828
rect 13127 5797 13139 5800
rect 13081 5791 13139 5797
rect 15746 5788 15752 5840
rect 15804 5828 15810 5840
rect 17218 5828 17224 5840
rect 15804 5800 17224 5828
rect 15804 5788 15810 5800
rect 17218 5788 17224 5800
rect 17276 5828 17282 5840
rect 17313 5831 17371 5837
rect 17313 5828 17325 5831
rect 17276 5800 17325 5828
rect 17276 5788 17282 5800
rect 17313 5797 17325 5800
rect 17359 5797 17371 5831
rect 17313 5791 17371 5797
rect 19058 5788 19064 5840
rect 19116 5828 19122 5840
rect 20257 5831 20315 5837
rect 20257 5828 20269 5831
rect 19116 5800 20269 5828
rect 19116 5788 19122 5800
rect 20257 5797 20269 5800
rect 20303 5797 20315 5831
rect 20257 5791 20315 5797
rect 20714 5788 20720 5840
rect 20772 5828 20778 5840
rect 22738 5828 22744 5840
rect 20772 5800 21496 5828
rect 22699 5800 22744 5828
rect 20772 5788 20778 5800
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5729 7067 5763
rect 7009 5723 7067 5729
rect 7368 5763 7426 5769
rect 7368 5729 7380 5763
rect 7414 5760 7426 5763
rect 8202 5760 8208 5772
rect 7414 5732 8208 5760
rect 7414 5729 7426 5732
rect 7368 5723 7426 5729
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 10134 5760 10140 5772
rect 9732 5732 10140 5760
rect 9732 5720 9738 5732
rect 10134 5720 10140 5732
rect 10192 5760 10198 5772
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10192 5732 10885 5760
rect 10192 5720 10198 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10873 5723 10931 5729
rect 10962 5720 10968 5772
rect 11020 5760 11026 5772
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 11020 5732 11529 5760
rect 11020 5720 11026 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11882 5760 11888 5772
rect 11843 5732 11888 5760
rect 11517 5723 11575 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12066 5760 12072 5772
rect 12027 5732 12072 5760
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 13446 5720 13452 5772
rect 13504 5760 13510 5772
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 13504 5732 13553 5760
rect 13504 5720 13510 5732
rect 13541 5729 13553 5732
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 13630 5720 13636 5772
rect 13688 5760 13694 5772
rect 13688 5732 13733 5760
rect 13688 5720 13694 5732
rect 14274 5720 14280 5772
rect 14332 5760 14338 5772
rect 15470 5760 15476 5772
rect 14332 5732 15476 5760
rect 14332 5720 14338 5732
rect 15470 5720 15476 5732
rect 15528 5760 15534 5772
rect 15637 5763 15695 5769
rect 15637 5760 15649 5763
rect 15528 5732 15649 5760
rect 15528 5720 15534 5732
rect 15637 5729 15649 5732
rect 15683 5729 15695 5763
rect 15637 5723 15695 5729
rect 18230 5720 18236 5772
rect 18288 5760 18294 5772
rect 18581 5763 18639 5769
rect 18581 5760 18593 5763
rect 18288 5732 18593 5760
rect 18288 5720 18294 5732
rect 18581 5729 18593 5732
rect 18627 5729 18639 5763
rect 18581 5723 18639 5729
rect 20806 5720 20812 5772
rect 20864 5760 20870 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20864 5732 21281 5760
rect 20864 5720 20870 5732
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4304 5664 4353 5692
rect 4304 5652 4310 5664
rect 4341 5661 4353 5664
rect 4387 5661 4399 5695
rect 7098 5692 7104 5704
rect 7059 5664 7104 5692
rect 4341 5655 4399 5661
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 2590 5556 2596 5568
rect 2464 5528 2596 5556
rect 2464 5516 2470 5528
rect 2590 5516 2596 5528
rect 2648 5556 2654 5568
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 2648 5528 2881 5556
rect 2648 5516 2654 5528
rect 2869 5525 2881 5528
rect 2915 5556 2927 5559
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 2915 5528 3433 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3421 5525 3433 5528
rect 3467 5556 3479 5559
rect 3602 5556 3608 5568
rect 3467 5528 3608 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 4356 5556 4384 5655
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 10410 5652 10416 5704
rect 10468 5692 10474 5704
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 10468 5664 11069 5692
rect 10468 5652 10474 5664
rect 11057 5661 11069 5664
rect 11103 5692 11115 5695
rect 11146 5692 11152 5704
rect 11103 5664 11152 5692
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 13722 5692 13728 5704
rect 13683 5664 13728 5692
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15252 5664 15393 5692
rect 15252 5652 15258 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 15381 5655 15439 5661
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5692 20775 5695
rect 21358 5692 21364 5704
rect 20763 5664 21364 5692
rect 20763 5661 20775 5664
rect 20717 5655 20775 5661
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 21468 5701 21496 5800
rect 22738 5788 22744 5800
rect 22796 5788 22802 5840
rect 23753 5831 23811 5837
rect 23753 5797 23765 5831
rect 23799 5828 23811 5831
rect 24210 5828 24216 5840
rect 23799 5800 24216 5828
rect 23799 5797 23811 5800
rect 23753 5791 23811 5797
rect 24210 5788 24216 5800
rect 24268 5788 24274 5840
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 22462 5720 22468 5732
rect 22520 5760 22526 5772
rect 23201 5763 23259 5769
rect 23201 5760 23213 5763
rect 22520 5732 23213 5760
rect 22520 5720 22526 5732
rect 23201 5729 23213 5732
rect 23247 5729 23259 5763
rect 23201 5723 23259 5729
rect 24026 5720 24032 5772
rect 24084 5760 24090 5772
rect 24397 5763 24455 5769
rect 24397 5760 24409 5763
rect 24084 5732 24409 5760
rect 24084 5720 24090 5732
rect 24397 5729 24409 5732
rect 24443 5760 24455 5763
rect 24670 5760 24676 5772
rect 24443 5732 24676 5760
rect 24443 5729 24455 5732
rect 24397 5723 24455 5729
rect 24670 5720 24676 5732
rect 24728 5720 24734 5772
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 23658 5652 23664 5704
rect 23716 5692 23722 5704
rect 24489 5695 24547 5701
rect 24489 5692 24501 5695
rect 23716 5664 24501 5692
rect 23716 5652 23722 5664
rect 24489 5661 24501 5664
rect 24535 5692 24547 5695
rect 24854 5692 24860 5704
rect 24535 5664 24860 5692
rect 24535 5661 24547 5664
rect 24489 5655 24547 5661
rect 24854 5652 24860 5664
rect 24912 5652 24918 5704
rect 6825 5627 6883 5633
rect 6825 5593 6837 5627
rect 6871 5624 6883 5627
rect 7006 5624 7012 5636
rect 6871 5596 7012 5624
rect 6871 5593 6883 5596
rect 6825 5587 6883 5593
rect 5258 5556 5264 5568
rect 4356 5528 5264 5556
rect 5258 5516 5264 5528
rect 5316 5556 5322 5568
rect 6840 5556 6868 5587
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 8478 5624 8484 5636
rect 8439 5596 8484 5624
rect 8478 5584 8484 5596
rect 8536 5584 8542 5636
rect 12710 5584 12716 5636
rect 12768 5624 12774 5636
rect 13354 5624 13360 5636
rect 12768 5596 13360 5624
rect 12768 5584 12774 5596
rect 13354 5584 13360 5596
rect 13412 5584 13418 5636
rect 5316 5528 6868 5556
rect 5316 5516 5322 5528
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 8628 5528 9413 5556
rect 8628 5516 8634 5528
rect 9401 5525 9413 5528
rect 9447 5525 9459 5559
rect 10042 5556 10048 5568
rect 10003 5528 10048 5556
rect 9401 5519 9459 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 12250 5556 12256 5568
rect 12211 5528 12256 5556
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 12618 5556 12624 5568
rect 12579 5528 12624 5556
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 14274 5556 14280 5568
rect 14235 5528 14280 5556
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 14550 5556 14556 5568
rect 14511 5528 14556 5556
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 15013 5559 15071 5565
rect 15013 5525 15025 5559
rect 15059 5556 15071 5559
rect 15378 5556 15384 5568
rect 15059 5528 15384 5556
rect 15059 5525 15071 5528
rect 15013 5519 15071 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19705 5559 19763 5565
rect 19705 5556 19717 5559
rect 19392 5528 19717 5556
rect 19392 5516 19398 5528
rect 19705 5525 19717 5528
rect 19751 5556 19763 5559
rect 20714 5556 20720 5568
rect 19751 5528 20720 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 1946 5352 1952 5364
rect 1535 5324 1952 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 1946 5312 1952 5324
rect 2004 5352 2010 5364
rect 2498 5352 2504 5364
rect 2004 5324 2504 5352
rect 2004 5312 2010 5324
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3142 5352 3148 5364
rect 3099 5324 3148 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 4338 5352 4344 5364
rect 4299 5324 4344 5352
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6454 5352 6460 5364
rect 6227 5324 6460 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7340 5324 7849 5352
rect 7340 5312 7346 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 8941 5355 8999 5361
rect 8941 5321 8953 5355
rect 8987 5352 8999 5355
rect 9674 5352 9680 5364
rect 8987 5324 9680 5352
rect 8987 5321 8999 5324
rect 8941 5315 8999 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 10410 5352 10416 5364
rect 10371 5324 10416 5352
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 10505 5355 10563 5361
rect 10505 5321 10517 5355
rect 10551 5352 10563 5355
rect 10962 5352 10968 5364
rect 10551 5324 10968 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 12066 5352 12072 5364
rect 11931 5324 12072 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 13780 5324 14933 5352
rect 13780 5312 13786 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 17218 5352 17224 5364
rect 17179 5324 17224 5352
rect 14921 5315 14979 5321
rect 17218 5312 17224 5324
rect 17276 5352 17282 5364
rect 17589 5355 17647 5361
rect 17589 5352 17601 5355
rect 17276 5324 17601 5352
rect 17276 5312 17282 5324
rect 17589 5321 17601 5324
rect 17635 5321 17647 5355
rect 21358 5352 21364 5364
rect 21319 5324 21364 5352
rect 17589 5315 17647 5321
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 22646 5312 22652 5364
rect 22704 5352 22710 5364
rect 23477 5355 23535 5361
rect 23477 5352 23489 5355
rect 22704 5324 23489 5352
rect 22704 5312 22710 5324
rect 2958 5284 2964 5296
rect 2919 5256 2964 5284
rect 2958 5244 2964 5256
rect 3016 5244 3022 5296
rect 6641 5287 6699 5293
rect 6641 5253 6653 5287
rect 6687 5284 6699 5287
rect 10045 5287 10103 5293
rect 6687 5256 7420 5284
rect 6687 5253 6699 5256
rect 6641 5247 6699 5253
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1820 5188 2053 5216
rect 1820 5176 1826 5188
rect 2041 5185 2053 5188
rect 2087 5216 2099 5219
rect 2406 5216 2412 5228
rect 2087 5188 2412 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4764 5188 4997 5216
rect 4764 5176 4770 5188
rect 4985 5185 4997 5188
rect 5031 5216 5043 5219
rect 5718 5216 5724 5228
rect 5031 5188 5724 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 6822 5216 6828 5228
rect 6783 5188 6828 5216
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7392 5225 7420 5256
rect 10045 5253 10057 5287
rect 10091 5284 10103 5287
rect 10870 5284 10876 5296
rect 10091 5256 10876 5284
rect 10091 5253 10103 5256
rect 10045 5247 10103 5253
rect 10870 5244 10876 5256
rect 10928 5284 10934 5296
rect 13909 5287 13967 5293
rect 10928 5256 11100 5284
rect 10928 5244 10934 5256
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 8202 5216 8208 5228
rect 7423 5188 8208 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 8202 5176 8208 5188
rect 8260 5216 8266 5228
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8260 5188 8401 5216
rect 8260 5176 8266 5188
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 11072 5225 11100 5256
rect 13909 5253 13921 5287
rect 13955 5284 13967 5287
rect 16485 5287 16543 5293
rect 16485 5284 16497 5287
rect 13955 5256 16497 5284
rect 13955 5253 13967 5256
rect 13909 5247 13967 5253
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10744 5188 10977 5216
rect 10744 5176 10750 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11057 5219 11115 5225
rect 11057 5185 11069 5219
rect 11103 5185 11115 5219
rect 11057 5179 11115 5185
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 15948 5225 15976 5256
rect 16485 5253 16497 5256
rect 16531 5253 16543 5287
rect 16485 5247 16543 5253
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14332 5188 14473 5216
rect 14332 5176 14338 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5216 16083 5219
rect 16114 5216 16120 5228
rect 16071 5188 16120 5216
rect 16071 5185 16083 5188
rect 16025 5179 16083 5185
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 2130 5148 2136 5160
rect 1903 5120 2136 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 2130 5108 2136 5120
rect 2188 5148 2194 5160
rect 3510 5148 3516 5160
rect 2188 5120 2728 5148
rect 3471 5120 3516 5148
rect 2188 5108 2194 5120
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 2038 5012 2044 5024
rect 1995 4984 2044 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 2038 4972 2044 4984
rect 2096 5012 2102 5024
rect 2222 5012 2228 5024
rect 2096 4984 2228 5012
rect 2096 4972 2102 4984
rect 2222 4972 2228 4984
rect 2280 5012 2286 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2280 4984 2513 5012
rect 2280 4972 2286 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2700 5012 2728 5120
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5500 5120 5549 5148
rect 5500 5108 5506 5120
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 9309 5151 9367 5157
rect 9309 5117 9321 5151
rect 9355 5148 9367 5151
rect 9398 5148 9404 5160
rect 9355 5120 9404 5148
rect 9355 5117 9367 5120
rect 9309 5111 9367 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10778 5148 10784 5160
rect 10100 5120 10784 5148
rect 10100 5108 10106 5120
rect 10778 5108 10784 5120
rect 10836 5148 10842 5160
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10836 5120 10885 5148
rect 10836 5108 10842 5120
rect 10873 5117 10885 5120
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12621 5151 12679 5157
rect 12621 5148 12633 5151
rect 12299 5120 12633 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12621 5117 12633 5120
rect 12667 5117 12679 5151
rect 14366 5148 14372 5160
rect 14327 5120 14372 5148
rect 12621 5111 12679 5117
rect 2774 5040 2780 5092
rect 2832 5080 2838 5092
rect 2832 5052 3464 5080
rect 2832 5040 2838 5052
rect 2958 5012 2964 5024
rect 2700 4984 2964 5012
rect 2501 4975 2559 4981
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 3436 5021 3464 5052
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 8297 5083 8355 5089
rect 8297 5080 8309 5083
rect 8076 5052 8309 5080
rect 8076 5040 8082 5052
rect 8297 5049 8309 5052
rect 8343 5049 8355 5083
rect 8297 5043 8355 5049
rect 12636 5024 12664 5111
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 15381 5151 15439 5157
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 16040 5148 16068 5179
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 18288 5188 18429 5216
rect 18288 5176 18294 5188
rect 18417 5185 18429 5188
rect 18463 5216 18475 5219
rect 21913 5219 21971 5225
rect 18463 5188 19012 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 18874 5148 18880 5160
rect 15427 5120 16068 5148
rect 18835 5120 18880 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 18874 5108 18880 5120
rect 18932 5108 18938 5160
rect 18984 5148 19012 5188
rect 21913 5185 21925 5219
rect 21959 5185 21971 5219
rect 21913 5179 21971 5185
rect 21928 5148 21956 5179
rect 18984 5120 21956 5148
rect 23400 5148 23428 5324
rect 23477 5321 23489 5324
rect 23523 5321 23535 5355
rect 23477 5315 23535 5321
rect 24670 5312 24676 5364
rect 24728 5352 24734 5364
rect 25593 5355 25651 5361
rect 25593 5352 25605 5355
rect 24728 5324 25605 5352
rect 24728 5312 24734 5324
rect 25593 5321 25605 5324
rect 25639 5321 25651 5355
rect 25958 5352 25964 5364
rect 25919 5324 25964 5352
rect 25593 5315 25651 5321
rect 25958 5312 25964 5324
rect 26016 5352 26022 5364
rect 26329 5355 26387 5361
rect 26329 5352 26341 5355
rect 26016 5324 26341 5352
rect 26016 5312 26022 5324
rect 26329 5321 26341 5324
rect 26375 5321 26387 5355
rect 26329 5315 26387 5321
rect 24854 5244 24860 5296
rect 24912 5284 24918 5296
rect 25041 5287 25099 5293
rect 25041 5284 25053 5287
rect 24912 5256 25053 5284
rect 24912 5244 24918 5256
rect 25041 5253 25053 5256
rect 25087 5253 25099 5287
rect 25041 5247 25099 5253
rect 23474 5176 23480 5228
rect 23532 5216 23538 5228
rect 23658 5216 23664 5228
rect 23532 5188 23664 5216
rect 23532 5176 23538 5188
rect 23658 5176 23664 5188
rect 23716 5176 23722 5228
rect 23917 5151 23975 5157
rect 23917 5148 23929 5151
rect 23400 5120 23929 5148
rect 12894 5080 12900 5092
rect 12855 5052 12900 5080
rect 12894 5040 12900 5052
rect 12952 5040 12958 5092
rect 13814 5080 13820 5092
rect 13727 5052 13820 5080
rect 13814 5040 13820 5052
rect 13872 5080 13878 5092
rect 14277 5083 14335 5089
rect 14277 5080 14289 5083
rect 13872 5052 14289 5080
rect 13872 5040 13878 5052
rect 14277 5049 14289 5052
rect 14323 5080 14335 5083
rect 14642 5080 14648 5092
rect 14323 5052 14648 5080
rect 14323 5049 14335 5052
rect 14277 5043 14335 5049
rect 14642 5040 14648 5052
rect 14700 5040 14706 5092
rect 18785 5083 18843 5089
rect 18785 5049 18797 5083
rect 18831 5080 18843 5083
rect 19144 5083 19202 5089
rect 19144 5080 19156 5083
rect 18831 5052 19156 5080
rect 18831 5049 18843 5052
rect 18785 5043 18843 5049
rect 19144 5049 19156 5052
rect 19190 5080 19202 5083
rect 19242 5080 19248 5092
rect 19190 5052 19248 5080
rect 19190 5049 19202 5052
rect 19144 5043 19202 5049
rect 19242 5040 19248 5052
rect 19300 5040 19306 5092
rect 20901 5083 20959 5089
rect 20901 5049 20913 5083
rect 20947 5080 20959 5083
rect 21726 5080 21732 5092
rect 20947 5052 21732 5080
rect 20947 5049 20959 5052
rect 20901 5043 20959 5049
rect 21726 5040 21732 5052
rect 21784 5040 21790 5092
rect 21928 5080 21956 5120
rect 23917 5117 23929 5120
rect 23963 5148 23975 5151
rect 24946 5148 24952 5160
rect 23963 5120 24952 5148
rect 23963 5117 23975 5120
rect 23917 5111 23975 5117
rect 24946 5108 24952 5120
rect 25004 5108 25010 5160
rect 22278 5080 22284 5092
rect 21928 5052 22284 5080
rect 22278 5040 22284 5052
rect 22336 5080 22342 5092
rect 22373 5083 22431 5089
rect 22373 5080 22385 5083
rect 22336 5052 22385 5080
rect 22336 5040 22342 5052
rect 22373 5049 22385 5052
rect 22419 5049 22431 5083
rect 22373 5043 22431 5049
rect 23109 5083 23167 5089
rect 23109 5049 23121 5083
rect 23155 5080 23167 5083
rect 23750 5080 23756 5092
rect 23155 5052 23756 5080
rect 23155 5049 23167 5052
rect 23109 5043 23167 5049
rect 23750 5040 23756 5052
rect 23808 5040 23814 5092
rect 24210 5040 24216 5092
rect 24268 5080 24274 5092
rect 25222 5080 25228 5092
rect 24268 5052 25228 5080
rect 24268 5040 24274 5052
rect 25222 5040 25228 5052
rect 25280 5040 25286 5092
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 4062 5012 4068 5024
rect 3467 4984 4068 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5350 5012 5356 5024
rect 5123 4984 5356 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 5012 5503 5015
rect 5994 5012 6000 5024
rect 5491 4984 6000 5012
rect 5491 4981 5503 4984
rect 5445 4975 5503 4981
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 7745 5015 7803 5021
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 8110 5012 8116 5024
rect 7791 4984 8116 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 8110 4972 8116 4984
rect 8168 5012 8174 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 8168 4984 8217 5012
rect 8168 4972 8174 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 9582 5012 9588 5024
rect 9543 4984 9588 5012
rect 8205 4975 8263 4981
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 12618 4972 12624 5024
rect 12676 4972 12682 5024
rect 13446 5012 13452 5024
rect 13407 4984 13452 5012
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 15470 5012 15476 5024
rect 15431 4984 15476 5012
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 15838 5012 15844 5024
rect 15751 4984 15844 5012
rect 15838 4972 15844 4984
rect 15896 5012 15902 5024
rect 16853 5015 16911 5021
rect 16853 5012 16865 5015
rect 15896 4984 16865 5012
rect 15896 4972 15902 4984
rect 16853 4981 16865 4984
rect 16899 4981 16911 5015
rect 16853 4975 16911 4981
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 20070 5012 20076 5024
rect 19392 4984 20076 5012
rect 19392 4972 19398 4984
rect 20070 4972 20076 4984
rect 20128 5012 20134 5024
rect 20257 5015 20315 5021
rect 20257 5012 20269 5015
rect 20128 4984 20269 5012
rect 20128 4972 20134 4984
rect 20257 4981 20269 4984
rect 20303 4981 20315 5015
rect 20257 4975 20315 4981
rect 21269 5015 21327 5021
rect 21269 4981 21281 5015
rect 21315 5012 21327 5015
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21315 4984 21833 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 21821 4981 21833 4984
rect 21867 5012 21879 5015
rect 22186 5012 22192 5024
rect 21867 4984 22192 5012
rect 21867 4981 21879 4984
rect 21821 4975 21879 4981
rect 22186 4972 22192 4984
rect 22244 5012 22250 5024
rect 22922 5012 22928 5024
rect 22244 4984 22928 5012
rect 22244 4972 22250 4984
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 1578 4808 1584 4820
rect 1443 4780 1584 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 1762 4808 1768 4820
rect 1723 4780 1768 4808
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 1946 4808 1952 4820
rect 1903 4780 1952 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 5776 4780 6745 4808
rect 5776 4768 5782 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 6733 4771 6791 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 9122 4808 9128 4820
rect 9035 4780 9128 4808
rect 9122 4768 9128 4780
rect 9180 4808 9186 4820
rect 9306 4808 9312 4820
rect 9180 4780 9312 4808
rect 9180 4768 9186 4780
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 11149 4811 11207 4817
rect 11149 4777 11161 4811
rect 11195 4808 11207 4811
rect 11330 4808 11336 4820
rect 11195 4780 11336 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11698 4808 11704 4820
rect 11659 4780 11704 4808
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12342 4808 12348 4820
rect 12303 4780 12348 4808
rect 12342 4768 12348 4780
rect 12400 4808 12406 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12400 4780 12909 4808
rect 12400 4768 12406 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 12897 4771 12955 4777
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 13078 4808 13084 4820
rect 13035 4780 13084 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 3510 4700 3516 4752
rect 3568 4740 3574 4752
rect 3789 4743 3847 4749
rect 3789 4740 3801 4743
rect 3568 4712 3801 4740
rect 3568 4700 3574 4712
rect 3789 4709 3801 4712
rect 3835 4709 3847 4743
rect 3789 4703 3847 4709
rect 5534 4700 5540 4752
rect 5592 4749 5598 4752
rect 5592 4743 5656 4749
rect 5592 4709 5610 4743
rect 5644 4709 5656 4743
rect 5592 4703 5656 4709
rect 8481 4743 8539 4749
rect 8481 4709 8493 4743
rect 8527 4740 8539 4743
rect 8846 4740 8852 4752
rect 8527 4712 8852 4740
rect 8527 4709 8539 4712
rect 8481 4703 8539 4709
rect 5592 4700 5598 4703
rect 8846 4700 8852 4712
rect 8904 4700 8910 4752
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 9732 4712 10180 4740
rect 9732 4700 9738 4712
rect 4246 4672 4252 4684
rect 4207 4644 4252 4672
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 5316 4644 5365 4672
rect 5316 4632 5322 4644
rect 5353 4641 5365 4644
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 9398 4672 9404 4684
rect 8435 4644 9404 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 10042 4681 10048 4684
rect 10036 4672 10048 4681
rect 10003 4644 10048 4672
rect 10036 4635 10048 4644
rect 10042 4632 10048 4635
rect 10100 4632 10106 4684
rect 10152 4672 10180 4712
rect 12802 4700 12808 4752
rect 12860 4740 12866 4752
rect 13004 4740 13032 4771
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 14366 4808 14372 4820
rect 14047 4780 14372 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15562 4808 15568 4820
rect 15344 4780 15568 4808
rect 15344 4768 15350 4780
rect 15562 4768 15568 4780
rect 15620 4808 15626 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15620 4780 15853 4808
rect 15620 4768 15626 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 15841 4771 15899 4777
rect 17589 4811 17647 4817
rect 17589 4777 17601 4811
rect 17635 4808 17647 4811
rect 17678 4808 17684 4820
rect 17635 4780 17684 4808
rect 17635 4777 17647 4780
rect 17589 4771 17647 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18230 4808 18236 4820
rect 18191 4780 18236 4808
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 18414 4768 18420 4820
rect 18472 4808 18478 4820
rect 18874 4808 18880 4820
rect 18472 4780 18880 4808
rect 18472 4768 18478 4780
rect 18874 4768 18880 4780
rect 18932 4808 18938 4820
rect 19337 4811 19395 4817
rect 19337 4808 19349 4811
rect 18932 4780 19349 4808
rect 18932 4768 18938 4780
rect 19337 4777 19349 4780
rect 19383 4777 19395 4811
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 19337 4771 19395 4777
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 21266 4808 21272 4820
rect 21227 4780 21272 4808
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 23106 4768 23112 4820
rect 23164 4808 23170 4820
rect 23477 4811 23535 4817
rect 23477 4808 23489 4811
rect 23164 4780 23489 4808
rect 23164 4768 23170 4780
rect 23477 4777 23489 4780
rect 23523 4808 23535 4811
rect 24029 4811 24087 4817
rect 23523 4780 23888 4808
rect 23523 4777 23535 4780
rect 23477 4771 23535 4777
rect 12860 4712 13032 4740
rect 22005 4743 22063 4749
rect 12860 4700 12866 4712
rect 22005 4709 22017 4743
rect 22051 4740 22063 4743
rect 22833 4743 22891 4749
rect 22833 4740 22845 4743
rect 22051 4712 22845 4740
rect 22051 4709 22063 4712
rect 22005 4703 22063 4709
rect 22833 4709 22845 4712
rect 22879 4740 22891 4743
rect 23750 4740 23756 4752
rect 22879 4712 23756 4740
rect 22879 4709 22891 4712
rect 22833 4703 22891 4709
rect 23750 4700 23756 4712
rect 23808 4700 23814 4752
rect 13906 4672 13912 4684
rect 10152 4644 13912 4672
rect 13906 4632 13912 4644
rect 13964 4632 13970 4684
rect 14090 4672 14096 4684
rect 14051 4644 14096 4672
rect 14090 4632 14096 4644
rect 14148 4672 14154 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 14148 4644 14657 4672
rect 14148 4632 14154 4644
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 16206 4672 16212 4684
rect 16167 4644 16212 4672
rect 14645 4635 14703 4641
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 16482 4681 16488 4684
rect 16476 4672 16488 4681
rect 16443 4644 16488 4672
rect 16476 4635 16488 4644
rect 16482 4632 16488 4635
rect 16540 4632 16546 4684
rect 19242 4672 19248 4684
rect 19203 4644 19248 4672
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 22373 4675 22431 4681
rect 22373 4641 22385 4675
rect 22419 4672 22431 4675
rect 22925 4675 22983 4681
rect 22925 4672 22937 4675
rect 22419 4644 22937 4672
rect 22419 4641 22431 4644
rect 22373 4635 22431 4641
rect 22925 4641 22937 4644
rect 22971 4672 22983 4675
rect 23382 4672 23388 4684
rect 22971 4644 23388 4672
rect 22971 4641 22983 4644
rect 22925 4635 22983 4641
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 23860 4672 23888 4780
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 24118 4808 24124 4820
rect 24075 4780 24124 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24489 4811 24547 4817
rect 24489 4777 24501 4811
rect 24535 4808 24547 4811
rect 24762 4808 24768 4820
rect 24535 4780 24768 4808
rect 24535 4777 24547 4780
rect 24489 4771 24547 4777
rect 23937 4743 23995 4749
rect 23937 4709 23949 4743
rect 23983 4740 23995 4743
rect 24504 4740 24532 4771
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 25038 4808 25044 4820
rect 24999 4780 25044 4808
rect 25038 4768 25044 4780
rect 25096 4808 25102 4820
rect 25409 4811 25467 4817
rect 25409 4808 25421 4811
rect 25096 4780 25421 4808
rect 25096 4768 25102 4780
rect 25409 4777 25421 4780
rect 25455 4777 25467 4811
rect 25409 4771 25467 4777
rect 23983 4712 24532 4740
rect 23983 4709 23995 4712
rect 23937 4703 23995 4709
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23860 4644 24409 4672
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 2038 4604 2044 4616
rect 1995 4576 2044 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4604 7987 4607
rect 8018 4604 8024 4616
rect 7975 4576 8024 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9766 4604 9772 4616
rect 9364 4576 9772 4604
rect 9364 4564 9370 4576
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 2056 4536 2084 4564
rect 2590 4536 2596 4548
rect 2056 4508 2596 4536
rect 2590 4496 2596 4508
rect 2648 4536 2654 4548
rect 3053 4539 3111 4545
rect 3053 4536 3065 4539
rect 2648 4508 3065 4536
rect 2648 4496 2654 4508
rect 3053 4505 3065 4508
rect 3099 4505 3111 4539
rect 4890 4536 4896 4548
rect 3053 4499 3111 4505
rect 3436 4508 4896 4536
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3436 4477 3464 4508
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 2832 4440 3433 4468
rect 2832 4428 2838 4440
rect 3421 4437 3433 4440
rect 3467 4437 3479 4471
rect 4430 4468 4436 4480
rect 4391 4440 4436 4468
rect 3421 4431 3479 4437
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 8294 4468 8300 4480
rect 8067 4440 8300 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 9674 4468 9680 4480
rect 9539 4440 9680 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9784 4468 9812 4564
rect 13188 4536 13216 4567
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19208 4576 19441 4604
rect 19208 4564 19214 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 20772 4576 21373 4604
rect 20772 4564 20778 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 23014 4604 23020 4616
rect 21508 4576 23020 4604
rect 21508 4564 21514 4576
rect 23014 4564 23020 4576
rect 23072 4564 23078 4616
rect 24673 4607 24731 4613
rect 24673 4573 24685 4607
rect 24719 4604 24731 4607
rect 24854 4604 24860 4616
rect 24719 4576 24860 4604
rect 24719 4573 24731 4576
rect 24673 4567 24731 4573
rect 24854 4564 24860 4576
rect 24912 4564 24918 4616
rect 14090 4536 14096 4548
rect 13188 4508 14096 4536
rect 14090 4496 14096 4508
rect 14148 4496 14154 4548
rect 20806 4536 20812 4548
rect 20272 4508 20812 4536
rect 20272 4480 20300 4508
rect 20806 4496 20812 4508
rect 20864 4496 20870 4548
rect 10502 4468 10508 4480
rect 9784 4440 10508 4468
rect 10502 4428 10508 4440
rect 10560 4428 10566 4480
rect 12526 4468 12532 4480
rect 12487 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 14274 4468 14280 4480
rect 14235 4440 14280 4468
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 14734 4428 14740 4480
rect 14792 4468 14798 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14792 4440 15025 4468
rect 14792 4428 14798 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15013 4431 15071 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 18785 4471 18843 4477
rect 18785 4437 18797 4471
rect 18831 4468 18843 4471
rect 18877 4471 18935 4477
rect 18877 4468 18889 4471
rect 18831 4440 18889 4468
rect 18831 4437 18843 4440
rect 18785 4431 18843 4437
rect 18877 4437 18889 4440
rect 18923 4468 18935 4471
rect 19058 4468 19064 4480
rect 18923 4440 19064 4468
rect 18923 4437 18935 4440
rect 18877 4431 18935 4437
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19886 4468 19892 4480
rect 19847 4440 19892 4468
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 20254 4468 20260 4480
rect 20215 4440 20260 4468
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 20901 4471 20959 4477
rect 20901 4468 20913 4471
rect 20772 4440 20913 4468
rect 20772 4428 20778 4440
rect 20901 4437 20913 4440
rect 20947 4437 20959 4471
rect 22462 4468 22468 4480
rect 22423 4440 22468 4468
rect 20901 4431 20959 4437
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 2041 4267 2099 4273
rect 2041 4264 2053 4267
rect 1719 4236 2053 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 2041 4233 2053 4236
rect 2087 4264 2099 4267
rect 2314 4264 2320 4276
rect 2087 4236 2320 4264
rect 2087 4233 2099 4236
rect 2041 4227 2099 4233
rect 2314 4224 2320 4236
rect 2372 4224 2378 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 4304 4236 4353 4264
rect 4304 4224 4310 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 6454 4264 6460 4276
rect 6319 4236 6460 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 9398 4264 9404 4276
rect 9359 4236 9404 4264
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 10778 4264 10784 4276
rect 10739 4236 10784 4264
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 15013 4267 15071 4273
rect 15013 4233 15025 4267
rect 15059 4264 15071 4267
rect 15286 4264 15292 4276
rect 15059 4236 15292 4264
rect 15059 4233 15071 4236
rect 15013 4227 15071 4233
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 15473 4267 15531 4273
rect 15473 4233 15485 4267
rect 15519 4264 15531 4267
rect 15838 4264 15844 4276
rect 15519 4236 15844 4264
rect 15519 4233 15531 4236
rect 15473 4227 15531 4233
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16482 4264 16488 4276
rect 16443 4236 16488 4264
rect 16482 4224 16488 4236
rect 16540 4224 16546 4276
rect 18874 4224 18880 4276
rect 18932 4264 18938 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 18932 4236 19073 4264
rect 18932 4224 18938 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19061 4227 19119 4233
rect 20901 4267 20959 4273
rect 20901 4233 20913 4267
rect 20947 4264 20959 4267
rect 21266 4264 21272 4276
rect 20947 4236 21272 4264
rect 20947 4233 20959 4236
rect 20901 4227 20959 4233
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 23014 4264 23020 4276
rect 22975 4236 23020 4264
rect 23014 4224 23020 4236
rect 23072 4224 23078 4276
rect 24854 4224 24860 4276
rect 24912 4264 24918 4276
rect 25593 4267 25651 4273
rect 25593 4264 25605 4267
rect 24912 4236 25605 4264
rect 24912 4224 24918 4236
rect 25593 4233 25605 4236
rect 25639 4233 25651 4267
rect 25958 4264 25964 4276
rect 25919 4236 25964 4264
rect 25593 4227 25651 4233
rect 25958 4224 25964 4236
rect 26016 4264 26022 4276
rect 26329 4267 26387 4273
rect 26329 4264 26341 4267
rect 26016 4236 26341 4264
rect 26016 4224 26022 4236
rect 26329 4233 26341 4236
rect 26375 4233 26387 4267
rect 26329 4227 26387 4233
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 1544 4100 2421 4128
rect 1544 4088 1550 4100
rect 2409 4097 2421 4100
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 2424 4060 2452 4091
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 5258 4128 5264 4140
rect 4948 4100 5264 4128
rect 4948 4088 4954 4100
rect 5258 4088 5264 4100
rect 5316 4128 5322 4140
rect 5445 4131 5503 4137
rect 5445 4128 5457 4131
rect 5316 4100 5457 4128
rect 5316 4088 5322 4100
rect 5445 4097 5457 4100
rect 5491 4097 5503 4131
rect 6472 4128 6500 4224
rect 8570 4196 8576 4208
rect 8220 4168 8576 4196
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6472 4100 7389 4128
rect 5445 4091 5503 4097
rect 7377 4097 7389 4100
rect 7423 4128 7435 4131
rect 7926 4128 7932 4140
rect 7423 4100 7932 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8220 4128 8248 4168
rect 8570 4156 8576 4168
rect 8628 4196 8634 4208
rect 15304 4196 15332 4224
rect 18049 4199 18107 4205
rect 8628 4168 9444 4196
rect 15304 4168 16068 4196
rect 8628 4156 8634 4168
rect 9416 4140 9444 4168
rect 8159 4100 8248 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8444 4100 8953 4128
rect 8444 4088 8450 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9398 4088 9404 4140
rect 9456 4088 9462 4140
rect 11330 4128 11336 4140
rect 11291 4100 11336 4128
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12710 4128 12716 4140
rect 12299 4100 12572 4128
rect 12671 4100 12716 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 2498 4060 2504 4072
rect 2424 4032 2504 4060
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 5534 4060 5540 4072
rect 4847 4032 5540 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 6880 4032 8861 4060
rect 6880 4020 6886 4032
rect 8849 4029 8861 4032
rect 8895 4060 8907 4063
rect 9030 4060 9036 4072
rect 8895 4032 9036 4060
rect 8895 4029 8907 4032
rect 8849 4023 8907 4029
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10229 4063 10287 4069
rect 10229 4060 10241 4063
rect 10192 4032 10241 4060
rect 10192 4020 10198 4032
rect 10229 4029 10241 4032
rect 10275 4060 10287 4063
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 10275 4032 11161 4060
rect 10275 4029 10287 4032
rect 10229 4023 10287 4029
rect 11149 4029 11161 4032
rect 11195 4060 11207 4063
rect 12544 4060 12572 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 16040 4137 16068 4168
rect 18049 4165 18061 4199
rect 18095 4165 18107 4199
rect 18049 4159 18107 4165
rect 15933 4131 15991 4137
rect 15933 4128 15945 4131
rect 15488 4100 15945 4128
rect 15488 4072 15516 4100
rect 15933 4097 15945 4100
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16816 4100 16865 4128
rect 16816 4088 16822 4100
rect 16853 4097 16865 4100
rect 16899 4128 16911 4131
rect 17221 4131 17279 4137
rect 17221 4128 17233 4131
rect 16899 4100 17233 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17221 4097 17233 4100
rect 17267 4097 17279 4131
rect 17221 4091 17279 4097
rect 12980 4063 13038 4069
rect 12980 4060 12992 4063
rect 11195 4032 12388 4060
rect 12544 4032 12992 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 2676 3995 2734 4001
rect 2676 3961 2688 3995
rect 2722 3992 2734 3995
rect 3050 3992 3056 4004
rect 2722 3964 3056 3992
rect 2722 3961 2734 3964
rect 2676 3955 2734 3961
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 5261 3995 5319 4001
rect 5261 3961 5273 3995
rect 5307 3992 5319 3995
rect 6546 3992 6552 4004
rect 5307 3964 6552 3992
rect 5307 3961 5319 3964
rect 5261 3955 5319 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 6641 3995 6699 4001
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 6687 3964 7328 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 7300 3936 7328 3964
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 10689 3995 10747 4001
rect 10689 3992 10701 3995
rect 10376 3964 10701 3992
rect 10376 3952 10382 3964
rect 10689 3961 10701 3964
rect 10735 3992 10747 3995
rect 11241 3995 11299 4001
rect 11241 3992 11253 3995
rect 10735 3964 11253 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 11241 3961 11253 3964
rect 11287 3992 11299 3995
rect 11422 3992 11428 4004
rect 11287 3964 11428 3992
rect 11287 3961 11299 3964
rect 11241 3955 11299 3961
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 11793 3995 11851 4001
rect 11793 3961 11805 3995
rect 11839 3992 11851 3995
rect 11882 3992 11888 4004
rect 11839 3964 11888 3992
rect 11839 3961 11851 3964
rect 11793 3955 11851 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 12360 3992 12388 4032
rect 12980 4029 12992 4032
rect 13026 4060 13038 4063
rect 14182 4060 14188 4072
rect 13026 4032 14188 4060
rect 13026 4029 13038 4032
rect 12980 4023 13038 4029
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 15470 4060 15476 4072
rect 15427 4032 15476 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 15838 4060 15844 4072
rect 15620 4032 15844 4060
rect 15620 4020 15626 4032
rect 15838 4020 15844 4032
rect 15896 4020 15902 4072
rect 18064 4060 18092 4159
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 20254 4196 20260 4208
rect 18288 4168 18644 4196
rect 18288 4156 18294 4168
rect 18616 4137 18644 4168
rect 19260 4168 20260 4196
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 19260 4128 19288 4168
rect 20254 4156 20260 4168
rect 20312 4156 20318 4208
rect 18601 4091 18659 4097
rect 19168 4100 19288 4128
rect 19168 4060 19196 4100
rect 19886 4088 19892 4140
rect 19944 4088 19950 4140
rect 20898 4088 20904 4140
rect 20956 4128 20962 4140
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20956 4100 21005 4128
rect 20956 4088 20962 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 23658 4128 23664 4140
rect 23619 4100 23664 4128
rect 20993 4091 21051 4097
rect 23658 4088 23664 4100
rect 23716 4088 23722 4140
rect 18064 4032 19196 4060
rect 19613 4063 19671 4069
rect 19613 4029 19625 4063
rect 19659 4060 19671 4063
rect 19904 4060 19932 4088
rect 21266 4069 21272 4072
rect 21260 4060 21272 4069
rect 19659 4032 19932 4060
rect 21179 4032 21272 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 21260 4023 21272 4032
rect 21324 4060 21330 4072
rect 21818 4060 21824 4072
rect 21324 4032 21824 4060
rect 21266 4020 21272 4023
rect 21324 4020 21330 4032
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 13814 3992 13820 4004
rect 12360 3964 13820 3992
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 18417 3995 18475 4001
rect 18417 3992 18429 3995
rect 17788 3964 18429 3992
rect 17788 3936 17816 3964
rect 18417 3961 18429 3964
rect 18463 3961 18475 3995
rect 18417 3955 18475 3961
rect 19889 3995 19947 4001
rect 19889 3961 19901 3995
rect 19935 3992 19947 3995
rect 19978 3992 19984 4004
rect 19935 3964 19984 3992
rect 19935 3961 19947 3964
rect 19889 3955 19947 3961
rect 19978 3952 19984 3964
rect 20036 3952 20042 4004
rect 22278 3952 22284 4004
rect 22336 3992 22342 4004
rect 23477 3995 23535 4001
rect 23477 3992 23489 3995
rect 22336 3964 23489 3992
rect 22336 3952 22342 3964
rect 23477 3961 23489 3964
rect 23523 3992 23535 3995
rect 23906 3995 23964 4001
rect 23906 3992 23918 3995
rect 23523 3964 23918 3992
rect 23523 3961 23535 3964
rect 23477 3955 23535 3961
rect 23906 3961 23918 3964
rect 23952 3961 23964 3995
rect 23906 3955 23964 3961
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 3789 3927 3847 3933
rect 3789 3924 3801 3927
rect 3292 3896 3801 3924
rect 3292 3884 3298 3896
rect 3789 3893 3801 3896
rect 3835 3893 3847 3927
rect 3789 3887 3847 3893
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4893 3927 4951 3933
rect 4893 3924 4905 3927
rect 4028 3896 4905 3924
rect 4028 3884 4034 3896
rect 4893 3893 4905 3896
rect 4939 3893 4951 3927
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 4893 3887 4951 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6788 3896 6837 3924
rect 6788 3884 6794 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 6825 3887 6883 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 7156 3896 7205 3924
rect 7156 3884 7162 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 8389 3927 8447 3933
rect 7340 3896 7385 3924
rect 7340 3884 7346 3896
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 8662 3924 8668 3936
rect 8435 3896 8668 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9861 3927 9919 3933
rect 8812 3896 8857 3924
rect 8812 3884 8818 3896
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 10042 3924 10048 3936
rect 9907 3896 10048 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 14090 3924 14096 3936
rect 14003 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3924 14154 3936
rect 16206 3924 16212 3936
rect 14148 3896 16212 3924
rect 14148 3884 14154 3896
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 18564 3896 18609 3924
rect 18564 3884 18570 3896
rect 19334 3884 19340 3936
rect 19392 3924 19398 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 19392 3896 19441 3924
rect 19392 3884 19398 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19429 3887 19487 3893
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20312 3896 20453 3924
rect 20312 3884 20318 3896
rect 20441 3893 20453 3896
rect 20487 3924 20499 3927
rect 20622 3924 20628 3936
rect 20487 3896 20628 3924
rect 20487 3893 20499 3896
rect 20441 3887 20499 3893
rect 20622 3884 20628 3896
rect 20680 3884 20686 3936
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22373 3927 22431 3933
rect 22373 3924 22385 3927
rect 21968 3896 22385 3924
rect 21968 3884 21974 3896
rect 22373 3893 22385 3896
rect 22419 3893 22431 3927
rect 22373 3887 22431 3893
rect 24946 3884 24952 3936
rect 25004 3924 25010 3936
rect 25041 3927 25099 3933
rect 25041 3924 25053 3927
rect 25004 3896 25053 3924
rect 25004 3884 25010 3896
rect 25041 3893 25053 3896
rect 25087 3893 25099 3927
rect 25041 3887 25099 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 1762 3720 1768 3732
rect 1443 3692 1768 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 2409 3723 2467 3729
rect 2409 3720 2421 3723
rect 2096 3692 2421 3720
rect 2096 3680 2102 3692
rect 2409 3689 2421 3692
rect 2455 3689 2467 3723
rect 4062 3720 4068 3732
rect 4023 3692 4068 3720
rect 2409 3683 2467 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 4212 3692 5089 3720
rect 4212 3680 4218 3692
rect 5077 3689 5089 3692
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5592 3692 5641 3720
rect 5592 3680 5598 3692
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 5629 3683 5687 3689
rect 5813 3723 5871 3729
rect 5813 3689 5825 3723
rect 5859 3720 5871 3723
rect 5994 3720 6000 3732
rect 5859 3692 6000 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 1857 3655 1915 3661
rect 1857 3652 1869 3655
rect 1636 3624 1869 3652
rect 1636 3612 1642 3624
rect 1857 3621 1869 3624
rect 1903 3621 1915 3655
rect 1857 3615 1915 3621
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 3694 3652 3700 3664
rect 3384 3624 3700 3652
rect 3384 3612 3390 3624
rect 3694 3612 3700 3624
rect 3752 3652 3758 3664
rect 4525 3655 4583 3661
rect 4525 3652 4537 3655
rect 3752 3624 4537 3652
rect 3752 3612 3758 3624
rect 4525 3621 4537 3624
rect 4571 3621 4583 3655
rect 5644 3652 5672 3683
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 6181 3723 6239 3729
rect 6181 3689 6193 3723
rect 6227 3720 6239 3723
rect 6362 3720 6368 3732
rect 6227 3692 6368 3720
rect 6227 3689 6239 3692
rect 6181 3683 6239 3689
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 7377 3723 7435 3729
rect 7377 3720 7389 3723
rect 7248 3692 7389 3720
rect 7248 3680 7254 3692
rect 7377 3689 7389 3692
rect 7423 3689 7435 3723
rect 7377 3683 7435 3689
rect 8294 3680 8300 3732
rect 8352 3720 8358 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 8352 3692 9413 3720
rect 8352 3680 8358 3692
rect 9401 3689 9413 3692
rect 9447 3720 9459 3723
rect 9490 3720 9496 3732
rect 9447 3692 9496 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 10100 3692 11069 3720
rect 10100 3680 10106 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11057 3683 11115 3689
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11609 3723 11667 3729
rect 11609 3720 11621 3723
rect 11388 3692 11621 3720
rect 11388 3680 11394 3692
rect 11609 3689 11621 3692
rect 11655 3689 11667 3723
rect 11609 3683 11667 3689
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12584 3692 13001 3720
rect 12584 3680 12590 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 12989 3683 13047 3689
rect 13081 3723 13139 3729
rect 13081 3689 13093 3723
rect 13127 3720 13139 3723
rect 15289 3723 15347 3729
rect 15289 3720 15301 3723
rect 13127 3692 15301 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 15289 3689 15301 3692
rect 15335 3689 15347 3723
rect 15654 3720 15660 3732
rect 15615 3692 15660 3720
rect 15289 3683 15347 3689
rect 8386 3652 8392 3664
rect 5644 3624 6408 3652
rect 8347 3624 8392 3652
rect 4525 3615 4583 3621
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 1452 3556 1777 3584
rect 1452 3544 1458 3556
rect 1765 3553 1777 3556
rect 1811 3584 1823 3587
rect 2222 3584 2228 3596
rect 1811 3556 2228 3584
rect 1811 3553 1823 3556
rect 1765 3547 1823 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3418 3584 3424 3596
rect 3007 3556 3424 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3418 3544 3424 3556
rect 3476 3584 3482 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 3476 3556 4445 3584
rect 3476 3544 3482 3556
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 4540 3556 4844 3584
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2314 3516 2320 3528
rect 2087 3488 2320 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 4540 3516 4568 3556
rect 4706 3516 4712 3528
rect 3436 3488 4568 3516
rect 4667 3488 4712 3516
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 3436 3448 3464 3488
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 1360 3420 3464 3448
rect 3513 3451 3571 3457
rect 1360 3408 1366 3420
rect 3513 3417 3525 3451
rect 3559 3448 3571 3451
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3559 3420 3893 3448
rect 3559 3417 3571 3420
rect 3513 3411 3571 3417
rect 3881 3417 3893 3420
rect 3927 3448 3939 3451
rect 4724 3448 4752 3476
rect 3927 3420 4752 3448
rect 4816 3448 4844 3556
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 6178 3584 6184 3596
rect 5592 3556 6184 3584
rect 5592 3544 5598 3556
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6270 3516 6276 3528
rect 6231 3488 6276 3516
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6380 3525 6408 3624
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 9858 3612 9864 3664
rect 9916 3661 9922 3664
rect 9916 3655 9980 3661
rect 9916 3621 9934 3655
rect 9968 3621 9980 3655
rect 9916 3615 9980 3621
rect 9916 3612 9922 3615
rect 7745 3587 7803 3593
rect 7745 3553 7757 3587
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 6825 3451 6883 3457
rect 6825 3448 6837 3451
rect 4816 3420 6837 3448
rect 3927 3417 3939 3420
rect 3881 3411 3939 3417
rect 6825 3417 6837 3420
rect 6871 3448 6883 3451
rect 7098 3448 7104 3460
rect 6871 3420 7104 3448
rect 6871 3417 6883 3420
rect 6825 3411 6883 3417
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 1854 3340 1860 3392
rect 1912 3380 1918 3392
rect 2314 3380 2320 3392
rect 1912 3352 2320 3380
rect 1912 3340 1918 3352
rect 2314 3340 2320 3352
rect 2372 3340 2378 3392
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3380 2927 3383
rect 3050 3380 3056 3392
rect 2915 3352 3056 3380
rect 2915 3349 2927 3352
rect 2869 3343 2927 3349
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 5074 3380 5080 3392
rect 4212 3352 5080 3380
rect 4212 3340 4218 3352
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 7190 3380 7196 3392
rect 7151 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 7760 3380 7788 3547
rect 7834 3544 7840 3596
rect 7892 3584 7898 3596
rect 7892 3556 7937 3584
rect 7892 3544 7898 3556
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8996 3556 9137 3584
rect 8996 3544 9002 3556
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 9398 3544 9404 3596
rect 9456 3584 9462 3596
rect 9876 3584 9904 3612
rect 9456 3556 9904 3584
rect 12529 3587 12587 3593
rect 9456 3544 9462 3556
rect 12529 3553 12541 3587
rect 12575 3584 12587 3587
rect 12802 3584 12808 3596
rect 12575 3556 12808 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 7926 3516 7932 3528
rect 7887 3488 7932 3516
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8846 3516 8852 3528
rect 8807 3488 8852 3516
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9306 3516 9312 3528
rect 8956 3488 9312 3516
rect 7926 3380 7932 3392
rect 7760 3352 7932 3380
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8956 3389 8984 3488
rect 9306 3476 9312 3488
rect 9364 3516 9370 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9364 3488 9689 3516
rect 9364 3476 9370 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 12161 3451 12219 3457
rect 12161 3417 12173 3451
rect 12207 3448 12219 3451
rect 13096 3448 13124 3683
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 16850 3720 16856 3732
rect 16811 3692 16856 3720
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 17313 3723 17371 3729
rect 17313 3720 17325 3723
rect 17092 3692 17325 3720
rect 17092 3680 17098 3692
rect 17313 3689 17325 3692
rect 17359 3689 17371 3723
rect 17313 3683 17371 3689
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18141 3723 18199 3729
rect 18141 3720 18153 3723
rect 18104 3692 18153 3720
rect 18104 3680 18110 3692
rect 18141 3689 18153 3692
rect 18187 3720 18199 3723
rect 18506 3720 18512 3732
rect 18187 3692 18512 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 19058 3720 19064 3732
rect 19019 3692 19064 3720
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 19153 3723 19211 3729
rect 19153 3689 19165 3723
rect 19199 3720 19211 3723
rect 20533 3723 20591 3729
rect 20533 3720 20545 3723
rect 19199 3692 20545 3720
rect 19199 3689 19211 3692
rect 19153 3683 19211 3689
rect 20533 3689 20545 3692
rect 20579 3720 20591 3723
rect 20622 3720 20628 3732
rect 20579 3692 20628 3720
rect 20579 3689 20591 3692
rect 20533 3683 20591 3689
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 21177 3723 21235 3729
rect 21177 3689 21189 3723
rect 21223 3720 21235 3723
rect 21266 3720 21272 3732
rect 21223 3692 21272 3720
rect 21223 3689 21235 3692
rect 21177 3683 21235 3689
rect 21266 3680 21272 3692
rect 21324 3680 21330 3732
rect 23014 3720 23020 3732
rect 22975 3692 23020 3720
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 24121 3723 24179 3729
rect 24121 3720 24133 3723
rect 23532 3692 24133 3720
rect 23532 3680 23538 3692
rect 24121 3689 24133 3692
rect 24167 3689 24179 3723
rect 24121 3683 24179 3689
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 24581 3723 24639 3729
rect 24581 3720 24593 3723
rect 24268 3692 24593 3720
rect 24268 3680 24274 3692
rect 24581 3689 24593 3692
rect 24627 3689 24639 3723
rect 24581 3683 24639 3689
rect 25038 3680 25044 3732
rect 25096 3720 25102 3732
rect 25133 3723 25191 3729
rect 25133 3720 25145 3723
rect 25096 3692 25145 3720
rect 25096 3680 25102 3692
rect 25133 3689 25145 3692
rect 25179 3689 25191 3723
rect 25133 3683 25191 3689
rect 25593 3723 25651 3729
rect 25593 3689 25605 3723
rect 25639 3720 25651 3723
rect 25958 3720 25964 3732
rect 25639 3692 25964 3720
rect 25639 3689 25651 3692
rect 25593 3683 25651 3689
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 14182 3652 14188 3664
rect 14143 3624 14188 3652
rect 14182 3612 14188 3624
rect 14240 3612 14246 3664
rect 14737 3655 14795 3661
rect 14737 3621 14749 3655
rect 14783 3652 14795 3655
rect 15672 3652 15700 3680
rect 14783 3624 15700 3652
rect 14783 3621 14795 3624
rect 14737 3615 14795 3621
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 17221 3655 17279 3661
rect 17221 3652 17233 3655
rect 17184 3624 17233 3652
rect 17184 3612 17190 3624
rect 17221 3621 17233 3624
rect 17267 3621 17279 3655
rect 17221 3615 17279 3621
rect 23934 3612 23940 3664
rect 23992 3652 23998 3664
rect 24762 3652 24768 3664
rect 23992 3624 24768 3652
rect 23992 3612 23998 3624
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 20990 3544 20996 3596
rect 21048 3584 21054 3596
rect 21910 3593 21916 3596
rect 21637 3587 21695 3593
rect 21637 3584 21649 3587
rect 21048 3556 21649 3584
rect 21048 3544 21054 3556
rect 21637 3553 21649 3556
rect 21683 3553 21695 3587
rect 21904 3584 21916 3593
rect 21871 3556 21916 3584
rect 21637 3547 21695 3553
rect 21904 3547 21916 3556
rect 21910 3544 21916 3547
rect 21968 3544 21974 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 24489 3587 24547 3593
rect 24489 3584 24501 3587
rect 22244 3556 24501 3584
rect 22244 3544 22250 3556
rect 24489 3553 24501 3556
rect 24535 3584 24547 3587
rect 24946 3584 24952 3596
rect 24535 3556 24952 3584
rect 24535 3553 24547 3556
rect 24489 3547 24547 3553
rect 24946 3544 24952 3556
rect 25004 3544 25010 3596
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3516 13323 3519
rect 13354 3516 13360 3528
rect 13311 3488 13360 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13630 3516 13636 3528
rect 13591 3488 13636 3516
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 15010 3516 15016 3528
rect 14971 3488 15016 3516
rect 15010 3476 15016 3488
rect 15068 3516 15074 3528
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 15068 3488 15761 3516
rect 15068 3476 15074 3488
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16206 3516 16212 3528
rect 15979 3488 16212 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 19334 3516 19340 3528
rect 17460 3488 17505 3516
rect 19295 3488 19340 3516
rect 17460 3476 17466 3488
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 24029 3519 24087 3525
rect 24029 3485 24041 3519
rect 24075 3516 24087 3519
rect 24670 3516 24676 3528
rect 24075 3488 24676 3516
rect 24075 3485 24087 3488
rect 24029 3479 24087 3485
rect 12207 3420 13124 3448
rect 12207 3417 12219 3420
rect 12161 3411 12219 3417
rect 15378 3408 15384 3460
rect 15436 3448 15442 3460
rect 16301 3451 16359 3457
rect 16301 3448 16313 3451
rect 15436 3420 16313 3448
rect 15436 3408 15442 3420
rect 16301 3417 16313 3420
rect 16347 3417 16359 3451
rect 19150 3448 19156 3460
rect 16301 3411 16359 3417
rect 18524 3420 19156 3448
rect 18524 3392 18552 3420
rect 19150 3408 19156 3420
rect 19208 3448 19214 3460
rect 19705 3451 19763 3457
rect 19705 3448 19717 3451
rect 19208 3420 19717 3448
rect 19208 3408 19214 3420
rect 19705 3417 19717 3420
rect 19751 3448 19763 3451
rect 21450 3448 21456 3460
rect 19751 3420 21456 3448
rect 19751 3417 19763 3420
rect 19705 3411 19763 3417
rect 21450 3408 21456 3420
rect 21508 3408 21514 3460
rect 22646 3408 22652 3460
rect 22704 3448 22710 3460
rect 24044 3448 24072 3479
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 22704 3420 24072 3448
rect 22704 3408 22710 3420
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 8352 3352 8953 3380
rect 8352 3340 8358 3352
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 8941 3343 8999 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 13998 3380 14004 3392
rect 13959 3352 14004 3380
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 16758 3380 16764 3392
rect 16719 3352 16764 3380
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 18506 3380 18512 3392
rect 18467 3352 18512 3380
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 18690 3380 18696 3392
rect 18651 3352 18696 3380
rect 18690 3340 18696 3352
rect 18748 3340 18754 3392
rect 20162 3380 20168 3392
rect 20123 3352 20168 3380
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 23566 3380 23572 3392
rect 23527 3352 23572 3380
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 3418 3176 3424 3188
rect 2096 3148 3004 3176
rect 3379 3148 3424 3176
rect 2096 3136 2102 3148
rect 2976 3108 3004 3148
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 5258 3176 5264 3188
rect 5219 3148 5264 3176
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6512 3148 6561 3176
rect 6512 3136 6518 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 7892 3148 8125 3176
rect 7892 3136 7898 3148
rect 8113 3145 8125 3148
rect 8159 3176 8171 3179
rect 8202 3176 8208 3188
rect 8159 3148 8208 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 9732 3148 10793 3176
rect 9732 3136 9738 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 10781 3139 10839 3145
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12434 3176 12440 3188
rect 12299 3148 12440 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12434 3136 12440 3148
rect 12492 3176 12498 3188
rect 13354 3176 13360 3188
rect 12492 3148 13360 3176
rect 12492 3136 12498 3148
rect 13354 3136 13360 3148
rect 13412 3176 13418 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13412 3148 14105 3176
rect 13412 3136 13418 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 16206 3176 16212 3188
rect 16167 3148 16212 3176
rect 14093 3139 14151 3145
rect 16206 3136 16212 3148
rect 16264 3136 16270 3188
rect 16666 3176 16672 3188
rect 16579 3148 16672 3176
rect 16666 3136 16672 3148
rect 16724 3176 16730 3188
rect 17402 3176 17408 3188
rect 16724 3148 17408 3176
rect 16724 3136 16730 3148
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19392 3148 19625 3176
rect 19392 3136 19398 3148
rect 19613 3145 19625 3148
rect 19659 3176 19671 3179
rect 20349 3179 20407 3185
rect 20349 3176 20361 3179
rect 19659 3148 20361 3176
rect 19659 3145 19671 3148
rect 19613 3139 19671 3145
rect 20349 3145 20361 3148
rect 20395 3176 20407 3179
rect 20438 3176 20444 3188
rect 20395 3148 20444 3176
rect 20395 3145 20407 3148
rect 20349 3139 20407 3145
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 20809 3179 20867 3185
rect 20809 3145 20821 3179
rect 20855 3176 20867 3179
rect 21910 3176 21916 3188
rect 20855 3148 21916 3176
rect 20855 3145 20867 3148
rect 20809 3139 20867 3145
rect 21910 3136 21916 3148
rect 21968 3136 21974 3188
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 22278 3176 22284 3188
rect 22060 3148 22284 3176
rect 22060 3136 22066 3148
rect 22278 3136 22284 3148
rect 22336 3136 22342 3188
rect 23014 3176 23020 3188
rect 22975 3148 23020 3176
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 23658 3176 23664 3188
rect 23619 3148 23664 3176
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 25958 3136 25964 3188
rect 26016 3176 26022 3188
rect 26329 3179 26387 3185
rect 26329 3176 26341 3179
rect 26016 3148 26341 3176
rect 26016 3136 26022 3148
rect 26329 3145 26341 3148
rect 26375 3145 26387 3179
rect 26329 3139 26387 3145
rect 3694 3108 3700 3120
rect 2976 3080 3700 3108
rect 3694 3068 3700 3080
rect 3752 3068 3758 3120
rect 16482 3068 16488 3120
rect 16540 3108 16546 3120
rect 16945 3111 17003 3117
rect 16945 3108 16957 3111
rect 16540 3080 16957 3108
rect 16540 3068 16546 3080
rect 16945 3077 16957 3080
rect 16991 3077 17003 3111
rect 16945 3071 17003 3077
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 17681 3111 17739 3117
rect 17681 3108 17693 3111
rect 17092 3080 17693 3108
rect 17092 3068 17098 3080
rect 17681 3077 17693 3080
rect 17727 3077 17739 3111
rect 21928 3108 21956 3136
rect 22646 3108 22652 3120
rect 21928 3080 22652 3108
rect 17681 3071 17739 3077
rect 22646 3068 22652 3080
rect 22704 3068 22710 3120
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 2648 3012 3893 3040
rect 2648 3000 2654 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 8294 3040 8300 3052
rect 8255 3012 8300 3040
rect 3881 3003 3939 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3040 10379 3043
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 10367 3012 10609 3040
rect 10367 3009 10379 3012
rect 10321 3003 10379 3009
rect 10597 3009 10609 3012
rect 10643 3040 10655 3043
rect 11333 3043 11391 3049
rect 11333 3040 11345 3043
rect 10643 3012 11345 3040
rect 10643 3009 10655 3012
rect 10597 3003 10655 3009
rect 11333 3009 11345 3012
rect 11379 3009 11391 3043
rect 12710 3040 12716 3052
rect 12671 3012 12716 3040
rect 11333 3003 11391 3009
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1664 2975 1722 2981
rect 1664 2941 1676 2975
rect 1710 2972 1722 2975
rect 2682 2972 2688 2984
rect 1710 2944 2688 2972
rect 1710 2941 1722 2944
rect 1664 2935 1722 2941
rect 1412 2904 1440 2935
rect 2682 2932 2688 2944
rect 2740 2932 2746 2984
rect 4148 2975 4206 2981
rect 4148 2941 4160 2975
rect 4194 2972 4206 2975
rect 4706 2972 4712 2984
rect 4194 2944 4712 2972
rect 4194 2941 4206 2944
rect 4148 2935 4206 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 6638 2972 6644 2984
rect 6420 2944 6644 2972
rect 6420 2932 6426 2944
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 7006 2972 7012 2984
rect 6919 2944 7012 2972
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 7190 2972 7196 2984
rect 7064 2944 7196 2972
rect 7064 2932 7070 2944
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 8386 2932 8392 2984
rect 8444 2972 8450 2984
rect 8570 2981 8576 2984
rect 8564 2972 8576 2981
rect 8444 2944 8576 2972
rect 8444 2932 8450 2944
rect 8564 2935 8576 2944
rect 8628 2972 8634 2984
rect 9398 2972 9404 2984
rect 8628 2944 9404 2972
rect 8570 2932 8576 2935
rect 8628 2932 8634 2944
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 2590 2904 2596 2916
rect 1412 2876 2596 2904
rect 2590 2864 2596 2876
rect 2648 2864 2654 2916
rect 4798 2864 4804 2916
rect 4856 2904 4862 2916
rect 5813 2907 5871 2913
rect 5813 2904 5825 2907
rect 4856 2876 5825 2904
rect 4856 2864 4862 2876
rect 5813 2873 5825 2876
rect 5859 2904 5871 2907
rect 6270 2904 6276 2916
rect 5859 2876 6276 2904
rect 5859 2873 5871 2876
rect 5813 2867 5871 2873
rect 6270 2864 6276 2876
rect 6328 2864 6334 2916
rect 7282 2904 7288 2916
rect 7243 2876 7288 2904
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 2777 2839 2835 2845
rect 2777 2805 2789 2839
rect 2823 2836 2835 2839
rect 3050 2836 3056 2848
rect 2823 2808 3056 2836
rect 2823 2805 2835 2808
rect 2777 2799 2835 2805
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6454 2836 6460 2848
rect 6227 2808 6460 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 7837 2839 7895 2845
rect 7837 2805 7849 2839
rect 7883 2836 7895 2839
rect 7926 2836 7932 2848
rect 7883 2808 7932 2836
rect 7883 2805 7895 2808
rect 7837 2799 7895 2805
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 9677 2839 9735 2845
rect 9677 2805 9689 2839
rect 9723 2836 9735 2839
rect 9858 2836 9864 2848
rect 9723 2808 9864 2836
rect 9723 2805 9735 2808
rect 9677 2799 9735 2805
rect 9858 2796 9864 2808
rect 9916 2836 9922 2848
rect 10336 2836 10364 3003
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 15105 3043 15163 3049
rect 15105 3040 15117 3043
rect 14700 3012 15117 3040
rect 14700 3000 14706 3012
rect 15105 3009 15117 3012
rect 15151 3040 15163 3043
rect 15654 3040 15660 3052
rect 15151 3012 15660 3040
rect 15151 3009 15163 3012
rect 15105 3003 15163 3009
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 16666 3040 16672 3052
rect 15887 3012 16672 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 17184 3012 17325 3040
rect 17184 3000 17190 3012
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 23032 3040 23060 3136
rect 24213 3043 24271 3049
rect 24213 3040 24225 3043
rect 23032 3012 24225 3040
rect 17313 3003 17371 3009
rect 24213 3009 24225 3012
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 25130 3000 25136 3052
rect 25188 3040 25194 3052
rect 25409 3043 25467 3049
rect 25409 3040 25421 3043
rect 25188 3012 25421 3040
rect 25188 3000 25194 3012
rect 25409 3009 25421 3012
rect 25455 3009 25467 3043
rect 25409 3003 25467 3009
rect 11882 2972 11888 2984
rect 11795 2944 11888 2972
rect 11882 2932 11888 2944
rect 11940 2972 11946 2984
rect 12980 2975 13038 2981
rect 12980 2972 12992 2975
rect 11940 2944 12992 2972
rect 11940 2932 11946 2944
rect 12980 2941 12992 2944
rect 13026 2972 13038 2975
rect 14090 2972 14096 2984
rect 13026 2944 14096 2972
rect 13026 2941 13038 2944
rect 12980 2935 13038 2941
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2972 18291 2975
rect 18322 2972 18328 2984
rect 18279 2944 18328 2972
rect 18279 2941 18291 2944
rect 18233 2935 18291 2941
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 18506 2981 18512 2984
rect 18500 2935 18512 2981
rect 18564 2972 18570 2984
rect 20901 2975 20959 2981
rect 18564 2944 18600 2972
rect 18506 2932 18512 2935
rect 18564 2932 18570 2944
rect 20901 2941 20913 2975
rect 20947 2972 20959 2975
rect 20990 2972 20996 2984
rect 20947 2944 20996 2972
rect 20947 2941 20959 2944
rect 20901 2935 20959 2941
rect 20990 2932 20996 2944
rect 21048 2932 21054 2984
rect 23658 2932 23664 2984
rect 23716 2972 23722 2984
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 23716 2944 24133 2972
rect 23716 2932 23722 2944
rect 24121 2941 24133 2944
rect 24167 2941 24179 2975
rect 25222 2972 25228 2984
rect 25183 2944 25228 2972
rect 24121 2935 24179 2941
rect 25222 2932 25228 2944
rect 25280 2972 25286 2984
rect 25961 2975 26019 2981
rect 25961 2972 25973 2975
rect 25280 2944 25973 2972
rect 25280 2932 25286 2944
rect 25961 2941 25973 2944
rect 26007 2941 26019 2975
rect 25961 2935 26019 2941
rect 14642 2864 14648 2916
rect 14700 2904 14706 2916
rect 14737 2907 14795 2913
rect 14737 2904 14749 2907
rect 14700 2876 14749 2904
rect 14700 2864 14706 2876
rect 14737 2873 14749 2876
rect 14783 2904 14795 2907
rect 15565 2907 15623 2913
rect 15565 2904 15577 2907
rect 14783 2876 15577 2904
rect 14783 2873 14795 2876
rect 14737 2867 14795 2873
rect 15565 2873 15577 2876
rect 15611 2873 15623 2907
rect 15565 2867 15623 2873
rect 20438 2864 20444 2916
rect 20496 2904 20502 2916
rect 21146 2907 21204 2913
rect 21146 2904 21158 2907
rect 20496 2876 21158 2904
rect 20496 2864 20502 2876
rect 21146 2873 21158 2876
rect 21192 2873 21204 2907
rect 21146 2867 21204 2873
rect 24210 2864 24216 2916
rect 24268 2904 24274 2916
rect 24765 2907 24823 2913
rect 24765 2904 24777 2907
rect 24268 2876 24777 2904
rect 24268 2864 24274 2876
rect 24765 2873 24777 2876
rect 24811 2904 24823 2907
rect 26050 2904 26056 2916
rect 24811 2876 26056 2904
rect 24811 2873 24823 2876
rect 24765 2867 24823 2873
rect 26050 2864 26056 2876
rect 26108 2864 26114 2916
rect 11146 2836 11152 2848
rect 9916 2808 10364 2836
rect 11107 2808 11152 2836
rect 9916 2796 9922 2808
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11296 2808 11341 2836
rect 11296 2796 11302 2808
rect 12986 2796 12992 2848
rect 13044 2836 13050 2848
rect 13630 2836 13636 2848
rect 13044 2808 13636 2836
rect 13044 2796 13050 2808
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 15194 2836 15200 2848
rect 15155 2808 15200 2836
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 23474 2836 23480 2848
rect 23387 2808 23480 2836
rect 23474 2796 23480 2808
rect 23532 2836 23538 2848
rect 24029 2839 24087 2845
rect 24029 2836 24041 2839
rect 23532 2808 24041 2836
rect 23532 2796 23538 2808
rect 24029 2805 24041 2808
rect 24075 2805 24087 2839
rect 24029 2799 24087 2805
rect 24946 2796 24952 2848
rect 25004 2836 25010 2848
rect 25133 2839 25191 2845
rect 25133 2836 25145 2839
rect 25004 2808 25145 2836
rect 25004 2796 25010 2808
rect 25133 2805 25145 2808
rect 25179 2836 25191 2839
rect 25222 2836 25228 2848
rect 25179 2808 25228 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 1857 2635 1915 2641
rect 1857 2632 1869 2635
rect 1636 2604 1869 2632
rect 1636 2592 1642 2604
rect 1857 2601 1869 2604
rect 1903 2601 1915 2635
rect 2222 2632 2228 2644
rect 2183 2604 2228 2632
rect 1857 2595 1915 2601
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2314 2592 2320 2644
rect 2372 2632 2378 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2372 2604 2421 2632
rect 2372 2592 2378 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 2958 2632 2964 2644
rect 2915 2604 2964 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 6822 2632 6828 2644
rect 4111 2604 6828 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 9732 2604 10149 2632
rect 9732 2592 9738 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 10137 2595 10195 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12069 2635 12127 2641
rect 12069 2601 12081 2635
rect 12115 2632 12127 2635
rect 12526 2632 12532 2644
rect 12115 2604 12532 2632
rect 12115 2601 12127 2604
rect 12069 2595 12127 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 19889 2635 19947 2641
rect 19889 2601 19901 2635
rect 19935 2632 19947 2635
rect 20162 2632 20168 2644
rect 19935 2604 20168 2632
rect 19935 2601 19947 2604
rect 19889 2595 19947 2601
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 20622 2632 20628 2644
rect 20583 2604 20628 2632
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 21266 2632 21272 2644
rect 21227 2604 21272 2632
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 21634 2632 21640 2644
rect 21595 2604 21640 2632
rect 21634 2592 21640 2604
rect 21692 2592 21698 2644
rect 21726 2592 21732 2644
rect 21784 2632 21790 2644
rect 22281 2635 22339 2641
rect 22281 2632 22293 2635
rect 21784 2604 22293 2632
rect 21784 2592 21790 2604
rect 22281 2601 22293 2604
rect 22327 2601 22339 2635
rect 22646 2632 22652 2644
rect 22607 2604 22652 2632
rect 22281 2595 22339 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 23750 2592 23756 2644
rect 23808 2632 23814 2644
rect 24029 2635 24087 2641
rect 24029 2632 24041 2635
rect 23808 2604 24041 2632
rect 23808 2592 23814 2604
rect 24029 2601 24041 2604
rect 24075 2601 24087 2635
rect 24029 2595 24087 2601
rect 24397 2635 24455 2641
rect 24397 2601 24409 2635
rect 24443 2632 24455 2635
rect 25501 2635 25559 2641
rect 25501 2632 25513 2635
rect 24443 2604 25513 2632
rect 24443 2601 24455 2604
rect 24397 2595 24455 2601
rect 25501 2601 25513 2604
rect 25547 2632 25559 2635
rect 25682 2632 25688 2644
rect 25547 2604 25688 2632
rect 25547 2601 25559 2604
rect 25501 2595 25559 2601
rect 25682 2592 25688 2604
rect 25740 2592 25746 2644
rect 1210 2524 1216 2576
rect 1268 2564 1274 2576
rect 3421 2567 3479 2573
rect 3421 2564 3433 2567
rect 1268 2536 3433 2564
rect 1268 2524 1274 2536
rect 3421 2533 3433 2536
rect 3467 2564 3479 2567
rect 4338 2564 4344 2576
rect 3467 2536 4344 2564
rect 3467 2533 3479 2536
rect 3421 2527 3479 2533
rect 4338 2524 4344 2536
rect 4396 2564 4402 2576
rect 4433 2567 4491 2573
rect 4433 2564 4445 2567
rect 4396 2536 4445 2564
rect 4396 2524 4402 2536
rect 4433 2533 4445 2536
rect 4479 2533 4491 2567
rect 4433 2527 4491 2533
rect 6178 2524 6184 2576
rect 6236 2564 6242 2576
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 6236 2536 7297 2564
rect 6236 2524 6242 2536
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 9490 2524 9496 2576
rect 9548 2564 9554 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9548 2536 10241 2564
rect 9548 2524 9554 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 12866 2567 12924 2573
rect 12866 2564 12878 2567
rect 12492 2536 12878 2564
rect 12492 2524 12498 2536
rect 12866 2533 12878 2536
rect 12912 2533 12924 2567
rect 12866 2527 12924 2533
rect 19981 2567 20039 2573
rect 19981 2533 19993 2567
rect 20027 2564 20039 2567
rect 20640 2564 20668 2592
rect 20027 2536 20668 2564
rect 24489 2567 24547 2573
rect 20027 2533 20039 2536
rect 19981 2527 20039 2533
rect 24489 2533 24501 2567
rect 24535 2564 24547 2567
rect 25133 2567 25191 2573
rect 25133 2564 25145 2567
rect 24535 2536 25145 2564
rect 24535 2533 24547 2536
rect 24489 2527 24547 2533
rect 25133 2533 25145 2536
rect 25179 2564 25191 2567
rect 25866 2564 25872 2576
rect 25179 2536 25872 2564
rect 25179 2533 25191 2536
rect 25133 2527 25191 2533
rect 25866 2524 25872 2536
rect 25924 2524 25930 2576
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 5721 2499 5779 2505
rect 2832 2468 2877 2496
rect 2832 2456 2838 2468
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6822 2496 6828 2508
rect 5767 2468 6828 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6822 2456 6828 2468
rect 6880 2456 6886 2508
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2496 7435 2499
rect 7742 2496 7748 2508
rect 7423 2468 7748 2496
rect 7423 2465 7435 2468
rect 7377 2459 7435 2465
rect 3050 2428 3056 2440
rect 2963 2400 3056 2428
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3510 2388 3516 2440
rect 3568 2428 3574 2440
rect 4525 2431 4583 2437
rect 4525 2428 4537 2431
rect 3568 2400 4537 2428
rect 3568 2388 3574 2400
rect 4525 2397 4537 2400
rect 4571 2397 4583 2431
rect 4706 2428 4712 2440
rect 4619 2400 4712 2428
rect 4525 2391 4583 2397
rect 4706 2388 4712 2400
rect 4764 2428 4770 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 4764 2400 5549 2428
rect 4764 2388 4770 2400
rect 5537 2397 5549 2400
rect 5583 2428 5595 2431
rect 6733 2431 6791 2437
rect 5583 2400 6040 2428
rect 5583 2397 5595 2400
rect 5537 2391 5595 2397
rect 3068 2360 3096 2388
rect 5077 2363 5135 2369
rect 5077 2360 5089 2363
rect 3068 2332 5089 2360
rect 5077 2329 5089 2332
rect 5123 2329 5135 2363
rect 5902 2360 5908 2372
rect 5863 2332 5908 2360
rect 5077 2323 5135 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 6012 2360 6040 2400
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7392 2428 7420 2459
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 9122 2496 9128 2508
rect 8619 2468 9128 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10781 2499 10839 2505
rect 10781 2496 10793 2499
rect 10008 2468 10793 2496
rect 10008 2456 10014 2468
rect 10781 2465 10793 2468
rect 10827 2496 10839 2499
rect 11238 2496 11244 2508
rect 10827 2468 11244 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 11238 2456 11244 2468
rect 11296 2456 11302 2508
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 11698 2496 11704 2508
rect 11471 2468 11704 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12710 2496 12716 2508
rect 12667 2468 12716 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 13170 2456 13176 2508
rect 13228 2496 13234 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 13228 2468 14841 2496
rect 13228 2456 13234 2468
rect 14829 2465 14841 2468
rect 14875 2496 14887 2499
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 14875 2468 15853 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 17034 2496 17040 2508
rect 16995 2468 17040 2496
rect 15841 2459 15899 2465
rect 17034 2456 17040 2468
rect 17092 2496 17098 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17092 2468 17601 2496
rect 17092 2456 17098 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2496 21051 2499
rect 25590 2496 25596 2508
rect 21039 2468 21956 2496
rect 25551 2468 25596 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 6779 2400 7420 2428
rect 7561 2431 7619 2437
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7607 2400 7941 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9306 2428 9312 2440
rect 9263 2400 9312 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 7576 2360 7604 2391
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 10042 2428 10048 2440
rect 9631 2400 10048 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10042 2388 10048 2400
rect 10100 2428 10106 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10100 2400 10333 2428
rect 10100 2388 10106 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 10321 2391 10379 2397
rect 15194 2388 15200 2400
rect 15252 2428 15258 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 15252 2400 15945 2428
rect 15252 2388 15258 2400
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2428 16083 2431
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16071 2400 16497 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 16485 2397 16497 2400
rect 16531 2428 16543 2431
rect 16666 2428 16672 2440
rect 16531 2400 16672 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 6012 2332 7604 2360
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 9858 2360 9864 2372
rect 9815 2332 9864 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 9858 2320 9864 2332
rect 9916 2320 9922 2372
rect 16040 2360 16068 2391
rect 16666 2388 16672 2400
rect 16724 2428 16730 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16724 2400 16865 2428
rect 16724 2388 16730 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 19061 2431 19119 2437
rect 19061 2397 19073 2431
rect 19107 2428 19119 2431
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19107 2400 19441 2428
rect 19107 2397 19119 2400
rect 19061 2391 19119 2397
rect 19429 2397 19441 2400
rect 19475 2428 19487 2431
rect 20165 2431 20223 2437
rect 20165 2428 20177 2431
rect 19475 2400 20177 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 20165 2397 20177 2400
rect 20211 2428 20223 2431
rect 20438 2428 20444 2440
rect 20211 2400 20444 2428
rect 20211 2397 20223 2400
rect 20165 2391 20223 2397
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 21726 2428 21732 2440
rect 21639 2400 21732 2428
rect 21726 2388 21732 2400
rect 21784 2388 21790 2440
rect 21928 2437 21956 2468
rect 25590 2456 25596 2468
rect 25648 2456 25654 2508
rect 21913 2431 21971 2437
rect 21913 2397 21925 2431
rect 21959 2428 21971 2431
rect 22002 2428 22008 2440
rect 21959 2400 22008 2428
rect 21959 2397 21971 2400
rect 21913 2391 21971 2397
rect 22002 2388 22008 2400
rect 22060 2388 22066 2440
rect 24670 2428 24676 2440
rect 24631 2400 24676 2428
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 14016 2332 16068 2360
rect 14016 2304 14044 2332
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 17221 2363 17279 2369
rect 17221 2360 17233 2363
rect 16172 2332 17233 2360
rect 16172 2320 16178 2332
rect 17221 2329 17233 2332
rect 17267 2329 17279 2363
rect 17221 2323 17279 2329
rect 19521 2363 19579 2369
rect 19521 2329 19533 2363
rect 19567 2360 19579 2363
rect 21744 2360 21772 2388
rect 19567 2332 21772 2360
rect 19567 2329 19579 2332
rect 19521 2323 19579 2329
rect 22738 2320 22744 2372
rect 22796 2360 22802 2372
rect 25958 2360 25964 2372
rect 22796 2332 25964 2360
rect 22796 2320 22802 2332
rect 25958 2320 25964 2332
rect 26016 2320 26022 2372
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3568 2264 3801 2292
rect 3568 2252 3574 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6273 2295 6331 2301
rect 6273 2292 6285 2295
rect 6236 2264 6285 2292
rect 6236 2252 6242 2264
rect 6273 2261 6285 2264
rect 6319 2261 6331 2295
rect 6273 2255 6331 2261
rect 6546 2252 6552 2304
rect 6604 2292 6610 2304
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 6604 2264 6929 2292
rect 6604 2252 6610 2264
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 8754 2292 8760 2304
rect 8715 2264 8760 2292
rect 6917 2255 6975 2261
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 13998 2292 14004 2304
rect 13959 2264 14004 2292
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 15470 2292 15476 2304
rect 15431 2264 15476 2292
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 17954 2292 17960 2304
rect 17915 2264 17960 2292
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 18598 2292 18604 2304
rect 18559 2264 18604 2292
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 23014 2292 23020 2304
rect 22975 2264 23020 2292
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 23658 2292 23664 2304
rect 23619 2264 23664 2292
rect 23658 2252 23664 2264
rect 23716 2252 23722 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 13722 2048 13728 2100
rect 13780 2088 13786 2100
rect 15378 2088 15384 2100
rect 13780 2060 15384 2088
rect 13780 2048 13786 2060
rect 15378 2048 15384 2060
rect 15436 2048 15442 2100
rect 15378 1912 15384 1964
rect 15436 1952 15442 1964
rect 16298 1952 16304 1964
rect 15436 1924 16304 1952
rect 15436 1912 15442 1924
rect 16298 1912 16304 1924
rect 16356 1912 16362 1964
rect 24302 1368 24308 1420
rect 24360 1408 24366 1420
rect 24762 1408 24768 1420
rect 24360 1380 24768 1408
rect 24360 1368 24366 1380
rect 24762 1368 24768 1380
rect 24820 1368 24826 1420
rect 4614 552 4620 604
rect 4672 592 4678 604
rect 5258 592 5264 604
rect 4672 564 5264 592
rect 4672 552 4678 564
rect 5258 552 5264 564
rect 5316 552 5322 604
<< via1 >>
rect 4068 26256 4120 26308
rect 22468 26256 22520 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 3332 24828 3384 24880
rect 7012 24828 7064 24880
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 22652 23851 22704 23860
rect 22652 23817 22661 23851
rect 22661 23817 22695 23851
rect 22695 23817 22704 23851
rect 22652 23808 22704 23817
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 1860 23604 1912 23656
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 24584 23647 24636 23656
rect 24584 23613 24593 23647
rect 24593 23613 24627 23647
rect 24627 23613 24636 23647
rect 24584 23604 24636 23613
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1492 23264 1544 23316
rect 20628 23196 20680 23248
rect 2504 23128 2556 23180
rect 19524 23171 19576 23180
rect 19524 23137 19533 23171
rect 19533 23137 19567 23171
rect 19567 23137 19576 23171
rect 19524 23128 19576 23137
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 2228 22516 2280 22568
rect 2504 22423 2556 22432
rect 2504 22389 2513 22423
rect 2513 22389 2547 22423
rect 2547 22389 2556 22423
rect 2504 22380 2556 22389
rect 19524 22423 19576 22432
rect 19524 22389 19533 22423
rect 19533 22389 19567 22423
rect 19567 22389 19576 22423
rect 19524 22380 19576 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2412 22040 2464 22092
rect 1400 21904 1452 21956
rect 2228 21836 2280 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 23940 21428 23992 21480
rect 2044 21335 2096 21344
rect 2044 21301 2053 21335
rect 2053 21301 2087 21335
rect 2087 21301 2096 21335
rect 2044 21292 2096 21301
rect 2412 21335 2464 21344
rect 2412 21301 2421 21335
rect 2421 21301 2455 21335
rect 2455 21301 2464 21335
rect 2412 21292 2464 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1492 21088 1544 21140
rect 4620 21131 4672 21140
rect 4620 21097 4629 21131
rect 4629 21097 4663 21131
rect 4663 21097 4672 21131
rect 4620 21088 4672 21097
rect 23940 21063 23992 21072
rect 23940 21029 23949 21063
rect 23949 21029 23983 21063
rect 23983 21029 23992 21063
rect 23940 21020 23992 21029
rect 2320 20952 2372 21004
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 23848 20952 23900 21004
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 24676 20544 24728 20596
rect 4436 20408 4488 20460
rect 2320 20340 2372 20392
rect 24584 20383 24636 20392
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 24584 20349 24593 20383
rect 24593 20349 24627 20383
rect 24627 20349 24636 20383
rect 24584 20340 24636 20349
rect 6092 20204 6144 20256
rect 23848 20247 23900 20256
rect 23848 20213 23857 20247
rect 23857 20213 23891 20247
rect 23891 20213 23900 20247
rect 23848 20204 23900 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 2688 20043 2740 20052
rect 2688 20009 2697 20043
rect 2697 20009 2731 20043
rect 2731 20009 2740 20043
rect 2688 20000 2740 20009
rect 24768 20043 24820 20052
rect 24768 20009 24777 20043
rect 24777 20009 24811 20043
rect 24811 20009 24820 20043
rect 24768 20000 24820 20009
rect 2412 19864 2464 19916
rect 2688 19864 2740 19916
rect 23940 19796 23992 19848
rect 23848 19728 23900 19780
rect 1952 19703 2004 19712
rect 1952 19669 1961 19703
rect 1961 19669 1995 19703
rect 1995 19669 2004 19703
rect 1952 19660 2004 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2504 19295 2556 19304
rect 2504 19261 2513 19295
rect 2513 19261 2547 19295
rect 2547 19261 2556 19295
rect 2504 19252 2556 19261
rect 2688 19252 2740 19304
rect 9220 19252 9272 19304
rect 17408 19252 17460 19304
rect 24584 19295 24636 19304
rect 24584 19261 24593 19295
rect 24593 19261 24627 19295
rect 24627 19261 24636 19295
rect 24584 19252 24636 19261
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2044 19159 2096 19168
rect 2044 19125 2053 19159
rect 2053 19125 2087 19159
rect 2087 19125 2096 19159
rect 2044 19116 2096 19125
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 2596 19116 2648 19168
rect 18328 19159 18380 19168
rect 18328 19125 18337 19159
rect 18337 19125 18371 19159
rect 18371 19125 18380 19159
rect 18328 19116 18380 19125
rect 23020 19116 23072 19168
rect 23848 19116 23900 19168
rect 24768 19159 24820 19168
rect 24768 19125 24777 19159
rect 24777 19125 24811 19159
rect 24811 19125 24820 19159
rect 24768 19116 24820 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 24676 18912 24728 18964
rect 17408 18887 17460 18896
rect 17408 18853 17417 18887
rect 17417 18853 17451 18887
rect 17451 18853 17460 18887
rect 17408 18844 17460 18853
rect 1676 18776 1728 18828
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 4068 18819 4120 18828
rect 2780 18776 2832 18785
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 17132 18819 17184 18828
rect 17132 18785 17141 18819
rect 17141 18785 17175 18819
rect 17175 18785 17184 18819
rect 17132 18776 17184 18785
rect 22376 18819 22428 18828
rect 22376 18785 22385 18819
rect 22385 18785 22419 18819
rect 22419 18785 22428 18819
rect 22376 18776 22428 18785
rect 23480 18819 23532 18828
rect 23480 18785 23489 18819
rect 23489 18785 23523 18819
rect 23523 18785 23532 18819
rect 23480 18776 23532 18785
rect 24584 18819 24636 18828
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 2872 18708 2924 18760
rect 25964 18640 26016 18692
rect 2596 18615 2648 18624
rect 2596 18581 2605 18615
rect 2605 18581 2639 18615
rect 2639 18581 2648 18615
rect 2596 18572 2648 18581
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 24768 18572 24820 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 24676 18368 24728 18420
rect 2780 18232 2832 18284
rect 4068 18232 4120 18284
rect 23848 18232 23900 18284
rect 24676 18232 24728 18284
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 1952 18164 2004 18216
rect 1676 18096 1728 18148
rect 2136 18071 2188 18080
rect 2136 18037 2145 18071
rect 2145 18037 2179 18071
rect 2179 18037 2188 18071
rect 2136 18028 2188 18037
rect 20720 18164 20772 18216
rect 22928 18164 22980 18216
rect 22376 18096 22428 18148
rect 23388 18096 23440 18148
rect 4068 18028 4120 18080
rect 16304 18028 16356 18080
rect 17132 18071 17184 18080
rect 17132 18037 17141 18071
rect 17141 18037 17175 18071
rect 17175 18037 17184 18071
rect 17132 18028 17184 18037
rect 19432 18028 19484 18080
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 22652 18071 22704 18080
rect 22652 18037 22661 18071
rect 22661 18037 22695 18071
rect 22695 18037 22704 18071
rect 22652 18028 22704 18037
rect 23480 18071 23532 18080
rect 23480 18037 23489 18071
rect 23489 18037 23523 18071
rect 23523 18037 23532 18071
rect 23480 18028 23532 18037
rect 23848 18028 23900 18080
rect 24492 18071 24544 18080
rect 24492 18037 24501 18071
rect 24501 18037 24535 18071
rect 24535 18037 24544 18071
rect 24492 18028 24544 18037
rect 25596 18071 25648 18080
rect 25596 18037 25605 18071
rect 25605 18037 25639 18071
rect 25639 18037 25648 18071
rect 25596 18028 25648 18037
rect 26148 18028 26200 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 4160 17824 4212 17876
rect 23756 17824 23808 17876
rect 2504 17756 2556 17808
rect 19524 17756 19576 17808
rect 20628 17756 20680 17808
rect 1860 17731 1912 17740
rect 1860 17697 1869 17731
rect 1869 17697 1903 17731
rect 1903 17697 1912 17731
rect 1860 17688 1912 17697
rect 2780 17688 2832 17740
rect 2872 17688 2924 17740
rect 3976 17688 4028 17740
rect 4988 17688 5040 17740
rect 19340 17688 19392 17740
rect 21272 17731 21324 17740
rect 21272 17697 21281 17731
rect 21281 17697 21315 17731
rect 21315 17697 21324 17731
rect 21272 17688 21324 17697
rect 22468 17688 22520 17740
rect 23572 17688 23624 17740
rect 25136 17688 25188 17740
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 17408 17663 17460 17672
rect 17408 17629 17417 17663
rect 17417 17629 17451 17663
rect 17451 17629 17460 17663
rect 17408 17620 17460 17629
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 19892 17663 19944 17672
rect 19892 17629 19901 17663
rect 19901 17629 19935 17663
rect 19935 17629 19944 17663
rect 19892 17620 19944 17629
rect 26516 17620 26568 17672
rect 22560 17595 22612 17604
rect 22560 17561 22569 17595
rect 22569 17561 22603 17595
rect 22603 17561 22612 17595
rect 22560 17552 22612 17561
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 1768 17484 1820 17536
rect 2412 17484 2464 17536
rect 2872 17484 2924 17536
rect 3332 17527 3384 17536
rect 3332 17493 3341 17527
rect 3341 17493 3375 17527
rect 3375 17493 3384 17527
rect 3332 17484 3384 17493
rect 3700 17527 3752 17536
rect 3700 17493 3709 17527
rect 3709 17493 3743 17527
rect 3743 17493 3752 17527
rect 3700 17484 3752 17493
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 19248 17527 19300 17536
rect 19248 17493 19257 17527
rect 19257 17493 19291 17527
rect 19291 17493 19300 17527
rect 19248 17484 19300 17493
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 21916 17527 21968 17536
rect 21916 17493 21925 17527
rect 21925 17493 21959 17527
rect 21959 17493 21968 17527
rect 21916 17484 21968 17493
rect 23848 17484 23900 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2780 17323 2832 17332
rect 2780 17289 2789 17323
rect 2789 17289 2823 17323
rect 2823 17289 2832 17323
rect 3976 17323 4028 17332
rect 2780 17280 2832 17289
rect 3976 17289 3985 17323
rect 3985 17289 4019 17323
rect 4019 17289 4028 17323
rect 3976 17280 4028 17289
rect 16028 17323 16080 17332
rect 16028 17289 16037 17323
rect 16037 17289 16071 17323
rect 16071 17289 16080 17323
rect 16028 17280 16080 17289
rect 17500 17280 17552 17332
rect 18604 17280 18656 17332
rect 19892 17280 19944 17332
rect 21272 17323 21324 17332
rect 21272 17289 21281 17323
rect 21281 17289 21315 17323
rect 21315 17289 21324 17323
rect 21272 17280 21324 17289
rect 24124 17280 24176 17332
rect 19708 17255 19760 17264
rect 19708 17221 19717 17255
rect 19717 17221 19751 17255
rect 19751 17221 19760 17255
rect 19708 17212 19760 17221
rect 20536 17212 20588 17264
rect 2136 17144 2188 17196
rect 2872 17144 2924 17196
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 21916 17187 21968 17196
rect 21916 17153 21925 17187
rect 21925 17153 21959 17187
rect 21959 17153 21968 17187
rect 21916 17144 21968 17153
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 1952 17008 2004 17060
rect 3148 17008 3200 17060
rect 5264 17076 5316 17128
rect 15844 17119 15896 17128
rect 15844 17085 15853 17119
rect 15853 17085 15887 17119
rect 15887 17085 15896 17119
rect 15844 17076 15896 17085
rect 19340 17119 19392 17128
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 20628 17076 20680 17128
rect 20996 17008 21048 17060
rect 2320 16940 2372 16992
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 2964 16983 3016 16992
rect 2964 16949 2973 16983
rect 2973 16949 3007 16983
rect 3007 16949 3016 16983
rect 2964 16940 3016 16949
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 4344 16983 4396 16992
rect 4344 16949 4353 16983
rect 4353 16949 4387 16983
rect 4387 16949 4396 16983
rect 4344 16940 4396 16949
rect 4988 16940 5040 16992
rect 16764 16940 16816 16992
rect 18880 16983 18932 16992
rect 18880 16949 18889 16983
rect 18889 16949 18923 16983
rect 18923 16949 18932 16983
rect 18880 16940 18932 16949
rect 20168 16940 20220 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 21364 16940 21416 16992
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 21824 16940 21876 16949
rect 22560 16983 22612 16992
rect 22560 16949 22569 16983
rect 22569 16949 22603 16983
rect 22603 16949 22612 16983
rect 22560 16940 22612 16949
rect 23572 16940 23624 16992
rect 25136 16983 25188 16992
rect 25136 16949 25145 16983
rect 25145 16949 25179 16983
rect 25179 16949 25188 16983
rect 25136 16940 25188 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1952 16736 2004 16788
rect 2136 16736 2188 16788
rect 2320 16736 2372 16788
rect 3148 16736 3200 16788
rect 5540 16779 5592 16788
rect 5540 16745 5549 16779
rect 5549 16745 5583 16779
rect 5583 16745 5592 16779
rect 5540 16736 5592 16745
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 2320 16600 2372 16652
rect 5172 16668 5224 16720
rect 7656 16736 7708 16788
rect 17500 16736 17552 16788
rect 19064 16736 19116 16788
rect 20352 16736 20404 16788
rect 20628 16736 20680 16788
rect 21824 16736 21876 16788
rect 24032 16736 24084 16788
rect 25688 16736 25740 16788
rect 7196 16668 7248 16720
rect 16212 16668 16264 16720
rect 22284 16711 22336 16720
rect 22284 16677 22293 16711
rect 22293 16677 22327 16711
rect 22327 16677 22336 16711
rect 22284 16668 22336 16677
rect 22560 16668 22612 16720
rect 5356 16643 5408 16652
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 2688 16532 2740 16584
rect 2596 16464 2648 16516
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 13360 16600 13412 16652
rect 19524 16600 19576 16652
rect 20444 16600 20496 16652
rect 21272 16643 21324 16652
rect 21272 16609 21281 16643
rect 21281 16609 21315 16643
rect 21315 16609 21324 16643
rect 21272 16600 21324 16609
rect 21548 16600 21600 16652
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 24124 16600 24176 16652
rect 25780 16600 25832 16652
rect 7564 16575 7616 16584
rect 7564 16541 7573 16575
rect 7573 16541 7607 16575
rect 7607 16541 7616 16575
rect 7564 16532 7616 16541
rect 9036 16532 9088 16584
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 19340 16532 19392 16584
rect 1952 16396 2004 16448
rect 3240 16396 3292 16448
rect 3700 16396 3752 16448
rect 6276 16396 6328 16448
rect 18788 16396 18840 16448
rect 20904 16532 20956 16584
rect 22376 16532 22428 16584
rect 22284 16464 22336 16516
rect 24216 16464 24268 16516
rect 19984 16396 20036 16448
rect 20904 16396 20956 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2320 16192 2372 16244
rect 3424 16192 3476 16244
rect 5356 16235 5408 16244
rect 5356 16201 5365 16235
rect 5365 16201 5399 16235
rect 5399 16201 5408 16235
rect 5356 16192 5408 16201
rect 6000 16192 6052 16244
rect 7564 16192 7616 16244
rect 9036 16235 9088 16244
rect 9036 16201 9045 16235
rect 9045 16201 9079 16235
rect 9079 16201 9088 16235
rect 9036 16192 9088 16201
rect 16212 16192 16264 16244
rect 22376 16235 22428 16244
rect 22376 16201 22385 16235
rect 22385 16201 22419 16235
rect 22419 16201 22428 16235
rect 22376 16192 22428 16201
rect 22744 16192 22796 16244
rect 23664 16235 23716 16244
rect 23664 16201 23673 16235
rect 23673 16201 23707 16235
rect 23707 16201 23716 16235
rect 23664 16192 23716 16201
rect 25412 16235 25464 16244
rect 25412 16201 25421 16235
rect 25421 16201 25455 16235
rect 25455 16201 25464 16235
rect 25412 16192 25464 16201
rect 2044 16124 2096 16176
rect 1860 16056 1912 16108
rect 2320 16056 2372 16108
rect 2872 16056 2924 16108
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 14280 16056 14332 16108
rect 15844 16056 15896 16108
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 19064 16056 19116 16108
rect 1676 15988 1728 16040
rect 2136 15988 2188 16040
rect 3240 15988 3292 16040
rect 3516 15920 3568 15972
rect 1492 15852 1544 15904
rect 1860 15895 1912 15904
rect 1860 15861 1869 15895
rect 1869 15861 1903 15895
rect 1903 15861 1912 15895
rect 1860 15852 1912 15861
rect 2136 15852 2188 15904
rect 2504 15852 2556 15904
rect 4344 15852 4396 15904
rect 13544 15988 13596 16040
rect 13820 15988 13872 16040
rect 19248 15988 19300 16040
rect 21548 16056 21600 16108
rect 21088 15988 21140 16040
rect 24032 16056 24084 16108
rect 24216 16099 24268 16108
rect 24216 16065 24225 16099
rect 24225 16065 24259 16099
rect 24259 16065 24268 16099
rect 24216 16056 24268 16065
rect 7104 15920 7156 15972
rect 20260 15920 20312 15972
rect 24676 15920 24728 15972
rect 6368 15852 6420 15904
rect 7196 15852 7248 15904
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 12716 15895 12768 15904
rect 12716 15861 12725 15895
rect 12725 15861 12759 15895
rect 12759 15861 12768 15895
rect 12716 15852 12768 15861
rect 13268 15852 13320 15904
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 16212 15852 16264 15904
rect 17040 15895 17092 15904
rect 17040 15861 17049 15895
rect 17049 15861 17083 15895
rect 17083 15861 17092 15895
rect 17040 15852 17092 15861
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 19156 15852 19208 15904
rect 19524 15852 19576 15904
rect 21180 15852 21232 15904
rect 24952 15852 25004 15904
rect 25780 15895 25832 15904
rect 25780 15861 25789 15895
rect 25789 15861 25823 15895
rect 25823 15861 25832 15895
rect 25780 15852 25832 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1860 15648 1912 15700
rect 4344 15691 4396 15700
rect 4344 15657 4353 15691
rect 4353 15657 4387 15691
rect 4387 15657 4396 15691
rect 4344 15648 4396 15657
rect 2688 15580 2740 15632
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 1952 15555 2004 15564
rect 1952 15521 1961 15555
rect 1961 15521 1995 15555
rect 1995 15521 2004 15555
rect 1952 15512 2004 15521
rect 2780 15512 2832 15564
rect 1952 15376 2004 15428
rect 2320 15444 2372 15496
rect 3700 15580 3752 15632
rect 5080 15648 5132 15700
rect 6276 15691 6328 15700
rect 6276 15657 6285 15691
rect 6285 15657 6319 15691
rect 6319 15657 6328 15691
rect 6276 15648 6328 15657
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 7656 15648 7708 15700
rect 10140 15648 10192 15700
rect 12532 15648 12584 15700
rect 13728 15580 13780 15632
rect 20076 15648 20128 15700
rect 21272 15648 21324 15700
rect 24216 15580 24268 15632
rect 5080 15512 5132 15564
rect 5540 15555 5592 15564
rect 5540 15521 5549 15555
rect 5549 15521 5583 15555
rect 5583 15521 5592 15555
rect 5540 15512 5592 15521
rect 6828 15512 6880 15564
rect 10968 15555 11020 15564
rect 10968 15521 11002 15555
rect 11002 15521 11020 15555
rect 10968 15512 11020 15521
rect 15292 15555 15344 15564
rect 3608 15376 3660 15428
rect 5448 15444 5500 15496
rect 7104 15444 7156 15496
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 6276 15376 6328 15428
rect 9036 15376 9088 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 2688 15308 2740 15360
rect 2872 15308 2924 15360
rect 3516 15308 3568 15360
rect 4344 15308 4396 15360
rect 10140 15351 10192 15360
rect 10140 15317 10149 15351
rect 10149 15317 10183 15351
rect 10183 15317 10192 15351
rect 13452 15444 13504 15496
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 16672 15512 16724 15564
rect 20352 15512 20404 15564
rect 21088 15512 21140 15564
rect 21272 15512 21324 15564
rect 14280 15444 14332 15496
rect 17040 15487 17092 15496
rect 12256 15376 12308 15428
rect 10140 15308 10192 15317
rect 12440 15308 12492 15360
rect 14832 15308 14884 15360
rect 16028 15351 16080 15360
rect 16028 15317 16037 15351
rect 16037 15317 16071 15351
rect 16071 15317 16080 15351
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 16028 15308 16080 15317
rect 18512 15308 18564 15360
rect 19340 15351 19392 15360
rect 19340 15317 19349 15351
rect 19349 15317 19383 15351
rect 19383 15317 19392 15351
rect 19340 15308 19392 15317
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 22100 15308 22152 15360
rect 22836 15308 22888 15360
rect 23664 15308 23716 15360
rect 24860 15308 24912 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 2596 15104 2648 15156
rect 3700 15147 3752 15156
rect 3700 15113 3709 15147
rect 3709 15113 3743 15147
rect 3743 15113 3752 15147
rect 3700 15104 3752 15113
rect 5448 15104 5500 15156
rect 6828 15104 6880 15156
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 15292 15104 15344 15156
rect 2320 14968 2372 15020
rect 2688 14968 2740 15020
rect 7656 14968 7708 15020
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 12440 14968 12492 15020
rect 18972 15104 19024 15156
rect 19524 15104 19576 15156
rect 20260 15036 20312 15088
rect 20076 14968 20128 15020
rect 21272 14968 21324 15020
rect 22468 15011 22520 15020
rect 22468 14977 22477 15011
rect 22477 14977 22511 15011
rect 22511 14977 22520 15011
rect 22468 14968 22520 14977
rect 22652 15011 22704 15020
rect 22652 14977 22661 15011
rect 22661 14977 22695 15011
rect 22695 14977 22704 15011
rect 22652 14968 22704 14977
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 25412 15011 25464 15020
rect 25412 14977 25421 15011
rect 25421 14977 25455 15011
rect 25455 14977 25464 15011
rect 25412 14968 25464 14977
rect 2872 14900 2924 14952
rect 3240 14900 3292 14952
rect 3700 14900 3752 14952
rect 4344 14900 4396 14952
rect 5080 14900 5132 14952
rect 1860 14832 1912 14884
rect 2596 14764 2648 14816
rect 4068 14764 4120 14816
rect 11060 14900 11112 14952
rect 12072 14900 12124 14952
rect 12808 14943 12860 14952
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 14832 14900 14884 14952
rect 18512 14943 18564 14952
rect 11980 14832 12032 14884
rect 14648 14832 14700 14884
rect 17868 14875 17920 14884
rect 17868 14841 17877 14875
rect 17877 14841 17911 14875
rect 17911 14841 17920 14875
rect 18512 14909 18546 14943
rect 18546 14909 18564 14943
rect 18512 14900 18564 14909
rect 23204 14900 23256 14952
rect 24768 14900 24820 14952
rect 25320 14900 25372 14952
rect 17868 14832 17920 14841
rect 19064 14832 19116 14884
rect 20996 14875 21048 14884
rect 5448 14764 5500 14816
rect 7472 14807 7524 14816
rect 7472 14773 7481 14807
rect 7481 14773 7515 14807
rect 7515 14773 7524 14807
rect 7472 14764 7524 14773
rect 7932 14807 7984 14816
rect 7932 14773 7941 14807
rect 7941 14773 7975 14807
rect 7975 14773 7984 14807
rect 7932 14764 7984 14773
rect 9956 14764 10008 14816
rect 10876 14764 10928 14816
rect 11060 14764 11112 14816
rect 12072 14764 12124 14816
rect 12348 14764 12400 14816
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 13820 14764 13872 14816
rect 14740 14764 14792 14816
rect 15476 14764 15528 14816
rect 16488 14764 16540 14816
rect 16672 14807 16724 14816
rect 16672 14773 16681 14807
rect 16681 14773 16715 14807
rect 16715 14773 16724 14807
rect 16672 14764 16724 14773
rect 17040 14807 17092 14816
rect 17040 14773 17049 14807
rect 17049 14773 17083 14807
rect 17083 14773 17092 14807
rect 17040 14764 17092 14773
rect 17316 14764 17368 14816
rect 20352 14764 20404 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 20996 14841 21005 14875
rect 21005 14841 21039 14875
rect 21039 14841 21048 14875
rect 20996 14832 21048 14841
rect 21916 14875 21968 14884
rect 21916 14841 21925 14875
rect 21925 14841 21959 14875
rect 21959 14841 21968 14875
rect 21916 14832 21968 14841
rect 24032 14875 24084 14884
rect 24032 14841 24041 14875
rect 24041 14841 24075 14875
rect 24075 14841 24084 14875
rect 24032 14832 24084 14841
rect 21456 14764 21508 14816
rect 22008 14807 22060 14816
rect 22008 14773 22017 14807
rect 22017 14773 22051 14807
rect 22051 14773 22060 14807
rect 22008 14764 22060 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14560 1636 14612
rect 2412 14560 2464 14612
rect 2872 14560 2924 14612
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 4712 14560 4764 14612
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 12808 14560 12860 14612
rect 14924 14560 14976 14612
rect 20536 14560 20588 14612
rect 21456 14560 21508 14612
rect 22468 14603 22520 14612
rect 22468 14569 22477 14603
rect 22477 14569 22511 14603
rect 22511 14569 22520 14603
rect 22468 14560 22520 14569
rect 23480 14560 23532 14612
rect 23940 14560 23992 14612
rect 25504 14560 25556 14612
rect 1952 14424 2004 14476
rect 3700 14492 3752 14544
rect 4620 14492 4672 14544
rect 4804 14492 4856 14544
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 6736 14424 6788 14476
rect 7748 14424 7800 14476
rect 8392 14467 8444 14476
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 2412 14356 2464 14408
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 4528 14399 4580 14408
rect 2320 14288 2372 14340
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 4068 14288 4120 14340
rect 6184 14356 6236 14408
rect 9588 14424 9640 14476
rect 9956 14467 10008 14476
rect 9956 14433 9990 14467
rect 9990 14433 10008 14467
rect 9956 14424 10008 14433
rect 10140 14492 10192 14544
rect 11704 14492 11756 14544
rect 12440 14535 12492 14544
rect 12440 14501 12474 14535
rect 12474 14501 12492 14535
rect 12440 14492 12492 14501
rect 15292 14492 15344 14544
rect 16396 14492 16448 14544
rect 20260 14492 20312 14544
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 18052 14424 18104 14476
rect 19616 14467 19668 14476
rect 19616 14433 19625 14467
rect 19625 14433 19659 14467
rect 19659 14433 19668 14467
rect 19616 14424 19668 14433
rect 20904 14424 20956 14476
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 14648 14356 14700 14408
rect 15752 14356 15804 14408
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 9312 14288 9364 14340
rect 19340 14288 19392 14340
rect 20076 14356 20128 14408
rect 22744 14492 22796 14544
rect 23664 14492 23716 14544
rect 22652 14424 22704 14476
rect 23388 14424 23440 14476
rect 24768 14424 24820 14476
rect 25228 14467 25280 14476
rect 25228 14433 25237 14467
rect 25237 14433 25271 14467
rect 25271 14433 25280 14467
rect 25228 14424 25280 14433
rect 21640 14356 21692 14408
rect 22744 14399 22796 14408
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 2044 14220 2096 14272
rect 2780 14220 2832 14272
rect 7012 14263 7064 14272
rect 7012 14229 7021 14263
rect 7021 14229 7055 14263
rect 7055 14229 7064 14263
rect 7012 14220 7064 14229
rect 7932 14263 7984 14272
rect 7932 14229 7941 14263
rect 7941 14229 7975 14263
rect 7975 14229 7984 14263
rect 7932 14220 7984 14229
rect 8300 14220 8352 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 11704 14263 11756 14272
rect 11704 14229 11713 14263
rect 11713 14229 11747 14263
rect 11747 14229 11756 14263
rect 11704 14220 11756 14229
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 12440 14220 12492 14272
rect 14832 14220 14884 14272
rect 15568 14220 15620 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 17224 14263 17276 14272
rect 17224 14229 17233 14263
rect 17233 14229 17267 14263
rect 17267 14229 17276 14263
rect 17224 14220 17276 14229
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 20720 14263 20772 14272
rect 20720 14229 20729 14263
rect 20729 14229 20763 14263
rect 20763 14229 20772 14263
rect 20720 14220 20772 14229
rect 24124 14263 24176 14272
rect 24124 14229 24133 14263
rect 24133 14229 24167 14263
rect 24167 14229 24176 14263
rect 24124 14220 24176 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2412 14016 2464 14068
rect 2780 14016 2832 14068
rect 3056 14016 3108 14068
rect 7748 14059 7800 14068
rect 7748 14025 7757 14059
rect 7757 14025 7791 14059
rect 7791 14025 7800 14059
rect 7748 14016 7800 14025
rect 9312 14059 9364 14068
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 11704 14016 11756 14068
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 19248 14016 19300 14068
rect 19616 14059 19668 14068
rect 19616 14025 19625 14059
rect 19625 14025 19659 14059
rect 19659 14025 19668 14059
rect 19616 14016 19668 14025
rect 20904 14059 20956 14068
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 21456 14016 21508 14068
rect 21640 14059 21692 14068
rect 21640 14025 21649 14059
rect 21649 14025 21683 14059
rect 21683 14025 21692 14059
rect 21640 14016 21692 14025
rect 23020 14059 23072 14068
rect 23020 14025 23029 14059
rect 23029 14025 23063 14059
rect 23063 14025 23072 14059
rect 23020 14016 23072 14025
rect 23480 14059 23532 14068
rect 23480 14025 23489 14059
rect 23489 14025 23523 14059
rect 23523 14025 23532 14059
rect 24768 14059 24820 14068
rect 23480 14016 23532 14025
rect 4804 13948 4856 14000
rect 5080 13948 5132 14000
rect 11980 13948 12032 14000
rect 15200 13948 15252 14000
rect 15752 13948 15804 14000
rect 17868 13991 17920 14000
rect 17868 13957 17877 13991
rect 17877 13957 17911 13991
rect 17911 13957 17920 13991
rect 17868 13948 17920 13957
rect 18512 13948 18564 14000
rect 5632 13923 5684 13932
rect 5632 13889 5641 13923
rect 5641 13889 5675 13923
rect 5675 13889 5684 13923
rect 5632 13880 5684 13889
rect 6276 13923 6328 13932
rect 1308 13812 1360 13864
rect 2688 13812 2740 13864
rect 2228 13744 2280 13796
rect 4804 13812 4856 13864
rect 5448 13812 5500 13864
rect 6276 13889 6285 13923
rect 6285 13889 6319 13923
rect 6319 13889 6328 13923
rect 6276 13880 6328 13889
rect 7288 13880 7340 13932
rect 6736 13812 6788 13864
rect 7656 13812 7708 13864
rect 11060 13880 11112 13932
rect 8208 13855 8260 13864
rect 8208 13821 8231 13855
rect 8231 13821 8260 13855
rect 8208 13812 8260 13821
rect 8760 13812 8812 13864
rect 9956 13812 10008 13864
rect 3700 13744 3752 13796
rect 4988 13744 5040 13796
rect 6000 13744 6052 13796
rect 11428 13812 11480 13864
rect 13176 13855 13228 13864
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 16488 13880 16540 13932
rect 18236 13880 18288 13932
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 22008 13880 22060 13932
rect 22468 13880 22520 13932
rect 22652 13923 22704 13932
rect 22652 13889 22661 13923
rect 22661 13889 22695 13923
rect 22695 13889 22704 13923
rect 22652 13880 22704 13889
rect 24124 13880 24176 13932
rect 14832 13812 14884 13864
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 16672 13812 16724 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17408 13812 17460 13864
rect 18512 13855 18564 13864
rect 16396 13744 16448 13796
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 19248 13812 19300 13864
rect 19432 13812 19484 13864
rect 20536 13812 20588 13864
rect 23020 13812 23072 13864
rect 24768 14025 24777 14059
rect 24777 14025 24811 14059
rect 24811 14025 24820 14059
rect 24768 14016 24820 14025
rect 25228 13948 25280 14000
rect 25136 13880 25188 13932
rect 24860 13812 24912 13864
rect 25044 13855 25096 13864
rect 25044 13821 25053 13855
rect 25053 13821 25087 13855
rect 25087 13821 25096 13855
rect 25044 13812 25096 13821
rect 2412 13676 2464 13728
rect 3516 13676 3568 13728
rect 4068 13719 4120 13728
rect 4068 13685 4077 13719
rect 4077 13685 4111 13719
rect 4111 13685 4120 13719
rect 4068 13676 4120 13685
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 12164 13676 12216 13728
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 14648 13719 14700 13728
rect 14648 13685 14657 13719
rect 14657 13685 14691 13719
rect 14691 13685 14700 13719
rect 14648 13676 14700 13685
rect 17132 13676 17184 13728
rect 18328 13676 18380 13728
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 22284 13676 22336 13728
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 23664 13719 23716 13728
rect 23664 13685 23673 13719
rect 23673 13685 23707 13719
rect 23707 13685 23716 13719
rect 23664 13676 23716 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2596 13472 2648 13524
rect 4528 13472 4580 13524
rect 4712 13515 4764 13524
rect 4712 13481 4721 13515
rect 4721 13481 4755 13515
rect 4755 13481 4764 13515
rect 4712 13472 4764 13481
rect 5448 13472 5500 13524
rect 6184 13472 6236 13524
rect 6920 13472 6972 13524
rect 8116 13472 8168 13524
rect 8300 13472 8352 13524
rect 9588 13472 9640 13524
rect 10048 13472 10100 13524
rect 11060 13472 11112 13524
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 12348 13472 12400 13524
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 18052 13472 18104 13524
rect 19248 13515 19300 13524
rect 19248 13481 19257 13515
rect 19257 13481 19291 13515
rect 19291 13481 19300 13515
rect 19248 13472 19300 13481
rect 20076 13515 20128 13524
rect 20076 13481 20085 13515
rect 20085 13481 20119 13515
rect 20119 13481 20128 13515
rect 20076 13472 20128 13481
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 22652 13472 22704 13524
rect 23388 13472 23440 13524
rect 23664 13515 23716 13524
rect 23664 13481 23673 13515
rect 23673 13481 23707 13515
rect 23707 13481 23716 13515
rect 23664 13472 23716 13481
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 2228 13336 2280 13345
rect 1216 13268 1268 13320
rect 3516 13404 3568 13456
rect 5356 13404 5408 13456
rect 9864 13404 9916 13456
rect 14648 13404 14700 13456
rect 4712 13268 4764 13320
rect 7748 13336 7800 13388
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 14372 13336 14424 13388
rect 15108 13336 15160 13388
rect 15292 13336 15344 13388
rect 8760 13268 8812 13320
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 11888 13311 11940 13320
rect 10232 13268 10284 13277
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 12440 13268 12492 13320
rect 12624 13268 12676 13320
rect 14096 13311 14148 13320
rect 8024 13243 8076 13252
rect 8024 13209 8033 13243
rect 8033 13209 8067 13243
rect 8067 13209 8076 13243
rect 8024 13200 8076 13209
rect 13636 13243 13688 13252
rect 13636 13209 13645 13243
rect 13645 13209 13679 13243
rect 13679 13209 13688 13243
rect 13636 13200 13688 13209
rect 3240 13175 3292 13184
rect 3240 13141 3249 13175
rect 3249 13141 3283 13175
rect 3283 13141 3292 13175
rect 3240 13132 3292 13141
rect 3700 13175 3752 13184
rect 3700 13141 3709 13175
rect 3709 13141 3743 13175
rect 3743 13141 3752 13175
rect 3700 13132 3752 13141
rect 4620 13132 4672 13184
rect 9404 13132 9456 13184
rect 10692 13132 10744 13184
rect 11060 13132 11112 13184
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 15476 13268 15528 13320
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 19432 13404 19484 13456
rect 19984 13404 20036 13456
rect 20168 13404 20220 13456
rect 21916 13404 21968 13456
rect 24124 13404 24176 13456
rect 17408 13336 17460 13388
rect 19340 13379 19392 13388
rect 19340 13345 19349 13379
rect 19349 13345 19383 13379
rect 19383 13345 19392 13379
rect 19340 13336 19392 13345
rect 22284 13336 22336 13388
rect 23020 13336 23072 13388
rect 14556 13132 14608 13184
rect 16396 13132 16448 13184
rect 20168 13268 20220 13320
rect 20904 13268 20956 13320
rect 21640 13268 21692 13320
rect 22192 13268 22244 13320
rect 22744 13268 22796 13320
rect 18236 13243 18288 13252
rect 18236 13209 18245 13243
rect 18245 13209 18279 13243
rect 18279 13209 18288 13243
rect 18236 13200 18288 13209
rect 17500 13132 17552 13184
rect 25136 13175 25188 13184
rect 25136 13141 25145 13175
rect 25145 13141 25179 13175
rect 25179 13141 25188 13175
rect 25136 13132 25188 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1308 12928 1360 12980
rect 2228 12860 2280 12912
rect 2320 12792 2372 12844
rect 1952 12724 2004 12776
rect 2688 12724 2740 12776
rect 3424 12928 3476 12980
rect 5356 12928 5408 12980
rect 6000 12928 6052 12980
rect 7748 12971 7800 12980
rect 7748 12937 7757 12971
rect 7757 12937 7791 12971
rect 7791 12937 7800 12971
rect 7748 12928 7800 12937
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9404 12928 9456 12980
rect 10232 12928 10284 12980
rect 10968 12928 11020 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12348 12928 12400 12980
rect 13636 12971 13688 12980
rect 13636 12937 13645 12971
rect 13645 12937 13679 12971
rect 13679 12937 13688 12971
rect 13636 12928 13688 12937
rect 14096 12928 14148 12980
rect 16212 12928 16264 12980
rect 17500 12928 17552 12980
rect 19340 12928 19392 12980
rect 19616 12928 19668 12980
rect 3148 12860 3200 12912
rect 7932 12860 7984 12912
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 9772 12792 9824 12844
rect 14648 12835 14700 12844
rect 14648 12801 14657 12835
rect 14657 12801 14691 12835
rect 14691 12801 14700 12835
rect 14648 12792 14700 12801
rect 18512 12860 18564 12912
rect 22468 12928 22520 12980
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 24124 12928 24176 12980
rect 4712 12724 4764 12776
rect 5264 12724 5316 12776
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 9036 12724 9088 12776
rect 9588 12724 9640 12776
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 13452 12724 13504 12776
rect 17132 12792 17184 12844
rect 17316 12792 17368 12844
rect 20076 12860 20128 12912
rect 23756 12860 23808 12912
rect 24952 12860 25004 12912
rect 22376 12792 22428 12844
rect 23480 12792 23532 12844
rect 15476 12767 15528 12776
rect 15476 12733 15510 12767
rect 15510 12733 15528 12767
rect 7932 12656 7984 12708
rect 9864 12656 9916 12708
rect 10048 12656 10100 12708
rect 10876 12656 10928 12708
rect 12072 12656 12124 12708
rect 15476 12724 15528 12733
rect 17500 12767 17552 12776
rect 17500 12733 17509 12767
rect 17509 12733 17543 12767
rect 17543 12733 17552 12767
rect 17500 12724 17552 12733
rect 17776 12724 17828 12776
rect 16396 12656 16448 12708
rect 19064 12656 19116 12708
rect 20444 12724 20496 12776
rect 20720 12656 20772 12708
rect 21272 12656 21324 12708
rect 25780 12656 25832 12708
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 1952 12588 2004 12597
rect 2964 12631 3016 12640
rect 2964 12597 2973 12631
rect 2973 12597 3007 12631
rect 3007 12597 3016 12631
rect 2964 12588 3016 12597
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 9404 12588 9456 12640
rect 10692 12588 10744 12640
rect 13728 12588 13780 12640
rect 14372 12588 14424 12640
rect 16580 12588 16632 12640
rect 17040 12588 17092 12640
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 18328 12588 18380 12640
rect 21640 12588 21692 12640
rect 23020 12588 23072 12640
rect 24124 12588 24176 12640
rect 24676 12588 24728 12640
rect 25412 12588 25464 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1216 12384 1268 12436
rect 2136 12384 2188 12436
rect 3516 12427 3568 12436
rect 3516 12393 3525 12427
rect 3525 12393 3559 12427
rect 3559 12393 3568 12427
rect 3516 12384 3568 12393
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 4528 12384 4580 12436
rect 4712 12384 4764 12436
rect 8300 12384 8352 12436
rect 9864 12384 9916 12436
rect 11520 12384 11572 12436
rect 11612 12384 11664 12436
rect 13636 12384 13688 12436
rect 13820 12384 13872 12436
rect 14004 12384 14056 12436
rect 15752 12384 15804 12436
rect 17408 12427 17460 12436
rect 17408 12393 17417 12427
rect 17417 12393 17451 12427
rect 17451 12393 17460 12427
rect 17408 12384 17460 12393
rect 19432 12384 19484 12436
rect 20444 12427 20496 12436
rect 20444 12393 20453 12427
rect 20453 12393 20487 12427
rect 20487 12393 20496 12427
rect 20444 12384 20496 12393
rect 20904 12427 20956 12436
rect 20904 12393 20913 12427
rect 20913 12393 20947 12427
rect 20947 12393 20956 12427
rect 20904 12384 20956 12393
rect 21916 12427 21968 12436
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 23940 12384 23992 12436
rect 24124 12384 24176 12436
rect 24860 12427 24912 12436
rect 24860 12393 24869 12427
rect 24869 12393 24903 12427
rect 24903 12393 24912 12427
rect 24860 12384 24912 12393
rect 1676 12248 1728 12300
rect 2596 12248 2648 12300
rect 3424 12316 3476 12368
rect 5356 12248 5408 12300
rect 8576 12316 8628 12368
rect 7380 12248 7432 12300
rect 9588 12316 9640 12368
rect 10416 12316 10468 12368
rect 10692 12316 10744 12368
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 3240 12180 3292 12232
rect 4528 12180 4580 12232
rect 5448 12180 5500 12232
rect 6828 12223 6880 12232
rect 6828 12189 6837 12223
rect 6837 12189 6871 12223
rect 6871 12189 6880 12223
rect 6828 12180 6880 12189
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 1492 12112 1544 12164
rect 2136 12112 2188 12164
rect 4712 12112 4764 12164
rect 4896 12112 4948 12164
rect 6276 12112 6328 12164
rect 9220 12112 9272 12164
rect 15200 12316 15252 12368
rect 15844 12316 15896 12368
rect 13728 12248 13780 12300
rect 14004 12291 14056 12300
rect 14004 12257 14013 12291
rect 14013 12257 14047 12291
rect 14047 12257 14056 12291
rect 14004 12248 14056 12257
rect 15476 12248 15528 12300
rect 16856 12291 16908 12300
rect 16856 12257 16865 12291
rect 16865 12257 16899 12291
rect 16899 12257 16908 12291
rect 16856 12248 16908 12257
rect 20076 12316 20128 12368
rect 22744 12316 22796 12368
rect 18604 12248 18656 12300
rect 19340 12248 19392 12300
rect 23204 12291 23256 12300
rect 23204 12257 23213 12291
rect 23213 12257 23247 12291
rect 23247 12257 23256 12291
rect 23204 12248 23256 12257
rect 13912 12180 13964 12232
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 14648 12180 14700 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 16028 12180 16080 12232
rect 20720 12180 20772 12232
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 22836 12180 22888 12232
rect 24584 12316 24636 12368
rect 23940 12248 23992 12300
rect 23388 12180 23440 12232
rect 23756 12180 23808 12232
rect 25136 12180 25188 12232
rect 22744 12155 22796 12164
rect 22744 12121 22753 12155
rect 22753 12121 22787 12155
rect 22787 12121 22796 12155
rect 22744 12112 22796 12121
rect 22928 12112 22980 12164
rect 2412 12044 2464 12096
rect 2596 12044 2648 12096
rect 5172 12044 5224 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 8852 12044 8904 12096
rect 9956 12087 10008 12096
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 11060 12044 11112 12096
rect 11796 12044 11848 12096
rect 13452 12044 13504 12096
rect 14372 12044 14424 12096
rect 16488 12044 16540 12096
rect 16856 12044 16908 12096
rect 17316 12044 17368 12096
rect 17776 12087 17828 12096
rect 17776 12053 17785 12087
rect 17785 12053 17819 12087
rect 17819 12053 17828 12087
rect 17776 12044 17828 12053
rect 17960 12044 18012 12096
rect 18696 12044 18748 12096
rect 22376 12087 22428 12096
rect 22376 12053 22385 12087
rect 22385 12053 22419 12087
rect 22419 12053 22428 12087
rect 22376 12044 22428 12053
rect 23112 12044 23164 12096
rect 24768 12044 24820 12096
rect 25412 12044 25464 12096
rect 25872 12044 25924 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1676 11840 1728 11892
rect 2412 11840 2464 11892
rect 2688 11840 2740 11892
rect 5540 11840 5592 11892
rect 7196 11840 7248 11892
rect 10784 11883 10836 11892
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 14096 11840 14148 11892
rect 15752 11840 15804 11892
rect 16948 11840 17000 11892
rect 18604 11883 18656 11892
rect 1124 11772 1176 11824
rect 1584 11772 1636 11824
rect 1308 11704 1360 11756
rect 1676 11704 1728 11756
rect 5080 11704 5132 11756
rect 9588 11772 9640 11824
rect 10416 11772 10468 11824
rect 11796 11772 11848 11824
rect 11888 11772 11940 11824
rect 15292 11772 15344 11824
rect 16672 11772 16724 11824
rect 17684 11815 17736 11824
rect 17684 11781 17693 11815
rect 17693 11781 17727 11815
rect 17727 11781 17736 11815
rect 17684 11772 17736 11781
rect 17776 11772 17828 11824
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 7012 11704 7064 11756
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 8852 11704 8904 11756
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 11428 11747 11480 11756
rect 11428 11713 11437 11747
rect 11437 11713 11471 11747
rect 11471 11713 11480 11747
rect 11428 11704 11480 11713
rect 16488 11704 16540 11756
rect 1584 11636 1636 11688
rect 2596 11636 2648 11688
rect 8300 11636 8352 11688
rect 9312 11636 9364 11688
rect 9588 11636 9640 11688
rect 10324 11636 10376 11688
rect 2412 11568 2464 11620
rect 2964 11568 3016 11620
rect 5356 11568 5408 11620
rect 6184 11568 6236 11620
rect 2136 11500 2188 11552
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 5172 11500 5224 11552
rect 7380 11500 7432 11552
rect 8852 11500 8904 11552
rect 9772 11568 9824 11620
rect 12532 11636 12584 11688
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 17776 11636 17828 11688
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 19340 11840 19392 11892
rect 20444 11840 20496 11892
rect 21456 11840 21508 11892
rect 22468 11840 22520 11892
rect 23204 11840 23256 11892
rect 23940 11883 23992 11892
rect 23940 11849 23949 11883
rect 23949 11849 23983 11883
rect 23983 11849 23992 11883
rect 23940 11840 23992 11849
rect 20628 11772 20680 11824
rect 18052 11679 18104 11688
rect 14556 11568 14608 11620
rect 14648 11568 14700 11620
rect 16028 11568 16080 11620
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 19432 11636 19484 11688
rect 22008 11704 22060 11756
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 22928 11636 22980 11688
rect 25412 11636 25464 11688
rect 20076 11568 20128 11620
rect 25044 11568 25096 11620
rect 9588 11543 9640 11552
rect 9588 11509 9597 11543
rect 9597 11509 9631 11543
rect 9631 11509 9640 11543
rect 9588 11500 9640 11509
rect 9864 11500 9916 11552
rect 11612 11500 11664 11552
rect 12532 11500 12584 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 16856 11500 16908 11552
rect 17776 11500 17828 11552
rect 18972 11500 19024 11552
rect 21916 11543 21968 11552
rect 21916 11509 21925 11543
rect 21925 11509 21959 11543
rect 21959 11509 21968 11543
rect 21916 11500 21968 11509
rect 22652 11500 22704 11552
rect 22744 11500 22796 11552
rect 25136 11500 25188 11552
rect 25872 11500 25924 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11296 1452 11348
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 5448 11296 5500 11348
rect 5632 11296 5684 11348
rect 8300 11339 8352 11348
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 9864 11296 9916 11348
rect 14004 11296 14056 11348
rect 14556 11339 14608 11348
rect 14556 11305 14565 11339
rect 14565 11305 14599 11339
rect 14599 11305 14608 11339
rect 14556 11296 14608 11305
rect 16120 11296 16172 11348
rect 16304 11296 16356 11348
rect 16672 11296 16724 11348
rect 19064 11339 19116 11348
rect 19064 11305 19073 11339
rect 19073 11305 19107 11339
rect 19107 11305 19116 11339
rect 19064 11296 19116 11305
rect 20720 11339 20772 11348
rect 20720 11305 20729 11339
rect 20729 11305 20763 11339
rect 20763 11305 20772 11339
rect 20720 11296 20772 11305
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 22008 11339 22060 11348
rect 22008 11305 22017 11339
rect 22017 11305 22051 11339
rect 22051 11305 22060 11339
rect 22008 11296 22060 11305
rect 24860 11339 24912 11348
rect 24860 11305 24869 11339
rect 24869 11305 24903 11339
rect 24903 11305 24912 11339
rect 24860 11296 24912 11305
rect 25044 11296 25096 11348
rect 2872 11228 2924 11280
rect 4804 11228 4856 11280
rect 5540 11228 5592 11280
rect 7840 11228 7892 11280
rect 9128 11228 9180 11280
rect 9588 11228 9640 11280
rect 1400 11160 1452 11212
rect 6276 11160 6328 11212
rect 8208 11160 8260 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 11428 11228 11480 11280
rect 13360 11228 13412 11280
rect 13728 11228 13780 11280
rect 10324 11160 10376 11212
rect 15384 11160 15436 11212
rect 15752 11160 15804 11212
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2044 11024 2096 11076
rect 2412 11024 2464 11076
rect 1492 10956 1544 11008
rect 1676 10956 1728 11008
rect 8024 11092 8076 11144
rect 9864 11092 9916 11144
rect 10140 11092 10192 11144
rect 7196 11067 7248 11076
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 4712 10956 4764 11008
rect 6460 10956 6512 11008
rect 7196 11033 7205 11067
rect 7205 11033 7239 11067
rect 7239 11033 7248 11067
rect 7196 11024 7248 11033
rect 11520 11024 11572 11076
rect 13360 11092 13412 11144
rect 13084 11067 13136 11076
rect 13084 11033 13093 11067
rect 13093 11033 13127 11067
rect 13127 11033 13136 11067
rect 13820 11092 13872 11144
rect 16028 11092 16080 11144
rect 17868 11228 17920 11280
rect 20260 11228 20312 11280
rect 21916 11228 21968 11280
rect 23388 11228 23440 11280
rect 17960 11160 18012 11212
rect 22928 11203 22980 11212
rect 14924 11067 14976 11076
rect 13084 11024 13136 11033
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 17684 11092 17736 11144
rect 18052 11092 18104 11144
rect 22928 11169 22937 11203
rect 22937 11169 22971 11203
rect 22971 11169 22980 11203
rect 22928 11160 22980 11169
rect 23204 11203 23256 11212
rect 23204 11169 23238 11203
rect 23238 11169 23256 11203
rect 23204 11160 23256 11169
rect 17868 11067 17920 11076
rect 17868 11033 17877 11067
rect 17877 11033 17911 11067
rect 17911 11033 17920 11067
rect 17868 11024 17920 11033
rect 18328 11024 18380 11076
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 13176 10956 13228 10965
rect 14832 10956 14884 11008
rect 16212 10956 16264 11008
rect 18144 10956 18196 11008
rect 18604 10956 18656 11008
rect 20352 11092 20404 11144
rect 20812 11092 20864 11144
rect 25412 11135 25464 11144
rect 20536 11024 20588 11076
rect 20904 11067 20956 11076
rect 20904 11033 20913 11067
rect 20913 11033 20947 11067
rect 20947 11033 20956 11067
rect 20904 11024 20956 11033
rect 25412 11101 25421 11135
rect 25421 11101 25455 11135
rect 25455 11101 25464 11135
rect 25412 11092 25464 11101
rect 20076 10956 20128 11008
rect 22468 11024 22520 11076
rect 22928 11024 22980 11076
rect 22652 10956 22704 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 4160 10752 4212 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 6460 10752 6512 10804
rect 4712 10684 4764 10736
rect 7104 10752 7156 10804
rect 9772 10752 9824 10804
rect 11336 10752 11388 10804
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 13728 10752 13780 10804
rect 15384 10752 15436 10804
rect 15660 10752 15712 10804
rect 16580 10752 16632 10804
rect 20076 10795 20128 10804
rect 20076 10761 20085 10795
rect 20085 10761 20119 10795
rect 20119 10761 20128 10795
rect 20076 10752 20128 10761
rect 21272 10752 21324 10804
rect 22284 10795 22336 10804
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 9680 10684 9732 10736
rect 17408 10727 17460 10736
rect 17408 10693 17417 10727
rect 17417 10693 17451 10727
rect 17451 10693 17460 10727
rect 17408 10684 17460 10693
rect 17960 10684 18012 10736
rect 10692 10659 10744 10668
rect 2964 10548 3016 10600
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 11612 10616 11664 10668
rect 22284 10761 22293 10795
rect 22293 10761 22327 10795
rect 22327 10761 22336 10795
rect 22284 10752 22336 10761
rect 22836 10752 22888 10804
rect 24032 10752 24084 10804
rect 25872 10795 25924 10804
rect 21916 10659 21968 10668
rect 21916 10625 21925 10659
rect 21925 10625 21959 10659
rect 21959 10625 21968 10659
rect 21916 10616 21968 10625
rect 6276 10548 6328 10600
rect 10140 10548 10192 10600
rect 16304 10548 16356 10600
rect 18144 10548 18196 10600
rect 1124 10480 1176 10532
rect 1676 10480 1728 10532
rect 4620 10480 4672 10532
rect 10324 10480 10376 10532
rect 10692 10480 10744 10532
rect 13084 10480 13136 10532
rect 13728 10480 13780 10532
rect 15844 10480 15896 10532
rect 17684 10480 17736 10532
rect 21088 10523 21140 10532
rect 21088 10489 21097 10523
rect 21097 10489 21131 10523
rect 21131 10489 21140 10523
rect 21088 10480 21140 10489
rect 25872 10761 25881 10795
rect 25881 10761 25915 10795
rect 25915 10761 25924 10795
rect 25872 10752 25924 10761
rect 24768 10616 24820 10668
rect 24308 10548 24360 10600
rect 25136 10616 25188 10668
rect 1584 10412 1636 10464
rect 6000 10412 6052 10464
rect 7288 10412 7340 10464
rect 8024 10412 8076 10464
rect 10784 10412 10836 10464
rect 11428 10412 11480 10464
rect 13360 10412 13412 10464
rect 13636 10412 13688 10464
rect 17408 10412 17460 10464
rect 18052 10412 18104 10464
rect 19340 10412 19392 10464
rect 20812 10455 20864 10464
rect 20812 10421 20821 10455
rect 20821 10421 20855 10455
rect 20855 10421 20864 10455
rect 20812 10412 20864 10421
rect 21824 10412 21876 10464
rect 23204 10412 23256 10464
rect 23664 10412 23716 10464
rect 24308 10412 24360 10464
rect 24676 10412 24728 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1952 10208 2004 10260
rect 2872 10208 2924 10260
rect 3240 10208 3292 10260
rect 6276 10251 6328 10260
rect 6276 10217 6285 10251
rect 6285 10217 6319 10251
rect 6319 10217 6328 10251
rect 6276 10208 6328 10217
rect 7840 10208 7892 10260
rect 2136 10072 2188 10124
rect 3608 10140 3660 10192
rect 4252 10183 4304 10192
rect 4252 10149 4261 10183
rect 4261 10149 4295 10183
rect 4295 10149 4304 10183
rect 4252 10140 4304 10149
rect 5448 10140 5500 10192
rect 7748 10140 7800 10192
rect 9588 10208 9640 10260
rect 11428 10251 11480 10260
rect 11428 10217 11437 10251
rect 11437 10217 11471 10251
rect 11471 10217 11480 10251
rect 11428 10208 11480 10217
rect 11520 10208 11572 10260
rect 12532 10208 12584 10260
rect 13176 10208 13228 10260
rect 13544 10208 13596 10260
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 15292 10251 15344 10260
rect 15292 10217 15301 10251
rect 15301 10217 15335 10251
rect 15335 10217 15344 10251
rect 15292 10208 15344 10217
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 19524 10208 19576 10260
rect 21916 10251 21968 10260
rect 21916 10217 21925 10251
rect 21925 10217 21959 10251
rect 21959 10217 21968 10251
rect 21916 10208 21968 10217
rect 22652 10251 22704 10260
rect 22652 10217 22661 10251
rect 22661 10217 22695 10251
rect 22695 10217 22704 10251
rect 22652 10208 22704 10217
rect 23020 10208 23072 10260
rect 24308 10208 24360 10260
rect 8484 10183 8536 10192
rect 8484 10149 8493 10183
rect 8493 10149 8527 10183
rect 8527 10149 8536 10183
rect 8484 10140 8536 10149
rect 10048 10140 10100 10192
rect 16580 10183 16632 10192
rect 16580 10149 16614 10183
rect 16614 10149 16632 10183
rect 16580 10140 16632 10149
rect 19432 10140 19484 10192
rect 21548 10140 21600 10192
rect 22376 10140 22428 10192
rect 4712 10072 4764 10124
rect 3056 10047 3108 10056
rect 2412 9979 2464 9988
rect 2412 9945 2421 9979
rect 2421 9945 2455 9979
rect 2455 9945 2464 9979
rect 2412 9936 2464 9945
rect 3056 10013 3065 10047
rect 3065 10013 3099 10047
rect 3099 10013 3108 10047
rect 3056 10004 3108 10013
rect 4068 10004 4120 10056
rect 8392 10072 8444 10124
rect 12532 10072 12584 10124
rect 15752 10072 15804 10124
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 22008 10072 22060 10124
rect 23480 10072 23532 10124
rect 25044 10072 25096 10124
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 9956 10004 10008 10056
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 3516 9936 3568 9988
rect 8944 9936 8996 9988
rect 9496 9936 9548 9988
rect 16120 9979 16172 9988
rect 16120 9945 16129 9979
rect 16129 9945 16163 9979
rect 16163 9945 16172 9979
rect 16120 9936 16172 9945
rect 3976 9868 4028 9920
rect 5080 9868 5132 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 8208 9868 8260 9920
rect 10968 9868 11020 9920
rect 13452 9868 13504 9920
rect 17224 9868 17276 9920
rect 17684 9868 17736 9920
rect 18420 9868 18472 9920
rect 18880 9868 18932 9920
rect 19340 10004 19392 10056
rect 20260 10004 20312 10056
rect 20996 10004 21048 10056
rect 20720 9936 20772 9988
rect 21916 10004 21968 10056
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 24860 10047 24912 10056
rect 23204 10004 23256 10013
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 24032 9936 24084 9988
rect 24584 9936 24636 9988
rect 19248 9911 19300 9920
rect 19248 9877 19257 9911
rect 19257 9877 19291 9911
rect 19291 9877 19300 9911
rect 19248 9868 19300 9877
rect 21732 9868 21784 9920
rect 22284 9868 22336 9920
rect 23664 9868 23716 9920
rect 24676 9868 24728 9920
rect 24860 9868 24912 9920
rect 26056 9868 26108 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 1400 9639 1452 9648
rect 1400 9605 1409 9639
rect 1409 9605 1443 9639
rect 1443 9605 1452 9639
rect 1400 9596 1452 9605
rect 3516 9664 3568 9716
rect 4252 9664 4304 9716
rect 4620 9707 4672 9716
rect 4620 9673 4629 9707
rect 4629 9673 4663 9707
rect 4663 9673 4672 9707
rect 4620 9664 4672 9673
rect 8668 9664 8720 9716
rect 10048 9707 10100 9716
rect 10048 9673 10057 9707
rect 10057 9673 10091 9707
rect 10091 9673 10100 9707
rect 10048 9664 10100 9673
rect 10692 9664 10744 9716
rect 11060 9664 11112 9716
rect 11520 9664 11572 9716
rect 12256 9664 12308 9716
rect 3884 9596 3936 9648
rect 1584 9528 1636 9580
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 5448 9596 5500 9648
rect 7748 9596 7800 9648
rect 8852 9596 8904 9648
rect 2320 9460 2372 9512
rect 3424 9460 3476 9512
rect 7380 9528 7432 9580
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 12440 9596 12492 9648
rect 16580 9664 16632 9716
rect 12900 9596 12952 9648
rect 12532 9528 12584 9580
rect 7656 9460 7708 9512
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 15936 9596 15988 9648
rect 17960 9596 18012 9648
rect 19524 9664 19576 9716
rect 23020 9664 23072 9716
rect 23940 9664 23992 9716
rect 15660 9528 15712 9580
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 23296 9596 23348 9648
rect 23388 9596 23440 9648
rect 24860 9664 24912 9716
rect 23664 9528 23716 9580
rect 16120 9460 16172 9512
rect 17132 9460 17184 9512
rect 17408 9460 17460 9512
rect 18328 9460 18380 9512
rect 18880 9460 18932 9512
rect 21456 9460 21508 9512
rect 22284 9460 22336 9512
rect 22468 9503 22520 9512
rect 22468 9469 22477 9503
rect 22477 9469 22511 9503
rect 22511 9469 22520 9503
rect 22468 9460 22520 9469
rect 24216 9460 24268 9512
rect 24952 9460 25004 9512
rect 2228 9392 2280 9444
rect 5356 9392 5408 9444
rect 7012 9392 7064 9444
rect 7840 9392 7892 9444
rect 13636 9392 13688 9444
rect 14924 9435 14976 9444
rect 14924 9401 14933 9435
rect 14933 9401 14967 9435
rect 14967 9401 14976 9435
rect 14924 9392 14976 9401
rect 20260 9392 20312 9444
rect 3240 9324 3292 9376
rect 5080 9367 5132 9376
rect 5080 9333 5089 9367
rect 5089 9333 5123 9367
rect 5123 9333 5132 9367
rect 5080 9324 5132 9333
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 6736 9324 6788 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 15292 9367 15344 9376
rect 15292 9333 15301 9367
rect 15301 9333 15335 9367
rect 15335 9333 15344 9367
rect 15292 9324 15344 9333
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 17040 9324 17092 9376
rect 18052 9324 18104 9376
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 21548 9367 21600 9376
rect 21548 9333 21557 9367
rect 21557 9333 21591 9367
rect 21591 9333 21600 9367
rect 21548 9324 21600 9333
rect 21916 9367 21968 9376
rect 21916 9333 21925 9367
rect 21925 9333 21959 9367
rect 21959 9333 21968 9367
rect 21916 9324 21968 9333
rect 23480 9367 23532 9376
rect 23480 9333 23489 9367
rect 23489 9333 23523 9367
rect 23523 9333 23532 9367
rect 23480 9324 23532 9333
rect 25504 9367 25556 9376
rect 25504 9333 25513 9367
rect 25513 9333 25547 9367
rect 25547 9333 25556 9367
rect 25504 9324 25556 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1860 9120 1912 9172
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2596 9120 2648 9172
rect 6092 9120 6144 9172
rect 7840 9120 7892 9172
rect 10140 9120 10192 9172
rect 10784 9120 10836 9172
rect 12348 9120 12400 9172
rect 14648 9120 14700 9172
rect 15384 9120 15436 9172
rect 16764 9120 16816 9172
rect 18328 9120 18380 9172
rect 18420 9120 18472 9172
rect 18788 9120 18840 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 21272 9163 21324 9172
rect 21272 9129 21281 9163
rect 21281 9129 21315 9163
rect 21315 9129 21324 9163
rect 21272 9120 21324 9129
rect 22100 9120 22152 9172
rect 23204 9120 23256 9172
rect 2780 9095 2832 9104
rect 2780 9061 2789 9095
rect 2789 9061 2823 9095
rect 2823 9061 2832 9095
rect 2780 9052 2832 9061
rect 3792 9052 3844 9104
rect 6000 9095 6052 9104
rect 6000 9061 6009 9095
rect 6009 9061 6043 9095
rect 6043 9061 6052 9095
rect 6000 9052 6052 9061
rect 8024 9052 8076 9104
rect 2136 8984 2188 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 6460 8984 6512 9036
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 11980 8984 12032 9036
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 4528 8959 4580 8968
rect 2596 8848 2648 8900
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 7012 8916 7064 8968
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 10876 8959 10928 8968
rect 7104 8916 7156 8925
rect 10876 8925 10885 8959
rect 10885 8925 10919 8959
rect 10919 8925 10928 8959
rect 10876 8916 10928 8925
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 12532 8959 12584 8968
rect 10968 8916 11020 8925
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 4896 8848 4948 8900
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 3516 8780 3568 8832
rect 4068 8780 4120 8832
rect 4988 8823 5040 8832
rect 4988 8789 4997 8823
rect 4997 8789 5031 8823
rect 5031 8789 5040 8823
rect 4988 8780 5040 8789
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 7104 8780 7156 8832
rect 9128 8780 9180 8832
rect 11152 8780 11204 8832
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 11704 8780 11756 8832
rect 15844 9052 15896 9104
rect 18052 9095 18104 9104
rect 18052 9061 18061 9095
rect 18061 9061 18095 9095
rect 18095 9061 18104 9095
rect 18052 9052 18104 9061
rect 18144 9095 18196 9104
rect 18144 9061 18153 9095
rect 18153 9061 18187 9095
rect 18187 9061 18196 9095
rect 19064 9095 19116 9104
rect 18144 9052 18196 9061
rect 19064 9061 19073 9095
rect 19073 9061 19107 9095
rect 19107 9061 19116 9095
rect 19064 9052 19116 9061
rect 13636 9027 13688 9036
rect 13636 8993 13670 9027
rect 13670 8993 13688 9027
rect 13636 8984 13688 8993
rect 15384 8984 15436 9036
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 19340 8984 19392 9036
rect 13176 8916 13228 8968
rect 16028 8916 16080 8968
rect 18604 8916 18656 8968
rect 19524 8916 19576 8968
rect 16856 8848 16908 8900
rect 20260 8984 20312 9036
rect 21088 8984 21140 9036
rect 23664 9052 23716 9104
rect 25596 9052 25648 9104
rect 20168 8916 20220 8968
rect 20996 8916 21048 8968
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 23388 9027 23440 9036
rect 23388 8993 23422 9027
rect 23422 8993 23440 9027
rect 23388 8984 23440 8993
rect 25780 8848 25832 8900
rect 25964 8848 26016 8900
rect 14004 8780 14056 8832
rect 14832 8780 14884 8832
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 20720 8823 20772 8832
rect 20720 8789 20729 8823
rect 20729 8789 20763 8823
rect 20763 8789 20772 8823
rect 20720 8780 20772 8789
rect 21272 8780 21324 8832
rect 25044 8823 25096 8832
rect 25044 8789 25053 8823
rect 25053 8789 25087 8823
rect 25087 8789 25096 8823
rect 25044 8780 25096 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2872 8576 2924 8628
rect 3608 8576 3660 8628
rect 3792 8619 3844 8628
rect 3792 8585 3801 8619
rect 3801 8585 3835 8619
rect 3835 8585 3844 8619
rect 3792 8576 3844 8585
rect 6092 8576 6144 8628
rect 6184 8576 6236 8628
rect 6368 8576 6420 8628
rect 3332 8508 3384 8560
rect 4344 8551 4396 8560
rect 4344 8517 4353 8551
rect 4353 8517 4387 8551
rect 4387 8517 4396 8551
rect 4344 8508 4396 8517
rect 8208 8576 8260 8628
rect 9588 8576 9640 8628
rect 10048 8576 10100 8628
rect 10692 8576 10744 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 13544 8619 13596 8628
rect 12440 8576 12492 8585
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 16856 8576 16908 8628
rect 18052 8576 18104 8628
rect 18144 8576 18196 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 20260 8576 20312 8628
rect 21364 8576 21416 8628
rect 21916 8576 21968 8628
rect 25596 8619 25648 8628
rect 25596 8585 25605 8619
rect 25605 8585 25639 8619
rect 25639 8585 25648 8619
rect 25596 8576 25648 8585
rect 8024 8508 8076 8560
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 10876 8440 10928 8492
rect 13820 8508 13872 8560
rect 14556 8508 14608 8560
rect 14832 8508 14884 8560
rect 12532 8440 12584 8492
rect 13728 8440 13780 8492
rect 20628 8508 20680 8560
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 18880 8440 18932 8492
rect 21272 8440 21324 8492
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 2136 8415 2188 8424
rect 2136 8381 2170 8415
rect 2170 8381 2188 8415
rect 2136 8372 2188 8381
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 7288 8415 7340 8424
rect 6644 8372 6696 8381
rect 7288 8381 7322 8415
rect 7322 8381 7340 8415
rect 7288 8372 7340 8381
rect 2320 8304 2372 8356
rect 4160 8304 4212 8356
rect 5448 8304 5500 8356
rect 9772 8372 9824 8424
rect 14004 8415 14056 8424
rect 6368 8236 6420 8288
rect 8484 8236 8536 8288
rect 10140 8304 10192 8356
rect 10784 8347 10836 8356
rect 10784 8313 10793 8347
rect 10793 8313 10827 8347
rect 10827 8313 10836 8347
rect 10784 8304 10836 8313
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 14832 8372 14884 8424
rect 16764 8415 16816 8424
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 16856 8415 16908 8424
rect 16856 8381 16865 8415
rect 16865 8381 16899 8415
rect 16899 8381 16908 8415
rect 16856 8372 16908 8381
rect 18420 8372 18472 8424
rect 13360 8304 13412 8356
rect 13912 8347 13964 8356
rect 13912 8313 13921 8347
rect 13921 8313 13955 8347
rect 13955 8313 13964 8347
rect 13912 8304 13964 8313
rect 15660 8304 15712 8356
rect 16488 8304 16540 8356
rect 22284 8372 22336 8424
rect 19340 8304 19392 8356
rect 22744 8372 22796 8424
rect 26240 8372 26292 8424
rect 11980 8279 12032 8288
rect 11980 8245 11989 8279
rect 11989 8245 12023 8279
rect 12023 8245 12032 8279
rect 11980 8236 12032 8245
rect 12716 8236 12768 8288
rect 14464 8236 14516 8288
rect 16764 8236 16816 8288
rect 22652 8236 22704 8288
rect 23388 8236 23440 8288
rect 23664 8236 23716 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2136 8032 2188 8084
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 4528 8032 4580 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 6276 8032 6328 8084
rect 7196 8032 7248 8084
rect 10140 8032 10192 8084
rect 10968 8032 11020 8084
rect 12532 8032 12584 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 2964 7896 3016 7948
rect 2872 7871 2924 7880
rect 2872 7837 2881 7871
rect 2881 7837 2915 7871
rect 2915 7837 2924 7871
rect 2872 7828 2924 7837
rect 4160 7964 4212 8016
rect 3884 7896 3936 7948
rect 3240 7828 3292 7880
rect 4436 7828 4488 7880
rect 5264 7896 5316 7948
rect 5540 7828 5592 7880
rect 6736 7828 6788 7880
rect 7380 7828 7432 7880
rect 8024 7964 8076 8016
rect 11152 7964 11204 8016
rect 11428 7964 11480 8016
rect 13912 8032 13964 8084
rect 14464 8075 14516 8084
rect 14464 8041 14473 8075
rect 14473 8041 14507 8075
rect 14507 8041 14516 8075
rect 14464 8032 14516 8041
rect 14740 8032 14792 8084
rect 16028 8032 16080 8084
rect 17500 8032 17552 8084
rect 19064 8075 19116 8084
rect 19064 8041 19073 8075
rect 19073 8041 19107 8075
rect 19107 8041 19116 8075
rect 19064 8032 19116 8041
rect 19156 8032 19208 8084
rect 19984 8032 20036 8084
rect 20168 8075 20220 8084
rect 20168 8041 20177 8075
rect 20177 8041 20211 8075
rect 20211 8041 20220 8075
rect 20168 8032 20220 8041
rect 20628 8032 20680 8084
rect 21088 8075 21140 8084
rect 21088 8041 21097 8075
rect 21097 8041 21131 8075
rect 21131 8041 21140 8075
rect 21088 8032 21140 8041
rect 21180 8032 21232 8084
rect 21640 8032 21692 8084
rect 22100 8032 22152 8084
rect 14832 8007 14884 8016
rect 14832 7973 14841 8007
rect 14841 7973 14875 8007
rect 14875 7973 14884 8007
rect 14832 7964 14884 7973
rect 19524 7964 19576 8016
rect 20720 7964 20772 8016
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9772 7896 9824 7948
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 13820 7939 13872 7948
rect 13820 7905 13829 7939
rect 13829 7905 13863 7939
rect 13863 7905 13872 7939
rect 13820 7896 13872 7905
rect 13912 7939 13964 7948
rect 13912 7905 13921 7939
rect 13921 7905 13955 7939
rect 13955 7905 13964 7939
rect 13912 7896 13964 7905
rect 15936 7896 15988 7948
rect 16948 7896 17000 7948
rect 17960 7896 18012 7948
rect 19064 7896 19116 7948
rect 19340 7896 19392 7948
rect 22560 7964 22612 8016
rect 23480 8032 23532 8084
rect 23296 7964 23348 8016
rect 23756 7964 23808 8016
rect 25412 8032 25464 8084
rect 27252 7964 27304 8016
rect 22652 7939 22704 7948
rect 8024 7828 8076 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 5356 7760 5408 7812
rect 6460 7803 6512 7812
rect 6460 7769 6469 7803
rect 6469 7769 6503 7803
rect 6503 7769 6512 7803
rect 6460 7760 6512 7769
rect 18604 7803 18656 7812
rect 18604 7769 18613 7803
rect 18613 7769 18647 7803
rect 18647 7769 18656 7803
rect 18604 7760 18656 7769
rect 19432 7760 19484 7812
rect 20444 7828 20496 7880
rect 21180 7828 21232 7880
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 23480 7939 23532 7948
rect 23480 7905 23489 7939
rect 23489 7905 23523 7939
rect 23523 7905 23532 7939
rect 23480 7896 23532 7905
rect 23480 7760 23532 7812
rect 23664 7871 23716 7880
rect 23664 7837 23673 7871
rect 23673 7837 23707 7871
rect 23707 7837 23716 7871
rect 25136 7871 25188 7880
rect 23664 7828 23716 7837
rect 25136 7837 25145 7871
rect 25145 7837 25179 7871
rect 25179 7837 25188 7871
rect 25136 7828 25188 7837
rect 25688 7828 25740 7880
rect 23756 7760 23808 7812
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 8116 7692 8168 7744
rect 8944 7692 8996 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 12716 7692 12768 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 15936 7692 15988 7744
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 22100 7692 22152 7744
rect 24216 7692 24268 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2504 7488 2556 7540
rect 3608 7531 3660 7540
rect 3608 7497 3617 7531
rect 3617 7497 3651 7531
rect 3651 7497 3660 7531
rect 3608 7488 3660 7497
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 6000 7488 6052 7540
rect 8668 7488 8720 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12532 7488 12584 7540
rect 13728 7488 13780 7540
rect 16120 7488 16172 7540
rect 19156 7531 19208 7540
rect 19156 7497 19165 7531
rect 19165 7497 19199 7531
rect 19199 7497 19208 7531
rect 19156 7488 19208 7497
rect 19524 7488 19576 7540
rect 20444 7488 20496 7540
rect 21272 7488 21324 7540
rect 21456 7488 21508 7540
rect 21640 7488 21692 7540
rect 22008 7531 22060 7540
rect 22008 7497 22017 7531
rect 22017 7497 22051 7531
rect 22051 7497 22060 7531
rect 22008 7488 22060 7497
rect 23664 7488 23716 7540
rect 23940 7488 23992 7540
rect 5264 7420 5316 7472
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 3884 7352 3936 7404
rect 5540 7352 5592 7404
rect 6368 7420 6420 7472
rect 9496 7420 9548 7472
rect 2872 7284 2924 7336
rect 3608 7284 3660 7336
rect 6828 7284 6880 7336
rect 7196 7352 7248 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 9220 7395 9272 7404
rect 7380 7352 7432 7361
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 10876 7352 10928 7404
rect 21180 7463 21232 7472
rect 21180 7429 21189 7463
rect 21189 7429 21223 7463
rect 21223 7429 21232 7463
rect 21180 7420 21232 7429
rect 17500 7352 17552 7404
rect 17776 7352 17828 7404
rect 20444 7395 20496 7404
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9496 7284 9548 7336
rect 13176 7284 13228 7336
rect 13636 7327 13688 7336
rect 13636 7293 13670 7327
rect 13670 7293 13688 7327
rect 3884 7216 3936 7268
rect 6460 7216 6512 7268
rect 13636 7284 13688 7293
rect 14556 7284 14608 7336
rect 16580 7284 16632 7336
rect 16764 7327 16816 7336
rect 16764 7293 16773 7327
rect 16773 7293 16807 7327
rect 16807 7293 16816 7327
rect 16764 7284 16816 7293
rect 18052 7284 18104 7336
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 21088 7352 21140 7404
rect 22652 7395 22704 7404
rect 22652 7361 22661 7395
rect 22661 7361 22695 7395
rect 22695 7361 22704 7395
rect 22652 7352 22704 7361
rect 13728 7216 13780 7268
rect 14280 7216 14332 7268
rect 17684 7216 17736 7268
rect 20628 7284 20680 7336
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 25136 7488 25188 7540
rect 25412 7488 25464 7540
rect 25688 7488 25740 7540
rect 24952 7352 25004 7404
rect 18604 7216 18656 7268
rect 20812 7216 20864 7268
rect 22376 7259 22428 7268
rect 22376 7225 22385 7259
rect 22385 7225 22419 7259
rect 22419 7225 22428 7259
rect 22376 7216 22428 7225
rect 1584 7148 1636 7200
rect 2596 7148 2648 7200
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3792 7148 3844 7200
rect 4436 7148 4488 7200
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7748 7148 7800 7200
rect 8024 7191 8076 7200
rect 8024 7157 8033 7191
rect 8033 7157 8067 7191
rect 8067 7157 8076 7191
rect 8024 7148 8076 7157
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 8944 7148 8996 7157
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 10048 7191 10100 7200
rect 9036 7148 9088 7157
rect 10048 7157 10057 7191
rect 10057 7157 10091 7191
rect 10091 7157 10100 7191
rect 10048 7148 10100 7157
rect 10140 7191 10192 7200
rect 10140 7157 10149 7191
rect 10149 7157 10183 7191
rect 10183 7157 10192 7191
rect 10140 7148 10192 7157
rect 10784 7148 10836 7200
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 14004 7148 14056 7200
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 16488 7148 16540 7200
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 17776 7148 17828 7157
rect 17960 7148 18012 7200
rect 19432 7191 19484 7200
rect 19432 7157 19441 7191
rect 19441 7157 19475 7191
rect 19475 7157 19484 7191
rect 19432 7148 19484 7157
rect 22468 7191 22520 7200
rect 22468 7157 22477 7191
rect 22477 7157 22511 7191
rect 22511 7157 22520 7191
rect 22468 7148 22520 7157
rect 24768 7148 24820 7200
rect 25228 7148 25280 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 2688 6876 2740 6928
rect 4528 6944 4580 6996
rect 4804 6944 4856 6996
rect 5540 6944 5592 6996
rect 6184 6944 6236 6996
rect 7288 6944 7340 6996
rect 7932 6944 7984 6996
rect 9220 6944 9272 6996
rect 11152 6944 11204 6996
rect 12624 6987 12676 6996
rect 12624 6953 12633 6987
rect 12633 6953 12667 6987
rect 12667 6953 12676 6987
rect 12624 6944 12676 6953
rect 12900 6944 12952 6996
rect 14004 6944 14056 6996
rect 15936 6944 15988 6996
rect 20444 6944 20496 6996
rect 20720 6987 20772 6996
rect 20720 6953 20729 6987
rect 20729 6953 20763 6987
rect 20763 6953 20772 6987
rect 20720 6944 20772 6953
rect 4068 6876 4120 6928
rect 9036 6876 9088 6928
rect 9956 6876 10008 6928
rect 13636 6876 13688 6928
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 6184 6851 6236 6860
rect 4712 6808 4764 6817
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 10048 6808 10100 6860
rect 10876 6851 10928 6860
rect 10876 6817 10899 6851
rect 10899 6817 10928 6851
rect 10876 6808 10928 6817
rect 13084 6808 13136 6860
rect 14280 6808 14332 6860
rect 14556 6808 14608 6860
rect 14832 6851 14884 6860
rect 14832 6817 14841 6851
rect 14841 6817 14875 6851
rect 14875 6817 14884 6851
rect 14832 6808 14884 6817
rect 15752 6808 15804 6860
rect 16580 6876 16632 6928
rect 20168 6876 20220 6928
rect 16396 6851 16448 6860
rect 16396 6817 16430 6851
rect 16430 6817 16448 6851
rect 16396 6808 16448 6817
rect 17868 6808 17920 6860
rect 18788 6851 18840 6860
rect 18788 6817 18797 6851
rect 18797 6817 18831 6851
rect 18831 6817 18840 6851
rect 18788 6808 18840 6817
rect 19248 6808 19300 6860
rect 21456 6944 21508 6996
rect 22376 6944 22428 6996
rect 23756 6944 23808 6996
rect 25596 6944 25648 6996
rect 22652 6876 22704 6928
rect 20904 6851 20956 6860
rect 1952 6740 2004 6792
rect 2780 6740 2832 6792
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6644 6740 6696 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8208 6740 8260 6792
rect 9772 6740 9824 6792
rect 13176 6740 13228 6792
rect 5356 6715 5408 6724
rect 5356 6681 5365 6715
rect 5365 6681 5399 6715
rect 5399 6681 5408 6715
rect 5356 6672 5408 6681
rect 2044 6604 2096 6656
rect 2688 6604 2740 6656
rect 2964 6604 3016 6656
rect 3792 6604 3844 6656
rect 5448 6604 5500 6656
rect 6644 6604 6696 6656
rect 6828 6604 6880 6656
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 10784 6604 10836 6656
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 16120 6783 16172 6792
rect 13636 6740 13688 6749
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 19156 6740 19208 6792
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 20996 6808 21048 6860
rect 23480 6808 23532 6860
rect 23664 6851 23716 6860
rect 23664 6817 23698 6851
rect 23698 6817 23716 6851
rect 23664 6808 23716 6817
rect 24216 6808 24268 6860
rect 13176 6604 13228 6656
rect 13912 6604 13964 6656
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 20720 6672 20772 6724
rect 17776 6604 17828 6656
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 18512 6604 18564 6656
rect 18604 6647 18656 6656
rect 18604 6613 18613 6647
rect 18613 6613 18647 6647
rect 18647 6613 18656 6647
rect 18604 6604 18656 6613
rect 19340 6604 19392 6656
rect 22284 6647 22336 6656
rect 22284 6613 22293 6647
rect 22293 6613 22327 6647
rect 22327 6613 22336 6647
rect 22284 6604 22336 6613
rect 23664 6604 23716 6656
rect 25688 6876 25740 6928
rect 24952 6604 25004 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1952 6443 2004 6452
rect 1952 6409 1961 6443
rect 1961 6409 1995 6443
rect 1995 6409 2004 6443
rect 1952 6400 2004 6409
rect 2044 6400 2096 6452
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 4528 6400 4580 6452
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 5080 6443 5132 6452
rect 5080 6409 5089 6443
rect 5089 6409 5123 6443
rect 5123 6409 5132 6443
rect 5080 6400 5132 6409
rect 7932 6443 7984 6452
rect 7932 6409 7941 6443
rect 7941 6409 7975 6443
rect 7975 6409 7984 6443
rect 7932 6400 7984 6409
rect 9220 6400 9272 6452
rect 4252 6332 4304 6384
rect 4620 6332 4672 6384
rect 6552 6332 6604 6384
rect 7840 6332 7892 6384
rect 1492 6264 1544 6316
rect 2320 6264 2372 6316
rect 5356 6264 5408 6316
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 7012 6264 7064 6316
rect 8484 6264 8536 6316
rect 12164 6400 12216 6452
rect 12992 6400 13044 6452
rect 14280 6400 14332 6452
rect 11336 6332 11388 6384
rect 4252 6196 4304 6248
rect 1308 6128 1360 6180
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 2412 6128 2464 6180
rect 8852 6171 8904 6180
rect 8852 6137 8861 6171
rect 8861 6137 8895 6171
rect 8895 6137 8904 6171
rect 8852 6128 8904 6137
rect 9772 6196 9824 6248
rect 12624 6264 12676 6316
rect 13636 6264 13688 6316
rect 19248 6400 19300 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 22008 6400 22060 6452
rect 22100 6400 22152 6452
rect 23480 6400 23532 6452
rect 25596 6400 25648 6452
rect 25964 6400 26016 6452
rect 18696 6332 18748 6384
rect 20812 6332 20864 6384
rect 22652 6332 22704 6384
rect 24124 6332 24176 6384
rect 24308 6332 24360 6384
rect 24492 6332 24544 6384
rect 25044 6332 25096 6384
rect 20076 6264 20128 6316
rect 21824 6264 21876 6316
rect 11336 6196 11388 6248
rect 11796 6196 11848 6248
rect 13820 6196 13872 6248
rect 15200 6196 15252 6248
rect 16120 6196 16172 6248
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 18512 6196 18564 6248
rect 21732 6196 21784 6248
rect 22100 6196 22152 6248
rect 12900 6128 12952 6180
rect 14004 6128 14056 6180
rect 16856 6171 16908 6180
rect 16856 6137 16865 6171
rect 16865 6137 16899 6171
rect 16899 6137 16908 6171
rect 16856 6128 16908 6137
rect 19524 6171 19576 6180
rect 19524 6137 19533 6171
rect 19533 6137 19567 6171
rect 19567 6137 19576 6171
rect 19524 6128 19576 6137
rect 23664 6264 23716 6316
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 24216 6264 24268 6273
rect 25412 6307 25464 6316
rect 25412 6273 25421 6307
rect 25421 6273 25455 6307
rect 25455 6273 25464 6307
rect 25412 6264 25464 6273
rect 24124 6239 24176 6248
rect 24124 6205 24133 6239
rect 24133 6205 24167 6239
rect 24167 6205 24176 6239
rect 24124 6196 24176 6205
rect 24860 6196 24912 6248
rect 23940 6128 23992 6180
rect 2596 6060 2648 6112
rect 3608 6060 3660 6112
rect 6000 6060 6052 6112
rect 6920 6103 6972 6112
rect 6920 6069 6929 6103
rect 6929 6069 6963 6103
rect 6963 6069 6972 6103
rect 6920 6060 6972 6069
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 8208 6060 8260 6112
rect 8576 6060 8628 6112
rect 9404 6103 9456 6112
rect 9404 6069 9413 6103
rect 9413 6069 9447 6103
rect 9447 6069 9456 6103
rect 9404 6060 9456 6069
rect 10876 6060 10928 6112
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 13084 6060 13136 6112
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 19340 6060 19392 6112
rect 20076 6103 20128 6112
rect 20076 6069 20085 6103
rect 20085 6069 20119 6103
rect 20119 6069 20128 6103
rect 20076 6060 20128 6069
rect 20720 6060 20772 6112
rect 22008 6060 22060 6112
rect 22376 6060 22428 6112
rect 25044 6103 25096 6112
rect 25044 6069 25053 6103
rect 25053 6069 25087 6103
rect 25087 6069 25096 6103
rect 25044 6060 25096 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1768 5856 1820 5908
rect 2136 5856 2188 5908
rect 4804 5856 4856 5908
rect 5540 5856 5592 5908
rect 6184 5856 6236 5908
rect 6828 5856 6880 5908
rect 7288 5856 7340 5908
rect 9404 5856 9456 5908
rect 13176 5899 13228 5908
rect 13176 5865 13185 5899
rect 13185 5865 13219 5899
rect 13219 5865 13228 5899
rect 13176 5856 13228 5865
rect 13636 5856 13688 5908
rect 16120 5856 16172 5908
rect 16396 5856 16448 5908
rect 17868 5899 17920 5908
rect 17868 5865 17877 5899
rect 17877 5865 17911 5899
rect 17911 5865 17920 5899
rect 17868 5856 17920 5865
rect 19340 5856 19392 5908
rect 19524 5856 19576 5908
rect 21824 5856 21876 5908
rect 22376 5899 22428 5908
rect 22376 5865 22385 5899
rect 22385 5865 22419 5899
rect 22419 5865 22428 5899
rect 22376 5856 22428 5865
rect 23940 5899 23992 5908
rect 23940 5865 23949 5899
rect 23949 5865 23983 5899
rect 23983 5865 23992 5899
rect 23940 5856 23992 5865
rect 24676 5856 24728 5908
rect 25044 5856 25096 5908
rect 3792 5788 3844 5840
rect 4344 5788 4396 5840
rect 6276 5831 6328 5840
rect 6276 5797 6285 5831
rect 6285 5797 6319 5831
rect 6319 5797 6328 5831
rect 6276 5788 6328 5797
rect 1492 5763 1544 5772
rect 1492 5729 1501 5763
rect 1501 5729 1535 5763
rect 1535 5729 1544 5763
rect 1492 5720 1544 5729
rect 1768 5763 1820 5772
rect 1768 5729 1802 5763
rect 1802 5729 1820 5763
rect 1768 5720 1820 5729
rect 8944 5788 8996 5840
rect 10784 5788 10836 5840
rect 15752 5788 15804 5840
rect 17224 5788 17276 5840
rect 19064 5788 19116 5840
rect 20720 5788 20772 5840
rect 22744 5831 22796 5840
rect 8208 5720 8260 5772
rect 9680 5720 9732 5772
rect 10140 5720 10192 5772
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 12072 5763 12124 5772
rect 12072 5729 12081 5763
rect 12081 5729 12115 5763
rect 12115 5729 12124 5763
rect 12072 5720 12124 5729
rect 13452 5720 13504 5772
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 14280 5720 14332 5772
rect 15476 5720 15528 5772
rect 18236 5720 18288 5772
rect 20812 5720 20864 5772
rect 4252 5652 4304 5704
rect 7104 5695 7156 5704
rect 2412 5516 2464 5568
rect 2596 5516 2648 5568
rect 3608 5516 3660 5568
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 10416 5652 10468 5704
rect 11152 5652 11204 5704
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 15200 5652 15252 5704
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 21364 5695 21416 5704
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 22744 5797 22753 5831
rect 22753 5797 22787 5831
rect 22787 5797 22796 5831
rect 22744 5788 22796 5797
rect 24216 5788 24268 5840
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 24032 5720 24084 5772
rect 24676 5720 24728 5772
rect 23664 5652 23716 5704
rect 24860 5652 24912 5704
rect 5264 5516 5316 5568
rect 7012 5584 7064 5636
rect 8484 5627 8536 5636
rect 8484 5593 8493 5627
rect 8493 5593 8527 5627
rect 8527 5593 8536 5627
rect 8484 5584 8536 5593
rect 12716 5584 12768 5636
rect 13360 5584 13412 5636
rect 8576 5516 8628 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 12256 5559 12308 5568
rect 12256 5525 12265 5559
rect 12265 5525 12299 5559
rect 12299 5525 12308 5559
rect 12256 5516 12308 5525
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 14280 5559 14332 5568
rect 14280 5525 14289 5559
rect 14289 5525 14323 5559
rect 14323 5525 14332 5559
rect 14280 5516 14332 5525
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 15384 5516 15436 5568
rect 19340 5516 19392 5568
rect 20720 5516 20772 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1952 5312 2004 5364
rect 2504 5312 2556 5364
rect 3148 5312 3200 5364
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 6460 5312 6512 5364
rect 7288 5312 7340 5364
rect 9680 5312 9732 5364
rect 10416 5355 10468 5364
rect 10416 5321 10425 5355
rect 10425 5321 10459 5355
rect 10459 5321 10468 5355
rect 10416 5312 10468 5321
rect 10968 5312 11020 5364
rect 12072 5312 12124 5364
rect 13728 5312 13780 5364
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 22652 5312 22704 5364
rect 2964 5287 3016 5296
rect 2964 5253 2973 5287
rect 2973 5253 3007 5287
rect 3007 5253 3016 5287
rect 2964 5244 3016 5253
rect 1768 5176 1820 5228
rect 2412 5176 2464 5228
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 4712 5176 4764 5228
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 10876 5244 10928 5296
rect 8208 5176 8260 5228
rect 10692 5176 10744 5228
rect 14280 5176 14332 5228
rect 2136 5108 2188 5160
rect 3516 5151 3568 5160
rect 2044 4972 2096 5024
rect 2228 4972 2280 5024
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 5448 5108 5500 5160
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 10048 5108 10100 5160
rect 10784 5108 10836 5160
rect 14372 5151 14424 5160
rect 2780 5040 2832 5092
rect 2964 4972 3016 5024
rect 8024 5040 8076 5092
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 16120 5176 16172 5228
rect 18236 5176 18288 5228
rect 18880 5151 18932 5160
rect 18880 5117 18889 5151
rect 18889 5117 18923 5151
rect 18923 5117 18932 5151
rect 18880 5108 18932 5117
rect 24676 5312 24728 5364
rect 25964 5355 26016 5364
rect 25964 5321 25973 5355
rect 25973 5321 26007 5355
rect 26007 5321 26016 5355
rect 25964 5312 26016 5321
rect 24860 5244 24912 5296
rect 23480 5176 23532 5228
rect 23664 5219 23716 5228
rect 23664 5185 23673 5219
rect 23673 5185 23707 5219
rect 23707 5185 23716 5219
rect 23664 5176 23716 5185
rect 12900 5083 12952 5092
rect 12900 5049 12909 5083
rect 12909 5049 12943 5083
rect 12943 5049 12952 5083
rect 12900 5040 12952 5049
rect 13820 5083 13872 5092
rect 13820 5049 13829 5083
rect 13829 5049 13863 5083
rect 13863 5049 13872 5083
rect 13820 5040 13872 5049
rect 14648 5040 14700 5092
rect 19248 5040 19300 5092
rect 21732 5083 21784 5092
rect 21732 5049 21741 5083
rect 21741 5049 21775 5083
rect 21775 5049 21784 5083
rect 21732 5040 21784 5049
rect 24952 5108 25004 5160
rect 22284 5040 22336 5092
rect 23756 5040 23808 5092
rect 24216 5040 24268 5092
rect 25228 5040 25280 5092
rect 4068 4972 4120 5024
rect 5356 4972 5408 5024
rect 6000 4972 6052 5024
rect 8116 4972 8168 5024
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 12624 4972 12676 5024
rect 13452 5015 13504 5024
rect 13452 4981 13461 5015
rect 13461 4981 13495 5015
rect 13495 4981 13504 5015
rect 13452 4972 13504 4981
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 19340 4972 19392 5024
rect 20076 4972 20128 5024
rect 22192 4972 22244 5024
rect 22928 4972 22980 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1584 4768 1636 4820
rect 1768 4811 1820 4820
rect 1768 4777 1777 4811
rect 1777 4777 1811 4811
rect 1811 4777 1820 4811
rect 1768 4768 1820 4777
rect 1952 4768 2004 4820
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 5724 4768 5776 4820
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 9128 4811 9180 4820
rect 9128 4777 9137 4811
rect 9137 4777 9171 4811
rect 9171 4777 9180 4811
rect 9128 4768 9180 4777
rect 9312 4768 9364 4820
rect 11336 4768 11388 4820
rect 11704 4811 11756 4820
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 3516 4700 3568 4752
rect 5540 4700 5592 4752
rect 8852 4700 8904 4752
rect 9680 4700 9732 4752
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 5264 4632 5316 4684
rect 9404 4632 9456 4684
rect 10048 4675 10100 4684
rect 10048 4641 10082 4675
rect 10082 4641 10100 4675
rect 10048 4632 10100 4641
rect 12808 4700 12860 4752
rect 13084 4768 13136 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14372 4768 14424 4820
rect 15292 4768 15344 4820
rect 15568 4768 15620 4820
rect 17684 4768 17736 4820
rect 18236 4811 18288 4820
rect 18236 4777 18245 4811
rect 18245 4777 18279 4811
rect 18279 4777 18288 4811
rect 18236 4768 18288 4777
rect 18420 4768 18472 4820
rect 18880 4768 18932 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 23112 4768 23164 4820
rect 23756 4700 23808 4752
rect 13912 4632 13964 4684
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 16488 4675 16540 4684
rect 16488 4641 16522 4675
rect 16522 4641 16540 4675
rect 16488 4632 16540 4641
rect 19248 4675 19300 4684
rect 19248 4641 19257 4675
rect 19257 4641 19291 4675
rect 19291 4641 19300 4675
rect 19248 4632 19300 4641
rect 23388 4632 23440 4684
rect 24124 4768 24176 4820
rect 24768 4768 24820 4820
rect 25044 4811 25096 4820
rect 25044 4777 25053 4811
rect 25053 4777 25087 4811
rect 25087 4777 25096 4811
rect 25044 4768 25096 4777
rect 2044 4564 2096 4616
rect 8024 4564 8076 4616
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 9312 4564 9364 4616
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 2596 4496 2648 4548
rect 4896 4539 4948 4548
rect 2780 4428 2832 4480
rect 4896 4505 4905 4539
rect 4905 4505 4939 4539
rect 4939 4505 4948 4539
rect 4896 4496 4948 4505
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 8300 4428 8352 4480
rect 9680 4428 9732 4480
rect 19156 4564 19208 4616
rect 20720 4564 20772 4616
rect 21456 4607 21508 4616
rect 21456 4573 21465 4607
rect 21465 4573 21499 4607
rect 21499 4573 21508 4607
rect 23020 4607 23072 4616
rect 21456 4564 21508 4573
rect 23020 4573 23029 4607
rect 23029 4573 23063 4607
rect 23063 4573 23072 4607
rect 23020 4564 23072 4573
rect 24860 4564 24912 4616
rect 14096 4496 14148 4548
rect 20812 4496 20864 4548
rect 10508 4428 10560 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 14280 4471 14332 4480
rect 14280 4437 14289 4471
rect 14289 4437 14323 4471
rect 14323 4437 14332 4471
rect 14280 4428 14332 4437
rect 14740 4428 14792 4480
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 19064 4428 19116 4480
rect 19892 4471 19944 4480
rect 19892 4437 19901 4471
rect 19901 4437 19935 4471
rect 19935 4437 19944 4471
rect 19892 4428 19944 4437
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 20720 4428 20772 4480
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2320 4224 2372 4276
rect 4252 4224 4304 4276
rect 6460 4224 6512 4276
rect 9404 4267 9456 4276
rect 9404 4233 9413 4267
rect 9413 4233 9447 4267
rect 9447 4233 9456 4267
rect 9404 4224 9456 4233
rect 10784 4267 10836 4276
rect 10784 4233 10793 4267
rect 10793 4233 10827 4267
rect 10827 4233 10836 4267
rect 10784 4224 10836 4233
rect 15292 4224 15344 4276
rect 15844 4224 15896 4276
rect 16488 4267 16540 4276
rect 16488 4233 16497 4267
rect 16497 4233 16531 4267
rect 16531 4233 16540 4267
rect 16488 4224 16540 4233
rect 18880 4224 18932 4276
rect 21272 4224 21324 4276
rect 23020 4267 23072 4276
rect 23020 4233 23029 4267
rect 23029 4233 23063 4267
rect 23063 4233 23072 4267
rect 23020 4224 23072 4233
rect 24860 4224 24912 4276
rect 25964 4267 26016 4276
rect 25964 4233 25973 4267
rect 25973 4233 26007 4267
rect 26007 4233 26016 4267
rect 25964 4224 26016 4233
rect 1492 4088 1544 4140
rect 4896 4088 4948 4140
rect 5264 4088 5316 4140
rect 7932 4088 7984 4140
rect 8576 4156 8628 4208
rect 8392 4088 8444 4140
rect 9404 4088 9456 4140
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 12716 4131 12768 4140
rect 2504 4020 2556 4072
rect 5540 4020 5592 4072
rect 6828 4020 6880 4072
rect 9036 4020 9088 4072
rect 10140 4020 10192 4072
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 16764 4088 16816 4140
rect 3056 3952 3108 4004
rect 6552 3952 6604 4004
rect 10324 3952 10376 4004
rect 11428 3952 11480 4004
rect 11888 3952 11940 4004
rect 14188 4020 14240 4072
rect 15476 4020 15528 4072
rect 15568 4020 15620 4072
rect 15844 4063 15896 4072
rect 15844 4029 15853 4063
rect 15853 4029 15887 4063
rect 15887 4029 15896 4063
rect 15844 4020 15896 4029
rect 18236 4156 18288 4208
rect 20260 4156 20312 4208
rect 19892 4088 19944 4140
rect 20904 4088 20956 4140
rect 23664 4131 23716 4140
rect 23664 4097 23673 4131
rect 23673 4097 23707 4131
rect 23707 4097 23716 4131
rect 23664 4088 23716 4097
rect 21272 4063 21324 4072
rect 21272 4029 21306 4063
rect 21306 4029 21324 4063
rect 21272 4020 21324 4029
rect 21824 4020 21876 4072
rect 13820 3952 13872 4004
rect 19984 3952 20036 4004
rect 22284 3952 22336 4004
rect 3240 3884 3292 3936
rect 3976 3884 4028 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 6736 3884 6788 3936
rect 7104 3884 7156 3936
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 8668 3884 8720 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 10048 3884 10100 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 16212 3884 16264 3936
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 18512 3927 18564 3936
rect 18512 3893 18521 3927
rect 18521 3893 18555 3927
rect 18555 3893 18564 3927
rect 18512 3884 18564 3893
rect 19340 3884 19392 3936
rect 20260 3884 20312 3936
rect 20628 3884 20680 3936
rect 21916 3884 21968 3936
rect 24952 3884 25004 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1768 3680 1820 3732
rect 2044 3680 2096 3732
rect 4068 3723 4120 3732
rect 4068 3689 4077 3723
rect 4077 3689 4111 3723
rect 4111 3689 4120 3723
rect 4068 3680 4120 3689
rect 4160 3680 4212 3732
rect 5540 3680 5592 3732
rect 1584 3612 1636 3664
rect 3332 3612 3384 3664
rect 3700 3612 3752 3664
rect 6000 3680 6052 3732
rect 6368 3680 6420 3732
rect 7196 3680 7248 3732
rect 8300 3680 8352 3732
rect 9496 3680 9548 3732
rect 10048 3680 10100 3732
rect 11336 3680 11388 3732
rect 12532 3680 12584 3732
rect 15660 3723 15712 3732
rect 8392 3655 8444 3664
rect 1400 3544 1452 3596
rect 2228 3544 2280 3596
rect 3424 3544 3476 3596
rect 2320 3476 2372 3528
rect 4712 3519 4764 3528
rect 1308 3408 1360 3460
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 5540 3544 5592 3596
rect 6184 3544 6236 3596
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 8392 3621 8401 3655
rect 8401 3621 8435 3655
rect 8435 3621 8444 3655
rect 8392 3612 8444 3621
rect 9864 3612 9916 3664
rect 7104 3408 7156 3460
rect 1860 3340 1912 3392
rect 2320 3340 2372 3392
rect 3056 3340 3108 3392
rect 4160 3340 4212 3392
rect 5080 3340 5132 3392
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 7840 3587 7892 3596
rect 7840 3553 7849 3587
rect 7849 3553 7883 3587
rect 7883 3553 7892 3587
rect 7840 3544 7892 3553
rect 8944 3544 8996 3596
rect 9404 3544 9456 3596
rect 12808 3544 12860 3596
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 7932 3340 7984 3392
rect 8300 3340 8352 3392
rect 9312 3476 9364 3528
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 16856 3723 16908 3732
rect 16856 3689 16865 3723
rect 16865 3689 16899 3723
rect 16899 3689 16908 3723
rect 16856 3680 16908 3689
rect 17040 3680 17092 3732
rect 18052 3680 18104 3732
rect 18512 3680 18564 3732
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 20628 3680 20680 3732
rect 21272 3680 21324 3732
rect 23020 3723 23072 3732
rect 23020 3689 23029 3723
rect 23029 3689 23063 3723
rect 23063 3689 23072 3723
rect 23020 3680 23072 3689
rect 23480 3680 23532 3732
rect 24216 3680 24268 3732
rect 25044 3680 25096 3732
rect 25964 3680 26016 3732
rect 14188 3655 14240 3664
rect 14188 3621 14197 3655
rect 14197 3621 14231 3655
rect 14231 3621 14240 3655
rect 14188 3612 14240 3621
rect 17132 3612 17184 3664
rect 23940 3612 23992 3664
rect 24768 3612 24820 3664
rect 20996 3544 21048 3596
rect 21916 3587 21968 3596
rect 21916 3553 21950 3587
rect 21950 3553 21968 3587
rect 21916 3544 21968 3553
rect 22192 3544 22244 3596
rect 24952 3544 25004 3596
rect 13360 3476 13412 3528
rect 13636 3519 13688 3528
rect 13636 3485 13645 3519
rect 13645 3485 13679 3519
rect 13679 3485 13688 3519
rect 13636 3476 13688 3485
rect 15016 3519 15068 3528
rect 15016 3485 15025 3519
rect 15025 3485 15059 3519
rect 15059 3485 15068 3519
rect 15016 3476 15068 3485
rect 16212 3476 16264 3528
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 19340 3519 19392 3528
rect 17408 3476 17460 3485
rect 19340 3485 19349 3519
rect 19349 3485 19383 3519
rect 19383 3485 19392 3519
rect 19340 3476 19392 3485
rect 24676 3519 24728 3528
rect 15384 3408 15436 3460
rect 19156 3408 19208 3460
rect 21456 3451 21508 3460
rect 21456 3417 21465 3451
rect 21465 3417 21499 3451
rect 21499 3417 21508 3451
rect 21456 3408 21508 3417
rect 22652 3408 22704 3460
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 14004 3383 14056 3392
rect 14004 3349 14013 3383
rect 14013 3349 14047 3383
rect 14047 3349 14056 3383
rect 14004 3340 14056 3349
rect 16764 3383 16816 3392
rect 16764 3349 16773 3383
rect 16773 3349 16807 3383
rect 16807 3349 16816 3383
rect 16764 3340 16816 3349
rect 18512 3383 18564 3392
rect 18512 3349 18521 3383
rect 18521 3349 18555 3383
rect 18555 3349 18564 3383
rect 18512 3340 18564 3349
rect 18696 3383 18748 3392
rect 18696 3349 18705 3383
rect 18705 3349 18739 3383
rect 18739 3349 18748 3383
rect 18696 3340 18748 3349
rect 20168 3383 20220 3392
rect 20168 3349 20177 3383
rect 20177 3349 20211 3383
rect 20211 3349 20220 3383
rect 20168 3340 20220 3349
rect 23572 3383 23624 3392
rect 23572 3349 23581 3383
rect 23581 3349 23615 3383
rect 23615 3349 23624 3383
rect 23572 3340 23624 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2044 3136 2096 3188
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 6460 3136 6512 3188
rect 7840 3136 7892 3188
rect 8208 3136 8260 3188
rect 9680 3136 9732 3188
rect 12440 3136 12492 3188
rect 13360 3136 13412 3188
rect 16212 3179 16264 3188
rect 16212 3145 16221 3179
rect 16221 3145 16255 3179
rect 16255 3145 16264 3179
rect 16212 3136 16264 3145
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 17408 3136 17460 3188
rect 19340 3136 19392 3188
rect 20444 3136 20496 3188
rect 21916 3136 21968 3188
rect 22008 3136 22060 3188
rect 22284 3179 22336 3188
rect 22284 3145 22293 3179
rect 22293 3145 22327 3179
rect 22327 3145 22336 3179
rect 22284 3136 22336 3145
rect 23020 3179 23072 3188
rect 23020 3145 23029 3179
rect 23029 3145 23063 3179
rect 23063 3145 23072 3179
rect 23020 3136 23072 3145
rect 23664 3179 23716 3188
rect 23664 3145 23673 3179
rect 23673 3145 23707 3179
rect 23707 3145 23716 3179
rect 23664 3136 23716 3145
rect 25964 3136 26016 3188
rect 3700 3111 3752 3120
rect 3700 3077 3709 3111
rect 3709 3077 3743 3111
rect 3743 3077 3752 3111
rect 3700 3068 3752 3077
rect 16488 3068 16540 3120
rect 17040 3068 17092 3120
rect 22652 3068 22704 3120
rect 2596 3000 2648 3052
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 12716 3043 12768 3052
rect 2688 2932 2740 2984
rect 4712 2932 4764 2984
rect 6368 2932 6420 2984
rect 6644 2932 6696 2984
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 7196 2932 7248 2984
rect 8392 2932 8444 2984
rect 8576 2975 8628 2984
rect 8576 2941 8610 2975
rect 8610 2941 8628 2975
rect 8576 2932 8628 2941
rect 9404 2932 9456 2984
rect 2596 2864 2648 2916
rect 4804 2864 4856 2916
rect 6276 2864 6328 2916
rect 7288 2907 7340 2916
rect 7288 2873 7297 2907
rect 7297 2873 7331 2907
rect 7331 2873 7340 2907
rect 7288 2864 7340 2873
rect 3056 2796 3108 2848
rect 6460 2796 6512 2848
rect 7932 2796 7984 2848
rect 9864 2796 9916 2848
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 14648 3000 14700 3052
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 16672 3000 16724 3052
rect 17132 3000 17184 3052
rect 25136 3000 25188 3052
rect 11888 2975 11940 2984
rect 11888 2941 11897 2975
rect 11897 2941 11931 2975
rect 11931 2941 11940 2975
rect 11888 2932 11940 2941
rect 14096 2932 14148 2984
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 18328 2932 18380 2984
rect 18512 2975 18564 2984
rect 18512 2941 18546 2975
rect 18546 2941 18564 2975
rect 18512 2932 18564 2941
rect 20996 2932 21048 2984
rect 23664 2932 23716 2984
rect 25228 2975 25280 2984
rect 25228 2941 25237 2975
rect 25237 2941 25271 2975
rect 25271 2941 25280 2975
rect 25228 2932 25280 2941
rect 14648 2864 14700 2916
rect 20444 2864 20496 2916
rect 24216 2864 24268 2916
rect 26056 2864 26108 2916
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 11244 2839 11296 2848
rect 11244 2805 11253 2839
rect 11253 2805 11287 2839
rect 11287 2805 11296 2839
rect 11244 2796 11296 2805
rect 12992 2796 13044 2848
rect 13636 2796 13688 2848
rect 15200 2839 15252 2848
rect 15200 2805 15209 2839
rect 15209 2805 15243 2839
rect 15243 2805 15252 2839
rect 15200 2796 15252 2805
rect 23480 2839 23532 2848
rect 23480 2805 23489 2839
rect 23489 2805 23523 2839
rect 23523 2805 23532 2839
rect 23480 2796 23532 2805
rect 24952 2796 25004 2848
rect 25228 2796 25280 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1584 2592 1636 2644
rect 2228 2635 2280 2644
rect 2228 2601 2237 2635
rect 2237 2601 2271 2635
rect 2271 2601 2280 2635
rect 2228 2592 2280 2601
rect 2320 2592 2372 2644
rect 2964 2592 3016 2644
rect 6828 2592 6880 2644
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 9680 2592 9732 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 12532 2592 12584 2644
rect 20168 2592 20220 2644
rect 20628 2635 20680 2644
rect 20628 2601 20637 2635
rect 20637 2601 20671 2635
rect 20671 2601 20680 2635
rect 20628 2592 20680 2601
rect 21272 2635 21324 2644
rect 21272 2601 21281 2635
rect 21281 2601 21315 2635
rect 21315 2601 21324 2635
rect 21272 2592 21324 2601
rect 21640 2635 21692 2644
rect 21640 2601 21649 2635
rect 21649 2601 21683 2635
rect 21683 2601 21692 2635
rect 21640 2592 21692 2601
rect 21732 2592 21784 2644
rect 22652 2635 22704 2644
rect 22652 2601 22661 2635
rect 22661 2601 22695 2635
rect 22695 2601 22704 2635
rect 22652 2592 22704 2601
rect 23756 2592 23808 2644
rect 25688 2592 25740 2644
rect 1216 2524 1268 2576
rect 4344 2524 4396 2576
rect 6184 2524 6236 2576
rect 9496 2524 9548 2576
rect 12440 2567 12492 2576
rect 12440 2533 12449 2567
rect 12449 2533 12483 2567
rect 12483 2533 12492 2567
rect 12440 2524 12492 2533
rect 25872 2524 25924 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 6828 2456 6880 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 3516 2388 3568 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 5908 2363 5960 2372
rect 5908 2329 5917 2363
rect 5917 2329 5951 2363
rect 5951 2329 5960 2363
rect 5908 2320 5960 2329
rect 7748 2456 7800 2508
rect 9128 2456 9180 2508
rect 9956 2456 10008 2508
rect 11244 2456 11296 2508
rect 11704 2456 11756 2508
rect 12716 2456 12768 2508
rect 13176 2456 13228 2508
rect 17040 2499 17092 2508
rect 17040 2465 17049 2499
rect 17049 2465 17083 2499
rect 17083 2465 17092 2499
rect 17040 2456 17092 2465
rect 25596 2499 25648 2508
rect 9312 2388 9364 2440
rect 10048 2388 10100 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 9864 2320 9916 2372
rect 16672 2388 16724 2440
rect 20444 2388 20496 2440
rect 21732 2431 21784 2440
rect 21732 2397 21741 2431
rect 21741 2397 21775 2431
rect 21775 2397 21784 2431
rect 21732 2388 21784 2397
rect 25596 2465 25605 2499
rect 25605 2465 25639 2499
rect 25639 2465 25648 2499
rect 25596 2456 25648 2465
rect 22008 2388 22060 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 16120 2320 16172 2372
rect 22744 2320 22796 2372
rect 25964 2320 26016 2372
rect 3516 2252 3568 2304
rect 6184 2252 6236 2304
rect 6552 2252 6604 2304
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 14004 2295 14056 2304
rect 14004 2261 14013 2295
rect 14013 2261 14047 2295
rect 14047 2261 14056 2295
rect 14004 2252 14056 2261
rect 15476 2295 15528 2304
rect 15476 2261 15485 2295
rect 15485 2261 15519 2295
rect 15519 2261 15528 2295
rect 15476 2252 15528 2261
rect 17960 2295 18012 2304
rect 17960 2261 17969 2295
rect 17969 2261 18003 2295
rect 18003 2261 18012 2295
rect 17960 2252 18012 2261
rect 18604 2295 18656 2304
rect 18604 2261 18613 2295
rect 18613 2261 18647 2295
rect 18647 2261 18656 2295
rect 18604 2252 18656 2261
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 23664 2295 23716 2304
rect 23664 2261 23673 2295
rect 23673 2261 23707 2295
rect 23707 2261 23716 2295
rect 23664 2252 23716 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 13728 2048 13780 2100
rect 15384 2048 15436 2100
rect 15384 1912 15436 1964
rect 16304 1912 16356 1964
rect 24308 1368 24360 1420
rect 24768 1368 24820 1420
rect 4620 552 4672 604
rect 5264 552 5316 604
<< metal2 >>
rect 3514 27520 3570 28000
rect 4066 27704 4122 27713
rect 4066 27639 4122 27648
rect 2686 26616 2742 26625
rect 2686 26551 2742 26560
rect 1582 24984 1638 24993
rect 1582 24919 1638 24928
rect 1490 24440 1546 24449
rect 1490 24375 1546 24384
rect 1398 23896 1454 23905
rect 1398 23831 1454 23840
rect 1412 21962 1440 23831
rect 1504 23322 1532 24375
rect 1596 23866 1624 24919
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1492 23316 1544 23322
rect 1492 23258 1544 23264
rect 1582 23216 1638 23225
rect 1582 23151 1638 23160
rect 1490 22128 1546 22137
rect 1490 22063 1546 22072
rect 1400 21956 1452 21962
rect 1400 21898 1452 21904
rect 1504 21146 1532 22063
rect 1596 21690 1624 23151
rect 1872 22642 1900 23598
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 2228 22568 2280 22574
rect 2228 22510 2280 22516
rect 2240 21894 2268 22510
rect 2516 22438 2544 23122
rect 2504 22432 2556 22438
rect 2502 22400 2504 22409
rect 2556 22400 2558 22409
rect 2502 22335 2558 22344
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1582 21584 1638 21593
rect 1582 21519 1638 21528
rect 1492 21140 1544 21146
rect 1492 21082 1544 21088
rect 1596 20602 1624 21519
rect 2044 21344 2096 21350
rect 2042 21312 2044 21321
rect 2096 21312 2098 21321
rect 2042 21247 2098 21256
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1596 19961 1624 19994
rect 1582 19952 1638 19961
rect 1582 19887 1638 19896
rect 1952 19712 2004 19718
rect 1952 19654 2004 19660
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1596 19174 1624 19343
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1676 18828 1728 18834
rect 1676 18770 1728 18776
rect 1582 18728 1638 18737
rect 1582 18663 1638 18672
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1216 13320 1268 13326
rect 1216 13262 1268 13268
rect 1228 12442 1256 13262
rect 1320 12986 1348 13806
rect 1308 12980 1360 12986
rect 1308 12922 1360 12928
rect 1216 12436 1268 12442
rect 1216 12378 1268 12384
rect 1124 11824 1176 11830
rect 1124 11766 1176 11772
rect 1136 10538 1164 11766
rect 1320 11762 1348 12922
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1412 11354 1440 18158
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 15910 1532 17478
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 12170 1532 15302
rect 1596 15162 1624 18663
rect 1688 18154 1716 18770
rect 1964 18222 1992 19654
rect 2044 19168 2096 19174
rect 2042 19136 2044 19145
rect 2096 19136 2098 19145
rect 2042 19071 2098 19080
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1676 18148 1728 18154
rect 1676 18090 1728 18096
rect 1688 16946 1716 18090
rect 2136 18080 2188 18086
rect 2240 18057 2268 21830
rect 2424 21350 2452 22034
rect 2412 21344 2464 21350
rect 2412 21286 2464 21292
rect 2424 21185 2452 21286
rect 2410 21176 2466 21185
rect 2410 21111 2466 21120
rect 2594 21040 2650 21049
rect 2320 21004 2372 21010
rect 2594 20975 2650 20984
rect 2320 20946 2372 20952
rect 2332 20398 2360 20946
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 2136 18022 2188 18028
rect 2226 18048 2282 18057
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1780 17134 1808 17478
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1688 16918 1808 16946
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1492 12164 1544 12170
rect 1492 12106 1544 12112
rect 1490 12064 1546 12073
rect 1490 11999 1546 12008
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1124 10532 1176 10538
rect 1124 10474 1176 10480
rect 1412 9654 1440 11154
rect 1504 11121 1532 11999
rect 1596 11830 1624 14554
rect 1688 12306 1716 15982
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1688 11898 1716 12242
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1584 11824 1636 11830
rect 1584 11766 1636 11772
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1490 11112 1546 11121
rect 1490 11047 1546 11056
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1400 9648 1452 9654
rect 1400 9590 1452 9596
rect 1398 7984 1454 7993
rect 1398 7919 1400 7928
rect 1452 7919 1454 7928
rect 1400 7890 1452 7896
rect 1504 7426 1532 10950
rect 1596 10470 1624 11630
rect 1688 11014 1716 11698
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10674 1716 10950
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 9586 1624 10406
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1688 7528 1716 10474
rect 1780 7698 1808 16918
rect 1872 16114 1900 17682
rect 2148 17678 2176 18022
rect 2226 17983 2282 17992
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2148 17202 2176 17614
rect 2332 17241 2360 20334
rect 2412 20256 2464 20262
rect 2410 20224 2412 20233
rect 2464 20224 2466 20233
rect 2410 20159 2466 20168
rect 2412 19916 2464 19922
rect 2412 19858 2464 19864
rect 2424 19174 2452 19858
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2424 19009 2452 19110
rect 2410 19000 2466 19009
rect 2410 18935 2466 18944
rect 2516 18714 2544 19246
rect 2608 19174 2636 20975
rect 2700 20058 2728 26551
rect 3330 25528 3386 25537
rect 3330 25463 3386 25472
rect 3344 24886 3372 25463
rect 3332 24880 3384 24886
rect 3528 24857 3556 27520
rect 3790 27160 3846 27169
rect 3790 27095 3846 27104
rect 3332 24822 3384 24828
rect 3514 24848 3570 24857
rect 3514 24783 3570 24792
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2700 19310 2728 19858
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2516 18686 2636 18714
rect 2608 18630 2636 18686
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2608 18465 2636 18566
rect 2594 18456 2650 18465
rect 2594 18391 2650 18400
rect 2792 18290 2820 18770
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2504 17808 2556 17814
rect 2504 17750 2556 17756
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2318 17232 2374 17241
rect 2136 17196 2188 17202
rect 2318 17167 2374 17176
rect 2136 17138 2188 17144
rect 2148 17082 2176 17138
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 2056 17054 2176 17082
rect 1964 16794 1992 17002
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2056 16590 2084 17054
rect 2320 16992 2372 16998
rect 2226 16960 2282 16969
rect 2320 16934 2372 16940
rect 2226 16895 2282 16904
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1872 15706 1900 15846
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1964 15570 1992 16390
rect 2044 16176 2096 16182
rect 2044 16118 2096 16124
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1872 14890 1900 15506
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 1860 14884 1912 14890
rect 1860 14826 1912 14832
rect 1872 9178 1900 14826
rect 1964 14482 1992 15370
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 2056 14362 2084 16118
rect 2148 16046 2176 16730
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 1964 14334 2084 14362
rect 1964 12782 1992 14334
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 10266 1992 12582
rect 2056 11354 2084 14214
rect 2148 12442 2176 15846
rect 2240 14498 2268 16895
rect 2332 16794 2360 16934
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 2332 16250 2360 16594
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2332 15502 2360 16050
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2332 14657 2360 14962
rect 2318 14648 2374 14657
rect 2424 14618 2452 17478
rect 2516 16998 2544 17750
rect 2884 17746 2912 18702
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2792 17338 2820 17682
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2884 17202 2912 17478
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2516 15910 2544 16934
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2608 15162 2636 16458
rect 2700 15638 2728 16526
rect 2884 16114 2912 17138
rect 2976 17105 3004 18566
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 2962 17096 3018 17105
rect 2962 17031 3018 17040
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2700 15026 2728 15302
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2318 14583 2374 14592
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2240 14470 2544 14498
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 2240 13546 2268 13738
rect 2332 13716 2360 14282
rect 2424 14074 2452 14350
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2412 13728 2464 13734
rect 2332 13688 2412 13716
rect 2412 13670 2464 13676
rect 2240 13518 2360 13546
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2240 12918 2268 13330
rect 2228 12912 2280 12918
rect 2226 12880 2228 12889
rect 2280 12880 2282 12889
rect 2332 12850 2360 13518
rect 2226 12815 2282 12824
rect 2320 12844 2372 12850
rect 2240 12789 2268 12815
rect 2320 12786 2372 12792
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2332 12238 2360 12786
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2148 11642 2176 12106
rect 2424 12102 2452 13670
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2424 11778 2452 11834
rect 2332 11750 2452 11778
rect 2148 11614 2268 11642
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2148 11150 2176 11494
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1964 9178 1992 9522
rect 2056 9330 2084 11018
rect 2148 10130 2176 11086
rect 2240 10169 2268 11614
rect 2226 10160 2282 10169
rect 2136 10124 2188 10130
rect 2226 10095 2282 10104
rect 2136 10066 2188 10072
rect 2240 9450 2268 10095
rect 2332 9518 2360 11750
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 11082 2452 11562
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2410 10024 2466 10033
rect 2410 9959 2412 9968
rect 2464 9959 2466 9968
rect 2412 9930 2464 9936
rect 2410 9752 2466 9761
rect 2410 9687 2466 9696
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2056 9302 2268 9330
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2148 8430 2176 8978
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2148 8090 2176 8366
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 1780 7670 1900 7698
rect 1688 7500 1808 7528
rect 1504 7398 1716 7426
rect 1582 7304 1638 7313
rect 1582 7239 1638 7248
rect 1596 7206 1624 7239
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1398 6896 1454 6905
rect 1398 6831 1400 6840
rect 1452 6831 1454 6840
rect 1400 6802 1452 6808
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1308 6180 1360 6186
rect 1308 6122 1360 6128
rect 1320 3466 1348 6122
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 3602 1440 6054
rect 1504 5778 1532 6258
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 1504 4146 1532 5714
rect 1596 4826 1624 7142
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1688 4298 1716 7398
rect 1780 5914 1808 7500
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1766 5808 1822 5817
rect 1766 5743 1768 5752
rect 1820 5743 1822 5752
rect 1768 5714 1820 5720
rect 1780 5234 1808 5714
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1766 4856 1822 4865
rect 1766 4791 1768 4800
rect 1820 4791 1822 4800
rect 1768 4762 1820 4768
rect 1596 4270 1716 4298
rect 1596 4185 1624 4270
rect 1582 4176 1638 4185
rect 1492 4140 1544 4146
rect 1582 4111 1638 4120
rect 1492 4082 1544 4088
rect 1596 3670 1624 4111
rect 1780 3738 1808 4762
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1584 3664 1636 3670
rect 1636 3612 1716 3618
rect 1584 3606 1716 3612
rect 1400 3596 1452 3602
rect 1596 3590 1716 3606
rect 1400 3538 1452 3544
rect 1582 3496 1638 3505
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 1504 3454 1582 3482
rect 846 3360 902 3369
rect 846 3295 902 3304
rect 570 1592 626 1601
rect 308 1550 570 1578
rect 308 480 336 1550
rect 570 1527 626 1536
rect 860 480 888 3295
rect 1216 2576 1268 2582
rect 1214 2544 1216 2553
rect 1268 2544 1270 2553
rect 1214 2479 1270 2488
rect 1320 921 1348 3402
rect 1398 2544 1454 2553
rect 1398 2479 1400 2488
rect 1452 2479 1454 2488
rect 1400 2450 1452 2456
rect 1504 1442 1532 3454
rect 1582 3431 1638 3440
rect 1688 3380 1716 3590
rect 1872 3398 1900 7670
rect 2042 7440 2098 7449
rect 2042 7375 2044 7384
rect 2096 7375 2098 7384
rect 2136 7404 2188 7410
rect 2044 7346 2096 7352
rect 2136 7346 2188 7352
rect 1952 6792 2004 6798
rect 2148 6780 2176 7346
rect 1952 6734 2004 6740
rect 2056 6752 2176 6780
rect 1964 6458 1992 6734
rect 2056 6662 2084 6752
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 6458 2084 6598
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1964 4826 1992 5306
rect 2148 5166 2176 5850
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2056 4706 2084 4966
rect 1964 4678 2084 4706
rect 1596 3352 1716 3380
rect 1860 3392 1912 3398
rect 1596 2650 1624 3352
rect 1860 3334 1912 3340
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1964 2009 1992 4678
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2056 3738 2084 4558
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2042 3632 2098 3641
rect 2042 3567 2098 3576
rect 2056 3194 2084 3567
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2148 3097 2176 5102
rect 2240 5030 2268 9302
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2332 6322 2360 8298
rect 2424 8090 2452 9687
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2516 7546 2544 14470
rect 2608 13530 2636 14758
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 13870 2728 14350
rect 2792 14278 2820 15506
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 14958 2912 15302
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2976 14804 3004 16934
rect 3160 16794 3188 17002
rect 3344 16998 3372 17478
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 2884 14776 3004 14804
rect 2884 14618 2912 14776
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2780 14068 2832 14074
rect 3056 14068 3108 14074
rect 2832 14028 2912 14056
rect 2780 14010 2832 14016
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2594 12336 2650 12345
rect 2594 12271 2596 12280
rect 2648 12271 2650 12280
rect 2596 12242 2648 12248
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11694 2636 12038
rect 2700 11898 2728 12718
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2792 11098 2820 12951
rect 2884 11506 2912 14028
rect 3056 14010 3108 14016
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 11626 3004 12582
rect 3068 11812 3096 14010
rect 3160 13025 3188 16730
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3252 16046 3280 16390
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3252 14958 3280 15982
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3238 14376 3294 14385
rect 3238 14311 3294 14320
rect 3252 13433 3280 14311
rect 3238 13424 3294 13433
rect 3238 13359 3294 13368
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3146 13016 3202 13025
rect 3146 12951 3202 12960
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 3160 11880 3188 12854
rect 3252 12238 3280 13126
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3160 11852 3280 11880
rect 3068 11784 3188 11812
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2884 11478 3004 11506
rect 2870 11384 2926 11393
rect 2870 11319 2926 11328
rect 2884 11286 2912 11319
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2608 11070 2820 11098
rect 2608 9178 2636 11070
rect 2884 10996 2912 11222
rect 2976 11014 3004 11478
rect 2792 10968 2912 10996
rect 2964 11008 3016 11014
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2792 9110 2820 10968
rect 2964 10950 3016 10956
rect 2976 10606 3004 10950
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2870 10296 2926 10305
rect 2870 10231 2872 10240
rect 2924 10231 2926 10240
rect 2872 10202 2924 10208
rect 2884 9722 2912 10202
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2608 7290 2636 8842
rect 2792 8106 2820 9046
rect 2872 8968 2924 8974
rect 2976 8945 3004 10542
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 8974 3096 9998
rect 3160 9353 3188 11784
rect 3252 10266 3280 11852
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3252 9382 3280 10202
rect 3344 9761 3372 16934
rect 3712 16454 3740 17478
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3436 12986 3464 16186
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3528 15366 3556 15914
rect 3700 15632 3752 15638
rect 3698 15600 3700 15609
rect 3752 15600 3754 15609
rect 3698 15535 3754 15544
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 13734 3556 15302
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3528 13462 3556 13670
rect 3516 13456 3568 13462
rect 3516 13398 3568 13404
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3528 12442 3556 13398
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3436 9518 3464 12310
rect 3514 10432 3570 10441
rect 3514 10367 3570 10376
rect 3528 9994 3556 10367
rect 3620 10198 3648 15370
rect 3712 15162 3740 15535
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14550 3740 14894
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3700 13796 3752 13802
rect 3700 13738 3752 13744
rect 3712 13190 3740 13738
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3712 12481 3740 13126
rect 3698 12472 3754 12481
rect 3698 12407 3754 12416
rect 3804 12345 3832 27095
rect 4080 26314 4108 27639
rect 10506 27520 10562 28000
rect 17498 27520 17554 28000
rect 24122 27704 24178 27713
rect 24122 27639 24178 27648
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4066 26072 4122 26081
rect 4122 26030 4200 26058
rect 4066 26007 4122 26016
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4080 18290 4108 18770
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3988 17338 4016 17682
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 4080 16572 4108 18022
rect 4172 17882 4200 26030
rect 10520 25786 10548 27520
rect 10520 25758 10824 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 7012 24880 7064 24886
rect 7012 24822 7064 24828
rect 9218 24848 9274 24857
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 4618 22672 4674 22681
rect 4618 22607 4674 22616
rect 4526 21176 4582 21185
rect 4632 21146 4660 22607
rect 4894 22400 4950 22409
rect 4894 22335 4950 22344
rect 4526 21111 4582 21120
rect 4620 21140 4672 21146
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4250 20496 4306 20505
rect 4448 20466 4476 20946
rect 4250 20431 4306 20440
rect 4436 20460 4488 20466
rect 4264 18970 4292 20431
rect 4436 20402 4488 20408
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4080 16544 4200 16572
rect 4264 16561 4292 17478
rect 4344 16992 4396 16998
rect 4342 16960 4344 16969
rect 4396 16960 4398 16969
rect 4342 16895 4398 16904
rect 3974 16008 4030 16017
rect 3974 15943 4030 15952
rect 3882 15736 3938 15745
rect 3882 15671 3938 15680
rect 3790 12336 3846 12345
rect 3790 12271 3846 12280
rect 3804 11393 3832 12271
rect 3790 11384 3846 11393
rect 3790 11319 3846 11328
rect 3698 11248 3754 11257
rect 3698 11183 3754 11192
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3528 9722 3556 9930
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3240 9376 3292 9382
rect 3146 9344 3202 9353
rect 3240 9318 3292 9324
rect 3146 9279 3202 9288
rect 3056 8968 3108 8974
rect 2872 8910 2924 8916
rect 2962 8936 3018 8945
rect 2884 8634 2912 8910
rect 3056 8910 3108 8916
rect 2962 8871 3018 8880
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3252 8412 3280 9318
rect 3330 8936 3386 8945
rect 3330 8871 3386 8880
rect 3344 8566 3372 8871
rect 3436 8838 3464 9454
rect 3606 9072 3662 9081
rect 3606 9007 3662 9016
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3252 8384 3372 8412
rect 2700 8078 2820 8106
rect 2700 7426 2728 8078
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2700 7398 2820 7426
rect 2516 7262 2636 7290
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2424 5574 2452 6122
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2516 5370 2544 7262
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2608 6882 2636 7142
rect 2688 6928 2740 6934
rect 2608 6876 2688 6882
rect 2608 6870 2740 6876
rect 2608 6854 2728 6870
rect 2608 6118 2636 6854
rect 2792 6798 2820 7398
rect 2884 7342 2912 7822
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2976 7206 3004 7890
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3146 7440 3202 7449
rect 3146 7375 3202 7384
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2870 7032 2926 7041
rect 2870 6967 2926 6976
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2688 6656 2740 6662
rect 2884 6644 2912 6967
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2688 6598 2740 6604
rect 2792 6616 2912 6644
rect 2964 6656 3016 6662
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2424 4826 2452 5170
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2424 4706 2452 4762
rect 2332 4678 2452 4706
rect 2332 4282 2360 4678
rect 2608 4554 2636 5510
rect 2700 5114 2728 6598
rect 2792 5545 2820 6616
rect 2964 6598 3016 6604
rect 2976 5794 3004 6598
rect 3068 6361 3096 6734
rect 3054 6352 3110 6361
rect 3054 6287 3110 6296
rect 3068 5817 3096 6287
rect 2884 5766 3004 5794
rect 3054 5808 3110 5817
rect 2778 5536 2834 5545
rect 2778 5471 2834 5480
rect 2700 5098 2820 5114
rect 2700 5092 2832 5098
rect 2700 5086 2780 5092
rect 2780 5034 2832 5040
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4298 2820 4422
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2700 4270 2820 4298
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2134 3088 2190 3097
rect 2134 3023 2190 3032
rect 2240 2650 2268 3538
rect 2332 3534 2360 4218
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2516 3754 2544 4014
rect 2516 3726 2636 3754
rect 2502 3632 2558 3641
rect 2502 3567 2558 3576
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 2650 2360 3334
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 1950 2000 2006 2009
rect 1950 1935 2006 1944
rect 1950 1864 2006 1873
rect 1950 1799 2006 1808
rect 1412 1414 1532 1442
rect 1306 912 1362 921
rect 1306 847 1362 856
rect 1412 480 1440 1414
rect 1964 480 1992 1799
rect 2516 480 2544 3567
rect 2608 3058 2636 3726
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 2922 2636 2994
rect 2700 2990 2728 4270
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2884 2825 2912 5766
rect 3054 5743 3110 5752
rect 3160 5370 3188 7375
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 2964 5296 3016 5302
rect 2962 5264 2964 5273
rect 3016 5264 3018 5273
rect 2962 5199 3018 5208
rect 2976 5030 3004 5199
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2962 3768 3018 3777
rect 2962 3703 3018 3712
rect 2870 2816 2926 2825
rect 2870 2751 2926 2760
rect 2976 2650 3004 3703
rect 3068 3398 3096 3946
rect 3252 3942 3280 7822
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3344 3670 3372 8384
rect 3436 4604 3464 8774
rect 3528 5953 3556 8774
rect 3620 8634 3648 9007
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3606 7848 3662 7857
rect 3606 7783 3662 7792
rect 3620 7546 3648 7783
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 6118 3648 7278
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3514 5944 3570 5953
rect 3514 5879 3570 5888
rect 3514 5672 3570 5681
rect 3514 5607 3570 5616
rect 3528 5166 3556 5607
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3620 5234 3648 5510
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3528 4758 3556 5102
rect 3516 4752 3568 4758
rect 3712 4729 3740 11183
rect 3896 9654 3924 15671
rect 3988 13705 4016 15943
rect 4066 15600 4122 15609
rect 4066 15535 4122 15544
rect 4080 14822 4108 15535
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4080 14618 4108 14758
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 4080 13734 4108 14282
rect 4068 13728 4120 13734
rect 3974 13696 4030 13705
rect 4068 13670 4120 13676
rect 3974 13631 4030 13640
rect 4066 13152 4122 13161
rect 4066 13087 4122 13096
rect 4080 12753 4108 13087
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4172 10810 4200 16544
rect 4250 16552 4306 16561
rect 4250 16487 4306 16496
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4356 15706 4384 15846
rect 4344 15700 4396 15706
rect 4396 15660 4476 15688
rect 4344 15642 4396 15648
rect 4344 15360 4396 15366
rect 4264 15320 4344 15348
rect 4264 12442 4292 15320
rect 4344 15302 4396 15308
rect 4344 14952 4396 14958
rect 4448 14940 4476 15660
rect 4396 14912 4476 14940
rect 4344 14894 4396 14900
rect 4540 14804 4568 21111
rect 4620 21082 4672 21088
rect 4802 18456 4858 18465
rect 4802 18391 4858 18400
rect 4618 17776 4674 17785
rect 4618 17711 4674 17720
rect 4448 14776 4568 14804
rect 4448 14770 4476 14776
rect 4356 14742 4476 14770
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4250 11792 4306 11801
rect 4250 11727 4306 11736
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4264 10282 4292 11727
rect 4172 10254 4292 10282
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3804 8634 3832 9046
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3882 8392 3938 8401
rect 3882 8327 3938 8336
rect 3896 7954 3924 8327
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3896 7410 3924 7890
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3804 6662 3832 7142
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3804 5846 3832 6394
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3516 4694 3568 4700
rect 3698 4720 3754 4729
rect 3698 4655 3754 4664
rect 3436 4576 3556 4604
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3068 2854 3096 3334
rect 3436 3194 3464 3538
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 1737 2820 2450
rect 3068 2446 3096 2790
rect 3528 2446 3556 4576
rect 3896 4049 3924 7210
rect 3882 4040 3938 4049
rect 3882 3975 3938 3984
rect 3988 3942 4016 9862
rect 4080 8838 4108 9998
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4066 8664 4122 8673
rect 4066 8599 4122 8608
rect 4080 6934 4108 8599
rect 4172 8362 4200 10254
rect 4252 10192 4304 10198
rect 4250 10160 4252 10169
rect 4304 10160 4306 10169
rect 4250 10095 4306 10104
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4172 8022 4200 8298
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4264 6390 4292 9658
rect 4356 8650 4384 14742
rect 4632 14634 4660 17711
rect 4448 14606 4660 14634
rect 4712 14612 4764 14618
rect 4448 11257 4476 14606
rect 4712 14554 4764 14560
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 13530 4568 14350
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4540 12442 4568 13466
rect 4632 13308 4660 14486
rect 4724 13530 4752 14554
rect 4816 14550 4844 18391
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 4816 14006 4844 14486
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4712 13320 4764 13326
rect 4632 13280 4712 13308
rect 4712 13262 4764 13268
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4632 12617 4660 13126
rect 4724 12782 4752 13262
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4618 12608 4674 12617
rect 4618 12543 4674 12552
rect 4724 12442 4752 12718
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4618 12336 4674 12345
rect 4618 12271 4674 12280
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4540 11354 4568 12174
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4434 11248 4490 11257
rect 4632 11234 4660 12271
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4434 11183 4490 11192
rect 4540 11206 4660 11234
rect 4540 9602 4568 11206
rect 4724 11132 4752 12106
rect 4816 11286 4844 13806
rect 4908 12170 4936 22335
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6458 20224 6514 20233
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5538 18184 5594 18193
rect 5538 18119 5594 18128
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5000 16998 5028 17682
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 13802 5028 16934
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 5078 16144 5134 16153
rect 5078 16079 5134 16088
rect 5092 15706 5120 16079
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5092 14958 5120 15506
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5080 14000 5132 14006
rect 5080 13942 5132 13948
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 5092 11762 5120 13942
rect 5184 12628 5212 16662
rect 5276 12782 5304 17070
rect 5552 16794 5580 18119
rect 5998 17640 6054 17649
rect 5998 17575 6054 17584
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5368 16250 5396 16594
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16250 6040 17575
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5538 15600 5594 15609
rect 5538 15535 5540 15544
rect 5592 15535 5594 15544
rect 5540 15506 5592 15512
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 15162 5488 15438
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5448 15156 5500 15162
rect 5368 15116 5448 15144
rect 5368 13462 5396 15116
rect 5448 15098 5500 15104
rect 5998 14920 6054 14929
rect 5998 14855 6054 14864
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5460 13870 5488 14758
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5630 13968 5686 13977
rect 5630 13903 5632 13912
rect 5684 13903 5686 13912
rect 5632 13874 5684 13880
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 6012 13802 6040 14855
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 5998 13696 6054 13705
rect 5998 13631 6054 13640
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5368 12986 5396 13398
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5184 12600 5304 12628
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5184 11558 5212 12038
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4724 11104 4844 11132
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4724 10742 4752 10950
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4632 9722 4660 10474
rect 4724 10130 4752 10678
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4540 9574 4660 9602
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4356 8622 4476 8650
rect 4344 8560 4396 8566
rect 4342 8528 4344 8537
rect 4396 8528 4398 8537
rect 4342 8463 4398 8472
rect 4448 7970 4476 8622
rect 4540 8090 4568 8910
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4448 7942 4568 7970
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7206 4476 7822
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 5710 4292 6190
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4356 5370 4384 5782
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4448 5250 4476 7142
rect 4540 7002 4568 7942
rect 4632 7018 4660 9574
rect 4710 8664 4766 8673
rect 4816 8650 4844 11104
rect 4908 10674 4936 11494
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9382 5120 9862
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4766 8622 4844 8650
rect 4710 8599 4766 8608
rect 4724 8430 4752 8599
rect 4908 8498 4936 8842
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 5000 7449 5028 8774
rect 4986 7440 5042 7449
rect 4986 7375 5042 7384
rect 4802 7168 4858 7177
rect 4802 7103 4858 7112
rect 4710 7032 4766 7041
rect 4528 6996 4580 7002
rect 4632 6990 4710 7018
rect 4816 7002 4844 7103
rect 4710 6967 4766 6976
rect 4804 6996 4856 7002
rect 4528 6938 4580 6944
rect 4540 6458 4568 6938
rect 4724 6866 4752 6967
rect 4804 6938 4856 6944
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4724 6458 4752 6802
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4356 5222 4476 5250
rect 4250 5128 4306 5137
rect 4250 5063 4306 5072
rect 4068 5024 4120 5030
rect 4120 4984 4200 5012
rect 4068 4966 4120 4972
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 4066 3904 4122 3913
rect 3988 3777 4016 3878
rect 4066 3839 4122 3848
rect 3974 3768 4030 3777
rect 4080 3738 4108 3839
rect 4172 3738 4200 4984
rect 4264 4690 4292 5063
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4264 4282 4292 4626
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 3974 3703 4030 3712
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3712 3126 3740 3606
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 3700 3120 3752 3126
rect 3606 3088 3662 3097
rect 3700 3062 3752 3068
rect 3606 3023 3662 3032
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3528 2310 3556 2382
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 2778 1728 2834 1737
rect 2778 1663 2834 1672
rect 3528 1465 3556 2246
rect 3514 1456 3570 1465
rect 3514 1391 3570 1400
rect 3054 1048 3110 1057
rect 3054 983 3110 992
rect 3068 480 3096 983
rect 3620 480 3648 3023
rect 4172 480 4200 3334
rect 4356 2582 4384 5222
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4448 105 4476 4422
rect 4632 610 4660 6326
rect 4816 5914 4844 6734
rect 5092 6458 5120 9318
rect 5184 7546 5212 11494
rect 5276 7954 5304 12600
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5368 11626 5396 12242
rect 5460 12238 5488 13466
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12986 6040 13631
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5538 12880 5594 12889
rect 5538 12815 5540 12824
rect 5592 12815 5594 12824
rect 5540 12786 5592 12792
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5552 11762 5580 11834
rect 5540 11756 5592 11762
rect 5592 11716 5672 11744
rect 5540 11698 5592 11704
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5644 11354 5672 11716
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5354 10976 5410 10985
rect 5354 10911 5410 10920
rect 5368 10577 5396 10911
rect 5354 10568 5410 10577
rect 5354 10503 5410 10512
rect 5460 10198 5488 11290
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5552 10810 5580 11222
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10192 5500 10198
rect 5354 10160 5410 10169
rect 5448 10134 5500 10140
rect 5354 10095 5410 10104
rect 5368 9897 5396 10095
rect 5354 9888 5410 9897
rect 5354 9823 5410 9832
rect 5460 9654 5488 10134
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 8838 5396 9386
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5368 7818 5396 8774
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5276 6497 5304 7414
rect 5460 7041 5488 8298
rect 5552 8090 5580 10746
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9110 6040 10406
rect 6104 9178 6132 20198
rect 6458 20159 6514 20168
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6288 15706 6316 16390
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6288 15434 6316 15642
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 13530 6224 14350
rect 6288 13938 6316 14418
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6196 11393 6224 11562
rect 6182 11384 6238 11393
rect 6182 11319 6238 11328
rect 6196 10146 6224 11319
rect 6288 11218 6316 12106
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6288 10266 6316 10542
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6196 10118 6316 10146
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5552 7886 5580 8026
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5552 7410 5580 7822
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6012 7546 6040 9046
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6104 8634 6132 8910
rect 6196 8634 6224 9318
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6288 8480 6316 10118
rect 6380 9160 6408 15846
rect 6472 13025 6500 20159
rect 6918 18048 6974 18057
rect 6918 17983 6974 17992
rect 6932 16794 6960 17983
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6642 15736 6698 15745
rect 6840 15706 6868 16594
rect 6642 15671 6644 15680
rect 6696 15671 6698 15680
rect 6828 15700 6880 15706
rect 6644 15642 6696 15648
rect 6828 15642 6880 15648
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6840 15162 6868 15506
rect 7024 15162 7052 24822
rect 9218 24783 9274 24792
rect 7378 21312 7434 21321
rect 7378 21247 7434 21256
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 7116 15502 7144 15914
rect 7208 15910 7236 16662
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6748 13870 6776 14418
rect 7012 14272 7064 14278
rect 7116 14260 7144 15438
rect 7064 14232 7144 14260
rect 7012 14214 7064 14220
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6458 13016 6514 13025
rect 6458 12951 6514 12960
rect 6472 11014 6500 12951
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6656 12481 6684 12582
rect 6642 12472 6698 12481
rect 6642 12407 6698 12416
rect 6748 12073 6776 13806
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13530 6960 13670
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 12232 6880 12238
rect 6826 12200 6828 12209
rect 6880 12200 6882 12209
rect 6826 12135 6882 12144
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 7024 11762 7052 14214
rect 7208 11898 7236 15846
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7300 12345 7328 13874
rect 7392 13852 7420 21247
rect 9232 19961 9260 24783
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10796 20913 10824 25758
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 17512 23497 17540 27520
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 22480 23662 22508 26250
rect 24136 24970 24164 27639
rect 24490 27520 24546 28000
rect 24504 25242 24532 27520
rect 25410 27160 25466 27169
rect 25410 27095 25466 27104
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24044 24942 24164 24970
rect 24228 25214 24532 25242
rect 23846 24304 23902 24313
rect 23846 24239 23902 24248
rect 22650 24168 22706 24177
rect 22650 24103 22706 24112
rect 22664 23866 22692 24103
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22742 23760 22798 23769
rect 22742 23695 22798 23704
rect 22468 23656 22520 23662
rect 20626 23624 20682 23633
rect 22468 23598 22520 23604
rect 20626 23559 20682 23568
rect 15290 23488 15346 23497
rect 15290 23423 15346 23432
rect 17498 23488 17554 23497
rect 17498 23423 17554 23432
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 10782 20904 10838 20913
rect 10782 20839 10838 20848
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9218 19952 9274 19961
rect 9218 19887 9274 19896
rect 12898 19952 12954 19961
rect 12898 19887 12954 19896
rect 9220 19304 9272 19310
rect 9034 19272 9090 19281
rect 9220 19246 9272 19252
rect 9034 19207 9090 19216
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7576 16250 7604 16526
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7668 16114 7696 16730
rect 9048 16590 9076 19207
rect 9126 17232 9182 17241
rect 9126 17167 9182 17176
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16250 9076 16526
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7668 15706 7696 16050
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 7668 15026 7696 15642
rect 8022 15464 8078 15473
rect 8022 15399 8078 15408
rect 9036 15428 9088 15434
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 13977 7512 14758
rect 7470 13968 7526 13977
rect 7470 13903 7526 13912
rect 7668 13870 7696 14962
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14074 7788 14418
rect 7944 14278 7972 14758
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7656 13864 7708 13870
rect 7392 13824 7512 13852
rect 7286 12336 7342 12345
rect 7286 12271 7342 12280
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7392 11558 7420 12242
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6472 10810 6500 10950
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6458 10432 6514 10441
rect 6458 10367 6514 10376
rect 6734 10432 6790 10441
rect 6734 10367 6790 10376
rect 6472 9897 6500 10367
rect 6458 9888 6514 9897
rect 6458 9823 6514 9832
rect 6748 9466 6776 10367
rect 6748 9438 6868 9466
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6380 9132 6592 9160
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6104 8452 6316 8480
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5446 7032 5502 7041
rect 5552 7002 5580 7346
rect 5446 6967 5502 6976
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5354 6760 5410 6769
rect 5354 6695 5356 6704
rect 5408 6695 5410 6704
rect 5356 6666 5408 6672
rect 5262 6488 5318 6497
rect 5080 6452 5132 6458
rect 5262 6423 5318 6432
rect 5080 6394 5132 6400
rect 5368 6322 5396 6666
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5460 5817 5488 6598
rect 5552 6304 5580 6938
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5632 6316 5684 6322
rect 5552 6276 5632 6304
rect 5632 6258 5684 6264
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5446 5808 5502 5817
rect 5446 5743 5502 5752
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5354 5536 5410 5545
rect 4802 5400 4858 5409
rect 4802 5335 4858 5344
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4724 3534 4752 5170
rect 4816 4593 4844 5335
rect 5078 4720 5134 4729
rect 5276 4690 5304 5510
rect 5354 5471 5410 5480
rect 5368 5137 5396 5471
rect 5460 5166 5488 5743
rect 5448 5160 5500 5166
rect 5354 5128 5410 5137
rect 5448 5102 5500 5108
rect 5354 5063 5410 5072
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5078 4655 5134 4664
rect 5264 4684 5316 4690
rect 4802 4584 4858 4593
rect 4802 4519 4858 4528
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4908 4146 4936 4490
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 2990 4752 3470
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4724 2446 4752 2926
rect 4816 2922 4844 3975
rect 5092 3398 5120 4655
rect 5264 4626 5316 4632
rect 5262 4176 5318 4185
rect 5262 4111 5264 4120
rect 5316 4111 5318 4120
rect 5264 4082 5316 4088
rect 5170 4040 5226 4049
rect 5170 3975 5226 3984
rect 5080 3392 5132 3398
rect 5184 3369 5212 3975
rect 5080 3334 5132 3340
rect 5170 3360 5226 3369
rect 5170 3295 5226 3304
rect 5276 3194 5304 4082
rect 5368 3942 5396 4966
rect 5552 4758 5580 5850
rect 6012 5624 6040 6054
rect 6104 5794 6132 8452
rect 6380 8378 6408 8570
rect 6288 8350 6408 8378
rect 6288 8090 6316 8350
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6276 8084 6328 8090
rect 6196 8044 6276 8072
rect 6196 7002 6224 8044
rect 6276 8026 6328 8032
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7313 6316 7686
rect 6380 7478 6408 8230
rect 6472 7818 6500 8978
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6274 7304 6330 7313
rect 6274 7239 6330 7248
rect 6458 7304 6514 7313
rect 6458 7239 6460 7248
rect 6512 7239 6514 7248
rect 6460 7210 6512 7216
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 5914 6224 6802
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6288 5846 6316 6734
rect 6276 5840 6328 5846
rect 6104 5766 6224 5794
rect 6276 5782 6328 5788
rect 6012 5596 6132 5624
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5998 5400 6054 5409
rect 5998 5335 6054 5344
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5736 4826 5764 5170
rect 6012 5030 6040 5335
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5552 4078 5580 4694
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5368 3097 5396 3878
rect 5552 3738 5580 4014
rect 6012 3738 6040 4966
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5354 3088 5410 3097
rect 5354 3023 5410 3032
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4816 1442 4844 2858
rect 4724 1414 4844 1442
rect 5552 1442 5580 3538
rect 6104 3482 6132 5596
rect 6196 3602 6224 5766
rect 6288 5273 6316 5782
rect 6472 5370 6500 6734
rect 6564 6390 6592 9132
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6656 6798 6684 8366
rect 6748 7886 6776 9318
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6274 5264 6330 5273
rect 6274 5199 6330 5208
rect 6472 4282 6500 5306
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6276 3528 6328 3534
rect 6104 3454 6224 3482
rect 6276 3470 6328 3476
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6196 2582 6224 3454
rect 6288 2922 6316 3470
rect 6380 3074 6408 3674
rect 6472 3194 6500 4218
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6380 3046 6500 3074
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 5906 2408 5962 2417
rect 5906 2343 5908 2352
rect 5960 2343 5962 2352
rect 5908 2314 5960 2320
rect 6196 2310 6224 2518
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5552 1414 5856 1442
rect 4620 604 4672 610
rect 4620 546 4672 552
rect 4724 480 4752 1414
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5276 480 5304 546
rect 5828 480 5856 1414
rect 4434 96 4490 105
rect 4434 31 4490 40
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6196 377 6224 2246
rect 6380 480 6408 2926
rect 6472 2854 6500 3046
rect 6564 2961 6592 3946
rect 6656 2990 6684 6598
rect 6748 3942 6776 7822
rect 6840 7342 6868 9438
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 7024 8974 7052 9386
rect 7116 8974 7144 10746
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 6662 6868 7278
rect 7024 6848 7052 8434
rect 7116 7188 7144 8774
rect 7208 8090 7236 11018
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7300 9602 7328 10406
rect 7291 9574 7328 9602
rect 7392 9586 7420 11494
rect 7484 9761 7512 13824
rect 7656 13806 7708 13812
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7760 12986 7788 13330
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7944 12918 7972 14214
rect 8036 13258 8064 15399
rect 9036 15370 9088 15376
rect 9048 14618 9076 15370
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8404 14385 8432 14418
rect 8390 14376 8446 14385
rect 8390 14311 8446 14320
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8208 13864 8260 13870
rect 8206 13832 8208 13841
rect 8260 13832 8262 13841
rect 8206 13767 8262 13776
rect 8312 13530 8340 14214
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 8128 12782 8156 13466
rect 8206 13424 8262 13433
rect 8206 13359 8262 13368
rect 7564 12776 7616 12782
rect 7562 12744 7564 12753
rect 8116 12776 8168 12782
rect 7616 12744 7618 12753
rect 8220 12753 8248 13359
rect 8116 12718 8168 12724
rect 8206 12744 8262 12753
rect 7562 12679 7618 12688
rect 7932 12708 7984 12714
rect 8206 12679 8262 12688
rect 7932 12650 7984 12656
rect 7654 12200 7710 12209
rect 7654 12135 7710 12144
rect 7562 10568 7618 10577
rect 7562 10503 7618 10512
rect 7470 9752 7526 9761
rect 7470 9687 7526 9696
rect 7576 9586 7604 10503
rect 7380 9580 7432 9586
rect 7291 9500 7319 9574
rect 7380 9522 7432 9528
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7668 9518 7696 12135
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7852 10266 7880 11222
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7760 9654 7788 10134
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9512 7708 9518
rect 7291 9472 7328 9500
rect 7300 8430 7328 9472
rect 7656 9454 7708 9460
rect 7852 9450 7880 9862
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7378 9344 7434 9353
rect 7378 9279 7434 9288
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7208 7410 7236 8026
rect 7392 7970 7420 9279
rect 7852 9178 7880 9386
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7300 7942 7420 7970
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7196 7200 7248 7206
rect 7116 7160 7196 7188
rect 7196 7142 7248 7148
rect 7024 6820 7144 6848
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6361 7052 6598
rect 7010 6352 7066 6361
rect 7010 6287 7012 6296
rect 7064 6287 7066 6296
rect 7012 6258 7064 6264
rect 7024 6227 7052 6258
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6840 5234 6868 5850
rect 6932 5681 6960 6054
rect 7116 5794 7144 6820
rect 7024 5766 7144 5794
rect 6918 5672 6974 5681
rect 7024 5642 7052 5766
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 6918 5607 6974 5616
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7116 5545 7144 5646
rect 7102 5536 7158 5545
rect 7102 5471 7158 5480
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 2984 6696 2990
rect 6550 2952 6606 2961
rect 6644 2926 6696 2932
rect 6550 2887 6606 2896
rect 6460 2848 6512 2854
rect 6458 2816 6460 2825
rect 6512 2816 6514 2825
rect 6458 2751 6514 2760
rect 6564 2310 6592 2887
rect 6840 2650 6868 4014
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7116 3466 7144 3878
rect 7208 3738 7236 7142
rect 7300 7002 7328 7942
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7410 7420 7822
rect 7944 7562 7972 12650
rect 8312 12442 8340 13466
rect 8390 13424 8446 13433
rect 8390 13359 8446 13368
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11762 8248 12038
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8312 11354 8340 11630
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8036 10470 8064 11086
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8220 9926 8248 11154
rect 8298 10976 8354 10985
rect 8298 10911 8354 10920
rect 8312 10305 8340 10911
rect 8298 10296 8354 10305
rect 8298 10231 8354 10240
rect 8404 10130 8432 13359
rect 8772 13326 8800 13806
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8772 12986 8800 13262
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 9048 12782 9076 14554
rect 9140 12986 9168 17167
rect 9232 14657 9260 19246
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 9402 17232 9458 17241
rect 9402 17167 9458 17176
rect 9218 14648 9274 14657
rect 9218 14583 9274 14592
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9232 12458 9260 14583
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9324 14074 9352 14282
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9416 13190 9444 17167
rect 9862 17096 9918 17105
rect 9862 17031 9918 17040
rect 9586 15600 9642 15609
rect 9508 15558 9586 15586
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9416 12646 9444 12922
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9140 12430 9260 12458
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8588 11354 8616 12310
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11762 8892 12038
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8864 11558 8892 11698
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8482 10568 8538 10577
rect 8482 10503 8538 10512
rect 8496 10198 8524 10503
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8036 9625 8064 9862
rect 8022 9616 8078 9625
rect 8022 9551 8078 9560
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8036 8566 8064 9046
rect 8220 8634 8248 9862
rect 8680 9722 8708 9998
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8864 9654 8892 11494
rect 9140 11286 9168 12430
rect 9218 12200 9274 12209
rect 9218 12135 9220 12144
rect 9272 12135 9274 12144
rect 9220 12106 9272 12112
rect 9324 11694 9352 12582
rect 9508 12458 9536 15558
rect 9586 15535 9642 15544
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 13530 9628 14418
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9416 12430 9536 12458
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8956 9994 8984 11154
rect 9310 10976 9366 10985
rect 9310 10911 9366 10920
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 9126 9480 9182 9489
rect 9126 9415 9182 9424
rect 9140 8838 9168 9415
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8036 8022 8064 8502
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7576 7534 7972 7562
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6118 7420 6598
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7300 5914 7328 6054
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7300 5370 7328 5850
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7392 4826 7420 6054
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7196 3392 7248 3398
rect 7300 3369 7328 3878
rect 7196 3334 7248 3340
rect 7286 3360 7342 3369
rect 7208 2990 7236 3334
rect 7286 3295 7342 3304
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7024 2689 7052 2926
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7010 2680 7066 2689
rect 6828 2644 6880 2650
rect 7010 2615 7066 2624
rect 6828 2586 6880 2592
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6840 2417 6868 2450
rect 6826 2408 6882 2417
rect 6826 2343 6882 2352
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 7300 1329 7328 2858
rect 7286 1320 7342 1329
rect 7286 1255 7342 1264
rect 6932 598 7052 626
rect 6932 480 6960 598
rect 6182 368 6238 377
rect 6182 303 6238 312
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7024 241 7052 598
rect 7576 480 7604 7534
rect 8036 7206 8064 7822
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7760 4729 7788 7142
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7852 6633 7880 6734
rect 7838 6624 7894 6633
rect 7838 6559 7894 6568
rect 7852 6390 7880 6559
rect 7944 6458 7972 6938
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7840 6384 7892 6390
rect 7944 6361 7972 6394
rect 7840 6326 7892 6332
rect 7930 6352 7986 6361
rect 7930 6287 7986 6296
rect 8128 5114 8156 7686
rect 8404 7342 8432 7890
rect 8496 7886 8524 8230
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8680 7546 8708 7822
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6118 8248 6734
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5778 8248 6054
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8220 5234 8248 5714
rect 8496 5642 8524 6258
rect 8574 6216 8630 6225
rect 8574 6151 8630 6160
rect 8588 6118 8616 6151
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8024 5092 8076 5098
rect 8128 5086 8248 5114
rect 8024 5034 8076 5040
rect 7746 4720 7802 4729
rect 7746 4655 7802 4664
rect 8036 4622 8064 5034
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7852 3194 7880 3538
rect 7944 3534 7972 4082
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7944 2854 7972 3334
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7760 2009 7788 2450
rect 7746 2000 7802 2009
rect 7746 1935 7802 1944
rect 7944 1193 7972 2790
rect 7930 1184 7986 1193
rect 7930 1119 7986 1128
rect 8036 649 8064 4558
rect 8128 3233 8156 4966
rect 8220 3777 8248 5086
rect 8588 4865 8616 5510
rect 8574 4856 8630 4865
rect 8574 4791 8630 4800
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8206 3768 8262 3777
rect 8312 3738 8340 4422
rect 8588 4214 8616 4558
rect 8576 4208 8628 4214
rect 8390 4176 8446 4185
rect 8576 4150 8628 4156
rect 8390 4111 8392 4120
rect 8444 4111 8446 4120
rect 8392 4082 8444 4088
rect 8206 3703 8262 3712
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8404 3670 8432 4082
rect 8680 4026 8708 7482
rect 8956 7206 8984 7686
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8956 6905 8984 7142
rect 9048 6934 9076 7142
rect 9036 6928 9088 6934
rect 8942 6896 8998 6905
rect 9036 6870 9088 6876
rect 9140 6866 9168 8774
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9232 7002 9260 7346
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8942 6831 8998 6840
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8864 5137 8892 6122
rect 8956 5846 8984 6598
rect 9232 6458 9260 6938
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9324 6338 9352 10911
rect 9232 6310 9352 6338
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8956 5681 8984 5782
rect 8942 5672 8998 5681
rect 8942 5607 8998 5616
rect 8850 5128 8906 5137
rect 8850 5063 8906 5072
rect 8852 4752 8904 4758
rect 8852 4694 8904 4700
rect 8588 3998 8708 4026
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8114 3224 8170 3233
rect 8114 3159 8170 3168
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8022 640 8078 649
rect 8078 598 8156 626
rect 8022 575 8078 584
rect 8128 480 8156 598
rect 7010 232 7066 241
rect 7010 167 7066 176
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8220 241 8248 3130
rect 8312 3058 8340 3334
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8588 2990 8616 3998
rect 8668 3936 8720 3942
rect 8760 3936 8812 3942
rect 8668 3878 8720 3884
rect 8758 3904 8760 3913
rect 8812 3904 8814 3913
rect 8680 3346 8708 3878
rect 8758 3839 8814 3848
rect 8864 3534 8892 4694
rect 8956 3602 8984 5607
rect 9034 5264 9090 5273
rect 9034 5199 9090 5208
rect 9048 4457 9076 5199
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9034 4448 9090 4457
rect 9034 4383 9090 4392
rect 9034 4312 9090 4321
rect 9034 4247 9090 4256
rect 9048 4078 9076 4247
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8852 3528 8904 3534
rect 8850 3496 8852 3505
rect 8904 3496 8906 3505
rect 8850 3431 8906 3440
rect 8680 3318 8892 3346
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8404 2650 8432 2926
rect 8666 2816 8722 2825
rect 8666 2751 8722 2760
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8680 480 8708 2751
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 785 8800 2246
rect 8864 1737 8892 3318
rect 9140 2514 9168 4762
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 8850 1728 8906 1737
rect 8850 1663 8906 1672
rect 8864 921 8892 1663
rect 8850 912 8906 921
rect 8850 847 8906 856
rect 8758 776 8814 785
rect 8758 711 8814 720
rect 9232 480 9260 6310
rect 9416 6202 9444 12430
rect 9600 12374 9628 12718
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9600 11694 9628 11766
rect 9588 11688 9640 11694
rect 9586 11656 9588 11665
rect 9640 11656 9642 11665
rect 9586 11591 9642 11600
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11286 9628 11494
rect 9588 11280 9640 11286
rect 9586 11248 9588 11257
rect 9640 11248 9642 11257
rect 9586 11183 9642 11192
rect 9600 11157 9628 11183
rect 9692 10826 9720 15438
rect 9876 13462 9904 17031
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 11610 16144 11666 16153
rect 11610 16079 11666 16088
rect 11334 16008 11390 16017
rect 11334 15943 11390 15952
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11242 15872 11298 15881
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10152 15366 10180 15642
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 14482 9996 14758
rect 10152 14550 10180 15302
rect 10598 15056 10654 15065
rect 10598 14991 10600 15000
rect 10652 14991 10654 15000
rect 10600 14962 10652 14968
rect 10876 14816 10928 14822
rect 10980 14804 11008 15506
rect 11072 14958 11100 15846
rect 11242 15807 11298 15816
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11060 14816 11112 14822
rect 10980 14776 11060 14804
rect 10876 14758 10928 14764
rect 11060 14758 11112 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 13870 9996 14418
rect 10046 14104 10102 14113
rect 10046 14039 10102 14048
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 10060 13530 10088 14039
rect 10888 13852 10916 14758
rect 11072 14278 11100 14758
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13938 11100 14214
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10138 13832 10194 13841
rect 10888 13824 11008 13852
rect 10980 13818 11008 13824
rect 10980 13790 11100 13818
rect 10138 13767 10194 13776
rect 10048 13524 10100 13530
rect 9968 13484 10048 13512
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9784 11762 9812 12786
rect 9876 12714 9904 13398
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9862 12472 9918 12481
rect 9862 12407 9864 12416
rect 9916 12407 9918 12416
rect 9864 12378 9916 12384
rect 9968 12102 9996 13484
rect 10048 13466 10100 13472
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10060 12714 10088 13330
rect 10152 13308 10180 13767
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 11072 13530 11100 13790
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10232 13320 10284 13326
rect 10152 13280 10232 13308
rect 10232 13262 10284 13268
rect 10244 12986 10272 13262
rect 10692 13184 10744 13190
rect 11060 13184 11112 13190
rect 10692 13126 10744 13132
rect 10782 13152 10838 13161
rect 10704 13025 10732 13126
rect 11060 13126 11112 13132
rect 10782 13087 10838 13096
rect 10690 13016 10746 13025
rect 10232 12980 10284 12986
rect 10690 12951 10746 12960
rect 10232 12922 10284 12928
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12481 10732 12582
rect 10690 12472 10746 12481
rect 10690 12407 10746 12416
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 9956 12096 10008 12102
rect 9862 12064 9918 12073
rect 9956 12038 10008 12044
rect 9862 11999 9918 12008
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9784 11393 9812 11562
rect 9876 11558 9904 11999
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9770 11384 9826 11393
rect 9876 11354 9904 11494
rect 9968 11393 9996 12038
rect 10336 11694 10364 12174
rect 10428 11830 10456 12310
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10324 11688 10376 11694
rect 10152 11648 10324 11676
rect 9954 11384 10010 11393
rect 9770 11319 9826 11328
rect 9864 11348 9916 11354
rect 9954 11319 10010 11328
rect 9864 11290 9916 11296
rect 10152 11150 10180 11648
rect 10324 11630 10376 11636
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 9864 11144 9916 11150
rect 10140 11144 10192 11150
rect 9864 11086 9916 11092
rect 9968 11104 10140 11132
rect 9600 10798 9720 10826
rect 9772 10804 9824 10810
rect 9600 10266 9628 10798
rect 9772 10746 9824 10752
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9489 9536 9930
rect 9494 9480 9550 9489
rect 9494 9415 9550 9424
rect 9588 8628 9640 8634
rect 9692 8616 9720 10678
rect 9640 8588 9720 8616
rect 9588 8570 9640 8576
rect 9692 7954 9720 8588
rect 9784 8430 9812 10746
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7478 9536 7686
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9508 7342 9536 7414
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9784 6798 9812 7890
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9784 6254 9812 6734
rect 9324 6174 9444 6202
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9324 4826 9352 6174
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5914 9444 6054
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9692 5370 9720 5714
rect 9784 5545 9812 6190
rect 9770 5536 9826 5545
rect 9770 5471 9826 5480
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9402 5264 9458 5273
rect 9402 5199 9458 5208
rect 9416 5166 9444 5199
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9600 4706 9628 4966
rect 9680 4752 9732 4758
rect 9600 4700 9680 4706
rect 9600 4694 9732 4700
rect 9404 4684 9456 4690
rect 9600 4678 9720 4694
rect 9404 4626 9456 4632
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9324 3534 9352 4558
rect 9416 4282 9444 4626
rect 9784 4622 9812 5471
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9404 4276 9456 4282
rect 9456 4236 9628 4264
rect 9404 4218 9456 4224
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9416 3602 9444 4082
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9312 2440 9364 2446
rect 9310 2408 9312 2417
rect 9364 2408 9366 2417
rect 9310 2343 9366 2352
rect 9416 2145 9444 2926
rect 9508 2582 9536 3674
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9402 2136 9458 2145
rect 9402 2071 9458 2080
rect 9600 1737 9628 4236
rect 9692 3194 9720 4422
rect 9876 3890 9904 11086
rect 9968 10062 9996 11104
rect 10140 11086 10192 11092
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 10060 9722 10088 10134
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10060 8634 10088 9658
rect 10152 9178 10180 10542
rect 10336 10538 10364 11154
rect 10704 10674 10732 12310
rect 10796 11898 10824 13087
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 12617 10916 12650
rect 10874 12608 10930 12617
rect 10874 12543 10930 12552
rect 10980 12084 11008 12922
rect 11072 12782 11100 13126
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11060 12096 11112 12102
rect 10980 12056 11060 12084
rect 11060 12038 11112 12044
rect 10874 11928 10930 11937
rect 10784 11892 10836 11898
rect 10874 11863 10930 11872
rect 10784 11834 10836 11840
rect 10888 11121 10916 11863
rect 11164 11529 11192 13670
rect 11256 11665 11284 15807
rect 11242 11656 11298 11665
rect 11242 11591 11298 11600
rect 11150 11520 11206 11529
rect 11150 11455 11206 11464
rect 10874 11112 10930 11121
rect 10874 11047 10930 11056
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 9722 10732 10474
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10598 9616 10654 9625
rect 10796 9586 10824 10406
rect 10980 9982 11192 10010
rect 10980 9926 11008 9982
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10598 9551 10654 9560
rect 10784 9580 10836 9586
rect 10612 9518 10640 9551
rect 10784 9522 10836 9528
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10704 8634 10732 9318
rect 10796 9178 10824 9522
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8945 10824 8978
rect 10876 8968 10928 8974
rect 10782 8936 10838 8945
rect 10876 8910 10928 8916
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10782 8871 10838 8880
rect 10782 8800 10838 8809
rect 10782 8735 10838 8744
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10796 8362 10824 8735
rect 10888 8498 10916 8910
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10152 8129 10180 8298
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10138 8120 10194 8129
rect 10289 8112 10585 8132
rect 10980 8090 11008 8910
rect 10138 8055 10140 8064
rect 10192 8055 10194 8064
rect 10968 8084 11020 8090
rect 10140 8026 10192 8032
rect 10968 8026 11020 8032
rect 11072 7970 11100 9658
rect 11164 8838 11192 9982
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10980 7954 11100 7970
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 10968 7948 11100 7954
rect 11020 7942 11100 7948
rect 10968 7890 11020 7896
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9968 7449 9996 7822
rect 9954 7440 10010 7449
rect 9954 7375 10010 7384
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10690 7304 10746 7313
rect 10690 7239 10746 7248
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 9954 7032 10010 7041
rect 9954 6967 10010 6976
rect 9968 6934 9996 6967
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 10060 6866 10088 7142
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10152 5778 10180 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 5166 10088 5510
rect 10428 5370 10456 5646
rect 10704 5522 10732 7239
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 6662 10824 7142
rect 10888 6866 10916 7346
rect 11164 7206 11192 7958
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 7002 11192 7142
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10888 6118 10916 6802
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10782 5944 10838 5953
rect 10782 5879 10838 5888
rect 10796 5846 10824 5879
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10612 5494 10732 5522
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10612 5012 10640 5494
rect 10796 5250 10824 5782
rect 10888 5302 10916 6054
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10980 5370 11008 5714
rect 11164 5710 11192 6938
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10704 5234 10824 5250
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10692 5228 10824 5234
rect 10744 5222 10824 5228
rect 10692 5170 10744 5176
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10612 4984 10732 5012
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10060 3942 10088 4626
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10520 4185 10548 4422
rect 10322 4176 10378 4185
rect 10322 4111 10378 4120
rect 10506 4176 10562 4185
rect 10506 4111 10562 4120
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 9784 3862 9904 3890
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9692 2650 9720 3130
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 9784 480 9812 3862
rect 9954 3768 10010 3777
rect 10060 3738 10088 3878
rect 9954 3703 10010 3712
rect 10048 3732 10100 3738
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9876 2854 9904 3606
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9862 2680 9918 2689
rect 9862 2615 9918 2624
rect 9876 2378 9904 2615
rect 9968 2514 9996 3703
rect 10048 3674 10100 3680
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 10060 2446 10088 3674
rect 10152 3641 10180 4014
rect 10336 4010 10364 4111
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10138 3632 10194 3641
rect 10704 3618 10732 4984
rect 10796 4282 10824 5102
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10138 3567 10194 3576
rect 10244 3590 10732 3618
rect 11256 3618 11284 11591
rect 11348 10810 11376 15943
rect 11624 13954 11652 16079
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12544 15609 12572 15642
rect 12530 15600 12586 15609
rect 12530 15535 12586 15544
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11716 14278 11744 14486
rect 11992 14278 12020 14826
rect 12084 14822 12112 14894
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11716 14074 11744 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11992 14006 12020 14214
rect 11980 14000 12032 14006
rect 11624 13926 11744 13954
rect 11980 13942 12032 13948
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 13025 11468 13806
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11426 13016 11482 13025
rect 11426 12951 11482 12960
rect 11624 12442 11652 13466
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11426 12200 11482 12209
rect 11426 12135 11482 12144
rect 11440 11762 11468 12135
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11440 11286 11468 11698
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11532 11082 11560 12378
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11532 10810 11560 11018
rect 11624 11014 11652 11494
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 10266 11468 10406
rect 11532 10266 11560 10746
rect 11624 10674 11652 10950
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11532 9722 11560 10202
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11716 8838 11744 13926
rect 12084 13852 12112 14758
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11992 13824 12112 13852
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 12986 11928 13262
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11808 11830 11836 12038
rect 11900 11830 11928 12922
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11992 10169 12020 13824
rect 12176 13734 12204 14350
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11348 6254 11376 6326
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 4826 11376 6190
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11348 4146 11376 4762
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11348 3738 11376 4082
rect 11440 4010 11468 7958
rect 11532 6905 11560 8774
rect 11992 8294 12020 8978
rect 11980 8288 12032 8294
rect 11978 8256 11980 8265
rect 12032 8256 12034 8265
rect 11978 8191 12034 8200
rect 11886 7712 11942 7721
rect 11886 7647 11942 7656
rect 11900 7546 11928 7647
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11518 6896 11574 6905
rect 11518 6831 11574 6840
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11702 5128 11758 5137
rect 11702 5063 11758 5072
rect 11716 4826 11744 5063
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11256 3590 11468 3618
rect 10244 3516 10272 3590
rect 10152 3488 10272 3516
rect 10506 3496 10562 3505
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 10152 1442 10180 3488
rect 10506 3431 10562 3440
rect 10520 3097 10548 3431
rect 10506 3088 10562 3097
rect 10506 3023 10562 3032
rect 11164 2854 11192 2885
rect 11152 2848 11204 2854
rect 11150 2816 11152 2825
rect 11244 2848 11296 2854
rect 11204 2816 11206 2825
rect 10289 2748 10585 2768
rect 11244 2790 11296 2796
rect 11150 2751 11206 2760
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11164 2650 11192 2751
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11256 2514 11284 2790
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 10152 1414 10364 1442
rect 10336 480 10364 1414
rect 10874 1184 10930 1193
rect 10874 1119 10930 1128
rect 11058 1184 11114 1193
rect 11058 1119 11114 1128
rect 10888 626 10916 1119
rect 11072 921 11100 1119
rect 11058 912 11114 921
rect 11058 847 11114 856
rect 10888 598 11008 626
rect 10888 480 10916 598
rect 8206 232 8262 241
rect 8206 167 8262 176
rect 8666 0 8722 480
rect 9218 0 9274 480
rect 9770 0 9826 480
rect 10322 0 10378 480
rect 10874 0 10930 480
rect 10980 377 11008 598
rect 11440 480 11468 3590
rect 11716 2514 11744 4762
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1601 11652 2246
rect 11610 1592 11666 1601
rect 11610 1527 11666 1536
rect 11808 1465 11836 6190
rect 11886 5808 11942 5817
rect 12084 5778 12112 12650
rect 12162 10160 12218 10169
rect 12162 10095 12218 10104
rect 12176 9897 12204 10095
rect 12162 9888 12218 9897
rect 12162 9823 12218 9832
rect 12268 9722 12296 15370
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 15026 12480 15302
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12360 13530 12388 14758
rect 12452 14550 12480 14962
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12360 12986 12388 13466
rect 12452 13326 12480 14214
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13326 12664 13670
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12438 12472 12494 12481
rect 12438 12407 12494 12416
rect 12346 11520 12402 11529
rect 12346 11455 12402 11464
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12162 9208 12218 9217
rect 12360 9178 12388 11455
rect 12452 10441 12480 12407
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12544 11558 12572 11630
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12544 10130 12572 10202
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12162 9143 12218 9152
rect 12348 9172 12400 9178
rect 12176 6458 12204 9143
rect 12348 9114 12400 9120
rect 12452 9024 12480 9590
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12360 8996 12480 9024
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12162 6352 12218 6361
rect 12162 6287 12218 6296
rect 12176 5817 12204 6287
rect 12162 5808 12218 5817
rect 11886 5743 11888 5752
rect 11940 5743 11942 5752
rect 12072 5772 12124 5778
rect 11888 5714 11940 5720
rect 12162 5743 12218 5752
rect 12072 5714 12124 5720
rect 11886 5400 11942 5409
rect 12084 5370 12112 5714
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 11886 5335 11942 5344
rect 12072 5364 12124 5370
rect 11900 5137 11928 5335
rect 12072 5306 12124 5312
rect 11886 5128 11942 5137
rect 11886 5063 11942 5072
rect 12268 5001 12296 5510
rect 12254 4992 12310 5001
rect 12254 4927 12310 4936
rect 12360 4826 12388 8996
rect 12544 8974 12572 9522
rect 12532 8968 12584 8974
rect 12438 8936 12494 8945
rect 12728 8945 12756 15846
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12820 14618 12848 14894
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12806 12336 12862 12345
rect 12806 12271 12862 12280
rect 12820 11801 12848 12271
rect 12806 11792 12862 11801
rect 12806 11727 12862 11736
rect 12532 8910 12584 8916
rect 12714 8936 12770 8945
rect 12438 8871 12494 8880
rect 12452 8634 12480 8871
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12544 8498 12572 8910
rect 12714 8871 12770 8880
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12714 8392 12770 8401
rect 12714 8327 12770 8336
rect 12728 8294 12756 8327
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12544 7546 12572 8026
rect 12728 7750 12756 8230
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12622 7168 12678 7177
rect 12622 7103 12678 7112
rect 12636 7002 12664 7103
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12636 6322 12664 6938
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5953 12480 6054
rect 12438 5944 12494 5953
rect 12438 5879 12494 5888
rect 12728 5642 12756 7686
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12820 5522 12848 11727
rect 12912 9654 12940 19887
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19281 15332 23423
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 20640 23254 20668 23559
rect 20628 23248 20680 23254
rect 20628 23190 20680 23196
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19536 22438 19564 23122
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19536 22137 19564 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 17958 22128 18014 22137
rect 17958 22063 18014 22072
rect 19522 22128 19578 22137
rect 19522 22063 19578 22072
rect 16210 20904 16266 20913
rect 16210 20839 16266 20848
rect 15290 19272 15346 19281
rect 15290 19207 15346 19216
rect 15934 18864 15990 18873
rect 15934 18799 15990 18808
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 12990 14512 13046 14521
rect 12990 14447 13046 14456
rect 13004 12617 13032 14447
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12990 12608 13046 12617
rect 12990 12543 13046 12552
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 7002 12940 7142
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13004 6610 13032 12543
rect 13188 12345 13216 13806
rect 13174 12336 13230 12345
rect 13174 12271 13230 12280
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 10538 13124 11018
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13188 10266 13216 10950
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13082 7576 13138 7585
rect 13082 7511 13138 7520
rect 13096 6866 13124 7511
rect 13188 7342 13216 8910
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13176 6792 13228 6798
rect 12912 6582 13032 6610
rect 13096 6740 13176 6746
rect 13096 6734 13228 6740
rect 13096 6718 13216 6734
rect 12912 6186 12940 6582
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 13004 5794 13032 6394
rect 13096 6118 13124 6718
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13188 5914 13216 6598
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13004 5766 13216 5794
rect 12636 5137 12664 5510
rect 12820 5494 13032 5522
rect 12622 5128 12678 5137
rect 12622 5063 12678 5072
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11900 2990 11928 3946
rect 12544 3738 12572 4422
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 11978 3224 12034 3233
rect 11978 3159 12034 3168
rect 12440 3188 12492 3194
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11992 1465 12020 3159
rect 12440 3130 12492 3136
rect 12452 2582 12480 3130
rect 12544 2650 12572 3674
rect 12636 3398 12664 4966
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 12714 4176 12770 4185
rect 12714 4111 12716 4120
rect 12768 4111 12770 4120
rect 12716 4082 12768 4088
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12728 3058 12756 4082
rect 12820 3602 12848 4694
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12728 2514 12756 2994
rect 12912 2689 12940 5034
rect 13004 2854 13032 5494
rect 13082 5128 13138 5137
rect 13082 5063 13138 5072
rect 13096 4826 13124 5063
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13188 3754 13216 5766
rect 13280 3777 13308 15846
rect 13372 11286 13400 16594
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14462 16144 14518 16153
rect 14280 16108 14332 16114
rect 15856 16114 15884 17070
rect 14462 16079 14518 16088
rect 15844 16108 15896 16114
rect 14280 16050 14332 16056
rect 13544 16040 13596 16046
rect 13820 16040 13872 16046
rect 13544 15982 13596 15988
rect 13648 15988 13820 15994
rect 13648 15982 13872 15988
rect 13556 15910 13584 15982
rect 13648 15966 13860 15982
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13450 15600 13506 15609
rect 13450 15535 13506 15544
rect 13464 15502 13492 15535
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13464 14822 13492 15438
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13464 13433 13492 14758
rect 13556 14521 13584 15846
rect 13542 14512 13598 14521
rect 13542 14447 13598 14456
rect 13450 13424 13506 13433
rect 13450 13359 13506 13368
rect 13648 13258 13676 15966
rect 14292 15910 14320 16050
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13740 15450 13768 15574
rect 14292 15502 14320 15846
rect 14280 15496 14332 15502
rect 13740 15422 13860 15450
rect 14280 15438 14332 15444
rect 13832 14822 13860 15422
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 14002 13696 14058 13705
rect 14002 13631 14058 13640
rect 13910 13560 13966 13569
rect 13910 13495 13966 13504
rect 13924 13297 13952 13495
rect 13910 13288 13966 13297
rect 13636 13252 13688 13258
rect 13910 13223 13966 13232
rect 13636 13194 13688 13200
rect 13452 13184 13504 13190
rect 13450 13152 13452 13161
rect 13504 13152 13506 13161
rect 13450 13087 13506 13096
rect 13464 12782 13492 13087
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13648 12442 13676 12922
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13740 12306 13768 12582
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13452 12096 13504 12102
rect 13504 12056 13584 12084
rect 13452 12038 13504 12044
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 10713 13400 11086
rect 13358 10704 13414 10713
rect 13358 10639 13414 10648
rect 13372 10470 13400 10639
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13372 9625 13400 10406
rect 13556 10266 13584 12056
rect 13832 11642 13860 12378
rect 13924 12238 13952 13223
rect 14016 12442 14044 13631
rect 14292 13376 14320 15438
rect 14372 13388 14424 13394
rect 14292 13348 14372 13376
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 12986 14136 13262
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13832 11614 13952 11642
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13740 10810 13768 11222
rect 13832 11150 13860 11494
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13648 10062 13676 10406
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13358 9616 13414 9625
rect 13358 9551 13414 9560
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13372 5760 13400 8298
rect 13464 7834 13492 9862
rect 13556 8634 13584 9998
rect 13648 9450 13676 9998
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13648 9042 13676 9386
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13740 8498 13768 10474
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13464 7806 13584 7834
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 6361 13492 7686
rect 13450 6352 13506 6361
rect 13450 6287 13506 6296
rect 13452 6112 13504 6118
rect 13450 6080 13452 6089
rect 13504 6080 13506 6089
rect 13450 6015 13506 6024
rect 13452 5772 13504 5778
rect 13372 5732 13452 5760
rect 13452 5714 13504 5720
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13096 3726 13216 3754
rect 13266 3768 13322 3777
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 12898 2680 12954 2689
rect 12898 2615 12954 2624
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12530 2000 12586 2009
rect 12530 1935 12586 1944
rect 11794 1456 11850 1465
rect 11794 1391 11850 1400
rect 11978 1456 12034 1465
rect 11978 1391 12034 1400
rect 11992 480 12020 1391
rect 12544 480 12572 1935
rect 13096 480 13124 3726
rect 13266 3703 13322 3712
rect 13372 3618 13400 5578
rect 13464 5030 13492 5714
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13188 3590 13400 3618
rect 13188 2514 13216 3590
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13372 3194 13400 3470
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13188 1057 13216 2450
rect 13464 2281 13492 4966
rect 13556 4729 13584 7806
rect 13740 7546 13768 8434
rect 13832 7954 13860 8502
rect 13924 8362 13952 11614
rect 14016 11354 14044 12242
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14108 11898 14136 12174
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14002 10432 14058 10441
rect 14002 10367 14058 10376
rect 14016 8838 14044 10367
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14016 8430 14044 8774
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13924 8090 13952 8298
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13832 7721 13860 7890
rect 13818 7712 13874 7721
rect 13818 7647 13874 7656
rect 13818 7576 13874 7585
rect 13728 7540 13780 7546
rect 13818 7511 13874 7520
rect 13728 7482 13780 7488
rect 13636 7336 13688 7342
rect 13832 7313 13860 7511
rect 13636 7278 13688 7284
rect 13818 7304 13874 7313
rect 13648 6934 13676 7278
rect 13728 7268 13780 7274
rect 13818 7239 13874 7248
rect 13728 7210 13780 7216
rect 13740 6984 13768 7210
rect 13740 6956 13860 6984
rect 13636 6928 13688 6934
rect 13688 6888 13768 6916
rect 13636 6870 13688 6876
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6322 13676 6734
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13648 5914 13676 6258
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13634 5808 13690 5817
rect 13634 5743 13636 5752
rect 13688 5743 13690 5752
rect 13636 5714 13688 5720
rect 13648 4826 13676 5714
rect 13740 5710 13768 6888
rect 13832 6254 13860 6956
rect 13924 6662 13952 7890
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14016 7206 14044 7822
rect 14094 7440 14150 7449
rect 14094 7375 14150 7384
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 7002 14044 7142
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 14016 6186 14044 6938
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5370 13768 5646
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13542 4720 13598 4729
rect 13542 4655 13598 4664
rect 13832 4010 13860 5034
rect 14108 4690 14136 7375
rect 14292 7274 14320 13348
rect 14372 13330 14424 13336
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12102 14412 12582
rect 14372 12096 14424 12102
rect 14476 12073 14504 16079
rect 15844 16050 15896 16056
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15304 15473 15332 15506
rect 15290 15464 15346 15473
rect 15290 15399 15346 15408
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 14958 14872 15302
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 15162 15332 15399
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14660 14414 14688 14826
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 13734 14688 14350
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14660 13462 14688 13670
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14372 12038 14424 12044
rect 14462 12064 14518 12073
rect 14384 11665 14412 12038
rect 14462 11999 14518 12008
rect 14370 11656 14426 11665
rect 14370 11591 14426 11600
rect 14476 8294 14504 11999
rect 14568 11626 14596 13126
rect 14660 12850 14688 13398
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14646 12336 14702 12345
rect 14646 12271 14702 12280
rect 14660 12238 14688 12271
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14660 11626 14688 12174
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14568 11354 14596 11562
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 8560 14608 8566
rect 14556 8502 14608 8508
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 8090 14504 8230
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 14568 7342 14596 8502
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14280 7268 14332 7274
rect 14200 7228 14280 7256
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13636 3528 13688 3534
rect 13634 3496 13636 3505
rect 13924 3505 13952 4626
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14108 3942 14136 4490
rect 14200 4078 14228 7228
rect 14280 7210 14332 7216
rect 14370 7168 14426 7177
rect 14370 7103 14426 7112
rect 14554 7168 14610 7177
rect 14554 7103 14610 7112
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14292 6458 14320 6802
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14292 5574 14320 5714
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14292 5234 14320 5510
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14384 5166 14412 7103
rect 14568 6866 14596 7103
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14462 6760 14518 6769
rect 14462 6695 14518 6704
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14384 4826 14412 5102
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4185 14320 4422
rect 14278 4176 14334 4185
rect 14278 4111 14334 4120
rect 14188 4072 14240 4078
rect 14476 4060 14504 6695
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14188 4014 14240 4020
rect 14292 4032 14504 4060
rect 14568 4049 14596 5510
rect 14660 5098 14688 9114
rect 14752 8090 14780 14758
rect 14844 14278 14872 14894
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 14922 14648 14978 14657
rect 14922 14583 14924 14592
rect 14976 14583 14978 14592
rect 14924 14554 14976 14560
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 13870 14872 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15200 14000 15252 14006
rect 15120 13960 15200 13988
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 15120 13394 15148 13960
rect 15200 13942 15252 13948
rect 15304 13870 15332 14486
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15304 13705 15332 13806
rect 15290 13696 15346 13705
rect 15290 13631 15346 13640
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12458 15332 13330
rect 15488 13326 15516 14758
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15476 13320 15528 13326
rect 15382 13288 15438 13297
rect 15476 13262 15528 13268
rect 15382 13223 15438 13232
rect 15212 12430 15332 12458
rect 15212 12374 15240 12430
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 14922 12200 14978 12209
rect 14844 12158 14922 12186
rect 14844 11529 14872 12158
rect 14922 12135 14978 12144
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14830 11520 14886 11529
rect 14830 11455 14886 11464
rect 14830 11248 14886 11257
rect 14830 11183 14886 11192
rect 14844 11014 14872 11183
rect 14936 11121 14964 11630
rect 15108 11552 15160 11558
rect 15106 11520 15108 11529
rect 15160 11520 15162 11529
rect 15106 11455 15162 11464
rect 14922 11112 14978 11121
rect 14922 11047 14924 11056
rect 14976 11047 14978 11056
rect 14924 11018 14976 11024
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10792 15332 11766
rect 15396 11218 15424 13223
rect 15488 12782 15516 13262
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15488 11558 15516 12242
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15120 10764 15332 10792
rect 15384 10804 15436 10810
rect 15120 10266 15148 10764
rect 15384 10746 15436 10752
rect 15290 10296 15346 10305
rect 15108 10260 15160 10266
rect 15290 10231 15292 10240
rect 15108 10202 15160 10208
rect 15344 10231 15346 10240
rect 15292 10202 15344 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14922 9480 14978 9489
rect 14922 9415 14924 9424
rect 14976 9415 14978 9424
rect 14924 9386 14976 9392
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 8566 14872 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14832 8560 14884 8566
rect 15304 8537 15332 9318
rect 15396 9178 15424 10746
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15488 9081 15516 11494
rect 15474 9072 15530 9081
rect 15384 9036 15436 9042
rect 15474 9007 15530 9016
rect 15384 8978 15436 8984
rect 15396 8634 15424 8978
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 14832 8502 14884 8508
rect 15290 8528 15346 8537
rect 15290 8463 15346 8472
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14844 8022 14872 8366
rect 14832 8016 14884 8022
rect 14830 7984 14832 7993
rect 14884 7984 14886 7993
rect 14830 7919 14886 7928
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14830 6896 14886 6905
rect 14830 6831 14832 6840
rect 14884 6831 14886 6840
rect 14832 6802 14884 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15580 6474 15608 14214
rect 15672 13870 15700 14418
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15764 14006 15792 14350
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15660 13864 15712 13870
rect 15948 13818 15976 18799
rect 16026 18320 16082 18329
rect 16026 18255 16082 18264
rect 16040 17338 16068 18255
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16224 16726 16252 20839
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17420 18902 17448 19246
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17144 18086 17172 18770
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16040 15366 16068 16526
rect 16224 16250 16252 16662
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 15660 13806 15712 13812
rect 15672 10810 15700 13806
rect 15856 13790 15976 13818
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 12442 15792 13262
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15856 12374 15884 13790
rect 16224 12986 16252 15846
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 15934 12880 15990 12889
rect 15934 12815 15990 12824
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11898 15792 12174
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15764 11801 15792 11834
rect 15750 11792 15806 11801
rect 15750 11727 15806 11736
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15764 10266 15792 11154
rect 15842 10840 15898 10849
rect 15842 10775 15898 10784
rect 15856 10538 15884 10775
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 9382 15700 9522
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 8945 15700 9318
rect 15658 8936 15714 8945
rect 15658 8871 15714 8880
rect 15658 8392 15714 8401
rect 15658 8327 15660 8336
rect 15712 8327 15714 8336
rect 15660 8298 15712 8304
rect 15764 6866 15792 10066
rect 15948 9654 15976 12815
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11626 16068 12174
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16040 11150 16068 11562
rect 16316 11354 16344 18022
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16684 14822 16712 15506
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16408 14074 16436 14486
rect 16500 14278 16528 14758
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16500 13938 16528 14214
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16672 13864 16724 13870
rect 16500 13812 16672 13818
rect 16500 13806 16724 13812
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16500 13790 16712 13806
rect 16408 13190 16436 13738
rect 16500 13530 16528 13790
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12714 16436 13126
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16132 11257 16160 11290
rect 16118 11248 16174 11257
rect 16118 11183 16174 11192
rect 16028 11144 16080 11150
rect 16026 11112 16028 11121
rect 16080 11112 16082 11121
rect 16026 11047 16082 11056
rect 16212 11008 16264 11014
rect 16026 10976 16082 10985
rect 16212 10950 16264 10956
rect 16026 10911 16082 10920
rect 16040 10441 16068 10911
rect 16026 10432 16082 10441
rect 16026 10367 16082 10376
rect 16118 10024 16174 10033
rect 16118 9959 16120 9968
rect 16172 9959 16174 9968
rect 16120 9930 16172 9936
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 16132 9518 16160 9930
rect 16224 9636 16252 10950
rect 16408 10792 16436 12650
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11762 16528 12038
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16316 10764 16436 10792
rect 16500 10792 16528 11698
rect 16592 11234 16620 12582
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16684 11354 16712 11766
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16592 11206 16712 11234
rect 16580 10804 16632 10810
rect 16500 10764 16580 10792
rect 16316 10606 16344 10764
rect 16580 10746 16632 10752
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16316 10441 16344 10542
rect 16302 10432 16358 10441
rect 16302 10367 16358 10376
rect 16316 10130 16344 10367
rect 16592 10198 16620 10746
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16592 9722 16620 10134
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16224 9608 16436 9636
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 15844 9104 15896 9110
rect 15844 9046 15896 9052
rect 16026 9072 16082 9081
rect 15856 7993 15884 9046
rect 16026 9007 16082 9016
rect 16040 8974 16068 9007
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15842 7984 15898 7993
rect 15948 7954 15976 8774
rect 16040 8537 16068 8910
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16026 8528 16082 8537
rect 16026 8463 16082 8472
rect 16040 8090 16068 8463
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 15842 7919 15898 7928
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15948 7750 15976 7890
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15948 7206 15976 7686
rect 16132 7546 16160 8774
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 15936 7200 15988 7206
rect 16316 7154 16344 7822
rect 15936 7142 15988 7148
rect 15948 7002 15976 7142
rect 16132 7126 16344 7154
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15580 6446 15700 6474
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 5710 15240 6190
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5778 15516 6054
rect 15476 5772 15528 5778
rect 15528 5732 15608 5760
rect 15476 5714 15528 5720
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15382 5672 15438 5681
rect 15382 5607 15438 5616
rect 15396 5574 15424 5607
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 14740 4480 14792 4486
rect 14646 4448 14702 4457
rect 14740 4422 14792 4428
rect 14646 4383 14702 4392
rect 14554 4040 14610 4049
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14186 3904 14242 3913
rect 13688 3496 13690 3505
rect 13634 3431 13690 3440
rect 13910 3496 13966 3505
rect 13910 3431 13966 3440
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 14016 2961 14044 3334
rect 14108 2990 14136 3878
rect 14186 3839 14242 3848
rect 14200 3670 14228 3839
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14096 2984 14148 2990
rect 14002 2952 14058 2961
rect 14096 2926 14148 2932
rect 14002 2887 14058 2896
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13450 2272 13506 2281
rect 13450 2207 13506 2216
rect 13174 1048 13230 1057
rect 13174 983 13230 992
rect 13648 480 13676 2790
rect 14094 2408 14150 2417
rect 14094 2343 14150 2352
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14016 2145 14044 2246
rect 14002 2136 14058 2145
rect 13728 2100 13780 2106
rect 14002 2071 14058 2080
rect 13728 2042 13780 2048
rect 13740 2009 13768 2042
rect 14108 2009 14136 2343
rect 13726 2000 13782 2009
rect 13726 1935 13782 1944
rect 14094 2000 14150 2009
rect 14094 1935 14150 1944
rect 14292 480 14320 4032
rect 14554 3975 14610 3984
rect 14554 3360 14610 3369
rect 14554 3295 14610 3304
rect 14568 3097 14596 3295
rect 14554 3088 14610 3097
rect 14660 3058 14688 4383
rect 14752 4321 14780 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14738 4312 14794 4321
rect 14956 4304 15252 4324
rect 15304 4282 15332 4762
rect 14738 4247 14794 4256
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15014 3768 15070 3777
rect 15014 3703 15070 3712
rect 15028 3534 15056 3703
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15396 3466 15424 5510
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15488 4729 15516 4966
rect 15580 4826 15608 5732
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15474 4720 15530 4729
rect 15474 4655 15530 4664
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4078 15608 4422
rect 15476 4072 15528 4078
rect 15474 4040 15476 4049
rect 15568 4072 15620 4078
rect 15528 4040 15530 4049
rect 15568 4014 15620 4020
rect 15474 3975 15530 3984
rect 15672 3738 15700 6446
rect 15764 5846 15792 6802
rect 16132 6798 16160 7126
rect 16408 6984 16436 9608
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16500 8362 16528 8978
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16316 6956 16436 6984
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16132 6633 16160 6734
rect 16118 6624 16174 6633
rect 16118 6559 16174 6568
rect 16132 6254 16160 6559
rect 16120 6248 16172 6254
rect 16172 6196 16252 6202
rect 16120 6190 16252 6196
rect 16132 6174 16252 6190
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5914 16160 6054
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 16132 5234 16160 5850
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15856 4282 15884 4966
rect 16224 4690 16252 6174
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15658 3360 15714 3369
rect 14956 3292 15252 3312
rect 15658 3295 15714 3304
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15672 3058 15700 3295
rect 14554 3023 14610 3032
rect 14648 3052 14700 3058
rect 14568 2258 14596 3023
rect 14648 2994 14700 3000
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14660 2553 14688 2858
rect 15200 2848 15252 2854
rect 15198 2816 15200 2825
rect 15252 2816 15254 2825
rect 15198 2751 15254 2760
rect 15856 2553 15884 4014
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16224 3534 16252 3878
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 3194 16252 3470
rect 16212 3188 16264 3194
rect 16212 3130 16264 3136
rect 14646 2544 14702 2553
rect 14646 2479 14702 2488
rect 15842 2544 15898 2553
rect 15842 2479 15898 2488
rect 15200 2440 15252 2446
rect 15198 2408 15200 2417
rect 15252 2408 15254 2417
rect 15198 2343 15254 2352
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 15476 2304 15528 2310
rect 15382 2272 15438 2281
rect 14568 2230 14872 2258
rect 14844 480 14872 2230
rect 14956 2204 15252 2224
rect 15476 2246 15528 2252
rect 15382 2207 15438 2216
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15396 2106 15424 2207
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 15396 480 15424 1906
rect 15488 1737 15516 2246
rect 15474 1728 15530 1737
rect 15474 1663 15530 1672
rect 16132 1170 16160 2314
rect 16316 1970 16344 6956
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16408 5914 16436 6802
rect 16500 6497 16528 7142
rect 16592 6934 16620 7278
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16486 6488 16542 6497
rect 16486 6423 16542 6432
rect 16578 6352 16634 6361
rect 16578 6287 16634 6296
rect 16592 6254 16620 6287
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16684 5545 16712 11206
rect 16776 9178 16804 16934
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15502 17080 15846
rect 17040 15496 17092 15502
rect 16946 15464 17002 15473
rect 17040 15438 17092 15444
rect 16946 15399 17002 15408
rect 16854 14376 16910 14385
rect 16960 14362 16988 15399
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 16910 14334 16988 14362
rect 16854 14311 16910 14320
rect 16854 13968 16910 13977
rect 16854 13903 16910 13912
rect 16868 13870 16896 13903
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16960 12322 16988 14334
rect 17052 12646 17080 14758
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13308 17172 13670
rect 17236 13433 17264 14214
rect 17222 13424 17278 13433
rect 17222 13359 17278 13368
rect 17144 13280 17264 13308
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16856 12300 16908 12306
rect 16960 12294 17080 12322
rect 16856 12242 16908 12248
rect 16868 12209 16896 12242
rect 16854 12200 16910 12209
rect 16910 12158 16988 12186
rect 16854 12135 16910 12144
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16868 11558 16896 12038
rect 16960 11898 16988 12158
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16946 11792 17002 11801
rect 16946 11727 17002 11736
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16776 8430 16804 9114
rect 16868 8906 16896 11494
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16854 8664 16910 8673
rect 16854 8599 16856 8608
rect 16908 8599 16910 8608
rect 16960 8616 16988 11727
rect 17052 9382 17080 12294
rect 17144 9518 17172 12786
rect 17236 9926 17264 13280
rect 17328 12850 17356 14758
rect 17420 14074 17448 17614
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17512 16794 17540 17274
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17776 15904 17828 15910
rect 17774 15872 17776 15881
rect 17828 15872 17830 15881
rect 17774 15807 17830 15816
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17880 14414 17908 14826
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17420 13870 17448 14010
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17880 13569 17908 13942
rect 17866 13560 17922 13569
rect 17866 13495 17922 13504
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17420 12442 17448 13330
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17512 12986 17540 13126
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17500 12776 17552 12782
rect 17498 12744 17500 12753
rect 17776 12776 17828 12782
rect 17552 12744 17554 12753
rect 17776 12718 17828 12724
rect 17498 12679 17554 12688
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17328 9874 17356 12038
rect 17420 10826 17448 12378
rect 17788 12186 17816 12718
rect 17696 12158 17816 12186
rect 17696 11830 17724 12158
rect 17972 12102 18000 22063
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 18326 20632 18382 20641
rect 18326 20567 18382 20576
rect 18340 19174 18368 20567
rect 20074 20224 20130 20233
rect 19996 20182 20074 20210
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 18694 19952 18750 19961
rect 18694 19887 18750 19896
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18512 15360 18564 15366
rect 18142 15328 18198 15337
rect 18512 15302 18564 15308
rect 18142 15263 18198 15272
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18064 14074 18092 14418
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18064 13530 18092 14010
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17788 11830 17816 12038
rect 18064 11914 18092 12582
rect 17880 11886 18092 11914
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17776 11688 17828 11694
rect 17880 11676 17908 11886
rect 18050 11792 18106 11801
rect 18050 11727 18106 11736
rect 18064 11694 18092 11727
rect 17828 11648 17908 11676
rect 17776 11630 17828 11636
rect 17776 11552 17828 11558
rect 17590 11520 17646 11529
rect 17776 11494 17828 11500
rect 17590 11455 17646 11464
rect 17420 10798 17540 10826
rect 17408 10736 17460 10742
rect 17406 10704 17408 10713
rect 17460 10704 17462 10713
rect 17406 10639 17462 10648
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 10169 17448 10406
rect 17406 10160 17462 10169
rect 17406 10095 17462 10104
rect 17328 9846 17448 9874
rect 17420 9704 17448 9846
rect 17328 9676 17448 9704
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16960 8588 17172 8616
rect 16856 8570 16908 8576
rect 16868 8430 16896 8570
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 7342 16804 8230
rect 16960 7954 16988 8434
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 17038 7032 17094 7041
rect 17038 6967 17094 6976
rect 16762 6896 16818 6905
rect 16762 6831 16818 6840
rect 16670 5536 16726 5545
rect 16670 5471 16726 5480
rect 16486 4992 16542 5001
rect 16486 4927 16542 4936
rect 16500 4690 16528 4927
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16500 4282 16528 4626
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16776 4146 16804 6831
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16868 5273 16896 6122
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 17052 3738 17080 6967
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16868 3641 16896 3674
rect 16854 3632 16910 3641
rect 16854 3567 16910 3576
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 15948 1142 16160 1170
rect 15948 480 15976 1142
rect 16500 480 16528 3062
rect 16684 3058 16712 3130
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16684 2446 16712 2994
rect 16776 2990 16804 3334
rect 17052 3126 17080 3674
rect 17144 3670 17172 8588
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17236 5370 17264 5782
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17132 3664 17184 3670
rect 17328 3641 17356 9676
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17420 5409 17448 9454
rect 17512 8090 17540 10798
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17512 7410 17540 8026
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17406 5400 17462 5409
rect 17406 5335 17462 5344
rect 17604 4321 17632 11455
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17696 10538 17724 11086
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 17696 10266 17724 10474
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17696 7392 17724 9862
rect 17788 9489 17816 11494
rect 17880 11286 17908 11648
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10554 17908 11018
rect 17972 10742 18000 11154
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17880 10526 18000 10554
rect 17972 9654 18000 10526
rect 18064 10470 18092 11086
rect 18156 11014 18184 15263
rect 18524 14958 18552 15302
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 13938 18276 14214
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18248 13258 18276 13874
rect 18524 13870 18552 13942
rect 18512 13864 18564 13870
rect 18510 13832 18512 13841
rect 18564 13832 18566 13841
rect 18510 13767 18566 13776
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18340 12753 18368 13670
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18326 12744 18382 12753
rect 18326 12679 18382 12688
rect 18340 12646 18368 12679
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18234 12336 18290 12345
rect 18234 12271 18290 12280
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18142 10704 18198 10713
rect 18142 10639 18198 10648
rect 18156 10606 18184 10639
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18052 10464 18104 10470
rect 18156 10441 18184 10542
rect 18052 10406 18104 10412
rect 18142 10432 18198 10441
rect 18142 10367 18198 10376
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17774 9480 17830 9489
rect 17774 9415 17830 9424
rect 17788 9330 17816 9415
rect 18052 9376 18104 9382
rect 17788 9302 18000 9330
rect 18052 9318 18104 9324
rect 17972 7954 18000 9302
rect 18064 9110 18092 9318
rect 18142 9208 18198 9217
rect 18142 9143 18198 9152
rect 18156 9110 18184 9143
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18064 8634 18092 9046
rect 18156 8634 18184 9046
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17776 7404 17828 7410
rect 17696 7364 17776 7392
rect 17776 7346 17828 7352
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17696 4826 17724 7210
rect 17788 7206 17816 7346
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17788 6662 17816 7142
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17880 5914 17908 6802
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17972 5273 18000 7142
rect 18064 6662 18092 7278
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 18064 4593 18092 6598
rect 18248 5930 18276 12271
rect 18524 11098 18552 12854
rect 18616 12306 18644 17274
rect 18708 15994 18736 19887
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18892 16697 18920 16934
rect 19076 16794 19104 17478
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 18878 16688 18934 16697
rect 18878 16623 18934 16632
rect 18878 16552 18934 16561
rect 18878 16487 18934 16496
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18800 16114 18828 16390
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18708 15966 18828 15994
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18616 11898 18644 12242
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18328 11076 18380 11082
rect 18524 11070 18644 11098
rect 18328 11018 18380 11024
rect 18340 9518 18368 11018
rect 18616 11014 18644 11070
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18616 10849 18644 10950
rect 18602 10840 18658 10849
rect 18602 10775 18658 10784
rect 18616 10266 18644 10775
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18340 9178 18368 9454
rect 18432 9178 18460 9862
rect 18510 9616 18566 9625
rect 18510 9551 18512 9560
rect 18564 9551 18566 9560
rect 18512 9522 18564 9528
rect 18510 9480 18566 9489
rect 18510 9415 18566 9424
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18432 8430 18460 9114
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18524 6662 18552 9415
rect 18616 8974 18644 10202
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18616 8634 18644 8910
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18602 7848 18658 7857
rect 18602 7783 18604 7792
rect 18656 7783 18658 7792
rect 18604 7754 18656 7760
rect 18616 7274 18644 7754
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18512 6656 18564 6662
rect 18604 6656 18656 6662
rect 18512 6598 18564 6604
rect 18602 6624 18604 6633
rect 18656 6624 18658 6633
rect 18524 6254 18552 6598
rect 18602 6559 18658 6568
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18248 5902 18460 5930
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18248 5234 18276 5714
rect 18328 5704 18380 5710
rect 18326 5672 18328 5681
rect 18380 5672 18382 5681
rect 18326 5607 18382 5616
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18248 4826 18276 5170
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18050 4584 18106 4593
rect 18050 4519 18106 4528
rect 17590 4312 17646 4321
rect 17590 4247 17646 4256
rect 18248 4214 18276 4762
rect 18236 4208 18288 4214
rect 17590 4176 17646 4185
rect 18236 4150 18288 4156
rect 17590 4111 17646 4120
rect 17132 3606 17184 3612
rect 17314 3632 17370 3641
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 17144 3058 17172 3606
rect 17314 3567 17370 3576
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17420 3194 17448 3470
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16776 1329 16804 2926
rect 17038 2680 17094 2689
rect 17038 2615 17094 2624
rect 17052 2514 17080 2615
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17038 1592 17094 1601
rect 17038 1527 17094 1536
rect 16762 1320 16818 1329
rect 16762 1255 16818 1264
rect 17052 480 17080 1527
rect 17604 480 17632 4111
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 1465 17816 3878
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17774 1456 17830 1465
rect 17774 1391 17830 1400
rect 17972 1193 18000 2246
rect 17958 1184 18014 1193
rect 17958 1119 18014 1128
rect 18064 649 18092 3674
rect 18340 2990 18368 5607
rect 18432 4826 18460 5902
rect 18616 5681 18644 6559
rect 18708 6390 18736 12038
rect 18800 9178 18828 15966
rect 18892 12345 18920 16487
rect 19076 16114 19104 16730
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19076 15178 19104 16050
rect 19260 16046 19288 17478
rect 19352 17134 19380 17682
rect 19340 17128 19392 17134
rect 19338 17096 19340 17105
rect 19392 17096 19394 17105
rect 19338 17031 19394 17040
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 18984 15162 19104 15178
rect 18972 15156 19104 15162
rect 19024 15150 19104 15156
rect 18972 15098 19024 15104
rect 19062 15056 19118 15065
rect 19062 14991 19118 15000
rect 19076 14890 19104 14991
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18878 12336 18934 12345
rect 18878 12271 18934 12280
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18880 9920 18932 9926
rect 18878 9888 18880 9897
rect 18932 9888 18934 9897
rect 18878 9823 18934 9832
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18892 8498 18920 9454
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 7449 18828 7686
rect 18786 7440 18842 7449
rect 18786 7375 18842 7384
rect 18800 6866 18828 7375
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18602 5672 18658 5681
rect 18602 5607 18658 5616
rect 18892 5166 18920 8434
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18432 4049 18460 4762
rect 18892 4282 18920 4762
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18984 4049 19012 11494
rect 19076 11354 19104 12650
rect 19168 12322 19196 15846
rect 19352 15366 19380 16526
rect 19340 15360 19392 15366
rect 19338 15328 19340 15337
rect 19392 15328 19394 15337
rect 19338 15263 19394 15272
rect 19444 14532 19472 18022
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19536 16658 19564 17750
rect 19708 17672 19760 17678
rect 19892 17672 19944 17678
rect 19708 17614 19760 17620
rect 19890 17640 19892 17649
rect 19944 17640 19946 17649
rect 19720 17270 19748 17614
rect 19890 17575 19946 17584
rect 19904 17338 19932 17575
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19708 17264 19760 17270
rect 19996 17241 20024 20182
rect 20074 20159 20130 20168
rect 20810 19272 20866 19281
rect 20810 19207 20866 19216
rect 20720 18216 20772 18222
rect 20640 18164 20720 18170
rect 20640 18158 20772 18164
rect 20640 18142 20760 18158
rect 20074 17912 20130 17921
rect 20074 17847 20130 17856
rect 19708 17206 19760 17212
rect 19982 17232 20038 17241
rect 19982 17167 20038 17176
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19536 15910 19564 16594
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19536 15609 19564 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19522 15600 19578 15609
rect 19522 15535 19578 15544
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19260 14504 19472 14532
rect 19260 14074 19288 14504
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19260 13870 19288 14010
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19352 13716 19380 14282
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13734 19472 13806
rect 19260 13688 19380 13716
rect 19432 13728 19484 13734
rect 19260 13530 19288 13688
rect 19432 13670 19484 13676
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19432 13456 19484 13462
rect 19338 13424 19394 13433
rect 19432 13398 19484 13404
rect 19536 13410 19564 15098
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19628 14074 19656 14418
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 13462 20024 16390
rect 20088 15706 20116 17847
rect 20640 17814 20668 18142
rect 20628 17808 20680 17814
rect 20628 17750 20680 17756
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20364 16998 20392 17478
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20088 14414 20116 14962
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20088 13530 20116 14350
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20180 13462 20208 16934
rect 20364 16794 20392 16934
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20456 16658 20484 17138
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20260 15972 20312 15978
rect 20260 15914 20312 15920
rect 20272 15366 20300 15914
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20272 15094 20300 15302
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20272 14550 20300 15030
rect 20364 14822 20392 15506
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20260 14544 20312 14550
rect 20260 14486 20312 14492
rect 20272 13938 20300 14486
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 19984 13456 20036 13462
rect 19338 13359 19340 13368
rect 19392 13359 19394 13368
rect 19340 13330 19392 13336
rect 19352 12986 19380 13330
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19444 12442 19472 13398
rect 19536 13382 19656 13410
rect 19984 13398 20036 13404
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 19628 12986 19656 13382
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 19982 13152 20038 13161
rect 19982 13087 20038 13096
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19168 12306 19380 12322
rect 19168 12300 19392 12306
rect 19168 12294 19340 12300
rect 19340 12242 19392 12248
rect 19444 11914 19472 12378
rect 19522 12336 19578 12345
rect 19522 12271 19578 12280
rect 19352 11898 19472 11914
rect 19340 11892 19472 11898
rect 19392 11886 19472 11892
rect 19340 11834 19392 11840
rect 19444 11694 19472 11886
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19062 10296 19118 10305
rect 19062 10231 19118 10240
rect 19076 9110 19104 10231
rect 19352 10062 19380 10406
rect 19430 10296 19486 10305
rect 19536 10266 19564 12271
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19430 10231 19486 10240
rect 19524 10260 19576 10266
rect 19444 10198 19472 10231
rect 19524 10202 19576 10208
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9761 19288 9862
rect 19246 9752 19302 9761
rect 19536 9722 19564 10202
rect 19246 9687 19302 9696
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 19340 9036 19392 9042
rect 19260 8996 19340 9024
rect 19062 8936 19118 8945
rect 19062 8871 19118 8880
rect 19076 8090 19104 8871
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19156 8084 19208 8090
rect 19156 8026 19208 8032
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19076 5846 19104 7890
rect 19168 7546 19196 8026
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19260 7426 19288 8996
rect 19340 8978 19392 8984
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 7954 19380 8298
rect 19536 8022 19564 8910
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 8090 20024 13087
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 20088 12374 20116 12854
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 20088 11626 20116 12310
rect 20180 12209 20208 13262
rect 20166 12200 20222 12209
rect 20166 12135 20222 12144
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 20260 11280 20312 11286
rect 20166 11248 20222 11257
rect 20260 11222 20312 11228
rect 20364 11234 20392 14758
rect 20456 12782 20484 16594
rect 20548 14906 20576 17206
rect 20640 17134 20668 17478
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20640 16794 20668 17070
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20548 14878 20668 14906
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14618 20576 14758
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20548 13569 20576 13806
rect 20534 13560 20590 13569
rect 20534 13495 20590 13504
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12442 20484 12718
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20456 11898 20484 12378
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20640 11830 20668 14878
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20732 12714 20760 14214
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20732 11354 20760 12174
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20824 11234 20852 19207
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 21546 18184 21602 18193
rect 22388 18154 22416 18770
rect 21546 18119 21602 18128
rect 22376 18148 22428 18154
rect 21560 18086 21588 18119
rect 22376 18090 22428 18096
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 21270 17776 21326 17785
rect 21270 17711 21272 17720
rect 21324 17711 21326 17720
rect 22468 17740 22520 17746
rect 21272 17682 21324 17688
rect 22468 17682 22520 17688
rect 20994 17504 21050 17513
rect 20994 17439 21050 17448
rect 21008 17066 21036 17439
rect 21284 17338 21312 17682
rect 22282 17640 22338 17649
rect 22282 17575 22338 17584
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21928 17202 21956 17478
rect 21916 17196 21968 17202
rect 21916 17138 21968 17144
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16590 20944 16934
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20916 16454 20944 16526
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20902 16008 20958 16017
rect 20902 15943 20958 15952
rect 20916 14482 20944 15943
rect 21008 15450 21036 17002
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21270 16688 21326 16697
rect 21270 16623 21272 16632
rect 21324 16623 21326 16632
rect 21272 16594 21324 16600
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21100 15570 21128 15982
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21192 15586 21220 15846
rect 21284 15706 21312 16594
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21192 15570 21312 15586
rect 21088 15564 21140 15570
rect 21192 15564 21324 15570
rect 21192 15558 21272 15564
rect 21088 15506 21140 15512
rect 21272 15506 21324 15512
rect 21008 15422 21220 15450
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20916 14074 20944 14418
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20902 13696 20958 13705
rect 20902 13631 20958 13640
rect 20916 13530 20944 13631
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20904 13320 20956 13326
rect 21008 13297 21036 14826
rect 20904 13262 20956 13268
rect 20994 13288 21050 13297
rect 20916 12442 20944 13262
rect 20994 13223 21050 13232
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20166 11183 20222 11192
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 20088 10810 20116 10950
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 20180 9058 20208 11183
rect 20272 10062 20300 11222
rect 20364 11206 20484 11234
rect 20824 11206 21036 11234
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 20272 9178 20300 9386
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20088 9030 20208 9058
rect 20272 9042 20300 9114
rect 20260 9036 20312 9042
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19338 7848 19394 7857
rect 19338 7783 19394 7792
rect 19432 7812 19484 7818
rect 19168 7398 19288 7426
rect 19168 6798 19196 7398
rect 19352 7177 19380 7783
rect 19432 7754 19484 7760
rect 19444 7206 19472 7754
rect 19536 7546 19564 7958
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19432 7200 19484 7206
rect 19338 7168 19394 7177
rect 19432 7142 19484 7148
rect 19338 7103 19394 7112
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19260 6458 19288 6802
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19352 6118 19380 6598
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5914 19380 6054
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19340 5568 19392 5574
rect 19260 5528 19340 5556
rect 19260 5098 19288 5528
rect 19340 5510 19392 5516
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19340 5024 19392 5030
rect 19338 4992 19340 5001
rect 19392 4992 19394 5001
rect 19338 4927 19394 4936
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 18418 4040 18474 4049
rect 18418 3975 18474 3984
rect 18970 4040 19026 4049
rect 18970 3975 19026 3984
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18524 3738 18552 3878
rect 19076 3738 19104 4422
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19168 3466 19196 4558
rect 19260 4026 19288 4626
rect 19260 3998 19380 4026
rect 19352 3942 19380 3998
rect 19340 3936 19392 3942
rect 19338 3904 19340 3913
rect 19392 3904 19394 3913
rect 19338 3839 19394 3848
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18524 2990 18552 3334
rect 18708 3097 18736 3334
rect 19352 3194 19380 3470
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 18694 3088 18750 3097
rect 18694 3023 18750 3032
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18694 2952 18750 2961
rect 18694 2887 18750 2896
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18616 2009 18644 2246
rect 18602 2000 18658 2009
rect 18602 1935 18658 1944
rect 18142 776 18198 785
rect 18142 711 18198 720
rect 18050 640 18106 649
rect 18050 575 18106 584
rect 18156 480 18184 711
rect 18708 480 18736 2887
rect 19444 2281 19472 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20088 6440 20116 9030
rect 20260 8978 20312 8984
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20180 8090 20208 8910
rect 20272 8634 20300 8978
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20180 6934 20208 8026
rect 20168 6928 20220 6934
rect 20168 6870 20220 6876
rect 20088 6412 20208 6440
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19536 5914 19564 6122
rect 20088 6118 20116 6258
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 20088 5030 20116 6054
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19892 4480 19944 4486
rect 19890 4448 19892 4457
rect 19944 4448 19946 4457
rect 19890 4383 19946 4392
rect 19904 4146 19932 4383
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19522 3496 19578 3505
rect 19522 3431 19578 3440
rect 19430 2272 19486 2281
rect 19430 2207 19486 2216
rect 19246 1864 19302 1873
rect 19246 1799 19302 1808
rect 19260 480 19288 1799
rect 19536 1442 19564 3431
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2145 20024 3946
rect 20180 3777 20208 6412
rect 20364 6361 20392 11086
rect 20456 7993 20484 11206
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20442 7984 20498 7993
rect 20442 7919 20498 7928
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20456 7546 20484 7822
rect 20444 7540 20496 7546
rect 20444 7482 20496 7488
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20456 7002 20484 7346
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20350 6352 20406 6361
rect 20350 6287 20406 6296
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20272 4214 20300 4422
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 20350 4040 20406 4049
rect 20350 3975 20406 3984
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20166 3768 20222 3777
rect 20166 3703 20222 3712
rect 20180 3398 20208 3429
rect 20168 3392 20220 3398
rect 20166 3360 20168 3369
rect 20220 3360 20222 3369
rect 20166 3295 20222 3304
rect 20180 2650 20208 3295
rect 20272 3233 20300 3878
rect 20258 3224 20314 3233
rect 20258 3159 20314 3168
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19982 2136 20038 2145
rect 19982 2071 20038 2080
rect 19536 1414 19840 1442
rect 19812 480 19840 1414
rect 20364 480 20392 3975
rect 20548 3618 20576 11018
rect 20824 10470 20852 11086
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20732 8838 20760 9930
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 20640 8090 20668 8502
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20640 7342 20668 8026
rect 20732 8022 20760 8774
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20732 7002 20760 7958
rect 20824 7274 20852 10406
rect 20916 9625 20944 11018
rect 21008 10146 21036 11206
rect 21086 10568 21142 10577
rect 21086 10503 21088 10512
rect 21140 10503 21142 10512
rect 21088 10474 21140 10480
rect 21008 10118 21128 10146
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 20902 9616 20958 9625
rect 20902 9551 20958 9560
rect 21008 9500 21036 9998
rect 20916 9472 21036 9500
rect 20812 7268 20864 7274
rect 20916 7256 20944 9472
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 21008 8974 21036 9318
rect 21100 9217 21128 10118
rect 21086 9208 21142 9217
rect 21086 9143 21142 9152
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 21100 8090 21128 8978
rect 21192 8809 21220 15422
rect 21284 15026 21312 15506
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21284 11354 21312 12650
rect 21376 12238 21404 16934
rect 21836 16794 21864 16934
rect 21928 16833 21956 17138
rect 21914 16824 21970 16833
rect 21824 16788 21876 16794
rect 21914 16759 21970 16768
rect 21824 16730 21876 16736
rect 22296 16726 22324 17575
rect 22480 16980 22508 17682
rect 22558 17640 22614 17649
rect 22558 17575 22560 17584
rect 22612 17575 22614 17584
rect 22560 17546 22612 17552
rect 22560 16992 22612 16998
rect 22480 16952 22560 16980
rect 22560 16934 22612 16940
rect 22572 16726 22600 16934
rect 22284 16720 22336 16726
rect 22560 16720 22612 16726
rect 22284 16662 22336 16668
rect 22466 16688 22522 16697
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21560 16153 21588 16594
rect 22296 16522 22324 16662
rect 22560 16662 22612 16668
rect 22466 16623 22522 16632
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22480 16538 22508 16623
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22388 16250 22416 16526
rect 22480 16510 22600 16538
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 21546 16144 21602 16153
rect 21546 16079 21548 16088
rect 21600 16079 21602 16088
rect 21548 16050 21600 16056
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14657 21496 14758
rect 21454 14648 21510 14657
rect 21454 14583 21456 14592
rect 21508 14583 21510 14592
rect 21456 14554 21508 14560
rect 21468 14074 21496 14554
rect 21928 14521 21956 14826
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 21914 14512 21970 14521
rect 21914 14447 21970 14456
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21652 14074 21680 14350
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 22020 13938 22048 14758
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21916 13456 21968 13462
rect 21916 13398 21968 13404
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21652 12646 21680 13262
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21468 11898 21496 12174
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21284 10810 21312 11290
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 21270 9752 21326 9761
rect 21270 9687 21326 9696
rect 21284 9178 21312 9687
rect 21456 9512 21508 9518
rect 21456 9454 21508 9460
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21364 8968 21416 8974
rect 21362 8936 21364 8945
rect 21416 8936 21418 8945
rect 21362 8871 21418 8880
rect 21272 8832 21324 8838
rect 21178 8800 21234 8809
rect 21272 8774 21324 8780
rect 21178 8735 21234 8744
rect 21192 8090 21220 8735
rect 21284 8498 21312 8774
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21100 7410 21128 8026
rect 21178 7984 21234 7993
rect 21178 7919 21234 7928
rect 21192 7886 21220 7919
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21192 7478 21220 7822
rect 21284 7546 21312 8434
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 20916 7228 21128 7256
rect 20812 7210 20864 7216
rect 20720 6996 20772 7002
rect 20772 6956 20852 6984
rect 20720 6938 20772 6944
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20732 6118 20760 6666
rect 20824 6390 20852 6956
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 5846 20760 6054
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20732 5574 20760 5782
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 4826 20760 5510
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20720 4616 20772 4622
rect 20640 4564 20720 4570
rect 20640 4558 20772 4564
rect 20640 4542 20760 4558
rect 20824 4554 20852 5714
rect 20812 4548 20864 4554
rect 20640 3942 20668 4542
rect 20812 4490 20864 4496
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20732 3754 20760 4422
rect 20916 4146 20944 6802
rect 21008 6458 21036 6802
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20994 5944 21050 5953
rect 21100 5930 21128 7228
rect 21270 6896 21326 6905
rect 21270 6831 21326 6840
rect 21050 5902 21128 5930
rect 20994 5879 21050 5888
rect 21008 5681 21036 5879
rect 20994 5672 21050 5681
rect 20994 5607 21050 5616
rect 21284 4826 21312 6831
rect 21376 6633 21404 8570
rect 21468 7546 21496 9454
rect 21560 9382 21588 10134
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21560 7585 21588 9318
rect 21652 8401 21680 12582
rect 21928 12442 21956 13398
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 21914 11656 21970 11665
rect 21914 11591 21970 11600
rect 21928 11558 21956 11591
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 22020 11354 22048 11698
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 21916 11280 21968 11286
rect 21916 11222 21968 11228
rect 21928 10674 21956 11222
rect 22020 11121 22048 11290
rect 22006 11112 22062 11121
rect 22006 11047 22062 11056
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21638 8392 21694 8401
rect 21638 8327 21694 8336
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21546 7576 21602 7585
rect 21456 7540 21508 7546
rect 21652 7546 21680 8026
rect 21546 7511 21602 7520
rect 21640 7540 21692 7546
rect 21456 7482 21508 7488
rect 21640 7482 21692 7488
rect 21468 7002 21496 7482
rect 21546 7440 21602 7449
rect 21546 7375 21602 7384
rect 21560 7342 21588 7375
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21468 6905 21496 6938
rect 21454 6896 21510 6905
rect 21454 6831 21510 6840
rect 21362 6624 21418 6633
rect 21362 6559 21418 6568
rect 21744 6254 21772 9862
rect 21836 6322 21864 10406
rect 21928 10266 21956 10610
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21928 10062 21956 10202
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 22020 9874 22048 10066
rect 21928 9846 22048 9874
rect 21928 9382 21956 9846
rect 21916 9376 21968 9382
rect 22112 9353 22140 15302
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22296 13394 22324 13670
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 21916 9318 21968 9324
rect 22098 9344 22154 9353
rect 21928 8634 21956 9318
rect 22098 9279 22154 9288
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 21914 8392 21970 8401
rect 21914 8327 21970 8336
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21836 5914 21864 6258
rect 21824 5908 21876 5914
rect 21824 5850 21876 5856
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21376 5370 21404 5646
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21744 4865 21772 5034
rect 21730 4856 21786 4865
rect 21272 4820 21324 4826
rect 21730 4791 21786 4800
rect 21272 4762 21324 4768
rect 21284 4282 21312 4762
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21284 4162 21312 4218
rect 20904 4140 20956 4146
rect 21192 4134 21312 4162
rect 20956 4100 21036 4128
rect 20904 4082 20956 4088
rect 20640 3738 20760 3754
rect 20628 3732 20760 3738
rect 20680 3726 20760 3732
rect 20628 3674 20680 3680
rect 20548 3590 20944 3618
rect 21008 3602 21036 4100
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20456 2922 20484 3130
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20456 2446 20484 2858
rect 20626 2816 20682 2825
rect 20626 2751 20682 2760
rect 20640 2650 20668 2751
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 20916 480 20944 3590
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21008 2990 21036 3538
rect 21192 3505 21220 4134
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 21284 3738 21312 4014
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21178 3496 21234 3505
rect 21468 3466 21496 4558
rect 21824 4072 21876 4078
rect 21928 4060 21956 8327
rect 22112 8090 22140 9114
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22006 7984 22062 7993
rect 22006 7919 22062 7928
rect 22020 7546 22048 7919
rect 22098 7848 22154 7857
rect 22098 7783 22154 7792
rect 22112 7750 22140 7783
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22020 6118 22048 6394
rect 22112 6254 22140 6394
rect 22100 6248 22152 6254
rect 22100 6190 22152 6196
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22204 5137 22232 13262
rect 22388 12850 22416 16186
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22480 14618 22508 14962
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22480 13734 22508 13874
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22480 12986 22508 13670
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22296 10810 22324 11630
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22388 10713 22416 12038
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22480 11082 22508 11834
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22374 10704 22430 10713
rect 22374 10639 22430 10648
rect 22388 10198 22416 10639
rect 22376 10192 22428 10198
rect 22376 10134 22428 10140
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22296 9518 22324 9862
rect 22284 9512 22336 9518
rect 22468 9512 22520 9518
rect 22284 9454 22336 9460
rect 22466 9480 22468 9489
rect 22520 9480 22522 9489
rect 22466 9415 22522 9424
rect 22282 9208 22338 9217
rect 22282 9143 22338 9152
rect 22296 8430 22324 9143
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22572 8022 22600 16510
rect 22664 16153 22692 18022
rect 22756 16250 22784 23695
rect 23478 22536 23534 22545
rect 23478 22471 23534 22480
rect 23492 20754 23520 22471
rect 23860 21162 23888 24239
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23308 20726 23520 20754
rect 23768 21134 23888 21162
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22650 16144 22706 16153
rect 22650 16079 22706 16088
rect 22848 15366 22876 16594
rect 22940 16561 22968 18158
rect 22926 16552 22982 16561
rect 22926 16487 22982 16496
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22664 14482 22692 14962
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22756 14414 22784 14486
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22664 13530 22692 13874
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22756 13326 22784 14350
rect 23032 14074 23060 19110
rect 23204 14952 23256 14958
rect 23202 14920 23204 14929
rect 23256 14920 23258 14929
rect 23202 14855 23258 14864
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23032 13870 23060 14010
rect 23020 13864 23072 13870
rect 23020 13806 23072 13812
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22756 12374 22784 13262
rect 23032 12986 23060 13330
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 22756 12170 22784 12310
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22744 11552 22796 11558
rect 22848 11540 22876 12174
rect 22928 12164 22980 12170
rect 22928 12106 22980 12112
rect 22940 11694 22968 12106
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22796 11512 22876 11540
rect 22744 11494 22796 11500
rect 22664 11014 22692 11494
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22664 10266 22692 10950
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22756 8430 22784 11494
rect 22940 11218 22968 11630
rect 22928 11212 22980 11218
rect 22928 11154 22980 11160
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22744 8424 22796 8430
rect 22744 8366 22796 8372
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22664 7954 22692 8230
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22664 7410 22692 7890
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22388 7002 22416 7210
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 22284 6656 22336 6662
rect 22480 6610 22508 7142
rect 22664 6934 22692 7346
rect 22652 6928 22704 6934
rect 22652 6870 22704 6876
rect 22284 6598 22336 6604
rect 22190 5128 22246 5137
rect 22296 5098 22324 6598
rect 22388 6582 22508 6610
rect 22388 6118 22416 6582
rect 22466 6488 22522 6497
rect 22466 6423 22522 6432
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22388 5914 22416 6054
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22480 5778 22508 6423
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22742 6352 22798 6361
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 22664 5370 22692 6326
rect 22742 6287 22798 6296
rect 22756 5846 22784 6287
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22848 5681 22876 10746
rect 22834 5672 22890 5681
rect 22834 5607 22890 5616
rect 22742 5536 22798 5545
rect 22742 5471 22798 5480
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22190 5063 22246 5072
rect 22284 5092 22336 5098
rect 22284 5034 22336 5040
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 21876 4032 21956 4060
rect 21824 4014 21876 4020
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21546 3632 21602 3641
rect 21928 3602 21956 3878
rect 22098 3768 22154 3777
rect 22098 3703 22154 3712
rect 21546 3567 21602 3576
rect 21916 3596 21968 3602
rect 21178 3431 21234 3440
rect 21456 3460 21508 3466
rect 21456 3402 21508 3408
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21270 2680 21326 2689
rect 21270 2615 21272 2624
rect 21324 2615 21326 2624
rect 21272 2586 21324 2592
rect 21560 480 21588 3567
rect 21916 3538 21968 3544
rect 21928 3194 21956 3538
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21638 3088 21694 3097
rect 21638 3023 21694 3032
rect 21652 2650 21680 3023
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21744 2446 21772 2586
rect 22020 2446 22048 3130
rect 21732 2440 21784 2446
rect 21732 2382 21784 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 22112 480 22140 3703
rect 22204 3602 22232 4966
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22296 3194 22324 3946
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22480 2825 22508 4422
rect 22652 3460 22704 3466
rect 22652 3402 22704 3408
rect 22664 3126 22692 3402
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22466 2816 22522 2825
rect 22466 2751 22522 2760
rect 22664 2650 22692 3062
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22756 2378 22784 5471
rect 22940 5030 22968 11018
rect 23032 10266 23060 12582
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23032 9722 23060 10202
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 23124 4826 23152 12038
rect 23216 11898 23244 12242
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23216 10470 23244 11154
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23216 10062 23244 10406
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23216 9178 23244 9998
rect 23308 9654 23336 20726
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23388 18148 23440 18154
rect 23388 18090 23440 18096
rect 23400 14804 23428 18090
rect 23492 18086 23520 18770
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23492 15065 23520 18022
rect 23768 17882 23796 21134
rect 23952 21078 23980 21422
rect 23940 21072 23992 21078
rect 23940 21014 23992 21020
rect 23848 21004 23900 21010
rect 23848 20946 23900 20952
rect 23860 20262 23888 20946
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23860 19961 23888 20198
rect 23846 19952 23902 19961
rect 23846 19887 23902 19896
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23860 19174 23888 19722
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23860 18290 23888 19110
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23860 17762 23888 18022
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23768 17734 23888 17762
rect 23584 16998 23612 17682
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23478 15056 23534 15065
rect 23478 14991 23534 15000
rect 23400 14776 23520 14804
rect 23492 14618 23520 14776
rect 23480 14612 23532 14618
rect 23480 14554 23532 14560
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23400 13530 23428 14418
rect 23478 14104 23534 14113
rect 23478 14039 23480 14048
rect 23532 14039 23534 14048
rect 23480 14010 23532 14016
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23480 12844 23532 12850
rect 23480 12786 23532 12792
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23400 11286 23428 12174
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23492 10130 23520 12786
rect 23480 10124 23532 10130
rect 23480 10066 23532 10072
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23400 9217 23428 9590
rect 23492 9382 23520 10066
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 23386 9208 23442 9217
rect 23204 9172 23256 9178
rect 23386 9143 23442 9152
rect 23204 9114 23256 9120
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23400 8294 23428 8978
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23492 8090 23520 9318
rect 23584 8945 23612 16934
rect 23662 16824 23718 16833
rect 23662 16759 23718 16768
rect 23676 16250 23704 16759
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23676 14550 23704 15302
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 23676 13530 23704 13670
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23768 13410 23796 17734
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23676 13382 23796 13410
rect 23676 11121 23704 13382
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23768 12238 23796 12854
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23754 11792 23810 11801
rect 23754 11727 23810 11736
rect 23662 11112 23718 11121
rect 23662 11047 23718 11056
rect 23664 10464 23716 10470
rect 23664 10406 23716 10412
rect 23676 9926 23704 10406
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23676 9586 23704 9862
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23676 9110 23704 9522
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23570 8936 23626 8945
rect 23570 8871 23626 8880
rect 23676 8498 23704 9046
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23296 8016 23348 8022
rect 23296 7958 23348 7964
rect 23478 7984 23534 7993
rect 23308 5817 23336 7958
rect 23478 7919 23480 7928
rect 23532 7919 23534 7928
rect 23480 7890 23532 7896
rect 23676 7886 23704 8230
rect 23768 8022 23796 11727
rect 23756 8016 23808 8022
rect 23756 7958 23808 7964
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23386 6896 23442 6905
rect 23492 6866 23520 7754
rect 23676 7546 23704 7822
rect 23756 7812 23808 7818
rect 23756 7754 23808 7760
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23768 7002 23796 7754
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23386 6831 23442 6840
rect 23480 6860 23532 6866
rect 23400 6798 23428 6831
rect 23480 6802 23532 6808
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23294 5808 23350 5817
rect 23294 5743 23350 5752
rect 23294 5536 23350 5545
rect 23294 5471 23350 5480
rect 23308 4865 23336 5471
rect 23400 5216 23428 6734
rect 23492 6458 23520 6802
rect 23676 6662 23704 6802
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23676 6322 23704 6598
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 5710 23704 6258
rect 23860 5794 23888 17478
rect 23952 14770 23980 19790
rect 24044 16794 24072 24942
rect 24122 24848 24178 24857
rect 24122 24783 24178 24792
rect 24136 17338 24164 24783
rect 24228 24177 24256 25214
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24214 24168 24270 24177
rect 24214 24103 24270 24112
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23866 24808 25327
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24584 23656 24636 23662
rect 24582 23624 24584 23633
rect 24636 23624 24638 23633
rect 24582 23559 24638 23568
rect 24766 23216 24822 23225
rect 24766 23151 24822 23160
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24674 21992 24730 22001
rect 24674 21927 24730 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 21927
rect 24780 21690 24808 23151
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24766 21448 24822 21457
rect 24766 21383 24822 21392
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24674 20360 24730 20369
rect 24596 20233 24624 20334
rect 24674 20295 24730 20304
rect 24582 20224 24638 20233
rect 24582 20159 24638 20168
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24214 19408 24270 19417
rect 24214 19343 24270 19352
rect 24228 17921 24256 19343
rect 24584 19304 24636 19310
rect 24582 19272 24584 19281
rect 24636 19272 24638 19281
rect 24582 19207 24638 19216
rect 24688 18970 24716 20295
rect 24780 20058 24808 21383
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24768 19168 24820 19174
rect 24766 19136 24768 19145
rect 24820 19136 24822 19145
rect 24766 19071 24822 19080
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24582 18864 24638 18873
rect 24582 18799 24584 18808
rect 24636 18799 24638 18808
rect 24584 18770 24636 18776
rect 24596 18714 24624 18770
rect 24596 18686 24716 18714
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24688 18426 24716 18686
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24492 18080 24544 18086
rect 24490 18048 24492 18057
rect 24544 18048 24546 18057
rect 24490 17983 24546 17992
rect 24214 17912 24270 17921
rect 24214 17847 24270 17856
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 24044 16114 24072 16730
rect 24122 16688 24178 16697
rect 24122 16623 24124 16632
rect 24176 16623 24178 16632
rect 24124 16594 24176 16600
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 24228 16114 24256 16458
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16130 24716 18226
rect 24780 16833 24808 18566
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25148 16998 25176 17682
rect 25136 16992 25188 16998
rect 25134 16960 25136 16969
rect 25188 16960 25190 16969
rect 25134 16895 25190 16904
rect 24766 16824 24822 16833
rect 24766 16759 24822 16768
rect 25134 16552 25190 16561
rect 25134 16487 25190 16496
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24596 16102 24716 16130
rect 24044 15858 24072 16050
rect 24044 15830 24164 15858
rect 24030 15736 24086 15745
rect 24030 15671 24086 15680
rect 24044 14890 24072 15671
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 23952 14742 24072 14770
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 23952 12442 23980 14554
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 23940 12300 23992 12306
rect 23940 12242 23992 12248
rect 23952 11937 23980 12242
rect 23938 11928 23994 11937
rect 23938 11863 23940 11872
rect 23992 11863 23994 11872
rect 23940 11834 23992 11840
rect 24044 10810 24072 14742
rect 24136 14362 24164 15830
rect 24216 15632 24268 15638
rect 24216 15574 24268 15580
rect 24228 15026 24256 15574
rect 24596 15473 24624 16102
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24582 15464 24638 15473
rect 24582 15399 24638 15408
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24136 14334 24256 14362
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 13938 24164 14214
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24136 13462 24164 13874
rect 24124 13456 24176 13462
rect 24124 13398 24176 13404
rect 24136 12986 24164 13398
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24228 12730 24256 14334
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12968 24716 15914
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24860 15360 24912 15366
rect 24860 15302 24912 15308
rect 24766 15192 24822 15201
rect 24766 15127 24822 15136
rect 24780 14958 24808 15127
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24872 14498 24900 15302
rect 24780 14482 24900 14498
rect 24768 14476 24900 14482
rect 24820 14470 24900 14476
rect 24768 14418 24820 14424
rect 24768 14068 24820 14074
rect 24872 14056 24900 14470
rect 24820 14028 24900 14056
rect 24768 14010 24820 14016
rect 24964 13954 24992 15846
rect 24872 13926 24992 13954
rect 25148 13938 25176 16487
rect 25424 16250 25452 27095
rect 25686 26616 25742 26625
rect 25686 26551 25742 26560
rect 25502 26072 25558 26081
rect 25502 26007 25558 26016
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25410 15056 25466 15065
rect 25410 14991 25412 15000
rect 25464 14991 25466 15000
rect 25412 14962 25464 14968
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25240 14006 25268 14418
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25136 13932 25188 13938
rect 24872 13870 24900 13926
rect 25136 13874 25188 13880
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 25044 13864 25096 13870
rect 25240 13841 25268 13942
rect 25044 13806 25096 13812
rect 25226 13832 25282 13841
rect 25056 13705 25084 13806
rect 25226 13767 25282 13776
rect 25042 13696 25098 13705
rect 25042 13631 25098 13640
rect 24858 13424 24914 13433
rect 24858 13359 24914 13368
rect 24136 12702 24256 12730
rect 24596 12940 24716 12968
rect 24136 12646 24164 12702
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 23940 9716 23992 9722
rect 23940 9658 23992 9664
rect 23952 7546 23980 9658
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23952 5914 23980 6122
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23860 5766 23980 5794
rect 24044 5778 24072 9930
rect 24136 6390 24164 12378
rect 24596 12374 24624 12940
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24308 10600 24360 10606
rect 24688 10554 24716 12582
rect 24872 12442 24900 13359
rect 25136 13184 25188 13190
rect 25136 13126 25188 13132
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 10674 24808 12038
rect 24872 11354 24900 12378
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24308 10542 24360 10548
rect 24320 10470 24348 10542
rect 24596 10526 24716 10554
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24320 10266 24348 10406
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24320 9908 24348 10202
rect 24596 9994 24624 10526
rect 24676 10464 24728 10470
rect 24728 10424 24808 10452
rect 24676 10406 24728 10412
rect 24584 9988 24636 9994
rect 24584 9930 24636 9936
rect 24228 9880 24348 9908
rect 24676 9920 24728 9926
rect 24228 9518 24256 9880
rect 24676 9862 24728 9868
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24228 7449 24256 7686
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24214 7440 24270 7449
rect 24214 7375 24270 7384
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24228 6322 24256 6802
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24492 6384 24544 6390
rect 24492 6326 24544 6332
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24124 6248 24176 6254
rect 24124 6190 24176 6196
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 23846 5672 23902 5681
rect 23676 5386 23704 5646
rect 23846 5607 23902 5616
rect 23676 5358 23796 5386
rect 23480 5228 23532 5234
rect 23400 5188 23480 5216
rect 23480 5170 23532 5176
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23294 4856 23350 4865
rect 23112 4820 23164 4826
rect 23294 4791 23350 4800
rect 23112 4762 23164 4768
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23032 4282 23060 4558
rect 23202 4312 23258 4321
rect 23020 4276 23072 4282
rect 23202 4247 23258 4256
rect 23020 4218 23072 4224
rect 23032 3738 23060 4218
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23032 3194 23060 3674
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 22744 2372 22796 2378
rect 22744 2314 22796 2320
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23032 1737 23060 2246
rect 23018 1728 23074 1737
rect 23018 1663 23074 1672
rect 22572 598 22692 626
rect 10966 368 11022 377
rect 10966 303 11022 312
rect 11426 0 11482 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 17038 0 17094 480
rect 17590 0 17646 480
rect 18142 0 18198 480
rect 18694 0 18750 480
rect 19246 0 19302 480
rect 19798 0 19854 480
rect 20350 0 20406 480
rect 20902 0 20958 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22572 105 22600 598
rect 22664 480 22692 598
rect 23216 480 23244 4247
rect 23308 3777 23336 4791
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23400 4570 23428 4626
rect 23400 4542 23520 4570
rect 23294 3768 23350 3777
rect 23492 3738 23520 4542
rect 23676 4146 23704 5170
rect 23768 5098 23796 5358
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 23756 4752 23808 4758
rect 23756 4694 23808 4700
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 23294 3703 23350 3712
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23662 3360 23718 3369
rect 23584 2961 23612 3334
rect 23662 3295 23718 3304
rect 23676 3194 23704 3295
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23664 2984 23716 2990
rect 23570 2952 23626 2961
rect 23664 2926 23716 2932
rect 23570 2887 23626 2896
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 22558 96 22614 105
rect 22558 31 22614 40
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23492 377 23520 2790
rect 23676 2310 23704 2926
rect 23768 2650 23796 4694
rect 23860 4593 23888 5607
rect 23846 4584 23902 4593
rect 23846 4519 23902 4528
rect 23846 4040 23902 4049
rect 23846 3975 23902 3984
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23664 2304 23716 2310
rect 23664 2246 23716 2252
rect 23478 368 23534 377
rect 23478 303 23534 312
rect 23676 241 23704 2246
rect 23860 1442 23888 3975
rect 23952 3670 23980 5766
rect 24032 5772 24084 5778
rect 24032 5714 24084 5720
rect 24136 4826 24164 6190
rect 24228 5846 24256 6258
rect 24216 5840 24268 5846
rect 24216 5782 24268 5788
rect 24320 5658 24348 6326
rect 24504 5681 24532 6326
rect 24688 5914 24716 9862
rect 24780 7290 24808 10424
rect 24964 10062 24992 12854
rect 25148 12238 25176 13126
rect 25136 12232 25188 12238
rect 25056 12192 25136 12220
rect 25056 11626 25084 12192
rect 25136 12174 25188 12180
rect 25226 11656 25282 11665
rect 25044 11620 25096 11626
rect 25226 11591 25282 11600
rect 25044 11562 25096 11568
rect 25056 11354 25084 11562
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25148 10674 25176 11494
rect 25136 10668 25188 10674
rect 25136 10610 25188 10616
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24872 9926 24900 9998
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9722 24900 9862
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24964 9518 24992 9998
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 25056 8838 25084 10066
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24780 7262 24900 7290
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24228 5630 24348 5658
rect 24490 5672 24546 5681
rect 24228 5273 24256 5630
rect 24490 5607 24546 5616
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5714
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24214 5264 24270 5273
rect 24214 5199 24270 5208
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24228 3738 24256 5034
rect 24780 4826 24808 7142
rect 24872 6254 24900 7262
rect 24964 6662 24992 7346
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24872 5302 24900 5646
rect 24860 5296 24912 5302
rect 24860 5238 24912 5244
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24872 4622 24900 5238
rect 24964 5166 24992 6598
rect 25056 6390 25084 8774
rect 25136 7880 25188 7886
rect 25134 7848 25136 7857
rect 25188 7848 25190 7857
rect 25134 7783 25190 7792
rect 25148 7546 25176 7783
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25240 7426 25268 11591
rect 25148 7398 25268 7426
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5953 25084 6054
rect 25042 5944 25098 5953
rect 25042 5879 25044 5888
rect 25096 5879 25098 5888
rect 25044 5850 25096 5856
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24860 4616 24912 4622
rect 24860 4558 24912 4564
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24872 4282 24900 4558
rect 24860 4276 24912 4282
rect 24860 4218 24912 4224
rect 24858 4176 24914 4185
rect 24858 4111 24914 4120
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 23940 3664 23992 3670
rect 23940 3606 23992 3612
rect 24228 2922 24256 3674
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24216 2916 24268 2922
rect 24216 2858 24268 2864
rect 24688 2446 24716 3470
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23768 1414 23888 1442
rect 24780 1426 24808 3606
rect 24308 1420 24360 1426
rect 23768 480 23796 1414
rect 24308 1362 24360 1368
rect 24768 1420 24820 1426
rect 24768 1362 24820 1368
rect 24320 480 24348 1362
rect 24872 480 24900 4111
rect 24964 3942 24992 5102
rect 25056 4826 25084 5850
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 24952 3936 25004 3942
rect 24952 3878 25004 3884
rect 25056 3738 25084 4762
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24964 2854 24992 3538
rect 25148 3058 25176 7398
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 5098 25268 7142
rect 25228 5092 25280 5098
rect 25228 5034 25280 5040
rect 25226 4720 25282 4729
rect 25226 4655 25282 4664
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 25240 2990 25268 4655
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 24952 2848 25004 2854
rect 24952 2790 25004 2796
rect 25228 2848 25280 2854
rect 25332 2825 25360 14894
rect 25516 14618 25544 26007
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25424 12102 25452 12582
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25424 11694 25452 12038
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25424 8090 25452 11086
rect 25608 9704 25636 18022
rect 25700 16794 25728 26551
rect 25964 18692 26016 18698
rect 25964 18634 26016 18640
rect 25688 16788 25740 16794
rect 25688 16730 25740 16736
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25792 15910 25820 16594
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25792 13569 25820 15846
rect 25778 13560 25834 13569
rect 25778 13495 25834 13504
rect 25780 12708 25832 12714
rect 25780 12650 25832 12656
rect 25792 10690 25820 12650
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25884 11558 25912 12038
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25884 10810 25912 11494
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25792 10662 25912 10690
rect 25608 9676 25728 9704
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25412 8084 25464 8090
rect 25412 8026 25464 8032
rect 25424 7546 25452 8026
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25410 6488 25466 6497
rect 25410 6423 25466 6432
rect 25424 6322 25452 6423
rect 25412 6316 25464 6322
rect 25412 6258 25464 6264
rect 25516 6225 25544 9318
rect 25596 9104 25648 9110
rect 25596 9046 25648 9052
rect 25608 8634 25636 9046
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25608 7002 25636 8570
rect 25700 7993 25728 9676
rect 25780 8900 25832 8906
rect 25780 8842 25832 8848
rect 25686 7984 25742 7993
rect 25686 7919 25742 7928
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25700 7546 25728 7822
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25608 6458 25636 6938
rect 25700 6934 25728 7482
rect 25688 6928 25740 6934
rect 25688 6870 25740 6876
rect 25596 6452 25648 6458
rect 25596 6394 25648 6400
rect 25502 6216 25558 6225
rect 25502 6151 25558 6160
rect 25792 4842 25820 8842
rect 25424 4814 25820 4842
rect 25228 2790 25280 2796
rect 25318 2816 25374 2825
rect 25240 1465 25268 2790
rect 25318 2751 25374 2760
rect 25226 1456 25282 1465
rect 25226 1391 25282 1400
rect 25424 480 25452 4814
rect 25686 3768 25742 3777
rect 25686 3703 25742 3712
rect 25700 2650 25728 3703
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 25884 2582 25912 10662
rect 25976 8906 26004 18634
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 25964 8900 26016 8906
rect 25964 8842 26016 8848
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 25976 5370 26004 6394
rect 25964 5364 26016 5370
rect 25964 5306 26016 5312
rect 25976 4282 26004 5306
rect 25964 4276 26016 4282
rect 25964 4218 26016 4224
rect 25976 3738 26004 4218
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 25976 3194 26004 3674
rect 26068 3233 26096 9862
rect 26160 6633 26188 18022
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26146 6624 26202 6633
rect 26146 6559 26202 6568
rect 26054 3224 26110 3233
rect 25964 3188 26016 3194
rect 26054 3159 26110 3168
rect 25964 3130 26016 3136
rect 26056 2916 26108 2922
rect 26056 2858 26108 2864
rect 25872 2576 25924 2582
rect 25594 2544 25650 2553
rect 25594 2479 25596 2488
rect 25648 2479 25650 2488
rect 25870 2544 25872 2553
rect 25924 2544 25926 2553
rect 25870 2479 25926 2488
rect 25596 2450 25648 2456
rect 25964 2372 26016 2378
rect 25964 2314 26016 2320
rect 25976 480 26004 2314
rect 23662 232 23718 241
rect 23662 167 23718 176
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26068 377 26096 2858
rect 26252 921 26280 8366
rect 26238 912 26294 921
rect 26238 847 26294 856
rect 26528 480 26556 17614
rect 27252 8016 27304 8022
rect 27252 7958 27304 7964
rect 27264 2009 27292 7958
rect 27066 2000 27122 2009
rect 27066 1935 27122 1944
rect 27250 2000 27306 2009
rect 27250 1935 27306 1944
rect 27080 480 27108 1935
rect 27618 1728 27674 1737
rect 27618 1663 27674 1672
rect 27632 480 27660 1663
rect 26054 368 26110 377
rect 26054 303 26110 312
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 4066 27648 4122 27704
rect 2686 26560 2742 26616
rect 1582 24928 1638 24984
rect 1490 24384 1546 24440
rect 1398 23840 1454 23896
rect 1582 23160 1638 23216
rect 1490 22072 1546 22128
rect 2502 22380 2504 22400
rect 2504 22380 2556 22400
rect 2556 22380 2558 22400
rect 2502 22344 2558 22380
rect 1582 21528 1638 21584
rect 2042 21292 2044 21312
rect 2044 21292 2096 21312
rect 2096 21292 2098 21312
rect 2042 21256 2098 21292
rect 1582 19896 1638 19952
rect 1582 19352 1638 19408
rect 1582 18672 1638 18728
rect 2042 19116 2044 19136
rect 2044 19116 2096 19136
rect 2096 19116 2098 19136
rect 2042 19080 2098 19116
rect 2410 21120 2466 21176
rect 2594 20984 2650 21040
rect 1490 12008 1546 12064
rect 1490 11056 1546 11112
rect 1398 7948 1454 7984
rect 1398 7928 1400 7948
rect 1400 7928 1452 7948
rect 1452 7928 1454 7948
rect 2226 17992 2282 18048
rect 2410 20204 2412 20224
rect 2412 20204 2464 20224
rect 2464 20204 2466 20224
rect 2410 20168 2466 20204
rect 2410 18944 2466 19000
rect 3330 25472 3386 25528
rect 3790 27104 3846 27160
rect 3514 24792 3570 24848
rect 2594 18400 2650 18456
rect 2318 17176 2374 17232
rect 2226 16904 2282 16960
rect 2318 14592 2374 14648
rect 2962 17040 3018 17096
rect 2226 12860 2228 12880
rect 2228 12860 2280 12880
rect 2280 12860 2282 12880
rect 2226 12824 2282 12860
rect 2226 10104 2282 10160
rect 2410 9988 2466 10024
rect 2410 9968 2412 9988
rect 2412 9968 2464 9988
rect 2464 9968 2466 9988
rect 2410 9696 2466 9752
rect 1582 7248 1638 7304
rect 1398 6860 1454 6896
rect 1398 6840 1400 6860
rect 1400 6840 1452 6860
rect 1452 6840 1454 6860
rect 1766 5772 1822 5808
rect 1766 5752 1768 5772
rect 1768 5752 1820 5772
rect 1820 5752 1822 5772
rect 1766 4820 1822 4856
rect 1766 4800 1768 4820
rect 1768 4800 1820 4820
rect 1820 4800 1822 4820
rect 1582 4120 1638 4176
rect 846 3304 902 3360
rect 570 1536 626 1592
rect 1214 2524 1216 2544
rect 1216 2524 1268 2544
rect 1268 2524 1270 2544
rect 1214 2488 1270 2524
rect 1398 2508 1454 2544
rect 1398 2488 1400 2508
rect 1400 2488 1452 2508
rect 1452 2488 1454 2508
rect 1582 3440 1638 3496
rect 2042 7404 2098 7440
rect 2042 7384 2044 7404
rect 2044 7384 2096 7404
rect 2096 7384 2098 7404
rect 2042 3576 2098 3632
rect 2778 12960 2834 13016
rect 2594 12300 2650 12336
rect 2594 12280 2596 12300
rect 2596 12280 2648 12300
rect 2648 12280 2650 12300
rect 3238 14320 3294 14376
rect 3238 13368 3294 13424
rect 3146 12960 3202 13016
rect 2870 11328 2926 11384
rect 2870 10260 2926 10296
rect 2870 10240 2872 10260
rect 2872 10240 2924 10260
rect 2924 10240 2926 10260
rect 3698 15580 3700 15600
rect 3700 15580 3752 15600
rect 3752 15580 3754 15600
rect 3698 15544 3754 15580
rect 3330 9696 3386 9752
rect 3514 10376 3570 10432
rect 3698 12416 3754 12472
rect 24122 27648 24178 27704
rect 4066 26016 4122 26072
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 4618 22616 4674 22672
rect 4526 21120 4582 21176
rect 4894 22344 4950 22400
rect 4250 20440 4306 20496
rect 4342 16940 4344 16960
rect 4344 16940 4396 16960
rect 4396 16940 4398 16960
rect 4342 16904 4398 16940
rect 3974 15952 4030 16008
rect 3882 15680 3938 15736
rect 3790 12280 3846 12336
rect 3790 11328 3846 11384
rect 3698 11192 3754 11248
rect 3146 9288 3202 9344
rect 2962 8880 3018 8936
rect 3330 8880 3386 8936
rect 3606 9016 3662 9072
rect 3146 7384 3202 7440
rect 2870 6976 2926 7032
rect 3054 6296 3110 6352
rect 2778 5480 2834 5536
rect 2134 3032 2190 3088
rect 2502 3576 2558 3632
rect 1950 1944 2006 2000
rect 1950 1808 2006 1864
rect 1306 856 1362 912
rect 3054 5752 3110 5808
rect 2962 5244 2964 5264
rect 2964 5244 3016 5264
rect 3016 5244 3018 5264
rect 2962 5208 3018 5244
rect 2962 3712 3018 3768
rect 2870 2760 2926 2816
rect 3606 7792 3662 7848
rect 3514 5888 3570 5944
rect 3514 5616 3570 5672
rect 4066 15544 4122 15600
rect 3974 13640 4030 13696
rect 4066 13096 4122 13152
rect 4066 12688 4122 12744
rect 4250 16496 4306 16552
rect 4802 18400 4858 18456
rect 4618 17720 4674 17776
rect 4250 11736 4306 11792
rect 3882 8336 3938 8392
rect 3698 4664 3754 4720
rect 3882 3984 3938 4040
rect 4066 8608 4122 8664
rect 4250 10140 4252 10160
rect 4252 10140 4304 10160
rect 4304 10140 4306 10160
rect 4250 10104 4306 10140
rect 4618 12552 4674 12608
rect 4618 12280 4674 12336
rect 4434 11192 4490 11248
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5538 18128 5594 18184
rect 5078 16088 5134 16144
rect 5998 17584 6054 17640
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5538 15564 5594 15600
rect 5538 15544 5540 15564
rect 5540 15544 5592 15564
rect 5592 15544 5594 15564
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5998 14864 6054 14920
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5630 13932 5686 13968
rect 5630 13912 5632 13932
rect 5632 13912 5684 13932
rect 5684 13912 5686 13932
rect 5998 13640 6054 13696
rect 4342 8508 4344 8528
rect 4344 8508 4396 8528
rect 4396 8508 4398 8528
rect 4342 8472 4398 8508
rect 4710 8608 4766 8664
rect 4986 7384 5042 7440
rect 4802 7112 4858 7168
rect 4710 6976 4766 7032
rect 4250 5072 4306 5128
rect 4066 3848 4122 3904
rect 3974 3712 4030 3768
rect 3606 3032 3662 3088
rect 2778 1672 2834 1728
rect 3514 1400 3570 1456
rect 3054 992 3110 1048
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5538 12844 5594 12880
rect 5538 12824 5540 12844
rect 5540 12824 5592 12844
rect 5592 12824 5594 12844
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5354 10920 5410 10976
rect 5354 10512 5410 10568
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5354 10104 5410 10160
rect 5354 9832 5410 9888
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6458 20168 6514 20224
rect 6182 11328 6238 11384
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6918 17992 6974 18048
rect 6642 15700 6698 15736
rect 6642 15680 6644 15700
rect 6644 15680 6696 15700
rect 6696 15680 6698 15700
rect 9218 24792 9274 24848
rect 7378 21256 7434 21312
rect 6458 12960 6514 13016
rect 6642 12416 6698 12472
rect 6826 12180 6828 12200
rect 6828 12180 6880 12200
rect 6880 12180 6882 12200
rect 6826 12144 6882 12180
rect 6734 12008 6790 12064
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 25410 27104 25466 27160
rect 24766 25336 24822 25392
rect 23846 24248 23902 24304
rect 22650 24112 22706 24168
rect 22742 23704 22798 23760
rect 20626 23568 20682 23624
rect 15290 23432 15346 23488
rect 17498 23432 17554 23488
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 10782 20848 10838 20904
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9218 19896 9274 19952
rect 12898 19896 12954 19952
rect 9034 19216 9090 19272
rect 9126 17176 9182 17232
rect 8022 15408 8078 15464
rect 7470 13912 7526 13968
rect 7286 12280 7342 12336
rect 6458 10376 6514 10432
rect 6734 10376 6790 10432
rect 6458 9832 6514 9888
rect 5446 6976 5502 7032
rect 5354 6724 5410 6760
rect 5354 6704 5356 6724
rect 5356 6704 5408 6724
rect 5408 6704 5410 6724
rect 5262 6432 5318 6488
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5446 5752 5502 5808
rect 4802 5344 4858 5400
rect 5078 4664 5134 4720
rect 5354 5480 5410 5536
rect 5354 5072 5410 5128
rect 4802 4528 4858 4584
rect 4802 3984 4858 4040
rect 5262 4140 5318 4176
rect 5262 4120 5264 4140
rect 5264 4120 5316 4140
rect 5316 4120 5318 4140
rect 5170 3984 5226 4040
rect 5170 3304 5226 3360
rect 6274 7248 6330 7304
rect 6458 7268 6514 7304
rect 6458 7248 6460 7268
rect 6460 7248 6512 7268
rect 6512 7248 6514 7268
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5998 5344 6054 5400
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5354 3032 5410 3088
rect 6274 5208 6330 5264
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5906 2372 5962 2408
rect 5906 2352 5908 2372
rect 5908 2352 5960 2372
rect 5960 2352 5962 2372
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 4434 40 4490 96
rect 8390 14320 8446 14376
rect 8206 13812 8208 13832
rect 8208 13812 8260 13832
rect 8260 13812 8262 13832
rect 8206 13776 8262 13812
rect 8206 13368 8262 13424
rect 7562 12724 7564 12744
rect 7564 12724 7616 12744
rect 7616 12724 7618 12744
rect 7562 12688 7618 12724
rect 8206 12688 8262 12744
rect 7654 12144 7710 12200
rect 7562 10512 7618 10568
rect 7470 9696 7526 9752
rect 7378 9288 7434 9344
rect 7010 6316 7066 6352
rect 7010 6296 7012 6316
rect 7012 6296 7064 6316
rect 7064 6296 7066 6316
rect 6918 5616 6974 5672
rect 7102 5480 7158 5536
rect 6550 2896 6606 2952
rect 6458 2796 6460 2816
rect 6460 2796 6512 2816
rect 6512 2796 6514 2816
rect 6458 2760 6514 2796
rect 8390 13368 8446 13424
rect 8298 10920 8354 10976
rect 8298 10240 8354 10296
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9402 17176 9458 17232
rect 9218 14592 9274 14648
rect 9862 17040 9918 17096
rect 8482 10512 8538 10568
rect 8022 9560 8078 9616
rect 9218 12164 9274 12200
rect 9218 12144 9220 12164
rect 9220 12144 9272 12164
rect 9272 12144 9274 12164
rect 9586 15544 9642 15600
rect 9310 10920 9366 10976
rect 9126 9424 9182 9480
rect 7286 3304 7342 3360
rect 7010 2624 7066 2680
rect 6826 2352 6882 2408
rect 7286 1264 7342 1320
rect 6182 312 6238 368
rect 7838 6568 7894 6624
rect 7930 6296 7986 6352
rect 8574 6160 8630 6216
rect 7746 4664 7802 4720
rect 7746 1944 7802 2000
rect 7930 1128 7986 1184
rect 8574 4800 8630 4856
rect 8206 3712 8262 3768
rect 8390 4140 8446 4176
rect 8390 4120 8392 4140
rect 8392 4120 8444 4140
rect 8444 4120 8446 4140
rect 8942 6840 8998 6896
rect 8942 5616 8998 5672
rect 8850 5072 8906 5128
rect 8114 3168 8170 3224
rect 8022 584 8078 640
rect 7010 176 7066 232
rect 8758 3884 8760 3904
rect 8760 3884 8812 3904
rect 8812 3884 8814 3904
rect 8758 3848 8814 3884
rect 9034 5208 9090 5264
rect 9034 4392 9090 4448
rect 9034 4256 9090 4312
rect 8850 3476 8852 3496
rect 8852 3476 8904 3496
rect 8904 3476 8906 3496
rect 8850 3440 8906 3476
rect 8666 2760 8722 2816
rect 8850 1672 8906 1728
rect 8850 856 8906 912
rect 8758 720 8814 776
rect 9586 11636 9588 11656
rect 9588 11636 9640 11656
rect 9640 11636 9642 11656
rect 9586 11600 9642 11636
rect 9586 11228 9588 11248
rect 9588 11228 9640 11248
rect 9640 11228 9642 11248
rect 9586 11192 9642 11228
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 11610 16088 11666 16144
rect 11334 15952 11390 16008
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10598 15020 10654 15056
rect 10598 15000 10600 15020
rect 10600 15000 10652 15020
rect 10652 15000 10654 15020
rect 11242 15816 11298 15872
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10046 14048 10102 14104
rect 10138 13776 10194 13832
rect 9862 12436 9918 12472
rect 9862 12416 9864 12436
rect 9864 12416 9916 12436
rect 9916 12416 9918 12436
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10782 13096 10838 13152
rect 10690 12960 10746 13016
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10690 12416 10746 12472
rect 9862 12008 9918 12064
rect 9770 11328 9826 11384
rect 9954 11328 10010 11384
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 9494 9424 9550 9480
rect 9770 5480 9826 5536
rect 9402 5208 9458 5264
rect 9310 2388 9312 2408
rect 9312 2388 9364 2408
rect 9364 2388 9366 2408
rect 9310 2352 9366 2388
rect 9402 2080 9458 2136
rect 10874 12552 10930 12608
rect 10874 11872 10930 11928
rect 11242 11600 11298 11656
rect 11150 11464 11206 11520
rect 10874 11056 10930 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10598 9560 10654 9616
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10782 8880 10838 8936
rect 10782 8744 10838 8800
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10138 8084 10194 8120
rect 10138 8064 10140 8084
rect 10140 8064 10192 8084
rect 10192 8064 10194 8084
rect 9954 7384 10010 7440
rect 10690 7248 10746 7304
rect 9954 6976 10010 7032
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10782 5888 10838 5944
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10322 4120 10378 4176
rect 10506 4120 10562 4176
rect 9586 1672 9642 1728
rect 9954 3712 10010 3768
rect 9862 2624 9918 2680
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3576 10194 3632
rect 12530 15544 12586 15600
rect 11426 12960 11482 13016
rect 11426 12144 11482 12200
rect 11978 10104 12034 10160
rect 11978 8236 11980 8256
rect 11980 8236 12032 8256
rect 12032 8236 12034 8256
rect 11978 8200 12034 8236
rect 11886 7656 11942 7712
rect 11518 6840 11574 6896
rect 11702 5072 11758 5128
rect 10506 3440 10562 3496
rect 10506 3032 10562 3088
rect 11150 2796 11152 2816
rect 11152 2796 11204 2816
rect 11204 2796 11206 2816
rect 11150 2760 11206 2796
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10874 1128 10930 1184
rect 11058 1128 11114 1184
rect 11058 856 11114 912
rect 8206 176 8262 232
rect 11610 1536 11666 1592
rect 11886 5772 11942 5808
rect 12162 10104 12218 10160
rect 12162 9832 12218 9888
rect 12438 12416 12494 12472
rect 12346 11464 12402 11520
rect 12162 9152 12218 9208
rect 12438 10376 12494 10432
rect 12162 6296 12218 6352
rect 11886 5752 11888 5772
rect 11888 5752 11940 5772
rect 11940 5752 11942 5772
rect 12162 5752 12218 5808
rect 11886 5344 11942 5400
rect 11886 5072 11942 5128
rect 12254 4936 12310 4992
rect 12438 8880 12494 8936
rect 12806 12280 12862 12336
rect 12806 11736 12862 11792
rect 12714 8880 12770 8936
rect 12714 8336 12770 8392
rect 12622 7112 12678 7168
rect 12438 5888 12494 5944
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 17958 22072 18014 22128
rect 19522 22072 19578 22128
rect 16210 20848 16266 20904
rect 15290 19216 15346 19272
rect 15934 18808 15990 18864
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 12990 14456 13046 14512
rect 12990 12552 13046 12608
rect 13174 12280 13230 12336
rect 13082 7520 13138 7576
rect 12622 5072 12678 5128
rect 11978 3168 12034 3224
rect 12714 4140 12770 4176
rect 12714 4120 12716 4140
rect 12716 4120 12768 4140
rect 12768 4120 12770 4140
rect 13082 5072 13138 5128
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14462 16088 14518 16144
rect 13450 15544 13506 15600
rect 13542 14456 13598 14512
rect 13450 13368 13506 13424
rect 14002 13640 14058 13696
rect 13910 13504 13966 13560
rect 13910 13232 13966 13288
rect 13450 13132 13452 13152
rect 13452 13132 13504 13152
rect 13504 13132 13506 13152
rect 13450 13096 13506 13132
rect 13358 10648 13414 10704
rect 13358 9560 13414 9616
rect 13450 6296 13506 6352
rect 13450 6060 13452 6080
rect 13452 6060 13504 6080
rect 13504 6060 13506 6080
rect 13450 6024 13506 6060
rect 12898 2624 12954 2680
rect 12530 1944 12586 2000
rect 11794 1400 11850 1456
rect 11978 1400 12034 1456
rect 13266 3712 13322 3768
rect 14002 10376 14058 10432
rect 13818 7656 13874 7712
rect 13818 7520 13874 7576
rect 13818 7248 13874 7304
rect 13634 5772 13690 5808
rect 13634 5752 13636 5772
rect 13636 5752 13688 5772
rect 13688 5752 13690 5772
rect 14094 7384 14150 7440
rect 13542 4664 13598 4720
rect 15290 15408 15346 15464
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14462 12008 14518 12064
rect 14370 11600 14426 11656
rect 14646 12280 14702 12336
rect 14370 7112 14426 7168
rect 14554 7112 14610 7168
rect 14462 6704 14518 6760
rect 14278 4120 14334 4176
rect 14922 14612 14978 14648
rect 14922 14592 14924 14612
rect 14924 14592 14976 14612
rect 14976 14592 14978 14612
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15290 13640 15346 13696
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15382 13232 15438 13288
rect 14922 12144 14978 12200
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14830 11464 14886 11520
rect 14830 11192 14886 11248
rect 15106 11500 15108 11520
rect 15108 11500 15160 11520
rect 15160 11500 15162 11520
rect 15106 11464 15162 11500
rect 14922 11076 14978 11112
rect 14922 11056 14924 11076
rect 14924 11056 14976 11076
rect 14976 11056 14978 11076
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15290 10260 15346 10296
rect 15290 10240 15292 10260
rect 15292 10240 15344 10260
rect 15344 10240 15346 10260
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14922 9444 14978 9480
rect 14922 9424 14924 9444
rect 14924 9424 14976 9444
rect 14976 9424 14978 9444
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15474 9016 15530 9072
rect 15290 8472 15346 8528
rect 14830 7964 14832 7984
rect 14832 7964 14884 7984
rect 14884 7964 14886 7984
rect 14830 7928 14886 7964
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14830 6860 14886 6896
rect 14830 6840 14832 6860
rect 14832 6840 14884 6860
rect 14884 6840 14886 6860
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 16026 18264 16082 18320
rect 15934 12824 15990 12880
rect 15750 11736 15806 11792
rect 15842 10784 15898 10840
rect 15658 8880 15714 8936
rect 15658 8356 15714 8392
rect 15658 8336 15660 8356
rect 15660 8336 15712 8356
rect 15712 8336 15714 8356
rect 16118 11192 16174 11248
rect 16026 11092 16028 11112
rect 16028 11092 16080 11112
rect 16080 11092 16082 11112
rect 16026 11056 16082 11092
rect 16026 10920 16082 10976
rect 16026 10376 16082 10432
rect 16118 9988 16174 10024
rect 16118 9968 16120 9988
rect 16120 9968 16172 9988
rect 16172 9968 16174 9988
rect 16302 10376 16358 10432
rect 16026 9016 16082 9072
rect 15842 7928 15898 7984
rect 16026 8472 16082 8528
rect 15382 5616 15438 5672
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14646 4392 14702 4448
rect 13634 3476 13636 3496
rect 13636 3476 13688 3496
rect 13688 3476 13690 3496
rect 13634 3440 13690 3476
rect 13910 3440 13966 3496
rect 14186 3848 14242 3904
rect 14002 2896 14058 2952
rect 13450 2216 13506 2272
rect 13174 992 13230 1048
rect 14094 2352 14150 2408
rect 14002 2080 14058 2136
rect 13726 1944 13782 2000
rect 14094 1944 14150 2000
rect 14554 3984 14610 4040
rect 14554 3304 14610 3360
rect 14554 3032 14610 3088
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14738 4256 14794 4312
rect 15014 3712 15070 3768
rect 15474 4664 15530 4720
rect 15474 4020 15476 4040
rect 15476 4020 15528 4040
rect 15528 4020 15530 4040
rect 15474 3984 15530 4020
rect 16118 6568 16174 6624
rect 15658 3304 15714 3360
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15198 2796 15200 2816
rect 15200 2796 15252 2816
rect 15252 2796 15254 2816
rect 15198 2760 15254 2796
rect 14646 2488 14702 2544
rect 15842 2488 15898 2544
rect 15198 2388 15200 2408
rect 15200 2388 15252 2408
rect 15252 2388 15254 2408
rect 15198 2352 15254 2388
rect 15382 2216 15438 2272
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15474 1672 15530 1728
rect 16486 6432 16542 6488
rect 16578 6296 16634 6352
rect 16946 15408 17002 15464
rect 16854 14320 16910 14376
rect 16854 13912 16910 13968
rect 17222 13368 17278 13424
rect 16854 12144 16910 12200
rect 16946 11736 17002 11792
rect 16854 8628 16910 8664
rect 16854 8608 16856 8628
rect 16856 8608 16908 8628
rect 16908 8608 16910 8628
rect 17774 15852 17776 15872
rect 17776 15852 17828 15872
rect 17828 15852 17830 15872
rect 17774 15816 17830 15852
rect 17866 13504 17922 13560
rect 17498 12724 17500 12744
rect 17500 12724 17552 12744
rect 17552 12724 17554 12744
rect 17498 12688 17554 12724
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 18326 20576 18382 20632
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 18694 19896 18750 19952
rect 18142 15272 18198 15328
rect 18050 11736 18106 11792
rect 17590 11464 17646 11520
rect 17406 10684 17408 10704
rect 17408 10684 17460 10704
rect 17460 10684 17462 10704
rect 17406 10648 17462 10684
rect 17406 10104 17462 10160
rect 17038 6976 17094 7032
rect 16762 6840 16818 6896
rect 16670 5480 16726 5536
rect 16486 4936 16542 4992
rect 16854 5208 16910 5264
rect 16854 3576 16910 3632
rect 17406 5344 17462 5400
rect 18510 13812 18512 13832
rect 18512 13812 18564 13832
rect 18564 13812 18566 13832
rect 18510 13776 18566 13812
rect 18326 12688 18382 12744
rect 18234 12280 18290 12336
rect 18142 10648 18198 10704
rect 18142 10376 18198 10432
rect 17774 9424 17830 9480
rect 18142 9152 18198 9208
rect 17958 5208 18014 5264
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 18878 16632 18934 16688
rect 18878 16496 18934 16552
rect 18602 10784 18658 10840
rect 18510 9580 18566 9616
rect 18510 9560 18512 9580
rect 18512 9560 18564 9580
rect 18564 9560 18566 9580
rect 18510 9424 18566 9480
rect 18602 7812 18658 7848
rect 18602 7792 18604 7812
rect 18604 7792 18656 7812
rect 18656 7792 18658 7812
rect 18602 6604 18604 6624
rect 18604 6604 18656 6624
rect 18656 6604 18658 6624
rect 18602 6568 18658 6604
rect 18326 5652 18328 5672
rect 18328 5652 18380 5672
rect 18380 5652 18382 5672
rect 18326 5616 18382 5652
rect 18050 4528 18106 4584
rect 17590 4256 17646 4312
rect 17590 4120 17646 4176
rect 17314 3576 17370 3632
rect 17038 2624 17094 2680
rect 17038 1536 17094 1592
rect 16762 1264 16818 1320
rect 17774 1400 17830 1456
rect 17958 1128 18014 1184
rect 19338 17076 19340 17096
rect 19340 17076 19392 17096
rect 19392 17076 19394 17096
rect 19338 17040 19394 17076
rect 19062 15000 19118 15056
rect 18878 12280 18934 12336
rect 18878 9868 18880 9888
rect 18880 9868 18932 9888
rect 18932 9868 18934 9888
rect 18878 9832 18934 9868
rect 18786 7384 18842 7440
rect 18602 5616 18658 5672
rect 19338 15308 19340 15328
rect 19340 15308 19392 15328
rect 19392 15308 19394 15328
rect 19338 15272 19394 15308
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19890 17620 19892 17640
rect 19892 17620 19944 17640
rect 19944 17620 19946 17640
rect 19890 17584 19946 17620
rect 20074 20168 20130 20224
rect 20810 19216 20866 19272
rect 20074 17856 20130 17912
rect 19982 17176 20038 17232
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19522 15544 19578 15600
rect 19338 13388 19394 13424
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19338 13368 19340 13388
rect 19340 13368 19392 13388
rect 19392 13368 19394 13388
rect 19982 13096 20038 13152
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19522 12280 19578 12336
rect 19062 10240 19118 10296
rect 19430 10240 19486 10296
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19246 9696 19302 9752
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19062 8880 19118 8936
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 20166 12144 20222 12200
rect 20166 11192 20222 11248
rect 20534 13504 20590 13560
rect 21546 18128 21602 18184
rect 21270 17740 21326 17776
rect 21270 17720 21272 17740
rect 21272 17720 21324 17740
rect 21324 17720 21326 17740
rect 20994 17448 21050 17504
rect 22282 17584 22338 17640
rect 20902 15952 20958 16008
rect 21270 16652 21326 16688
rect 21270 16632 21272 16652
rect 21272 16632 21324 16652
rect 21324 16632 21326 16652
rect 20902 13640 20958 13696
rect 20994 13232 21050 13288
rect 19338 7792 19394 7848
rect 19338 7112 19394 7168
rect 19338 4972 19340 4992
rect 19340 4972 19392 4992
rect 19392 4972 19394 4992
rect 19338 4936 19394 4972
rect 18418 3984 18474 4040
rect 18970 3984 19026 4040
rect 19338 3884 19340 3904
rect 19340 3884 19392 3904
rect 19392 3884 19394 3904
rect 19338 3848 19394 3884
rect 18694 3032 18750 3088
rect 18694 2896 18750 2952
rect 18602 1944 18658 2000
rect 18142 720 18198 776
rect 18050 584 18106 640
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19890 4428 19892 4448
rect 19892 4428 19944 4448
rect 19944 4428 19946 4448
rect 19890 4392 19946 4428
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19522 3440 19578 3496
rect 19430 2216 19486 2272
rect 19246 1808 19302 1864
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20442 7928 20498 7984
rect 20350 6296 20406 6352
rect 20350 3984 20406 4040
rect 20166 3712 20222 3768
rect 20166 3340 20168 3360
rect 20168 3340 20220 3360
rect 20220 3340 20222 3360
rect 20166 3304 20222 3340
rect 20258 3168 20314 3224
rect 19982 2080 20038 2136
rect 21086 10532 21142 10568
rect 21086 10512 21088 10532
rect 21088 10512 21140 10532
rect 21140 10512 21142 10532
rect 20902 9560 20958 9616
rect 21086 9152 21142 9208
rect 21914 16768 21970 16824
rect 22558 17604 22614 17640
rect 22558 17584 22560 17604
rect 22560 17584 22612 17604
rect 22612 17584 22614 17604
rect 22466 16632 22522 16688
rect 21546 16108 21602 16144
rect 21546 16088 21548 16108
rect 21548 16088 21600 16108
rect 21600 16088 21602 16108
rect 21454 14612 21510 14648
rect 21454 14592 21456 14612
rect 21456 14592 21508 14612
rect 21508 14592 21510 14612
rect 21914 14456 21970 14512
rect 21270 9696 21326 9752
rect 21362 8916 21364 8936
rect 21364 8916 21416 8936
rect 21416 8916 21418 8936
rect 21362 8880 21418 8916
rect 21178 8744 21234 8800
rect 21178 7928 21234 7984
rect 20994 5888 21050 5944
rect 21270 6840 21326 6896
rect 20994 5616 21050 5672
rect 21914 11600 21970 11656
rect 22006 11056 22062 11112
rect 21638 8336 21694 8392
rect 21546 7520 21602 7576
rect 21546 7384 21602 7440
rect 21454 6840 21510 6896
rect 21362 6568 21418 6624
rect 22098 9288 22154 9344
rect 21914 8336 21970 8392
rect 21730 4800 21786 4856
rect 20626 2760 20682 2816
rect 21178 3440 21234 3496
rect 22006 7928 22062 7984
rect 22098 7792 22154 7848
rect 22374 10648 22430 10704
rect 22466 9460 22468 9480
rect 22468 9460 22520 9480
rect 22520 9460 22522 9480
rect 22466 9424 22522 9460
rect 22282 9152 22338 9208
rect 23478 22480 23534 22536
rect 22650 16088 22706 16144
rect 22926 16496 22982 16552
rect 23202 14900 23204 14920
rect 23204 14900 23256 14920
rect 23256 14900 23258 14920
rect 23202 14864 23258 14900
rect 22190 5072 22246 5128
rect 22466 6432 22522 6488
rect 22742 6296 22798 6352
rect 22834 5616 22890 5672
rect 22742 5480 22798 5536
rect 21546 3576 21602 3632
rect 22098 3712 22154 3768
rect 21270 2644 21326 2680
rect 21270 2624 21272 2644
rect 21272 2624 21324 2644
rect 21324 2624 21326 2644
rect 21638 3032 21694 3088
rect 22466 2760 22522 2816
rect 23846 19896 23902 19952
rect 23478 15000 23534 15056
rect 23478 14068 23534 14104
rect 23478 14048 23480 14068
rect 23480 14048 23532 14068
rect 23532 14048 23534 14068
rect 23386 9152 23442 9208
rect 23662 16768 23718 16824
rect 23754 11736 23810 11792
rect 23662 11056 23718 11112
rect 23570 8880 23626 8936
rect 23478 7948 23534 7984
rect 23478 7928 23480 7948
rect 23480 7928 23532 7948
rect 23532 7928 23534 7948
rect 23386 6840 23442 6896
rect 23294 5752 23350 5808
rect 23294 5480 23350 5536
rect 24122 24792 24178 24848
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24112 24270 24168
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24582 23604 24584 23624
rect 24584 23604 24636 23624
rect 24636 23604 24638 23624
rect 24582 23568 24638 23604
rect 24766 23160 24822 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24674 21936 24730 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24766 21392 24822 21448
rect 24674 20304 24730 20360
rect 24582 20168 24638 20224
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24214 19352 24270 19408
rect 24582 19252 24584 19272
rect 24584 19252 24636 19272
rect 24636 19252 24638 19272
rect 24582 19216 24638 19252
rect 24766 19116 24768 19136
rect 24768 19116 24820 19136
rect 24820 19116 24822 19136
rect 24766 19080 24822 19116
rect 24582 18828 24638 18864
rect 24582 18808 24584 18828
rect 24584 18808 24636 18828
rect 24636 18808 24638 18828
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24490 18028 24492 18048
rect 24492 18028 24544 18048
rect 24544 18028 24546 18048
rect 24490 17992 24546 18028
rect 24214 17856 24270 17912
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24122 16652 24178 16688
rect 24122 16632 24124 16652
rect 24124 16632 24176 16652
rect 24176 16632 24178 16652
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25134 16940 25136 16960
rect 25136 16940 25188 16960
rect 25188 16940 25190 16960
rect 25134 16904 25190 16940
rect 24766 16768 24822 16824
rect 25134 16496 25190 16552
rect 24030 15680 24086 15736
rect 23938 11892 23994 11928
rect 23938 11872 23940 11892
rect 23940 11872 23992 11892
rect 23992 11872 23994 11892
rect 24582 15408 24638 15464
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24766 15136 24822 15192
rect 25686 26560 25742 26616
rect 25502 26016 25558 26072
rect 25410 15020 25466 15056
rect 25410 15000 25412 15020
rect 25412 15000 25464 15020
rect 25464 15000 25466 15020
rect 25226 13776 25282 13832
rect 25042 13640 25098 13696
rect 24858 13368 24914 13424
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24214 7384 24270 7440
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23846 5616 23902 5672
rect 23294 4800 23350 4856
rect 23202 4256 23258 4312
rect 23018 1672 23074 1728
rect 10966 312 11022 368
rect 23294 3712 23350 3768
rect 23662 3304 23718 3360
rect 23570 2896 23626 2952
rect 22558 40 22614 96
rect 23846 4528 23902 4584
rect 23846 3984 23902 4040
rect 23478 312 23534 368
rect 25226 11600 25282 11656
rect 24490 5616 24546 5672
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24214 5208 24270 5264
rect 25134 7828 25136 7848
rect 25136 7828 25188 7848
rect 25188 7828 25190 7848
rect 25134 7792 25190 7828
rect 25042 5908 25098 5944
rect 25042 5888 25044 5908
rect 25044 5888 25096 5908
rect 25096 5888 25098 5908
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24858 4120 24914 4176
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25226 4664 25282 4720
rect 25778 13504 25834 13560
rect 25410 6432 25466 6488
rect 25686 7928 25742 7984
rect 25502 6160 25558 6216
rect 25318 2760 25374 2816
rect 25226 1400 25282 1456
rect 25686 3712 25742 3768
rect 26146 6568 26202 6624
rect 26054 3168 26110 3224
rect 25594 2508 25650 2544
rect 25594 2488 25596 2508
rect 25596 2488 25648 2508
rect 25648 2488 25650 2508
rect 25870 2524 25872 2544
rect 25872 2524 25924 2544
rect 25924 2524 25926 2544
rect 25870 2488 25926 2524
rect 23662 176 23718 232
rect 26238 856 26294 912
rect 27066 1944 27122 2000
rect 27250 1944 27306 2000
rect 27618 1672 27674 1728
rect 26054 312 26110 368
<< metal3 >>
rect 0 27706 480 27736
rect 4061 27706 4127 27709
rect 0 27704 4127 27706
rect 0 27648 4066 27704
rect 4122 27648 4127 27704
rect 0 27646 4127 27648
rect 0 27616 480 27646
rect 4061 27643 4127 27646
rect 24117 27706 24183 27709
rect 27520 27706 28000 27736
rect 24117 27704 28000 27706
rect 24117 27648 24122 27704
rect 24178 27648 28000 27704
rect 24117 27646 28000 27648
rect 24117 27643 24183 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 3785 27162 3851 27165
rect 0 27160 3851 27162
rect 0 27104 3790 27160
rect 3846 27104 3851 27160
rect 0 27102 3851 27104
rect 0 27072 480 27102
rect 3785 27099 3851 27102
rect 25405 27162 25471 27165
rect 27520 27162 28000 27192
rect 25405 27160 28000 27162
rect 25405 27104 25410 27160
rect 25466 27104 28000 27160
rect 25405 27102 28000 27104
rect 25405 27099 25471 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 2681 26618 2747 26621
rect 0 26616 2747 26618
rect 0 26560 2686 26616
rect 2742 26560 2747 26616
rect 0 26558 2747 26560
rect 0 26528 480 26558
rect 2681 26555 2747 26558
rect 25681 26618 25747 26621
rect 27520 26618 28000 26648
rect 25681 26616 28000 26618
rect 25681 26560 25686 26616
rect 25742 26560 28000 26616
rect 25681 26558 28000 26560
rect 25681 26555 25747 26558
rect 27520 26528 28000 26558
rect 0 26074 480 26104
rect 4061 26074 4127 26077
rect 0 26072 4127 26074
rect 0 26016 4066 26072
rect 4122 26016 4127 26072
rect 0 26014 4127 26016
rect 0 25984 480 26014
rect 4061 26011 4127 26014
rect 25497 26074 25563 26077
rect 27520 26074 28000 26104
rect 25497 26072 28000 26074
rect 25497 26016 25502 26072
rect 25558 26016 28000 26072
rect 25497 26014 28000 26016
rect 25497 26011 25563 26014
rect 27520 25984 28000 26014
rect 10277 25600 10597 25601
rect 0 25530 480 25560
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 3325 25530 3391 25533
rect 0 25528 3391 25530
rect 0 25472 3330 25528
rect 3386 25472 3391 25528
rect 0 25470 3391 25472
rect 0 25440 480 25470
rect 3325 25467 3391 25470
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 24761 25392 28000 25394
rect 24761 25336 24766 25392
rect 24822 25336 28000 25392
rect 24761 25334 28000 25336
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 0 24986 480 25016
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 1577 24986 1643 24989
rect 0 24984 1643 24986
rect 0 24928 1582 24984
rect 1638 24928 1643 24984
rect 0 24926 1643 24928
rect 0 24896 480 24926
rect 1577 24923 1643 24926
rect 3509 24850 3575 24853
rect 9213 24850 9279 24853
rect 3509 24848 9279 24850
rect 3509 24792 3514 24848
rect 3570 24792 9218 24848
rect 9274 24792 9279 24848
rect 3509 24790 9279 24792
rect 3509 24787 3575 24790
rect 9213 24787 9279 24790
rect 24117 24850 24183 24853
rect 27520 24850 28000 24880
rect 24117 24848 28000 24850
rect 24117 24792 24122 24848
rect 24178 24792 28000 24848
rect 24117 24790 28000 24792
rect 24117 24787 24183 24790
rect 27520 24760 28000 24790
rect 10277 24512 10597 24513
rect 0 24442 480 24472
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 1485 24442 1551 24445
rect 0 24440 1551 24442
rect 0 24384 1490 24440
rect 1546 24384 1551 24440
rect 0 24382 1551 24384
rect 0 24352 480 24382
rect 1485 24379 1551 24382
rect 23841 24306 23907 24309
rect 27520 24306 28000 24336
rect 23841 24304 28000 24306
rect 23841 24248 23846 24304
rect 23902 24248 28000 24304
rect 23841 24246 28000 24248
rect 23841 24243 23907 24246
rect 27520 24216 28000 24246
rect 22645 24170 22711 24173
rect 24209 24170 24275 24173
rect 22645 24168 24275 24170
rect 22645 24112 22650 24168
rect 22706 24112 24214 24168
rect 24270 24112 24275 24168
rect 22645 24110 24275 24112
rect 22645 24107 22711 24110
rect 24209 24107 24275 24110
rect 5610 23968 5930 23969
rect 0 23898 480 23928
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 1393 23898 1459 23901
rect 0 23896 1459 23898
rect 0 23840 1398 23896
rect 1454 23840 1459 23896
rect 0 23838 1459 23840
rect 0 23808 480 23838
rect 1393 23835 1459 23838
rect 22737 23762 22803 23765
rect 27520 23762 28000 23792
rect 22737 23760 28000 23762
rect 22737 23704 22742 23760
rect 22798 23704 28000 23760
rect 22737 23702 28000 23704
rect 22737 23699 22803 23702
rect 27520 23672 28000 23702
rect 20621 23626 20687 23629
rect 24577 23626 24643 23629
rect 20621 23624 24643 23626
rect 20621 23568 20626 23624
rect 20682 23568 24582 23624
rect 24638 23568 24643 23624
rect 20621 23566 24643 23568
rect 20621 23563 20687 23566
rect 24577 23563 24643 23566
rect 15285 23490 15351 23493
rect 17493 23490 17559 23493
rect 15285 23488 17559 23490
rect 15285 23432 15290 23488
rect 15346 23432 17498 23488
rect 17554 23432 17559 23488
rect 15285 23430 17559 23432
rect 15285 23427 15351 23430
rect 17493 23427 17559 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23218 480 23248
rect 1577 23218 1643 23221
rect 0 23216 1643 23218
rect 0 23160 1582 23216
rect 1638 23160 1643 23216
rect 0 23158 1643 23160
rect 0 23128 480 23158
rect 1577 23155 1643 23158
rect 24761 23218 24827 23221
rect 27520 23218 28000 23248
rect 24761 23216 28000 23218
rect 24761 23160 24766 23216
rect 24822 23160 28000 23216
rect 24761 23158 28000 23160
rect 24761 23155 24827 23158
rect 27520 23128 28000 23158
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22674 480 22704
rect 4613 22674 4679 22677
rect 0 22672 4679 22674
rect 0 22616 4618 22672
rect 4674 22616 4679 22672
rect 0 22614 4679 22616
rect 0 22584 480 22614
rect 4613 22611 4679 22614
rect 23473 22538 23539 22541
rect 27520 22538 28000 22568
rect 23473 22536 28000 22538
rect 23473 22480 23478 22536
rect 23534 22480 28000 22536
rect 23473 22478 28000 22480
rect 23473 22475 23539 22478
rect 27520 22448 28000 22478
rect 2497 22402 2563 22405
rect 4889 22402 4955 22405
rect 2497 22400 4955 22402
rect 2497 22344 2502 22400
rect 2558 22344 4894 22400
rect 4950 22344 4955 22400
rect 2497 22342 4955 22344
rect 2497 22339 2563 22342
rect 4889 22339 4955 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 0 22130 480 22160
rect 1485 22130 1551 22133
rect 0 22128 1551 22130
rect 0 22072 1490 22128
rect 1546 22072 1551 22128
rect 0 22070 1551 22072
rect 0 22040 480 22070
rect 1485 22067 1551 22070
rect 17953 22130 18019 22133
rect 19517 22130 19583 22133
rect 17953 22128 19583 22130
rect 17953 22072 17958 22128
rect 18014 22072 19522 22128
rect 19578 22072 19583 22128
rect 17953 22070 19583 22072
rect 17953 22067 18019 22070
rect 19517 22067 19583 22070
rect 24669 21994 24735 21997
rect 27520 21994 28000 22024
rect 24669 21992 28000 21994
rect 24669 21936 24674 21992
rect 24730 21936 28000 21992
rect 24669 21934 28000 21936
rect 24669 21931 24735 21934
rect 27520 21904 28000 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21586 480 21616
rect 1577 21586 1643 21589
rect 0 21584 1643 21586
rect 0 21528 1582 21584
rect 1638 21528 1643 21584
rect 0 21526 1643 21528
rect 0 21496 480 21526
rect 1577 21523 1643 21526
rect 24761 21450 24827 21453
rect 27520 21450 28000 21480
rect 24761 21448 28000 21450
rect 24761 21392 24766 21448
rect 24822 21392 28000 21448
rect 24761 21390 28000 21392
rect 24761 21387 24827 21390
rect 27520 21360 28000 21390
rect 2037 21314 2103 21317
rect 7373 21314 7439 21317
rect 2037 21312 7439 21314
rect 2037 21256 2042 21312
rect 2098 21256 7378 21312
rect 7434 21256 7439 21312
rect 2037 21254 7439 21256
rect 2037 21251 2103 21254
rect 7373 21251 7439 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 2405 21178 2471 21181
rect 4521 21178 4587 21181
rect 2405 21176 4587 21178
rect 2405 21120 2410 21176
rect 2466 21120 4526 21176
rect 4582 21120 4587 21176
rect 2405 21118 4587 21120
rect 2405 21115 2471 21118
rect 4521 21115 4587 21118
rect 0 21042 480 21072
rect 2589 21042 2655 21045
rect 0 21040 2655 21042
rect 0 20984 2594 21040
rect 2650 20984 2655 21040
rect 0 20982 2655 20984
rect 0 20952 480 20982
rect 2589 20979 2655 20982
rect 10777 20906 10843 20909
rect 16205 20906 16271 20909
rect 27520 20906 28000 20936
rect 10777 20904 16271 20906
rect 10777 20848 10782 20904
rect 10838 20848 16210 20904
rect 16266 20848 16271 20904
rect 10777 20846 16271 20848
rect 10777 20843 10843 20846
rect 16205 20843 16271 20846
rect 23982 20846 28000 20906
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 18321 20634 18387 20637
rect 23982 20634 24042 20846
rect 27520 20816 28000 20846
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 18321 20632 24042 20634
rect 18321 20576 18326 20632
rect 18382 20576 24042 20632
rect 18321 20574 24042 20576
rect 18321 20571 18387 20574
rect 0 20498 480 20528
rect 4245 20498 4311 20501
rect 0 20496 4311 20498
rect 0 20440 4250 20496
rect 4306 20440 4311 20496
rect 0 20438 4311 20440
rect 0 20408 480 20438
rect 4245 20435 4311 20438
rect 24669 20362 24735 20365
rect 27520 20362 28000 20392
rect 24669 20360 28000 20362
rect 24669 20304 24674 20360
rect 24730 20304 28000 20360
rect 24669 20302 28000 20304
rect 24669 20299 24735 20302
rect 27520 20272 28000 20302
rect 2405 20226 2471 20229
rect 6453 20226 6519 20229
rect 2405 20224 6519 20226
rect 2405 20168 2410 20224
rect 2466 20168 6458 20224
rect 6514 20168 6519 20224
rect 2405 20166 6519 20168
rect 2405 20163 2471 20166
rect 6453 20163 6519 20166
rect 20069 20226 20135 20229
rect 24577 20226 24643 20229
rect 20069 20224 24643 20226
rect 20069 20168 20074 20224
rect 20130 20168 24582 20224
rect 24638 20168 24643 20224
rect 20069 20166 24643 20168
rect 20069 20163 20135 20166
rect 24577 20163 24643 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19954 480 19984
rect 1577 19954 1643 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 480 19894
rect 1577 19891 1643 19894
rect 9213 19954 9279 19957
rect 12893 19954 12959 19957
rect 9213 19952 12959 19954
rect 9213 19896 9218 19952
rect 9274 19896 12898 19952
rect 12954 19896 12959 19952
rect 9213 19894 12959 19896
rect 9213 19891 9279 19894
rect 12893 19891 12959 19894
rect 18689 19954 18755 19957
rect 23841 19954 23907 19957
rect 18689 19952 23907 19954
rect 18689 19896 18694 19952
rect 18750 19896 23846 19952
rect 23902 19896 23907 19952
rect 18689 19894 23907 19896
rect 18689 19891 18755 19894
rect 23841 19891 23907 19894
rect 27520 19682 28000 19712
rect 24718 19622 28000 19682
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19410 480 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 480 19350
rect 1577 19347 1643 19350
rect 24209 19410 24275 19413
rect 24718 19410 24778 19622
rect 27520 19592 28000 19622
rect 24209 19408 24778 19410
rect 24209 19352 24214 19408
rect 24270 19352 24778 19408
rect 24209 19350 24778 19352
rect 24209 19347 24275 19350
rect 9029 19274 9095 19277
rect 15285 19274 15351 19277
rect 9029 19272 15351 19274
rect 9029 19216 9034 19272
rect 9090 19216 15290 19272
rect 15346 19216 15351 19272
rect 9029 19214 15351 19216
rect 9029 19211 9095 19214
rect 15285 19211 15351 19214
rect 20805 19274 20871 19277
rect 24577 19274 24643 19277
rect 20805 19272 24643 19274
rect 20805 19216 20810 19272
rect 20866 19216 24582 19272
rect 24638 19216 24643 19272
rect 20805 19214 24643 19216
rect 20805 19211 20871 19214
rect 24577 19211 24643 19214
rect 2037 19138 2103 19141
rect 2814 19138 2820 19140
rect 2037 19136 2820 19138
rect 2037 19080 2042 19136
rect 2098 19080 2820 19136
rect 2037 19078 2820 19080
rect 2037 19075 2103 19078
rect 2814 19076 2820 19078
rect 2884 19076 2890 19140
rect 24761 19138 24827 19141
rect 27520 19138 28000 19168
rect 24761 19136 28000 19138
rect 24761 19080 24766 19136
rect 24822 19080 28000 19136
rect 24761 19078 28000 19080
rect 24761 19075 24827 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 2405 19002 2471 19005
rect 3366 19002 3372 19004
rect 2405 19000 3372 19002
rect 2405 18944 2410 19000
rect 2466 18944 3372 19000
rect 2405 18942 3372 18944
rect 2405 18939 2471 18942
rect 3366 18940 3372 18942
rect 3436 18940 3442 19004
rect 15929 18866 15995 18869
rect 24577 18866 24643 18869
rect 15929 18864 24643 18866
rect 15929 18808 15934 18864
rect 15990 18808 24582 18864
rect 24638 18808 24643 18864
rect 15929 18806 24643 18808
rect 15929 18803 15995 18806
rect 24577 18803 24643 18806
rect 0 18730 480 18760
rect 1577 18730 1643 18733
rect 0 18728 1643 18730
rect 0 18672 1582 18728
rect 1638 18672 1643 18728
rect 0 18670 1643 18672
rect 0 18640 480 18670
rect 1577 18667 1643 18670
rect 27520 18594 28000 18624
rect 24902 18534 28000 18594
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 2589 18458 2655 18461
rect 4797 18458 4863 18461
rect 2589 18456 4863 18458
rect 2589 18400 2594 18456
rect 2650 18400 4802 18456
rect 4858 18400 4863 18456
rect 2589 18398 4863 18400
rect 2589 18395 2655 18398
rect 4797 18395 4863 18398
rect 16021 18322 16087 18325
rect 24902 18322 24962 18534
rect 27520 18504 28000 18534
rect 16021 18320 24962 18322
rect 16021 18264 16026 18320
rect 16082 18264 24962 18320
rect 16021 18262 24962 18264
rect 16021 18259 16087 18262
rect 0 18186 480 18216
rect 5533 18186 5599 18189
rect 0 18184 5599 18186
rect 0 18128 5538 18184
rect 5594 18128 5599 18184
rect 0 18126 5599 18128
rect 0 18096 480 18126
rect 5533 18123 5599 18126
rect 21541 18186 21607 18189
rect 21541 18184 24962 18186
rect 21541 18128 21546 18184
rect 21602 18128 24962 18184
rect 21541 18126 24962 18128
rect 21541 18123 21607 18126
rect 2221 18050 2287 18053
rect 6913 18050 6979 18053
rect 2221 18048 6979 18050
rect 2221 17992 2226 18048
rect 2282 17992 6918 18048
rect 6974 17992 6979 18048
rect 2221 17990 6979 17992
rect 2221 17987 2287 17990
rect 6913 17987 6979 17990
rect 24485 18050 24551 18053
rect 24710 18050 24716 18052
rect 24485 18048 24716 18050
rect 24485 17992 24490 18048
rect 24546 17992 24716 18048
rect 24485 17990 24716 17992
rect 24485 17987 24551 17990
rect 24710 17988 24716 17990
rect 24780 17988 24786 18052
rect 24902 18050 24962 18126
rect 27520 18050 28000 18080
rect 24902 17990 28000 18050
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 20069 17914 20135 17917
rect 24209 17914 24275 17917
rect 20069 17912 24275 17914
rect 20069 17856 20074 17912
rect 20130 17856 24214 17912
rect 24270 17856 24275 17912
rect 20069 17854 24275 17856
rect 20069 17851 20135 17854
rect 24209 17851 24275 17854
rect 4613 17778 4679 17781
rect 21265 17778 21331 17781
rect 4613 17776 21331 17778
rect 4613 17720 4618 17776
rect 4674 17720 21270 17776
rect 21326 17720 21331 17776
rect 4613 17718 21331 17720
rect 4613 17715 4679 17718
rect 21265 17715 21331 17718
rect 0 17642 480 17672
rect 5993 17642 6059 17645
rect 0 17640 6059 17642
rect 0 17584 5998 17640
rect 6054 17584 6059 17640
rect 0 17582 6059 17584
rect 0 17552 480 17582
rect 5993 17579 6059 17582
rect 19885 17642 19951 17645
rect 22277 17642 22343 17645
rect 19885 17640 22343 17642
rect 19885 17584 19890 17640
rect 19946 17584 22282 17640
rect 22338 17584 22343 17640
rect 19885 17582 22343 17584
rect 19885 17579 19951 17582
rect 22277 17579 22343 17582
rect 22553 17642 22619 17645
rect 22553 17640 25146 17642
rect 22553 17584 22558 17640
rect 22614 17584 25146 17640
rect 22553 17582 25146 17584
rect 22553 17579 22619 17582
rect 20989 17506 21055 17509
rect 15334 17504 21055 17506
rect 15334 17448 20994 17504
rect 21050 17448 21055 17504
rect 15334 17446 21055 17448
rect 25086 17506 25146 17582
rect 27520 17506 28000 17536
rect 25086 17446 28000 17506
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 2313 17234 2379 17237
rect 9121 17234 9187 17237
rect 2313 17232 9187 17234
rect 2313 17176 2318 17232
rect 2374 17176 9126 17232
rect 9182 17176 9187 17232
rect 2313 17174 9187 17176
rect 2313 17171 2379 17174
rect 9121 17171 9187 17174
rect 9397 17234 9463 17237
rect 15334 17234 15394 17446
rect 20989 17443 21055 17446
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 9397 17232 15394 17234
rect 9397 17176 9402 17232
rect 9458 17176 15394 17232
rect 9397 17174 15394 17176
rect 9397 17171 9463 17174
rect 17902 17172 17908 17236
rect 17972 17234 17978 17236
rect 19977 17234 20043 17237
rect 17972 17232 20043 17234
rect 17972 17176 19982 17232
rect 20038 17176 20043 17232
rect 17972 17174 20043 17176
rect 17972 17172 17978 17174
rect 19977 17171 20043 17174
rect 0 17098 480 17128
rect 2957 17098 3023 17101
rect 0 17096 3023 17098
rect 0 17040 2962 17096
rect 3018 17040 3023 17096
rect 0 17038 3023 17040
rect 0 17008 480 17038
rect 2957 17035 3023 17038
rect 9857 17098 9923 17101
rect 19333 17098 19399 17101
rect 9857 17096 19399 17098
rect 9857 17040 9862 17096
rect 9918 17040 19338 17096
rect 19394 17040 19399 17096
rect 9857 17038 19399 17040
rect 9857 17035 9923 17038
rect 19333 17035 19399 17038
rect 2221 16962 2287 16965
rect 4337 16962 4403 16965
rect 25129 16962 25195 16965
rect 2221 16960 4403 16962
rect 2221 16904 2226 16960
rect 2282 16904 4342 16960
rect 4398 16904 4403 16960
rect 2221 16902 4403 16904
rect 2221 16899 2287 16902
rect 4337 16899 4403 16902
rect 21406 16960 25195 16962
rect 21406 16904 25134 16960
rect 25190 16904 25195 16960
rect 21406 16902 25195 16904
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 18873 16690 18939 16693
rect 21265 16690 21331 16693
rect 18873 16688 21331 16690
rect 18873 16632 18878 16688
rect 18934 16632 21270 16688
rect 21326 16632 21331 16688
rect 18873 16630 21331 16632
rect 18873 16627 18939 16630
rect 21265 16627 21331 16630
rect 0 16554 480 16584
rect 4245 16554 4311 16557
rect 0 16552 4311 16554
rect 0 16496 4250 16552
rect 4306 16496 4311 16552
rect 0 16494 4311 16496
rect 0 16464 480 16494
rect 4245 16491 4311 16494
rect 18873 16554 18939 16557
rect 21406 16554 21466 16902
rect 25129 16899 25195 16902
rect 21909 16826 21975 16829
rect 23657 16826 23723 16829
rect 21909 16824 23723 16826
rect 21909 16768 21914 16824
rect 21970 16768 23662 16824
rect 23718 16768 23723 16824
rect 21909 16766 23723 16768
rect 21909 16763 21975 16766
rect 23657 16763 23723 16766
rect 24761 16826 24827 16829
rect 27520 16826 28000 16856
rect 24761 16824 28000 16826
rect 24761 16768 24766 16824
rect 24822 16768 28000 16824
rect 24761 16766 28000 16768
rect 24761 16763 24827 16766
rect 27520 16736 28000 16766
rect 22461 16690 22527 16693
rect 24117 16690 24183 16693
rect 22461 16688 24183 16690
rect 22461 16632 22466 16688
rect 22522 16632 24122 16688
rect 24178 16632 24183 16688
rect 22461 16630 24183 16632
rect 22461 16627 22527 16630
rect 24117 16627 24183 16630
rect 18873 16552 21466 16554
rect 18873 16496 18878 16552
rect 18934 16496 21466 16552
rect 18873 16494 21466 16496
rect 22921 16554 22987 16557
rect 25129 16554 25195 16557
rect 22921 16552 25195 16554
rect 22921 16496 22926 16552
rect 22982 16496 25134 16552
rect 25190 16496 25195 16552
rect 22921 16494 25195 16496
rect 18873 16491 18939 16494
rect 22921 16491 22987 16494
rect 25129 16491 25195 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 27520 16282 28000 16312
rect 27478 16192 28000 16282
rect 5073 16146 5139 16149
rect 11605 16146 11671 16149
rect 5073 16144 11671 16146
rect 5073 16088 5078 16144
rect 5134 16088 11610 16144
rect 11666 16088 11671 16144
rect 5073 16086 11671 16088
rect 5073 16083 5139 16086
rect 11605 16083 11671 16086
rect 14457 16146 14523 16149
rect 21541 16146 21607 16149
rect 14457 16144 21607 16146
rect 14457 16088 14462 16144
rect 14518 16088 21546 16144
rect 21602 16088 21607 16144
rect 14457 16086 21607 16088
rect 14457 16083 14523 16086
rect 21541 16083 21607 16086
rect 22645 16146 22711 16149
rect 27478 16146 27538 16192
rect 22645 16144 27538 16146
rect 22645 16088 22650 16144
rect 22706 16088 27538 16144
rect 22645 16086 27538 16088
rect 22645 16083 22711 16086
rect 0 16010 480 16040
rect 3969 16010 4035 16013
rect 0 16008 4035 16010
rect 0 15952 3974 16008
rect 4030 15952 4035 16008
rect 0 15950 4035 15952
rect 0 15920 480 15950
rect 3969 15947 4035 15950
rect 11329 16010 11395 16013
rect 20897 16010 20963 16013
rect 11329 16008 20963 16010
rect 11329 15952 11334 16008
rect 11390 15952 20902 16008
rect 20958 15952 20963 16008
rect 11329 15950 20963 15952
rect 11329 15947 11395 15950
rect 20897 15947 20963 15950
rect 11237 15874 11303 15877
rect 17769 15874 17835 15877
rect 11237 15872 17835 15874
rect 11237 15816 11242 15872
rect 11298 15816 17774 15872
rect 17830 15816 17835 15872
rect 11237 15814 17835 15816
rect 11237 15811 11303 15814
rect 17769 15811 17835 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 3877 15738 3943 15741
rect 6637 15738 6703 15741
rect 3877 15736 6703 15738
rect 3877 15680 3882 15736
rect 3938 15680 6642 15736
rect 6698 15680 6703 15736
rect 3877 15678 6703 15680
rect 3877 15675 3943 15678
rect 6637 15675 6703 15678
rect 24025 15738 24091 15741
rect 27520 15738 28000 15768
rect 24025 15736 28000 15738
rect 24025 15680 24030 15736
rect 24086 15680 28000 15736
rect 24025 15678 28000 15680
rect 24025 15675 24091 15678
rect 27520 15648 28000 15678
rect 3366 15540 3372 15604
rect 3436 15602 3442 15604
rect 3693 15602 3759 15605
rect 3436 15600 3759 15602
rect 3436 15544 3698 15600
rect 3754 15544 3759 15600
rect 3436 15542 3759 15544
rect 3436 15540 3442 15542
rect 3693 15539 3759 15542
rect 4061 15602 4127 15605
rect 5533 15602 5599 15605
rect 4061 15600 5599 15602
rect 4061 15544 4066 15600
rect 4122 15544 5538 15600
rect 5594 15544 5599 15600
rect 4061 15542 5599 15544
rect 4061 15539 4127 15542
rect 5533 15539 5599 15542
rect 9581 15602 9647 15605
rect 12525 15602 12591 15605
rect 9581 15600 12591 15602
rect 9581 15544 9586 15600
rect 9642 15544 12530 15600
rect 12586 15544 12591 15600
rect 9581 15542 12591 15544
rect 9581 15539 9647 15542
rect 12525 15539 12591 15542
rect 13445 15602 13511 15605
rect 19517 15602 19583 15605
rect 13445 15600 19583 15602
rect 13445 15544 13450 15600
rect 13506 15544 19522 15600
rect 19578 15544 19583 15600
rect 13445 15542 19583 15544
rect 13445 15539 13511 15542
rect 19517 15539 19583 15542
rect 0 15466 480 15496
rect 8017 15466 8083 15469
rect 15285 15466 15351 15469
rect 0 15406 4906 15466
rect 0 15376 480 15406
rect 4846 15058 4906 15406
rect 8017 15464 15351 15466
rect 8017 15408 8022 15464
rect 8078 15408 15290 15464
rect 15346 15408 15351 15464
rect 8017 15406 15351 15408
rect 8017 15403 8083 15406
rect 15285 15403 15351 15406
rect 16941 15466 17007 15469
rect 24577 15466 24643 15469
rect 16941 15464 19580 15466
rect 16941 15408 16946 15464
rect 17002 15408 19580 15464
rect 16941 15406 19580 15408
rect 16941 15403 17007 15406
rect 18137 15330 18203 15333
rect 19333 15330 19399 15333
rect 18137 15328 19399 15330
rect 18137 15272 18142 15328
rect 18198 15272 19338 15328
rect 19394 15272 19399 15328
rect 18137 15270 19399 15272
rect 19520 15330 19580 15406
rect 23982 15464 24643 15466
rect 23982 15408 24582 15464
rect 24638 15408 24643 15464
rect 23982 15406 24643 15408
rect 23982 15330 24042 15406
rect 24577 15403 24643 15406
rect 19520 15270 24042 15330
rect 18137 15267 18203 15270
rect 19333 15267 19399 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 24761 15194 24827 15197
rect 27520 15194 28000 15224
rect 24761 15192 28000 15194
rect 24761 15136 24766 15192
rect 24822 15136 28000 15192
rect 24761 15134 28000 15136
rect 24761 15131 24827 15134
rect 27520 15104 28000 15134
rect 10593 15058 10659 15061
rect 19057 15058 19123 15061
rect 4846 15056 10659 15058
rect 4846 15000 10598 15056
rect 10654 15000 10659 15056
rect 4846 14998 10659 15000
rect 10593 14995 10659 14998
rect 14460 15056 19123 15058
rect 14460 15000 19062 15056
rect 19118 15000 19123 15056
rect 14460 14998 19123 15000
rect 0 14922 480 14952
rect 5390 14922 5396 14924
rect 0 14862 5396 14922
rect 0 14832 480 14862
rect 5390 14860 5396 14862
rect 5460 14860 5466 14924
rect 5993 14922 6059 14925
rect 14460 14922 14520 14998
rect 19057 14995 19123 14998
rect 23473 15058 23539 15061
rect 25405 15058 25471 15061
rect 23473 15056 25471 15058
rect 23473 15000 23478 15056
rect 23534 15000 25410 15056
rect 25466 15000 25471 15056
rect 23473 14998 25471 15000
rect 23473 14995 23539 14998
rect 25405 14995 25471 14998
rect 23197 14922 23263 14925
rect 5993 14920 14520 14922
rect 5993 14864 5998 14920
rect 6054 14864 14520 14920
rect 5993 14862 14520 14864
rect 14598 14920 23263 14922
rect 14598 14864 23202 14920
rect 23258 14864 23263 14920
rect 14598 14862 23263 14864
rect 5993 14859 6059 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 2313 14650 2379 14653
rect 4654 14650 4660 14652
rect 2313 14648 4660 14650
rect 2313 14592 2318 14648
rect 2374 14592 4660 14648
rect 2313 14590 4660 14592
rect 2313 14587 2379 14590
rect 4654 14588 4660 14590
rect 4724 14588 4730 14652
rect 9213 14650 9279 14653
rect 14598 14650 14658 14862
rect 23197 14859 23263 14862
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 9213 14648 9506 14650
rect 9213 14592 9218 14648
rect 9274 14616 9506 14648
rect 9274 14592 9552 14616
rect 9213 14590 9552 14592
rect 9213 14587 9279 14590
rect 9446 14556 9552 14590
rect 9492 14548 9552 14556
rect 12804 14590 14658 14650
rect 14917 14650 14983 14653
rect 17902 14650 17908 14652
rect 14917 14648 17908 14650
rect 14917 14592 14922 14648
rect 14978 14592 17908 14648
rect 14917 14590 17908 14592
rect 9492 14514 9644 14548
rect 12804 14514 12864 14590
rect 14917 14587 14983 14590
rect 17902 14588 17908 14590
rect 17972 14588 17978 14652
rect 21449 14650 21515 14653
rect 27520 14650 28000 14680
rect 21449 14648 28000 14650
rect 21449 14592 21454 14648
rect 21510 14592 28000 14648
rect 21449 14590 28000 14592
rect 21449 14587 21515 14590
rect 27520 14560 28000 14590
rect 9492 14488 12864 14514
rect 9584 14454 12864 14488
rect 12985 14514 13051 14517
rect 13537 14514 13603 14517
rect 21909 14514 21975 14517
rect 12985 14512 21975 14514
rect 12985 14456 12990 14512
rect 13046 14456 13542 14512
rect 13598 14456 21914 14512
rect 21970 14456 21975 14512
rect 12985 14454 21975 14456
rect 12985 14451 13051 14454
rect 13537 14451 13603 14454
rect 21909 14451 21975 14454
rect 0 14378 480 14408
rect 3233 14378 3299 14381
rect 0 14376 3299 14378
rect 0 14320 3238 14376
rect 3294 14320 3299 14376
rect 0 14318 3299 14320
rect 0 14288 480 14318
rect 3233 14315 3299 14318
rect 8385 14378 8451 14381
rect 16849 14378 16915 14381
rect 8385 14376 9092 14378
rect 8385 14320 8390 14376
rect 8446 14320 9092 14376
rect 8385 14318 9092 14320
rect 8385 14315 8451 14318
rect 9032 14276 9092 14318
rect 9584 14376 16915 14378
rect 9584 14320 16854 14376
rect 16910 14320 16915 14376
rect 9584 14318 16915 14320
rect 9584 14276 9644 14318
rect 16849 14315 16915 14318
rect 9032 14216 9644 14276
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 10041 14106 10107 14109
rect 7284 14104 10107 14106
rect 7284 14048 10046 14104
rect 10102 14048 10107 14104
rect 7284 14046 10107 14048
rect 5625 13970 5691 13973
rect 7284 13970 7344 14046
rect 10041 14043 10107 14046
rect 19374 14044 19380 14108
rect 19444 14106 19450 14108
rect 23473 14106 23539 14109
rect 19444 14104 23539 14106
rect 19444 14048 23478 14104
rect 23534 14048 23539 14104
rect 19444 14046 23539 14048
rect 19444 14044 19450 14046
rect 23473 14043 23539 14046
rect 5625 13968 7344 13970
rect 5625 13912 5630 13968
rect 5686 13912 7344 13968
rect 5625 13910 7344 13912
rect 7465 13970 7531 13973
rect 16849 13970 16915 13973
rect 27520 13970 28000 14000
rect 7465 13968 28000 13970
rect 7465 13912 7470 13968
rect 7526 13912 16854 13968
rect 16910 13912 28000 13968
rect 7465 13910 28000 13912
rect 5625 13907 5691 13910
rect 7465 13907 7531 13910
rect 16849 13907 16915 13910
rect 27520 13880 28000 13910
rect 8201 13834 8267 13837
rect 10133 13834 10199 13837
rect 8201 13832 10199 13834
rect 8201 13776 8206 13832
rect 8262 13776 10138 13832
rect 10194 13776 10199 13832
rect 8201 13774 10199 13776
rect 8201 13771 8267 13774
rect 10133 13771 10199 13774
rect 18505 13834 18571 13837
rect 25221 13834 25287 13837
rect 18505 13832 25287 13834
rect 18505 13776 18510 13832
rect 18566 13776 25226 13832
rect 25282 13776 25287 13832
rect 18505 13774 25287 13776
rect 18505 13771 18571 13774
rect 25221 13771 25287 13774
rect 0 13698 480 13728
rect 3969 13698 4035 13701
rect 5993 13698 6059 13701
rect 0 13638 3112 13698
rect 0 13608 480 13638
rect 3052 13290 3112 13638
rect 3969 13696 6059 13698
rect 3969 13640 3974 13696
rect 4030 13640 5998 13696
rect 6054 13640 6059 13696
rect 3969 13638 6059 13640
rect 3969 13635 4035 13638
rect 5993 13635 6059 13638
rect 13997 13698 14063 13701
rect 15285 13698 15351 13701
rect 13997 13696 15351 13698
rect 13997 13640 14002 13696
rect 14058 13640 15290 13696
rect 15346 13640 15351 13696
rect 13997 13638 15351 13640
rect 13997 13635 14063 13638
rect 15285 13635 15351 13638
rect 20897 13698 20963 13701
rect 25037 13698 25103 13701
rect 20897 13696 25103 13698
rect 20897 13640 20902 13696
rect 20958 13640 25042 13696
rect 25098 13640 25103 13696
rect 20897 13638 25103 13640
rect 20897 13635 20963 13638
rect 25037 13635 25103 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 13905 13562 13971 13565
rect 17861 13562 17927 13565
rect 13905 13560 17927 13562
rect 13905 13504 13910 13560
rect 13966 13504 17866 13560
rect 17922 13504 17927 13560
rect 13905 13502 17927 13504
rect 13905 13499 13971 13502
rect 17861 13499 17927 13502
rect 20529 13562 20595 13565
rect 25773 13562 25839 13565
rect 20529 13560 25839 13562
rect 20529 13504 20534 13560
rect 20590 13504 25778 13560
rect 25834 13504 25839 13560
rect 20529 13502 25839 13504
rect 20529 13499 20595 13502
rect 25773 13499 25839 13502
rect 3233 13426 3299 13429
rect 8201 13426 8267 13429
rect 3233 13424 8267 13426
rect 3233 13368 3238 13424
rect 3294 13368 8206 13424
rect 8262 13368 8267 13424
rect 3233 13366 8267 13368
rect 3233 13363 3299 13366
rect 8201 13363 8267 13366
rect 8385 13426 8451 13429
rect 13445 13426 13511 13429
rect 8385 13424 13511 13426
rect 8385 13368 8390 13424
rect 8446 13368 13450 13424
rect 13506 13368 13511 13424
rect 8385 13366 13511 13368
rect 8385 13363 8451 13366
rect 13445 13363 13511 13366
rect 17217 13426 17283 13429
rect 19333 13426 19399 13429
rect 17217 13424 19399 13426
rect 17217 13368 17222 13424
rect 17278 13368 19338 13424
rect 19394 13368 19399 13424
rect 17217 13366 19399 13368
rect 17217 13363 17283 13366
rect 19333 13363 19399 13366
rect 24853 13426 24919 13429
rect 27520 13426 28000 13456
rect 24853 13424 28000 13426
rect 24853 13368 24858 13424
rect 24914 13368 28000 13424
rect 24853 13366 28000 13368
rect 24853 13363 24919 13366
rect 27520 13336 28000 13366
rect 13905 13290 13971 13293
rect 3052 13288 13971 13290
rect 3052 13232 13910 13288
rect 13966 13232 13971 13288
rect 3052 13230 13971 13232
rect 13905 13227 13971 13230
rect 15377 13290 15443 13293
rect 20989 13290 21055 13293
rect 15377 13288 21055 13290
rect 15377 13232 15382 13288
rect 15438 13232 20994 13288
rect 21050 13232 21055 13288
rect 15377 13230 21055 13232
rect 15377 13227 15443 13230
rect 20989 13227 21055 13230
rect 0 13154 480 13184
rect 4061 13154 4127 13157
rect 0 13152 4127 13154
rect 0 13096 4066 13152
rect 4122 13096 4127 13152
rect 0 13094 4127 13096
rect 0 13064 480 13094
rect 4061 13091 4127 13094
rect 10777 13154 10843 13157
rect 13445 13154 13511 13157
rect 10777 13152 13511 13154
rect 10777 13096 10782 13152
rect 10838 13096 13450 13152
rect 13506 13096 13511 13152
rect 10777 13094 13511 13096
rect 10777 13091 10843 13094
rect 13445 13091 13511 13094
rect 17902 13092 17908 13156
rect 17972 13154 17978 13156
rect 19977 13154 20043 13157
rect 17972 13152 20043 13154
rect 17972 13096 19982 13152
rect 20038 13096 20043 13152
rect 17972 13094 20043 13096
rect 17972 13092 17978 13094
rect 19977 13091 20043 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 2773 13018 2839 13021
rect 3141 13018 3207 13021
rect 2773 13016 3207 13018
rect 2773 12960 2778 13016
rect 2834 12960 3146 13016
rect 3202 12960 3207 13016
rect 2773 12958 3207 12960
rect 2773 12955 2839 12958
rect 3141 12955 3207 12958
rect 6453 13018 6519 13021
rect 10685 13018 10751 13021
rect 11094 13018 11100 13020
rect 6453 13016 11100 13018
rect 6453 12960 6458 13016
rect 6514 12960 10690 13016
rect 10746 12960 11100 13016
rect 6453 12958 11100 12960
rect 6453 12955 6519 12958
rect 10685 12955 10751 12958
rect 11094 12956 11100 12958
rect 11164 13018 11170 13020
rect 11421 13018 11487 13021
rect 11164 13016 11487 13018
rect 11164 12960 11426 13016
rect 11482 12960 11487 13016
rect 11164 12958 11487 12960
rect 11164 12956 11170 12958
rect 11421 12955 11487 12958
rect 2221 12882 2287 12885
rect 5533 12882 5599 12885
rect 15929 12882 15995 12885
rect 2221 12880 5599 12882
rect 2221 12824 2226 12880
rect 2282 12824 5538 12880
rect 5594 12824 5599 12880
rect 2221 12822 5599 12824
rect 2221 12819 2287 12822
rect 5533 12819 5599 12822
rect 7790 12880 15995 12882
rect 7790 12824 15934 12880
rect 15990 12824 15995 12880
rect 7790 12822 15995 12824
rect 4061 12746 4127 12749
rect 7557 12746 7623 12749
rect 4061 12744 7623 12746
rect 4061 12688 4066 12744
rect 4122 12688 7562 12744
rect 7618 12688 7623 12744
rect 4061 12686 7623 12688
rect 4061 12683 4127 12686
rect 7557 12683 7623 12686
rect 0 12610 480 12640
rect 4613 12610 4679 12613
rect 7790 12610 7850 12822
rect 15929 12819 15995 12822
rect 23606 12820 23612 12884
rect 23676 12882 23682 12884
rect 27520 12882 28000 12912
rect 23676 12822 28000 12882
rect 23676 12820 23682 12822
rect 27520 12792 28000 12822
rect 8201 12746 8267 12749
rect 17493 12746 17559 12749
rect 18321 12746 18387 12749
rect 8201 12744 18387 12746
rect 8201 12688 8206 12744
rect 8262 12688 17498 12744
rect 17554 12688 18326 12744
rect 18382 12688 18387 12744
rect 8201 12686 18387 12688
rect 8201 12683 8267 12686
rect 17493 12683 17559 12686
rect 18321 12683 18387 12686
rect 0 12608 4679 12610
rect 0 12552 4618 12608
rect 4674 12552 4679 12608
rect 0 12550 4679 12552
rect 0 12520 480 12550
rect 4613 12547 4679 12550
rect 4800 12550 7850 12610
rect 10869 12610 10935 12613
rect 12985 12610 13051 12613
rect 10869 12608 13051 12610
rect 10869 12552 10874 12608
rect 10930 12552 12990 12608
rect 13046 12552 13051 12608
rect 10869 12550 13051 12552
rect 3693 12474 3759 12477
rect 4800 12474 4860 12550
rect 10869 12547 10935 12550
rect 12985 12547 13051 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 3693 12472 4860 12474
rect 3693 12416 3698 12472
rect 3754 12416 4860 12472
rect 3693 12414 4860 12416
rect 6637 12474 6703 12477
rect 9857 12474 9923 12477
rect 6637 12472 9923 12474
rect 6637 12416 6642 12472
rect 6698 12416 9862 12472
rect 9918 12416 9923 12472
rect 6637 12414 9923 12416
rect 3693 12411 3759 12414
rect 6637 12411 6703 12414
rect 9857 12411 9923 12414
rect 10685 12474 10751 12477
rect 12433 12474 12499 12477
rect 10685 12472 12499 12474
rect 10685 12416 10690 12472
rect 10746 12416 12438 12472
rect 12494 12416 12499 12472
rect 10685 12414 12499 12416
rect 10685 12411 10751 12414
rect 12433 12411 12499 12414
rect 2589 12338 2655 12341
rect 3785 12338 3851 12341
rect 2589 12336 3851 12338
rect 2589 12280 2594 12336
rect 2650 12280 3790 12336
rect 3846 12280 3851 12336
rect 2589 12278 3851 12280
rect 2589 12275 2655 12278
rect 3785 12275 3851 12278
rect 4613 12340 4679 12341
rect 4613 12336 4660 12340
rect 4724 12338 4730 12340
rect 7281 12338 7347 12341
rect 12801 12338 12867 12341
rect 13169 12338 13235 12341
rect 14641 12338 14707 12341
rect 18229 12338 18295 12341
rect 18873 12338 18939 12341
rect 4613 12280 4618 12336
rect 4613 12276 4660 12280
rect 4724 12278 4770 12338
rect 7281 12336 12867 12338
rect 7281 12280 7286 12336
rect 7342 12280 12806 12336
rect 12862 12280 12867 12336
rect 7281 12278 12867 12280
rect 4724 12276 4730 12278
rect 4613 12275 4679 12276
rect 7281 12275 7347 12278
rect 12801 12275 12867 12278
rect 13126 12336 14707 12338
rect 13126 12280 13174 12336
rect 13230 12280 14646 12336
rect 14702 12280 14707 12336
rect 13126 12278 14707 12280
rect 13126 12275 13235 12278
rect 14641 12275 14707 12278
rect 14782 12336 18939 12338
rect 14782 12280 18234 12336
rect 18290 12280 18878 12336
rect 18934 12280 18939 12336
rect 14782 12278 18939 12280
rect 6821 12202 6887 12205
rect 7649 12202 7715 12205
rect 9213 12202 9279 12205
rect 6821 12200 9279 12202
rect 6821 12144 6826 12200
rect 6882 12144 7654 12200
rect 7710 12144 9218 12200
rect 9274 12144 9279 12200
rect 6821 12142 9279 12144
rect 6821 12139 6887 12142
rect 7649 12139 7715 12142
rect 9213 12139 9279 12142
rect 11421 12202 11487 12205
rect 13126 12202 13186 12275
rect 11421 12200 13186 12202
rect 11421 12144 11426 12200
rect 11482 12144 13186 12200
rect 11421 12142 13186 12144
rect 11421 12139 11487 12142
rect 0 12066 480 12096
rect 1485 12066 1551 12069
rect 0 12064 1551 12066
rect 0 12008 1490 12064
rect 1546 12008 1551 12064
rect 0 12006 1551 12008
rect 0 11976 480 12006
rect 1485 12003 1551 12006
rect 6729 12066 6795 12069
rect 9857 12066 9923 12069
rect 14457 12066 14523 12069
rect 6729 12064 9923 12066
rect 6729 12008 6734 12064
rect 6790 12008 9862 12064
rect 9918 12008 9923 12064
rect 6729 12006 9923 12008
rect 6729 12003 6795 12006
rect 9857 12003 9923 12006
rect 10734 12064 14523 12066
rect 10734 12008 14462 12064
rect 14518 12008 14523 12064
rect 10734 12006 14523 12008
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 2814 11732 2820 11796
rect 2884 11794 2890 11796
rect 4245 11794 4311 11797
rect 10734 11794 10794 12006
rect 14457 12003 14523 12006
rect 10869 11930 10935 11933
rect 14782 11930 14842 12278
rect 18229 12275 18295 12278
rect 18873 12275 18939 12278
rect 19374 12276 19380 12340
rect 19444 12338 19450 12340
rect 19517 12338 19583 12341
rect 19444 12336 19583 12338
rect 19444 12280 19522 12336
rect 19578 12280 19583 12336
rect 19444 12278 19583 12280
rect 19444 12276 19450 12278
rect 19517 12275 19583 12278
rect 23422 12276 23428 12340
rect 23492 12338 23498 12340
rect 27520 12338 28000 12368
rect 23492 12278 28000 12338
rect 23492 12276 23498 12278
rect 27520 12248 28000 12278
rect 14917 12202 14983 12205
rect 16849 12202 16915 12205
rect 20161 12202 20227 12205
rect 14917 12200 15394 12202
rect 14917 12144 14922 12200
rect 14978 12144 15394 12200
rect 14917 12142 15394 12144
rect 14917 12139 14983 12142
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 10869 11928 14842 11930
rect 10869 11872 10874 11928
rect 10930 11872 14842 11928
rect 10869 11870 14842 11872
rect 15334 11930 15394 12142
rect 16849 12200 20227 12202
rect 16849 12144 16854 12200
rect 16910 12144 20166 12200
rect 20222 12144 20227 12200
rect 16849 12142 20227 12144
rect 16849 12139 16915 12142
rect 20161 12139 20227 12142
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 23933 11930 23999 11933
rect 15334 11928 23999 11930
rect 15334 11872 23938 11928
rect 23994 11872 23999 11928
rect 15334 11870 23999 11872
rect 10869 11867 10935 11870
rect 16990 11797 17050 11870
rect 23933 11867 23999 11870
rect 2884 11792 4311 11794
rect 2884 11736 4250 11792
rect 4306 11736 4311 11792
rect 2884 11734 4311 11736
rect 2884 11732 2890 11734
rect 4245 11731 4311 11734
rect 7560 11734 10794 11794
rect 12801 11794 12867 11797
rect 15745 11794 15811 11797
rect 12801 11792 15811 11794
rect 12801 11736 12806 11792
rect 12862 11736 15750 11792
rect 15806 11736 15811 11792
rect 12801 11734 15811 11736
rect 0 11522 480 11552
rect 7560 11522 7620 11734
rect 12801 11731 12867 11734
rect 15745 11731 15811 11734
rect 16941 11792 17050 11797
rect 16941 11736 16946 11792
rect 17002 11736 17050 11792
rect 16941 11734 17050 11736
rect 18045 11794 18111 11797
rect 23749 11794 23815 11797
rect 27520 11794 28000 11824
rect 18045 11792 22340 11794
rect 18045 11736 18050 11792
rect 18106 11736 22340 11792
rect 18045 11734 22340 11736
rect 16941 11731 17007 11734
rect 18045 11731 18111 11734
rect 9581 11658 9647 11661
rect 11237 11658 11303 11661
rect 9581 11656 11303 11658
rect 9581 11600 9586 11656
rect 9642 11600 11242 11656
rect 11298 11600 11303 11656
rect 9581 11598 11303 11600
rect 9581 11595 9647 11598
rect 11237 11595 11303 11598
rect 14365 11658 14431 11661
rect 21909 11658 21975 11661
rect 14365 11656 21975 11658
rect 14365 11600 14370 11656
rect 14426 11600 21914 11656
rect 21970 11600 21975 11656
rect 14365 11598 21975 11600
rect 22280 11658 22340 11734
rect 23749 11792 28000 11794
rect 23749 11736 23754 11792
rect 23810 11736 28000 11792
rect 23749 11734 28000 11736
rect 23749 11731 23815 11734
rect 27520 11704 28000 11734
rect 25221 11658 25287 11661
rect 22280 11656 25287 11658
rect 22280 11600 25226 11656
rect 25282 11600 25287 11656
rect 22280 11598 25287 11600
rect 14365 11595 14431 11598
rect 21909 11595 21975 11598
rect 25221 11595 25287 11598
rect 0 11462 7620 11522
rect 11145 11522 11211 11525
rect 12341 11522 12407 11525
rect 14825 11522 14891 11525
rect 11145 11520 14891 11522
rect 11145 11464 11150 11520
rect 11206 11464 12346 11520
rect 12402 11464 14830 11520
rect 14886 11464 14891 11520
rect 11145 11462 14891 11464
rect 0 11432 480 11462
rect 11145 11459 11211 11462
rect 12341 11459 12407 11462
rect 14825 11459 14891 11462
rect 15101 11522 15167 11525
rect 17585 11522 17651 11525
rect 15101 11520 17651 11522
rect 15101 11464 15106 11520
rect 15162 11464 17590 11520
rect 17646 11464 17651 11520
rect 15101 11462 17651 11464
rect 15101 11459 15167 11462
rect 17585 11459 17651 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 2865 11386 2931 11389
rect 3785 11386 3851 11389
rect 2865 11384 3851 11386
rect 2865 11328 2870 11384
rect 2926 11328 3790 11384
rect 3846 11328 3851 11384
rect 2865 11326 3851 11328
rect 2865 11323 2931 11326
rect 3785 11323 3851 11326
rect 6177 11386 6243 11389
rect 9765 11386 9831 11389
rect 9949 11388 10015 11389
rect 9949 11386 9996 11388
rect 6177 11384 9831 11386
rect 6177 11328 6182 11384
rect 6238 11328 9770 11384
rect 9826 11328 9831 11384
rect 6177 11326 9831 11328
rect 9904 11384 9996 11386
rect 9904 11328 9954 11384
rect 9904 11326 9996 11328
rect 6177 11323 6243 11326
rect 9765 11323 9831 11326
rect 9949 11324 9996 11326
rect 10060 11324 10066 11388
rect 9949 11323 10015 11324
rect 3693 11250 3759 11253
rect 4429 11250 4495 11253
rect 3693 11248 4495 11250
rect 3693 11192 3698 11248
rect 3754 11192 4434 11248
rect 4490 11192 4495 11248
rect 3693 11190 4495 11192
rect 3693 11187 3759 11190
rect 4429 11187 4495 11190
rect 9581 11250 9647 11253
rect 14825 11250 14891 11253
rect 9581 11248 14891 11250
rect 9581 11192 9586 11248
rect 9642 11192 14830 11248
rect 14886 11192 14891 11248
rect 9581 11190 14891 11192
rect 9581 11187 9647 11190
rect 14825 11187 14891 11190
rect 16113 11250 16179 11253
rect 20161 11250 20227 11253
rect 16113 11248 20227 11250
rect 16113 11192 16118 11248
rect 16174 11192 20166 11248
rect 20222 11192 20227 11248
rect 16113 11190 20227 11192
rect 16113 11187 16179 11190
rect 20161 11187 20227 11190
rect 1485 11114 1551 11117
rect 10869 11114 10935 11117
rect 1485 11112 10935 11114
rect 1485 11056 1490 11112
rect 1546 11056 10874 11112
rect 10930 11056 10935 11112
rect 1485 11054 10935 11056
rect 1485 11051 1551 11054
rect 10869 11051 10935 11054
rect 14774 11052 14780 11116
rect 14844 11114 14850 11116
rect 14917 11114 14983 11117
rect 14844 11112 14983 11114
rect 14844 11056 14922 11112
rect 14978 11056 14983 11112
rect 14844 11054 14983 11056
rect 14844 11052 14850 11054
rect 14917 11051 14983 11054
rect 16021 11114 16087 11117
rect 22001 11114 22067 11117
rect 16021 11112 22067 11114
rect 16021 11056 16026 11112
rect 16082 11056 22006 11112
rect 22062 11056 22067 11112
rect 16021 11054 22067 11056
rect 16021 11051 16087 11054
rect 22001 11051 22067 11054
rect 23657 11114 23723 11117
rect 27520 11114 28000 11144
rect 23657 11112 28000 11114
rect 23657 11056 23662 11112
rect 23718 11056 28000 11112
rect 23657 11054 28000 11056
rect 23657 11051 23723 11054
rect 27520 11024 28000 11054
rect 0 10978 480 11008
rect 5349 10978 5415 10981
rect 0 10976 5415 10978
rect 0 10920 5354 10976
rect 5410 10920 5415 10976
rect 0 10918 5415 10920
rect 0 10888 480 10918
rect 5349 10915 5415 10918
rect 8293 10978 8359 10981
rect 9305 10978 9371 10981
rect 16021 10978 16087 10981
rect 8293 10976 14842 10978
rect 8293 10920 8298 10976
rect 8354 10920 9310 10976
rect 9366 10920 14842 10976
rect 8293 10918 14842 10920
rect 8293 10915 8359 10918
rect 9305 10915 9371 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 13353 10706 13419 10709
rect 3374 10704 13419 10706
rect 3374 10648 13358 10704
rect 13414 10648 13419 10704
rect 3374 10646 13419 10648
rect 14782 10706 14842 10918
rect 16021 10976 24042 10978
rect 16021 10920 16026 10976
rect 16082 10920 24042 10976
rect 16021 10918 24042 10920
rect 16021 10915 16087 10918
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 15837 10842 15903 10845
rect 18597 10842 18663 10845
rect 15837 10840 18663 10842
rect 15837 10784 15842 10840
rect 15898 10784 18602 10840
rect 18658 10784 18663 10840
rect 15837 10782 18663 10784
rect 15837 10779 15903 10782
rect 18597 10779 18663 10782
rect 17401 10706 17467 10709
rect 14782 10704 17467 10706
rect 14782 10648 17406 10704
rect 17462 10648 17467 10704
rect 14782 10646 17467 10648
rect 0 10434 480 10464
rect 3374 10434 3434 10646
rect 13353 10643 13419 10646
rect 17401 10643 17467 10646
rect 18137 10706 18203 10709
rect 22369 10706 22435 10709
rect 18137 10704 22435 10706
rect 18137 10648 18142 10704
rect 18198 10648 22374 10704
rect 22430 10648 22435 10704
rect 18137 10646 22435 10648
rect 18137 10643 18203 10646
rect 22369 10643 22435 10646
rect 5349 10570 5415 10573
rect 7557 10570 7623 10573
rect 8477 10570 8543 10573
rect 21081 10570 21147 10573
rect 5349 10568 8543 10570
rect 5349 10512 5354 10568
rect 5410 10512 7562 10568
rect 7618 10512 8482 10568
rect 8538 10512 8543 10568
rect 5349 10510 8543 10512
rect 5349 10507 5415 10510
rect 7557 10507 7623 10510
rect 8477 10507 8543 10510
rect 8710 10568 21147 10570
rect 8710 10512 21086 10568
rect 21142 10512 21147 10568
rect 8710 10510 21147 10512
rect 23982 10570 24042 10918
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 27520 10570 28000 10600
rect 23982 10510 28000 10570
rect 0 10374 3434 10434
rect 3509 10434 3575 10437
rect 6453 10434 6519 10437
rect 3509 10432 6519 10434
rect 3509 10376 3514 10432
rect 3570 10376 6458 10432
rect 6514 10376 6519 10432
rect 3509 10374 6519 10376
rect 0 10344 480 10374
rect 3509 10371 3575 10374
rect 6453 10371 6519 10374
rect 6729 10434 6795 10437
rect 8710 10434 8770 10510
rect 21081 10507 21147 10510
rect 27520 10480 28000 10510
rect 6729 10432 8770 10434
rect 6729 10376 6734 10432
rect 6790 10376 8770 10432
rect 6729 10374 8770 10376
rect 12433 10434 12499 10437
rect 13997 10434 14063 10437
rect 16021 10434 16087 10437
rect 12433 10432 16087 10434
rect 12433 10376 12438 10432
rect 12494 10376 14002 10432
rect 14058 10376 16026 10432
rect 16082 10376 16087 10432
rect 12433 10374 16087 10376
rect 6729 10371 6795 10374
rect 12433 10371 12499 10374
rect 13997 10371 14063 10374
rect 16021 10371 16087 10374
rect 16297 10434 16363 10437
rect 18137 10434 18203 10437
rect 16297 10432 18203 10434
rect 16297 10376 16302 10432
rect 16358 10376 18142 10432
rect 18198 10376 18203 10432
rect 16297 10374 18203 10376
rect 16297 10371 16363 10374
rect 18137 10371 18203 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 2865 10298 2931 10301
rect 8293 10298 8359 10301
rect 2865 10296 8359 10298
rect 2865 10240 2870 10296
rect 2926 10240 8298 10296
rect 8354 10240 8359 10296
rect 2865 10238 8359 10240
rect 2865 10235 2931 10238
rect 8293 10235 8359 10238
rect 15285 10298 15351 10301
rect 19057 10298 19123 10301
rect 19425 10298 19491 10301
rect 15285 10296 19491 10298
rect 15285 10240 15290 10296
rect 15346 10240 19062 10296
rect 19118 10240 19430 10296
rect 19486 10240 19491 10296
rect 15285 10238 19491 10240
rect 15285 10235 15351 10238
rect 19057 10235 19123 10238
rect 19425 10235 19491 10238
rect 2221 10162 2287 10165
rect 4245 10162 4311 10165
rect 2221 10160 4311 10162
rect 2221 10104 2226 10160
rect 2282 10104 4250 10160
rect 4306 10104 4311 10160
rect 2221 10102 4311 10104
rect 2221 10099 2287 10102
rect 4245 10099 4311 10102
rect 5349 10162 5415 10165
rect 11973 10162 12039 10165
rect 5349 10160 12039 10162
rect 5349 10104 5354 10160
rect 5410 10104 11978 10160
rect 12034 10104 12039 10160
rect 5349 10102 12039 10104
rect 5349 10099 5415 10102
rect 11973 10099 12039 10102
rect 12157 10162 12223 10165
rect 17401 10162 17467 10165
rect 12157 10160 17467 10162
rect 12157 10104 12162 10160
rect 12218 10104 17406 10160
rect 17462 10104 17467 10160
rect 12157 10102 17467 10104
rect 12157 10099 12223 10102
rect 17401 10099 17467 10102
rect 2405 10026 2471 10029
rect 16113 10026 16179 10029
rect 2405 10024 16179 10026
rect 2405 9968 2410 10024
rect 2466 9968 16118 10024
rect 16174 9968 16179 10024
rect 2405 9966 16179 9968
rect 2405 9963 2471 9966
rect 16113 9963 16179 9966
rect 23974 9964 23980 10028
rect 24044 10026 24050 10028
rect 27520 10026 28000 10056
rect 24044 9966 28000 10026
rect 24044 9964 24050 9966
rect 27520 9936 28000 9966
rect 0 9890 480 9920
rect 5349 9890 5415 9893
rect 0 9888 5415 9890
rect 0 9832 5354 9888
rect 5410 9832 5415 9888
rect 0 9830 5415 9832
rect 0 9800 480 9830
rect 5349 9827 5415 9830
rect 6453 9890 6519 9893
rect 12157 9890 12223 9893
rect 18873 9892 18939 9893
rect 6453 9888 12223 9890
rect 6453 9832 6458 9888
rect 6514 9832 12162 9888
rect 12218 9832 12223 9888
rect 6453 9830 12223 9832
rect 6453 9827 6519 9830
rect 12157 9827 12223 9830
rect 18822 9828 18828 9892
rect 18892 9890 18939 9892
rect 18892 9888 18984 9890
rect 18934 9832 18984 9888
rect 18892 9830 18984 9832
rect 18892 9828 18939 9830
rect 18873 9827 18939 9828
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 2405 9754 2471 9757
rect 3325 9754 3391 9757
rect 7465 9754 7531 9757
rect 2405 9752 3391 9754
rect 2405 9696 2410 9752
rect 2466 9696 3330 9752
rect 3386 9696 3391 9752
rect 2405 9694 3391 9696
rect 2405 9691 2471 9694
rect 3325 9691 3391 9694
rect 7422 9752 7531 9754
rect 7422 9696 7470 9752
rect 7526 9696 7531 9752
rect 7422 9691 7531 9696
rect 19241 9754 19307 9757
rect 21265 9754 21331 9757
rect 19241 9752 21331 9754
rect 19241 9696 19246 9752
rect 19302 9696 21270 9752
rect 21326 9696 21331 9752
rect 19241 9694 21331 9696
rect 19241 9691 19307 9694
rect 21265 9691 21331 9694
rect 7422 9349 7482 9691
rect 8017 9618 8083 9621
rect 10593 9618 10659 9621
rect 8017 9616 10659 9618
rect 8017 9560 8022 9616
rect 8078 9560 10598 9616
rect 10654 9560 10659 9616
rect 8017 9558 10659 9560
rect 8017 9555 8083 9558
rect 10593 9555 10659 9558
rect 13353 9618 13419 9621
rect 18505 9618 18571 9621
rect 20897 9618 20963 9621
rect 13353 9616 18154 9618
rect 13353 9560 13358 9616
rect 13414 9560 18154 9616
rect 13353 9558 18154 9560
rect 13353 9555 13419 9558
rect 9121 9482 9187 9485
rect 9489 9482 9555 9485
rect 14917 9482 14983 9485
rect 17769 9482 17835 9485
rect 9121 9480 17835 9482
rect 9121 9424 9126 9480
rect 9182 9424 9494 9480
rect 9550 9424 14922 9480
rect 14978 9424 17774 9480
rect 17830 9424 17835 9480
rect 9121 9422 17835 9424
rect 18094 9482 18154 9558
rect 18505 9616 20963 9618
rect 18505 9560 18510 9616
rect 18566 9560 20902 9616
rect 20958 9560 20963 9616
rect 18505 9558 20963 9560
rect 18505 9555 18571 9558
rect 20897 9555 20963 9558
rect 18505 9482 18571 9485
rect 22461 9482 22527 9485
rect 18094 9480 22527 9482
rect 18094 9424 18510 9480
rect 18566 9424 22466 9480
rect 22522 9424 22527 9480
rect 18094 9422 22527 9424
rect 9121 9419 9187 9422
rect 9489 9419 9555 9422
rect 14917 9419 14983 9422
rect 17769 9419 17835 9422
rect 18505 9419 18571 9422
rect 22461 9419 22527 9422
rect 23974 9420 23980 9484
rect 24044 9482 24050 9484
rect 27520 9482 28000 9512
rect 24044 9422 28000 9482
rect 24044 9420 24050 9422
rect 27520 9392 28000 9422
rect 3141 9346 3207 9349
rect 1396 9344 3207 9346
rect 1396 9288 3146 9344
rect 3202 9288 3207 9344
rect 1396 9286 3207 9288
rect 0 9210 480 9240
rect 1396 9210 1456 9286
rect 3141 9283 3207 9286
rect 7373 9344 7482 9349
rect 7373 9288 7378 9344
rect 7434 9288 7482 9344
rect 7373 9286 7482 9288
rect 22093 9346 22159 9349
rect 22093 9344 22202 9346
rect 22093 9288 22098 9344
rect 22154 9288 22202 9344
rect 7373 9283 7439 9286
rect 22093 9283 22202 9288
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 12157 9210 12223 9213
rect 18137 9210 18203 9213
rect 0 9150 1456 9210
rect 10688 9208 18203 9210
rect 10688 9152 12162 9208
rect 12218 9152 18142 9208
rect 18198 9152 18203 9208
rect 10688 9150 18203 9152
rect 0 9120 480 9150
rect 3601 9074 3667 9077
rect 10688 9074 10748 9150
rect 12157 9147 12223 9150
rect 18137 9147 18203 9150
rect 21081 9210 21147 9213
rect 21214 9210 21220 9212
rect 21081 9208 21220 9210
rect 21081 9152 21086 9208
rect 21142 9152 21220 9208
rect 21081 9150 21220 9152
rect 21081 9147 21147 9150
rect 21214 9148 21220 9150
rect 21284 9148 21290 9212
rect 22142 9210 22202 9283
rect 22277 9210 22343 9213
rect 23381 9210 23447 9213
rect 22142 9208 23447 9210
rect 22142 9152 22282 9208
rect 22338 9152 23386 9208
rect 23442 9152 23447 9208
rect 22142 9150 23447 9152
rect 22277 9147 22343 9150
rect 23381 9147 23447 9150
rect 15469 9074 15535 9077
rect 3601 9072 10748 9074
rect 3601 9016 3606 9072
rect 3662 9016 10748 9072
rect 3601 9014 10748 9016
rect 14644 9072 15535 9074
rect 14644 9016 15474 9072
rect 15530 9016 15535 9072
rect 14644 9014 15535 9016
rect 3601 9011 3667 9014
rect 2957 8938 3023 8941
rect 3325 8938 3391 8941
rect 10777 8938 10843 8941
rect 12433 8938 12499 8941
rect 2957 8936 6194 8938
rect 2957 8880 2962 8936
rect 3018 8880 3330 8936
rect 3386 8880 6194 8936
rect 2957 8878 6194 8880
rect 2957 8875 3023 8878
rect 3325 8875 3391 8878
rect 5610 8736 5930 8737
rect 0 8666 480 8696
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 4061 8666 4127 8669
rect 0 8664 4127 8666
rect 0 8608 4066 8664
rect 4122 8608 4127 8664
rect 0 8606 4127 8608
rect 0 8576 480 8606
rect 4061 8603 4127 8606
rect 4705 8666 4771 8669
rect 4838 8666 4844 8668
rect 4705 8664 4844 8666
rect 4705 8608 4710 8664
rect 4766 8608 4844 8664
rect 4705 8606 4844 8608
rect 4705 8603 4771 8606
rect 4838 8604 4844 8606
rect 4908 8604 4914 8668
rect 6134 8666 6194 8878
rect 10777 8936 12499 8938
rect 10777 8880 10782 8936
rect 10838 8880 12438 8936
rect 12494 8880 12499 8936
rect 10777 8878 12499 8880
rect 10777 8875 10843 8878
rect 12433 8875 12499 8878
rect 12709 8940 12775 8941
rect 12709 8936 12756 8940
rect 12820 8938 12826 8940
rect 12709 8880 12714 8936
rect 12709 8876 12756 8880
rect 12820 8878 12866 8938
rect 12820 8876 12826 8878
rect 12709 8875 12775 8876
rect 10777 8802 10843 8805
rect 14644 8802 14704 9014
rect 15469 9011 15535 9014
rect 16021 9074 16087 9077
rect 23606 9074 23612 9076
rect 16021 9072 23612 9074
rect 16021 9016 16026 9072
rect 16082 9016 23612 9072
rect 16021 9014 23612 9016
rect 16021 9011 16087 9014
rect 23606 9012 23612 9014
rect 23676 9012 23682 9076
rect 15653 8938 15719 8941
rect 10777 8800 14704 8802
rect 10777 8744 10782 8800
rect 10838 8744 14704 8800
rect 10777 8742 14704 8744
rect 14782 8936 15719 8938
rect 14782 8880 15658 8936
rect 15714 8880 15719 8936
rect 14782 8878 15719 8880
rect 10777 8739 10843 8742
rect 14782 8666 14842 8878
rect 15653 8875 15719 8878
rect 19057 8938 19123 8941
rect 21357 8938 21423 8941
rect 19057 8936 21423 8938
rect 19057 8880 19062 8936
rect 19118 8880 21362 8936
rect 21418 8880 21423 8936
rect 19057 8878 21423 8880
rect 19057 8875 19123 8878
rect 21357 8875 21423 8878
rect 23565 8938 23631 8941
rect 27520 8938 28000 8968
rect 23565 8936 28000 8938
rect 23565 8880 23570 8936
rect 23626 8880 28000 8936
rect 23565 8878 28000 8880
rect 23565 8875 23631 8878
rect 27520 8848 28000 8878
rect 21173 8800 21239 8805
rect 21173 8744 21178 8800
rect 21234 8744 21239 8800
rect 21173 8739 21239 8744
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 6134 8606 14842 8666
rect 16849 8666 16915 8669
rect 21176 8666 21236 8739
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 16849 8664 21236 8666
rect 16849 8608 16854 8664
rect 16910 8608 21236 8664
rect 16849 8606 21236 8608
rect 16849 8603 16915 8606
rect 4337 8530 4403 8533
rect 15285 8530 15351 8533
rect 4337 8528 15351 8530
rect 4337 8472 4342 8528
rect 4398 8472 15290 8528
rect 15346 8472 15351 8528
rect 4337 8470 15351 8472
rect 4337 8467 4403 8470
rect 15285 8467 15351 8470
rect 15878 8468 15884 8532
rect 15948 8530 15954 8532
rect 16021 8530 16087 8533
rect 15948 8528 16087 8530
rect 15948 8472 16026 8528
rect 16082 8472 16087 8528
rect 15948 8470 16087 8472
rect 15948 8468 15954 8470
rect 16021 8467 16087 8470
rect 3877 8394 3943 8397
rect 6862 8394 6868 8396
rect 3877 8392 6868 8394
rect 3877 8336 3882 8392
rect 3938 8336 6868 8392
rect 3877 8334 6868 8336
rect 3877 8331 3943 8334
rect 6862 8332 6868 8334
rect 6932 8332 6938 8396
rect 12709 8394 12775 8397
rect 15653 8394 15719 8397
rect 12709 8392 15719 8394
rect 12709 8336 12714 8392
rect 12770 8336 15658 8392
rect 15714 8336 15719 8392
rect 12709 8334 15719 8336
rect 12709 8331 12775 8334
rect 15653 8331 15719 8334
rect 21633 8394 21699 8397
rect 21909 8394 21975 8397
rect 21633 8392 21975 8394
rect 21633 8336 21638 8392
rect 21694 8336 21914 8392
rect 21970 8336 21975 8392
rect 21633 8334 21975 8336
rect 21633 8331 21699 8334
rect 21909 8331 21975 8334
rect 11646 8196 11652 8260
rect 11716 8258 11722 8260
rect 11973 8258 12039 8261
rect 27520 8258 28000 8288
rect 11716 8256 12039 8258
rect 11716 8200 11978 8256
rect 12034 8200 12039 8256
rect 11716 8198 12039 8200
rect 11716 8196 11722 8198
rect 11973 8195 12039 8198
rect 20164 8198 28000 8258
rect 10277 8192 10597 8193
rect 0 8122 480 8152
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 10133 8122 10199 8125
rect 0 8120 10199 8122
rect 0 8064 10138 8120
rect 10194 8064 10199 8120
rect 0 8062 10199 8064
rect 0 8032 480 8062
rect 10133 8059 10199 8062
rect 14774 8060 14780 8124
rect 14844 8122 14850 8124
rect 16614 8122 16620 8124
rect 14844 8062 16620 8122
rect 14844 8060 14850 8062
rect 16614 8060 16620 8062
rect 16684 8060 16690 8124
rect 1393 7986 1459 7989
rect 14825 7986 14891 7989
rect 1393 7984 14891 7986
rect 1393 7928 1398 7984
rect 1454 7928 14830 7984
rect 14886 7928 14891 7984
rect 1393 7926 14891 7928
rect 1393 7923 1459 7926
rect 14825 7923 14891 7926
rect 15837 7986 15903 7989
rect 20164 7986 20224 8198
rect 27520 8168 28000 8198
rect 20437 7986 20503 7989
rect 21173 7986 21239 7989
rect 15837 7984 20224 7986
rect 15837 7928 15842 7984
rect 15898 7928 20224 7984
rect 15837 7926 20224 7928
rect 20302 7984 21239 7986
rect 20302 7928 20442 7984
rect 20498 7928 21178 7984
rect 21234 7928 21239 7984
rect 20302 7926 21239 7928
rect 15837 7923 15903 7926
rect 3601 7850 3667 7853
rect 18597 7850 18663 7853
rect 3601 7848 18663 7850
rect 3601 7792 3606 7848
rect 3662 7792 18602 7848
rect 18658 7792 18663 7848
rect 3601 7790 18663 7792
rect 3601 7787 3667 7790
rect 18597 7787 18663 7790
rect 19333 7850 19399 7853
rect 20302 7850 20362 7926
rect 20437 7923 20503 7926
rect 21173 7923 21239 7926
rect 22001 7986 22067 7989
rect 23473 7986 23539 7989
rect 22001 7984 23539 7986
rect 22001 7928 22006 7984
rect 22062 7928 23478 7984
rect 23534 7928 23539 7984
rect 22001 7926 23539 7928
rect 22001 7923 22067 7926
rect 23473 7923 23539 7926
rect 25446 7924 25452 7988
rect 25516 7986 25522 7988
rect 25681 7986 25747 7989
rect 25516 7984 25747 7986
rect 25516 7928 25686 7984
rect 25742 7928 25747 7984
rect 25516 7926 25747 7928
rect 25516 7924 25522 7926
rect 25681 7923 25747 7926
rect 19333 7848 20362 7850
rect 19333 7792 19338 7848
rect 19394 7792 20362 7848
rect 19333 7790 20362 7792
rect 22093 7850 22159 7853
rect 25129 7850 25195 7853
rect 22093 7848 25195 7850
rect 22093 7792 22098 7848
rect 22154 7792 25134 7848
rect 25190 7792 25195 7848
rect 22093 7790 25195 7792
rect 19333 7787 19399 7790
rect 22093 7787 22159 7790
rect 25129 7787 25195 7790
rect 11881 7714 11947 7717
rect 13813 7714 13879 7717
rect 27520 7714 28000 7744
rect 11881 7712 13879 7714
rect 11881 7656 11886 7712
rect 11942 7656 13818 7712
rect 13874 7656 13879 7712
rect 11881 7654 13879 7656
rect 11881 7651 11947 7654
rect 13813 7651 13879 7654
rect 24902 7654 28000 7714
rect 5610 7648 5930 7649
rect 0 7578 480 7608
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 13077 7578 13143 7581
rect 0 7518 5458 7578
rect 0 7488 480 7518
rect 2037 7442 2103 7445
rect 3141 7442 3207 7445
rect 4981 7442 5047 7445
rect 2037 7440 5047 7442
rect 2037 7384 2042 7440
rect 2098 7384 3146 7440
rect 3202 7384 4986 7440
rect 5042 7384 5047 7440
rect 2037 7382 5047 7384
rect 5398 7442 5458 7518
rect 6134 7576 13143 7578
rect 6134 7520 13082 7576
rect 13138 7520 13143 7576
rect 6134 7518 13143 7520
rect 6134 7442 6194 7518
rect 13077 7515 13143 7518
rect 13813 7578 13879 7581
rect 21541 7578 21607 7581
rect 13813 7576 14842 7578
rect 13813 7520 13818 7576
rect 13874 7520 14842 7576
rect 13813 7518 14842 7520
rect 13813 7515 13879 7518
rect 5398 7382 6194 7442
rect 9949 7442 10015 7445
rect 14089 7442 14155 7445
rect 9949 7440 14155 7442
rect 9949 7384 9954 7440
rect 10010 7384 14094 7440
rect 14150 7384 14155 7440
rect 9949 7382 14155 7384
rect 14782 7442 14842 7518
rect 18646 7576 21607 7578
rect 18646 7520 21546 7576
rect 21602 7520 21607 7576
rect 18646 7518 21607 7520
rect 18646 7442 18706 7518
rect 21541 7515 21607 7518
rect 14782 7382 18706 7442
rect 18781 7442 18847 7445
rect 21541 7442 21607 7445
rect 24209 7442 24275 7445
rect 18781 7440 24275 7442
rect 18781 7384 18786 7440
rect 18842 7384 21546 7440
rect 21602 7384 24214 7440
rect 24270 7384 24275 7440
rect 18781 7382 24275 7384
rect 2037 7379 2103 7382
rect 3141 7379 3207 7382
rect 4981 7379 5047 7382
rect 9949 7379 10015 7382
rect 14089 7379 14155 7382
rect 18781 7379 18847 7382
rect 21541 7379 21607 7382
rect 24209 7379 24275 7382
rect 1577 7306 1643 7309
rect 6269 7306 6335 7309
rect 1577 7304 6335 7306
rect 1577 7248 1582 7304
rect 1638 7248 6274 7304
rect 6330 7248 6335 7304
rect 1577 7246 6335 7248
rect 1577 7243 1643 7246
rect 6269 7243 6335 7246
rect 6453 7306 6519 7309
rect 10685 7306 10751 7309
rect 13813 7306 13879 7309
rect 24902 7306 24962 7654
rect 27520 7624 28000 7654
rect 6453 7304 13879 7306
rect 6453 7248 6458 7304
rect 6514 7248 10690 7304
rect 10746 7248 13818 7304
rect 13874 7248 13879 7304
rect 6453 7246 13879 7248
rect 6453 7243 6519 7246
rect 10685 7243 10751 7246
rect 13813 7243 13879 7246
rect 14000 7246 24962 7306
rect 4797 7170 4863 7173
rect 5206 7170 5212 7172
rect 4797 7168 5212 7170
rect 4797 7112 4802 7168
rect 4858 7112 5212 7168
rect 4797 7110 5212 7112
rect 4797 7107 4863 7110
rect 5206 7108 5212 7110
rect 5276 7108 5282 7172
rect 12617 7170 12683 7173
rect 14000 7170 14060 7246
rect 14365 7172 14431 7173
rect 14365 7170 14412 7172
rect 12617 7168 14060 7170
rect 12617 7112 12622 7168
rect 12678 7112 14060 7168
rect 12617 7110 14060 7112
rect 14320 7168 14412 7170
rect 14320 7112 14370 7168
rect 14320 7110 14412 7112
rect 12617 7107 12683 7110
rect 14365 7108 14412 7110
rect 14476 7108 14482 7172
rect 14549 7170 14615 7173
rect 19333 7170 19399 7173
rect 27520 7170 28000 7200
rect 14549 7168 19399 7170
rect 14549 7112 14554 7168
rect 14610 7112 19338 7168
rect 19394 7112 19399 7168
rect 14549 7110 19399 7112
rect 14365 7107 14431 7108
rect 14549 7107 14615 7110
rect 19333 7107 19399 7110
rect 24902 7110 28000 7170
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2865 7034 2931 7037
rect 0 7032 2931 7034
rect 0 6976 2870 7032
rect 2926 6976 2931 7032
rect 0 6974 2931 6976
rect 0 6944 480 6974
rect 2865 6971 2931 6974
rect 4705 7034 4771 7037
rect 4838 7034 4844 7036
rect 4705 7032 4844 7034
rect 4705 6976 4710 7032
rect 4766 6976 4844 7032
rect 4705 6974 4844 6976
rect 4705 6971 4771 6974
rect 4838 6972 4844 6974
rect 4908 6972 4914 7036
rect 5441 7034 5507 7037
rect 9949 7034 10015 7037
rect 17033 7036 17099 7037
rect 5441 7032 10015 7034
rect 5441 6976 5446 7032
rect 5502 6976 9954 7032
rect 10010 6976 10015 7032
rect 5441 6974 10015 6976
rect 5441 6971 5507 6974
rect 9949 6971 10015 6974
rect 16982 6972 16988 7036
rect 17052 7034 17099 7036
rect 24902 7034 24962 7110
rect 27520 7080 28000 7110
rect 17052 7032 19442 7034
rect 17094 6976 19442 7032
rect 17052 6974 19442 6976
rect 17052 6972 17099 6974
rect 17033 6971 17099 6972
rect 1393 6898 1459 6901
rect 8937 6898 9003 6901
rect 1393 6896 9003 6898
rect 1393 6840 1398 6896
rect 1454 6840 8942 6896
rect 8998 6840 9003 6896
rect 1393 6838 9003 6840
rect 1393 6835 1459 6838
rect 8937 6835 9003 6838
rect 11513 6898 11579 6901
rect 14825 6898 14891 6901
rect 16757 6898 16823 6901
rect 11513 6896 16823 6898
rect 11513 6840 11518 6896
rect 11574 6840 14830 6896
rect 14886 6840 16762 6896
rect 16818 6840 16823 6896
rect 11513 6838 16823 6840
rect 19382 6898 19442 6974
rect 20118 6974 24962 7034
rect 20118 6898 20178 6974
rect 21265 6900 21331 6901
rect 19382 6838 20178 6898
rect 11513 6835 11579 6838
rect 14825 6835 14891 6838
rect 16757 6835 16823 6838
rect 21214 6836 21220 6900
rect 21284 6898 21331 6900
rect 21449 6898 21515 6901
rect 23381 6898 23447 6901
rect 21284 6896 21376 6898
rect 21326 6840 21376 6896
rect 21284 6838 21376 6840
rect 21449 6896 23447 6898
rect 21449 6840 21454 6896
rect 21510 6840 23386 6896
rect 23442 6840 23447 6896
rect 21449 6838 23447 6840
rect 21284 6836 21331 6838
rect 21265 6835 21331 6836
rect 21449 6835 21515 6838
rect 23381 6835 23447 6838
rect 5349 6762 5415 6765
rect 14457 6762 14523 6765
rect 5349 6760 18844 6762
rect 5349 6704 5354 6760
rect 5410 6704 14462 6760
rect 14518 6704 18844 6760
rect 5349 6702 18844 6704
rect 5349 6699 5415 6702
rect 14457 6699 14523 6702
rect 7833 6626 7899 6629
rect 7966 6626 7972 6628
rect 7833 6624 7972 6626
rect 7833 6568 7838 6624
rect 7894 6568 7972 6624
rect 7833 6566 7972 6568
rect 7833 6563 7899 6566
rect 7966 6564 7972 6566
rect 8036 6564 8042 6628
rect 16113 6626 16179 6629
rect 18597 6626 18663 6629
rect 16113 6624 18663 6626
rect 16113 6568 16118 6624
rect 16174 6568 18602 6624
rect 18658 6568 18663 6624
rect 16113 6566 18663 6568
rect 18784 6626 18844 6702
rect 21357 6626 21423 6629
rect 18784 6624 21423 6626
rect 18784 6568 21362 6624
rect 21418 6568 21423 6624
rect 18784 6566 21423 6568
rect 16113 6563 16179 6566
rect 18597 6563 18663 6566
rect 21357 6563 21423 6566
rect 26141 6626 26207 6629
rect 27520 6626 28000 6656
rect 26141 6624 28000 6626
rect 26141 6568 26146 6624
rect 26202 6568 28000 6624
rect 26141 6566 28000 6568
rect 26141 6563 26207 6566
rect 5610 6560 5930 6561
rect 0 6490 480 6520
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 5257 6490 5323 6493
rect 0 6488 5323 6490
rect 0 6432 5262 6488
rect 5318 6432 5323 6488
rect 0 6430 5323 6432
rect 0 6400 480 6430
rect 5257 6427 5323 6430
rect 16481 6490 16547 6493
rect 22461 6490 22527 6493
rect 16481 6488 22527 6490
rect 16481 6432 16486 6488
rect 16542 6432 22466 6488
rect 22522 6432 22527 6488
rect 16481 6430 22527 6432
rect 16481 6427 16547 6430
rect 22461 6427 22527 6430
rect 25078 6428 25084 6492
rect 25148 6490 25154 6492
rect 25405 6490 25471 6493
rect 25148 6488 25471 6490
rect 25148 6432 25410 6488
rect 25466 6432 25471 6488
rect 25148 6430 25471 6432
rect 25148 6428 25154 6430
rect 25405 6427 25471 6430
rect 3049 6354 3115 6357
rect 7005 6354 7071 6357
rect 3049 6352 7071 6354
rect 3049 6296 3054 6352
rect 3110 6296 7010 6352
rect 7066 6296 7071 6352
rect 3049 6294 7071 6296
rect 3049 6291 3115 6294
rect 7005 6291 7071 6294
rect 7925 6354 7991 6357
rect 12157 6354 12223 6357
rect 7925 6352 12223 6354
rect 7925 6296 7930 6352
rect 7986 6296 12162 6352
rect 12218 6296 12223 6352
rect 7925 6294 12223 6296
rect 7925 6291 7991 6294
rect 12157 6291 12223 6294
rect 13445 6354 13511 6357
rect 16573 6354 16639 6357
rect 13445 6352 16639 6354
rect 13445 6296 13450 6352
rect 13506 6296 16578 6352
rect 16634 6296 16639 6352
rect 13445 6294 16639 6296
rect 13445 6291 13511 6294
rect 16573 6291 16639 6294
rect 20345 6354 20411 6357
rect 22737 6354 22803 6357
rect 20345 6352 22803 6354
rect 20345 6296 20350 6352
rect 20406 6296 22742 6352
rect 22798 6296 22803 6352
rect 20345 6294 22803 6296
rect 20345 6291 20411 6294
rect 22737 6291 22803 6294
rect 8569 6218 8635 6221
rect 25497 6218 25563 6221
rect 8569 6216 25563 6218
rect 8569 6160 8574 6216
rect 8630 6160 25502 6216
rect 25558 6160 25563 6216
rect 8569 6158 25563 6160
rect 8569 6155 8635 6158
rect 25497 6155 25563 6158
rect 13302 6020 13308 6084
rect 13372 6082 13378 6084
rect 13445 6082 13511 6085
rect 13372 6080 13511 6082
rect 13372 6024 13450 6080
rect 13506 6024 13511 6080
rect 13372 6022 13511 6024
rect 13372 6020 13378 6022
rect 13445 6019 13511 6022
rect 23974 6020 23980 6084
rect 24044 6082 24050 6084
rect 27520 6082 28000 6112
rect 24044 6022 28000 6082
rect 24044 6020 24050 6022
rect 10277 6016 10597 6017
rect 0 5946 480 5976
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 3509 5946 3575 5949
rect 0 5944 3575 5946
rect 0 5888 3514 5944
rect 3570 5888 3575 5944
rect 0 5886 3575 5888
rect 0 5856 480 5886
rect 3509 5883 3575 5886
rect 10777 5946 10843 5949
rect 12433 5946 12499 5949
rect 10777 5944 12499 5946
rect 10777 5888 10782 5944
rect 10838 5888 12438 5944
rect 12494 5888 12499 5944
rect 10777 5886 12499 5888
rect 10777 5883 10843 5886
rect 12433 5883 12499 5886
rect 20989 5946 21055 5949
rect 25037 5946 25103 5949
rect 20989 5944 25103 5946
rect 20989 5888 20994 5944
rect 21050 5888 25042 5944
rect 25098 5888 25103 5944
rect 20989 5886 25103 5888
rect 20989 5883 21055 5886
rect 25037 5883 25103 5886
rect 1761 5810 1827 5813
rect 3049 5810 3115 5813
rect 1761 5808 3115 5810
rect 1761 5752 1766 5808
rect 1822 5752 3054 5808
rect 3110 5752 3115 5808
rect 1761 5750 3115 5752
rect 1761 5747 1827 5750
rect 3049 5747 3115 5750
rect 5441 5810 5507 5813
rect 11881 5810 11947 5813
rect 5441 5808 11947 5810
rect 5441 5752 5446 5808
rect 5502 5752 11886 5808
rect 11942 5752 11947 5808
rect 5441 5750 11947 5752
rect 5441 5747 5507 5750
rect 11881 5747 11947 5750
rect 12157 5810 12223 5813
rect 13629 5810 13695 5813
rect 23289 5810 23355 5813
rect 12157 5808 23355 5810
rect 12157 5752 12162 5808
rect 12218 5752 13634 5808
rect 13690 5752 23294 5808
rect 23350 5752 23355 5808
rect 12157 5750 23355 5752
rect 12157 5747 12223 5750
rect 13629 5747 13695 5750
rect 23289 5747 23355 5750
rect 3509 5674 3575 5677
rect 6913 5674 6979 5677
rect 3509 5672 6979 5674
rect 3509 5616 3514 5672
rect 3570 5616 6918 5672
rect 6974 5616 6979 5672
rect 3509 5614 6979 5616
rect 3509 5611 3575 5614
rect 6913 5611 6979 5614
rect 8937 5674 9003 5677
rect 15377 5674 15443 5677
rect 8937 5672 15443 5674
rect 8937 5616 8942 5672
rect 8998 5616 15382 5672
rect 15438 5616 15443 5672
rect 8937 5614 15443 5616
rect 8937 5611 9003 5614
rect 15377 5611 15443 5614
rect 18321 5674 18387 5677
rect 18597 5674 18663 5677
rect 20989 5674 21055 5677
rect 18321 5672 21055 5674
rect 18321 5616 18326 5672
rect 18382 5616 18602 5672
rect 18658 5616 20994 5672
rect 21050 5616 21055 5672
rect 18321 5614 21055 5616
rect 18321 5611 18387 5614
rect 18597 5611 18663 5614
rect 20989 5611 21055 5614
rect 22829 5674 22895 5677
rect 23841 5674 23907 5677
rect 24485 5674 24551 5677
rect 22829 5672 23907 5674
rect 22829 5616 22834 5672
rect 22890 5616 23846 5672
rect 23902 5616 23907 5672
rect 22829 5614 23907 5616
rect 22829 5611 22895 5614
rect 23841 5611 23907 5614
rect 23982 5672 24551 5674
rect 23982 5616 24490 5672
rect 24546 5616 24551 5672
rect 23982 5614 24551 5616
rect 2773 5538 2839 5541
rect 5349 5538 5415 5541
rect 2773 5536 5415 5538
rect 2773 5480 2778 5536
rect 2834 5480 5354 5536
rect 5410 5480 5415 5536
rect 2773 5478 5415 5480
rect 2773 5475 2839 5478
rect 5349 5475 5415 5478
rect 7097 5538 7163 5541
rect 9765 5538 9831 5541
rect 7097 5536 9831 5538
rect 7097 5480 7102 5536
rect 7158 5480 9770 5536
rect 9826 5480 9831 5536
rect 7097 5478 9831 5480
rect 7097 5475 7163 5478
rect 9765 5475 9831 5478
rect 16665 5538 16731 5541
rect 22737 5538 22803 5541
rect 16665 5536 22803 5538
rect 16665 5480 16670 5536
rect 16726 5480 22742 5536
rect 22798 5480 22803 5536
rect 16665 5478 22803 5480
rect 16665 5475 16731 5478
rect 22737 5475 22803 5478
rect 23289 5538 23355 5541
rect 23982 5538 24042 5614
rect 24485 5611 24551 5614
rect 23289 5536 24042 5538
rect 23289 5480 23294 5536
rect 23350 5480 24042 5536
rect 23289 5478 24042 5480
rect 23289 5475 23355 5478
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 4797 5402 4863 5405
rect 0 5400 4863 5402
rect 0 5344 4802 5400
rect 4858 5344 4863 5400
rect 0 5342 4863 5344
rect 0 5312 480 5342
rect 4797 5339 4863 5342
rect 5993 5402 6059 5405
rect 11881 5402 11947 5405
rect 5993 5400 11947 5402
rect 5993 5344 5998 5400
rect 6054 5344 11886 5400
rect 11942 5344 11947 5400
rect 5993 5342 11947 5344
rect 5993 5339 6059 5342
rect 11881 5339 11947 5342
rect 17401 5402 17467 5405
rect 27520 5402 28000 5432
rect 17401 5400 24042 5402
rect 17401 5344 17406 5400
rect 17462 5344 24042 5400
rect 17401 5342 24042 5344
rect 17401 5339 17467 5342
rect 2957 5266 3023 5269
rect 6269 5266 6335 5269
rect 9029 5266 9095 5269
rect 2957 5264 6335 5266
rect 2957 5208 2962 5264
rect 3018 5208 6274 5264
rect 6330 5208 6335 5264
rect 2957 5206 6335 5208
rect 2957 5203 3023 5206
rect 6269 5203 6335 5206
rect 6502 5264 9095 5266
rect 6502 5208 9034 5264
rect 9090 5208 9095 5264
rect 6502 5206 9095 5208
rect 4245 5132 4311 5133
rect 4245 5130 4292 5132
rect 4200 5128 4292 5130
rect 4200 5072 4250 5128
rect 4200 5070 4292 5072
rect 4245 5068 4292 5070
rect 4356 5068 4362 5132
rect 5349 5130 5415 5133
rect 6502 5130 6562 5206
rect 9029 5203 9095 5206
rect 9397 5266 9463 5269
rect 16849 5266 16915 5269
rect 17953 5266 18019 5269
rect 9397 5264 16915 5266
rect 9397 5208 9402 5264
rect 9458 5208 16854 5264
rect 16910 5208 16915 5264
rect 9397 5206 16915 5208
rect 9397 5203 9463 5206
rect 16849 5203 16915 5206
rect 16990 5264 18019 5266
rect 16990 5208 17958 5264
rect 18014 5208 18019 5264
rect 16990 5206 18019 5208
rect 5349 5128 6562 5130
rect 5349 5072 5354 5128
rect 5410 5072 6562 5128
rect 5349 5070 6562 5072
rect 8845 5130 8911 5133
rect 11697 5130 11763 5133
rect 8845 5128 11763 5130
rect 8845 5072 8850 5128
rect 8906 5072 11702 5128
rect 11758 5072 11763 5128
rect 8845 5070 11763 5072
rect 4245 5067 4311 5068
rect 5349 5067 5415 5070
rect 8845 5067 8911 5070
rect 11697 5067 11763 5070
rect 11881 5130 11947 5133
rect 12617 5130 12683 5133
rect 11881 5128 12683 5130
rect 11881 5072 11886 5128
rect 11942 5072 12622 5128
rect 12678 5072 12683 5128
rect 11881 5070 12683 5072
rect 11881 5067 11947 5070
rect 12617 5067 12683 5070
rect 13077 5130 13143 5133
rect 16990 5130 17050 5206
rect 17953 5203 18019 5206
rect 13077 5128 17050 5130
rect 13077 5072 13082 5128
rect 13138 5072 17050 5128
rect 13077 5070 17050 5072
rect 13077 5067 13143 5070
rect 17166 5068 17172 5132
rect 17236 5130 17242 5132
rect 22185 5130 22251 5133
rect 17236 5128 22251 5130
rect 17236 5072 22190 5128
rect 22246 5072 22251 5128
rect 17236 5070 22251 5072
rect 17236 5068 17242 5070
rect 22185 5067 22251 5070
rect 12249 4994 12315 4997
rect 15510 4994 15516 4996
rect 12249 4992 15516 4994
rect 12249 4936 12254 4992
rect 12310 4936 15516 4992
rect 12249 4934 15516 4936
rect 12249 4931 12315 4934
rect 15510 4932 15516 4934
rect 15580 4932 15586 4996
rect 16481 4994 16547 4997
rect 19333 4994 19399 4997
rect 16481 4992 19399 4994
rect 16481 4936 16486 4992
rect 16542 4936 19338 4992
rect 19394 4936 19399 4992
rect 16481 4934 19399 4936
rect 16481 4931 16547 4934
rect 19333 4931 19399 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 1761 4858 1827 4861
rect 8569 4858 8635 4861
rect 1761 4856 8635 4858
rect 1761 4800 1766 4856
rect 1822 4800 8574 4856
rect 8630 4800 8635 4856
rect 1761 4798 8635 4800
rect 1761 4795 1827 4798
rect 8569 4795 8635 4798
rect 21725 4858 21791 4861
rect 23289 4858 23355 4861
rect 21725 4856 23355 4858
rect 21725 4800 21730 4856
rect 21786 4800 23294 4856
rect 23350 4800 23355 4856
rect 21725 4798 23355 4800
rect 23982 4858 24042 5342
rect 24718 5342 28000 5402
rect 24209 5266 24275 5269
rect 24718 5266 24778 5342
rect 27520 5312 28000 5342
rect 24209 5264 24778 5266
rect 24209 5208 24214 5264
rect 24270 5208 24778 5264
rect 24209 5206 24778 5208
rect 24209 5203 24275 5206
rect 27520 4858 28000 4888
rect 23982 4798 28000 4858
rect 21725 4795 21791 4798
rect 23289 4795 23355 4798
rect 27520 4768 28000 4798
rect 0 4722 480 4752
rect 3693 4722 3759 4725
rect 0 4720 3759 4722
rect 0 4664 3698 4720
rect 3754 4664 3759 4720
rect 0 4662 3759 4664
rect 0 4632 480 4662
rect 3693 4659 3759 4662
rect 5073 4722 5139 4725
rect 7741 4722 7807 4725
rect 5073 4720 7807 4722
rect 5073 4664 5078 4720
rect 5134 4664 7746 4720
rect 7802 4664 7807 4720
rect 5073 4662 7807 4664
rect 5073 4659 5139 4662
rect 7741 4659 7807 4662
rect 13537 4722 13603 4725
rect 15326 4722 15332 4724
rect 13537 4720 15332 4722
rect 13537 4664 13542 4720
rect 13598 4664 15332 4720
rect 13537 4662 15332 4664
rect 13537 4659 13603 4662
rect 15326 4660 15332 4662
rect 15396 4660 15402 4724
rect 15469 4722 15535 4725
rect 25221 4722 25287 4725
rect 15469 4720 25287 4722
rect 15469 4664 15474 4720
rect 15530 4664 25226 4720
rect 25282 4664 25287 4720
rect 15469 4662 25287 4664
rect 15469 4659 15535 4662
rect 25221 4659 25287 4662
rect 4797 4586 4863 4589
rect 18045 4586 18111 4589
rect 4797 4584 18111 4586
rect 4797 4528 4802 4584
rect 4858 4528 18050 4584
rect 18106 4528 18111 4584
rect 4797 4526 18111 4528
rect 4797 4523 4863 4526
rect 18045 4523 18111 4526
rect 23841 4586 23907 4589
rect 23841 4584 24778 4586
rect 23841 4528 23846 4584
rect 23902 4528 24778 4584
rect 23841 4526 24778 4528
rect 23841 4523 23907 4526
rect 9029 4450 9095 4453
rect 14641 4450 14707 4453
rect 9029 4448 14707 4450
rect 9029 4392 9034 4448
rect 9090 4392 14646 4448
rect 14702 4392 14707 4448
rect 9029 4390 14707 4392
rect 9029 4387 9095 4390
rect 14641 4387 14707 4390
rect 15326 4388 15332 4452
rect 15396 4450 15402 4452
rect 19885 4450 19951 4453
rect 15396 4448 19951 4450
rect 15396 4392 19890 4448
rect 19946 4392 19951 4448
rect 15396 4390 19951 4392
rect 15396 4388 15402 4390
rect 19885 4387 19951 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 9029 4314 9095 4317
rect 14733 4314 14799 4317
rect 9029 4312 14799 4314
rect 9029 4256 9034 4312
rect 9090 4256 14738 4312
rect 14794 4256 14799 4312
rect 9029 4254 14799 4256
rect 9029 4251 9095 4254
rect 14733 4251 14799 4254
rect 17585 4314 17651 4317
rect 23197 4314 23263 4317
rect 17585 4312 23263 4314
rect 17585 4256 17590 4312
rect 17646 4256 23202 4312
rect 23258 4256 23263 4312
rect 17585 4254 23263 4256
rect 24718 4314 24778 4526
rect 27520 4314 28000 4344
rect 24718 4254 28000 4314
rect 17585 4251 17651 4254
rect 23197 4251 23263 4254
rect 27520 4224 28000 4254
rect 0 4178 480 4208
rect 1577 4178 1643 4181
rect 0 4176 1643 4178
rect 0 4120 1582 4176
rect 1638 4120 1643 4176
rect 0 4118 1643 4120
rect 0 4088 480 4118
rect 1577 4115 1643 4118
rect 5257 4178 5323 4181
rect 8385 4178 8451 4181
rect 10317 4178 10383 4181
rect 5257 4176 8451 4178
rect 5257 4120 5262 4176
rect 5318 4120 8390 4176
rect 8446 4120 8451 4176
rect 5257 4118 8451 4120
rect 5257 4115 5323 4118
rect 8385 4115 8451 4118
rect 8710 4176 10383 4178
rect 8710 4120 10322 4176
rect 10378 4120 10383 4176
rect 8710 4118 10383 4120
rect 3877 4042 3943 4045
rect 4797 4042 4863 4045
rect 3877 4040 4863 4042
rect 3877 3984 3882 4040
rect 3938 3984 4802 4040
rect 4858 3984 4863 4040
rect 3877 3982 4863 3984
rect 3877 3979 3943 3982
rect 4797 3979 4863 3982
rect 5165 4042 5231 4045
rect 8710 4042 8770 4118
rect 10317 4115 10383 4118
rect 10501 4178 10567 4181
rect 12709 4178 12775 4181
rect 10501 4176 12775 4178
rect 10501 4120 10506 4176
rect 10562 4120 12714 4176
rect 12770 4120 12775 4176
rect 10501 4118 12775 4120
rect 10501 4115 10567 4118
rect 12709 4115 12775 4118
rect 14273 4178 14339 4181
rect 17585 4178 17651 4181
rect 14273 4176 17651 4178
rect 14273 4120 14278 4176
rect 14334 4120 17590 4176
rect 17646 4120 17651 4176
rect 14273 4118 17651 4120
rect 14273 4115 14339 4118
rect 17585 4115 17651 4118
rect 24853 4178 24919 4181
rect 25446 4178 25452 4180
rect 24853 4176 25452 4178
rect 24853 4120 24858 4176
rect 24914 4120 25452 4176
rect 24853 4118 25452 4120
rect 24853 4115 24919 4118
rect 25446 4116 25452 4118
rect 25516 4116 25522 4180
rect 14549 4042 14615 4045
rect 5165 4040 8770 4042
rect 5165 3984 5170 4040
rect 5226 3984 8770 4040
rect 5165 3982 8770 3984
rect 8894 4040 14615 4042
rect 8894 3984 14554 4040
rect 14610 3984 14615 4040
rect 8894 3982 14615 3984
rect 5165 3979 5231 3982
rect 4061 3906 4127 3909
rect 8753 3906 8819 3909
rect 8894 3906 8954 3982
rect 14549 3979 14615 3982
rect 15469 4042 15535 4045
rect 18413 4042 18479 4045
rect 15469 4040 18479 4042
rect 15469 3984 15474 4040
rect 15530 3984 18418 4040
rect 18474 3984 18479 4040
rect 15469 3982 18479 3984
rect 15469 3979 15535 3982
rect 18413 3979 18479 3982
rect 18965 4042 19031 4045
rect 20345 4042 20411 4045
rect 18965 4040 20411 4042
rect 18965 3984 18970 4040
rect 19026 3984 20350 4040
rect 20406 3984 20411 4040
rect 18965 3982 20411 3984
rect 18965 3979 19031 3982
rect 20345 3979 20411 3982
rect 23841 4042 23907 4045
rect 24710 4042 24716 4044
rect 23841 4040 24716 4042
rect 23841 3984 23846 4040
rect 23902 3984 24716 4040
rect 23841 3982 24716 3984
rect 23841 3979 23907 3982
rect 24710 3980 24716 3982
rect 24780 3980 24786 4044
rect 4061 3904 8954 3906
rect 4061 3848 4066 3904
rect 4122 3848 8758 3904
rect 8814 3848 8954 3904
rect 4061 3846 8954 3848
rect 14181 3906 14247 3909
rect 19333 3906 19399 3909
rect 14181 3904 19399 3906
rect 14181 3848 14186 3904
rect 14242 3848 19338 3904
rect 19394 3848 19399 3904
rect 14181 3846 19399 3848
rect 4061 3843 4127 3846
rect 8753 3843 8819 3846
rect 14181 3843 14247 3846
rect 19333 3843 19399 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 2957 3770 3023 3773
rect 3969 3770 4035 3773
rect 2957 3768 4035 3770
rect 2957 3712 2962 3768
rect 3018 3712 3974 3768
rect 4030 3712 4035 3768
rect 2957 3710 4035 3712
rect 2957 3707 3023 3710
rect 3969 3707 4035 3710
rect 8201 3770 8267 3773
rect 9949 3770 10015 3773
rect 8201 3768 10015 3770
rect 8201 3712 8206 3768
rect 8262 3712 9954 3768
rect 10010 3712 10015 3768
rect 8201 3710 10015 3712
rect 8201 3707 8267 3710
rect 9949 3707 10015 3710
rect 13261 3770 13327 3773
rect 15009 3770 15075 3773
rect 13261 3768 15075 3770
rect 13261 3712 13266 3768
rect 13322 3712 15014 3768
rect 15070 3712 15075 3768
rect 13261 3710 15075 3712
rect 13261 3707 13327 3710
rect 15009 3707 15075 3710
rect 20161 3770 20227 3773
rect 22093 3770 22159 3773
rect 20161 3768 22159 3770
rect 20161 3712 20166 3768
rect 20222 3712 22098 3768
rect 22154 3712 22159 3768
rect 20161 3710 22159 3712
rect 20161 3707 20227 3710
rect 22093 3707 22159 3710
rect 23289 3770 23355 3773
rect 25681 3770 25747 3773
rect 27520 3770 28000 3800
rect 23289 3768 28000 3770
rect 23289 3712 23294 3768
rect 23350 3712 25686 3768
rect 25742 3712 28000 3768
rect 23289 3710 28000 3712
rect 23289 3707 23355 3710
rect 25681 3707 25747 3710
rect 27520 3680 28000 3710
rect 0 3634 480 3664
rect 2037 3634 2103 3637
rect 0 3632 2103 3634
rect 0 3576 2042 3632
rect 2098 3576 2103 3632
rect 0 3574 2103 3576
rect 0 3544 480 3574
rect 2037 3571 2103 3574
rect 2497 3634 2563 3637
rect 10133 3634 10199 3637
rect 16849 3634 16915 3637
rect 2497 3632 10199 3634
rect 2497 3576 2502 3632
rect 2558 3576 10138 3632
rect 10194 3576 10199 3632
rect 2497 3574 10199 3576
rect 2497 3571 2563 3574
rect 10133 3571 10199 3574
rect 10366 3632 16915 3634
rect 10366 3576 16854 3632
rect 16910 3576 16915 3632
rect 10366 3574 16915 3576
rect 1577 3498 1643 3501
rect 8845 3498 8911 3501
rect 10366 3498 10426 3574
rect 16849 3571 16915 3574
rect 17309 3634 17375 3637
rect 21541 3634 21607 3637
rect 17309 3632 21607 3634
rect 17309 3576 17314 3632
rect 17370 3576 21546 3632
rect 21602 3576 21607 3632
rect 17309 3574 21607 3576
rect 17309 3571 17375 3574
rect 21541 3571 21607 3574
rect 1577 3496 3250 3498
rect 1577 3440 1582 3496
rect 1638 3440 3250 3496
rect 1577 3438 3250 3440
rect 1577 3435 1643 3438
rect 841 3362 907 3365
rect 974 3362 980 3364
rect 841 3360 980 3362
rect 841 3304 846 3360
rect 902 3304 980 3360
rect 841 3302 980 3304
rect 841 3299 907 3302
rect 974 3300 980 3302
rect 1044 3300 1050 3364
rect 3190 3362 3250 3438
rect 8845 3496 10426 3498
rect 8845 3440 8850 3496
rect 8906 3440 10426 3496
rect 8845 3438 10426 3440
rect 10501 3498 10567 3501
rect 13629 3498 13695 3501
rect 10501 3496 13695 3498
rect 10501 3440 10506 3496
rect 10562 3440 13634 3496
rect 13690 3440 13695 3496
rect 10501 3438 13695 3440
rect 8845 3435 8911 3438
rect 10501 3435 10567 3438
rect 13629 3435 13695 3438
rect 13905 3498 13971 3501
rect 19517 3498 19583 3501
rect 21173 3498 21239 3501
rect 13905 3496 19583 3498
rect 13905 3440 13910 3496
rect 13966 3440 19522 3496
rect 19578 3440 19583 3496
rect 13905 3438 19583 3440
rect 13905 3435 13971 3438
rect 19517 3435 19583 3438
rect 19750 3496 21239 3498
rect 19750 3440 21178 3496
rect 21234 3440 21239 3496
rect 19750 3438 21239 3440
rect 5165 3362 5231 3365
rect 3190 3360 5231 3362
rect 3190 3304 5170 3360
rect 5226 3304 5231 3360
rect 3190 3302 5231 3304
rect 5165 3299 5231 3302
rect 7281 3362 7347 3365
rect 14549 3362 14615 3365
rect 7281 3360 14615 3362
rect 7281 3304 7286 3360
rect 7342 3304 14554 3360
rect 14610 3304 14615 3360
rect 7281 3302 14615 3304
rect 7281 3299 7347 3302
rect 14549 3299 14615 3302
rect 15653 3362 15719 3365
rect 19750 3362 19810 3438
rect 21173 3435 21239 3438
rect 15653 3360 19810 3362
rect 15653 3304 15658 3360
rect 15714 3304 19810 3360
rect 15653 3302 19810 3304
rect 20161 3362 20227 3365
rect 23657 3362 23723 3365
rect 20161 3360 23723 3362
rect 20161 3304 20166 3360
rect 20222 3304 23662 3360
rect 23718 3304 23723 3360
rect 20161 3302 23723 3304
rect 15653 3299 15719 3302
rect 20161 3299 20227 3302
rect 23657 3299 23723 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 8109 3226 8175 3229
rect 11973 3226 12039 3229
rect 20253 3226 20319 3229
rect 8109 3224 12039 3226
rect 8109 3168 8114 3224
rect 8170 3168 11978 3224
rect 12034 3168 12039 3224
rect 8109 3166 12039 3168
rect 8109 3163 8175 3166
rect 11973 3163 12039 3166
rect 15334 3224 20319 3226
rect 15334 3168 20258 3224
rect 20314 3168 20319 3224
rect 15334 3166 20319 3168
rect 0 3090 480 3120
rect 2129 3090 2195 3093
rect 0 3088 2195 3090
rect 0 3032 2134 3088
rect 2190 3032 2195 3088
rect 0 3030 2195 3032
rect 0 3000 480 3030
rect 2129 3027 2195 3030
rect 3601 3090 3667 3093
rect 3734 3090 3740 3092
rect 3601 3088 3740 3090
rect 3601 3032 3606 3088
rect 3662 3032 3740 3088
rect 3601 3030 3740 3032
rect 3601 3027 3667 3030
rect 3734 3028 3740 3030
rect 3804 3028 3810 3092
rect 5349 3090 5415 3093
rect 10501 3090 10567 3093
rect 5349 3088 10567 3090
rect 5349 3032 5354 3088
rect 5410 3032 10506 3088
rect 10562 3032 10567 3088
rect 5349 3030 10567 3032
rect 5349 3027 5415 3030
rect 10501 3027 10567 3030
rect 14549 3090 14615 3093
rect 15334 3090 15394 3166
rect 20253 3163 20319 3166
rect 26049 3226 26115 3229
rect 27520 3226 28000 3256
rect 26049 3224 28000 3226
rect 26049 3168 26054 3224
rect 26110 3168 28000 3224
rect 26049 3166 28000 3168
rect 26049 3163 26115 3166
rect 27520 3136 28000 3166
rect 14549 3088 15394 3090
rect 14549 3032 14554 3088
rect 14610 3032 15394 3088
rect 14549 3030 15394 3032
rect 18689 3090 18755 3093
rect 21633 3090 21699 3093
rect 18689 3088 21834 3090
rect 18689 3032 18694 3088
rect 18750 3032 21638 3088
rect 21694 3032 21834 3088
rect 18689 3030 21834 3032
rect 14549 3027 14615 3030
rect 18689 3027 18755 3030
rect 21633 3027 21699 3030
rect 6545 2954 6611 2957
rect 13997 2954 14063 2957
rect 6545 2952 14063 2954
rect 6545 2896 6550 2952
rect 6606 2896 14002 2952
rect 14058 2896 14063 2952
rect 6545 2894 14063 2896
rect 6545 2891 6611 2894
rect 13997 2891 14063 2894
rect 15510 2892 15516 2956
rect 15580 2954 15586 2956
rect 18689 2954 18755 2957
rect 15580 2952 18755 2954
rect 15580 2896 18694 2952
rect 18750 2896 18755 2952
rect 15580 2894 18755 2896
rect 21774 2954 21834 3030
rect 23565 2954 23631 2957
rect 21774 2952 23631 2954
rect 21774 2896 23570 2952
rect 23626 2896 23631 2952
rect 21774 2894 23631 2896
rect 15580 2892 15586 2894
rect 18689 2891 18755 2894
rect 23565 2891 23631 2894
rect 2865 2818 2931 2821
rect 6453 2818 6519 2821
rect 8661 2818 8727 2821
rect 2865 2816 8727 2818
rect 2865 2760 2870 2816
rect 2926 2760 6458 2816
rect 6514 2760 8666 2816
rect 8722 2760 8727 2816
rect 2865 2758 8727 2760
rect 2865 2755 2931 2758
rect 6453 2755 6519 2758
rect 8661 2755 8727 2758
rect 11145 2818 11211 2821
rect 15193 2818 15259 2821
rect 11145 2816 15259 2818
rect 11145 2760 11150 2816
rect 11206 2760 15198 2816
rect 15254 2760 15259 2816
rect 11145 2758 15259 2760
rect 11145 2755 11211 2758
rect 15193 2755 15259 2758
rect 20621 2818 20687 2821
rect 22461 2818 22527 2821
rect 25313 2818 25379 2821
rect 20621 2816 22527 2818
rect 20621 2760 20626 2816
rect 20682 2760 22466 2816
rect 22522 2760 22527 2816
rect 20621 2758 22527 2760
rect 20621 2755 20687 2758
rect 22461 2755 22527 2758
rect 23430 2816 25379 2818
rect 23430 2760 25318 2816
rect 25374 2760 25379 2816
rect 23430 2758 25379 2760
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 7005 2682 7071 2685
rect 9857 2682 9923 2685
rect 7005 2680 9923 2682
rect 7005 2624 7010 2680
rect 7066 2624 9862 2680
rect 9918 2624 9923 2680
rect 7005 2622 9923 2624
rect 7005 2619 7071 2622
rect 9857 2619 9923 2622
rect 12893 2682 12959 2685
rect 17033 2682 17099 2685
rect 12893 2680 17099 2682
rect 12893 2624 12898 2680
rect 12954 2624 17038 2680
rect 17094 2624 17099 2680
rect 12893 2622 17099 2624
rect 12893 2619 12959 2622
rect 17033 2619 17099 2622
rect 21265 2682 21331 2685
rect 23430 2682 23490 2758
rect 25313 2755 25379 2758
rect 21265 2680 23490 2682
rect 21265 2624 21270 2680
rect 21326 2624 23490 2680
rect 21265 2622 23490 2624
rect 21265 2619 21331 2622
rect 0 2546 480 2576
rect 1209 2546 1275 2549
rect 0 2544 1275 2546
rect 0 2488 1214 2544
rect 1270 2488 1275 2544
rect 0 2486 1275 2488
rect 0 2456 480 2486
rect 1209 2483 1275 2486
rect 1393 2546 1459 2549
rect 14641 2546 14707 2549
rect 1393 2544 14707 2546
rect 1393 2488 1398 2544
rect 1454 2488 14646 2544
rect 14702 2488 14707 2544
rect 1393 2486 14707 2488
rect 1393 2483 1459 2486
rect 14641 2483 14707 2486
rect 15837 2546 15903 2549
rect 25589 2546 25655 2549
rect 15837 2544 25655 2546
rect 15837 2488 15842 2544
rect 15898 2488 25594 2544
rect 25650 2488 25655 2544
rect 15837 2486 25655 2488
rect 15837 2483 15903 2486
rect 25589 2483 25655 2486
rect 25865 2546 25931 2549
rect 27520 2546 28000 2576
rect 25865 2544 28000 2546
rect 25865 2488 25870 2544
rect 25926 2488 28000 2544
rect 25865 2486 28000 2488
rect 25865 2483 25931 2486
rect 27520 2456 28000 2486
rect 5901 2410 5967 2413
rect 6678 2410 6684 2412
rect 5901 2408 6684 2410
rect 5901 2352 5906 2408
rect 5962 2352 6684 2408
rect 5901 2350 6684 2352
rect 5901 2347 5967 2350
rect 6678 2348 6684 2350
rect 6748 2348 6754 2412
rect 6821 2410 6887 2413
rect 9305 2410 9371 2413
rect 14089 2410 14155 2413
rect 15193 2410 15259 2413
rect 6821 2408 14155 2410
rect 6821 2352 6826 2408
rect 6882 2352 9310 2408
rect 9366 2352 14094 2408
rect 14150 2352 14155 2408
rect 6821 2350 14155 2352
rect 6821 2347 6887 2350
rect 9305 2347 9371 2350
rect 14089 2347 14155 2350
rect 14230 2408 15259 2410
rect 14230 2352 15198 2408
rect 15254 2352 15259 2408
rect 14230 2350 15259 2352
rect 13445 2274 13511 2277
rect 14230 2274 14290 2350
rect 15193 2347 15259 2350
rect 7606 2272 14290 2274
rect 7606 2216 13450 2272
rect 13506 2216 14290 2272
rect 7606 2214 14290 2216
rect 15377 2274 15443 2277
rect 19425 2274 19491 2277
rect 15377 2272 19491 2274
rect 15377 2216 15382 2272
rect 15438 2216 19430 2272
rect 19486 2216 19491 2272
rect 15377 2214 19491 2216
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 0 2002 480 2032
rect 1945 2002 2011 2005
rect 0 2000 2011 2002
rect 0 1944 1950 2000
rect 2006 1944 2011 2000
rect 0 1942 2011 1944
rect 0 1912 480 1942
rect 1945 1939 2011 1942
rect 1945 1866 2011 1869
rect 7606 1866 7666 2214
rect 13445 2211 13511 2214
rect 15377 2211 15443 2214
rect 19425 2211 19491 2214
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 9397 2138 9463 2141
rect 13997 2138 14063 2141
rect 19977 2138 20043 2141
rect 9397 2136 14063 2138
rect 9397 2080 9402 2136
rect 9458 2080 14002 2136
rect 14058 2080 14063 2136
rect 9397 2078 14063 2080
rect 9397 2075 9463 2078
rect 13997 2075 14063 2078
rect 15334 2136 20043 2138
rect 15334 2080 19982 2136
rect 20038 2080 20043 2136
rect 15334 2078 20043 2080
rect 7741 2002 7807 2005
rect 12525 2002 12591 2005
rect 13721 2002 13787 2005
rect 7741 2000 13787 2002
rect 7741 1944 7746 2000
rect 7802 1944 12530 2000
rect 12586 1944 13726 2000
rect 13782 1944 13787 2000
rect 7741 1942 13787 1944
rect 7741 1939 7807 1942
rect 12525 1939 12591 1942
rect 13721 1939 13787 1942
rect 14089 2002 14155 2005
rect 15334 2002 15394 2078
rect 19977 2075 20043 2078
rect 14089 2000 15394 2002
rect 14089 1944 14094 2000
rect 14150 1944 15394 2000
rect 14089 1942 15394 1944
rect 18597 2002 18663 2005
rect 27061 2002 27127 2005
rect 18597 2000 27127 2002
rect 18597 1944 18602 2000
rect 18658 1944 27066 2000
rect 27122 1944 27127 2000
rect 18597 1942 27127 1944
rect 14089 1939 14155 1942
rect 18597 1939 18663 1942
rect 27061 1939 27127 1942
rect 27245 2002 27311 2005
rect 27520 2002 28000 2032
rect 27245 2000 28000 2002
rect 27245 1944 27250 2000
rect 27306 1944 28000 2000
rect 27245 1942 28000 1944
rect 27245 1939 27311 1942
rect 27520 1912 28000 1942
rect 1945 1864 7666 1866
rect 1945 1808 1950 1864
rect 2006 1808 7666 1864
rect 1945 1806 7666 1808
rect 1945 1803 2011 1806
rect 14590 1804 14596 1868
rect 14660 1866 14666 1868
rect 19241 1866 19307 1869
rect 14660 1864 19307 1866
rect 14660 1808 19246 1864
rect 19302 1808 19307 1864
rect 14660 1806 19307 1808
rect 14660 1804 14666 1806
rect 19241 1803 19307 1806
rect 2773 1730 2839 1733
rect 8845 1730 8911 1733
rect 2773 1728 8911 1730
rect 2773 1672 2778 1728
rect 2834 1672 8850 1728
rect 8906 1672 8911 1728
rect 2773 1670 8911 1672
rect 2773 1667 2839 1670
rect 8845 1667 8911 1670
rect 9581 1730 9647 1733
rect 15469 1730 15535 1733
rect 9581 1728 15535 1730
rect 9581 1672 9586 1728
rect 9642 1672 15474 1728
rect 15530 1672 15535 1728
rect 9581 1670 15535 1672
rect 9581 1667 9647 1670
rect 15469 1667 15535 1670
rect 23013 1730 23079 1733
rect 27613 1730 27679 1733
rect 23013 1728 27679 1730
rect 23013 1672 23018 1728
rect 23074 1672 27618 1728
rect 27674 1672 27679 1728
rect 23013 1670 27679 1672
rect 23013 1667 23079 1670
rect 27613 1667 27679 1670
rect 565 1594 631 1597
rect 11605 1594 11671 1597
rect 17033 1594 17099 1597
rect 565 1592 7298 1594
rect 565 1536 570 1592
rect 626 1536 7298 1592
rect 565 1534 7298 1536
rect 565 1531 631 1534
rect 0 1458 480 1488
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 7238 1458 7298 1534
rect 11605 1592 17099 1594
rect 11605 1536 11610 1592
rect 11666 1536 17038 1592
rect 17094 1536 17099 1592
rect 11605 1534 17099 1536
rect 11605 1531 11671 1534
rect 17033 1531 17099 1534
rect 11789 1458 11855 1461
rect 7238 1456 11855 1458
rect 7238 1400 11794 1456
rect 11850 1400 11855 1456
rect 7238 1398 11855 1400
rect 0 1368 480 1398
rect 3509 1395 3575 1398
rect 11789 1395 11855 1398
rect 11973 1458 12039 1461
rect 17769 1458 17835 1461
rect 11973 1456 17835 1458
rect 11973 1400 11978 1456
rect 12034 1400 17774 1456
rect 17830 1400 17835 1456
rect 11973 1398 17835 1400
rect 11973 1395 12039 1398
rect 17769 1395 17835 1398
rect 25221 1458 25287 1461
rect 27520 1458 28000 1488
rect 25221 1456 28000 1458
rect 25221 1400 25226 1456
rect 25282 1400 28000 1456
rect 25221 1398 28000 1400
rect 25221 1395 25287 1398
rect 27520 1368 28000 1398
rect 7281 1322 7347 1325
rect 16757 1322 16823 1325
rect 7281 1320 16823 1322
rect 7281 1264 7286 1320
rect 7342 1264 16762 1320
rect 16818 1264 16823 1320
rect 7281 1262 16823 1264
rect 7281 1259 7347 1262
rect 16757 1259 16823 1262
rect 7925 1186 7991 1189
rect 10869 1186 10935 1189
rect 7925 1184 10935 1186
rect 7925 1128 7930 1184
rect 7986 1128 10874 1184
rect 10930 1128 10935 1184
rect 7925 1126 10935 1128
rect 7925 1123 7991 1126
rect 10869 1123 10935 1126
rect 11053 1186 11119 1189
rect 17953 1186 18019 1189
rect 11053 1184 18019 1186
rect 11053 1128 11058 1184
rect 11114 1128 17958 1184
rect 18014 1128 18019 1184
rect 11053 1126 18019 1128
rect 11053 1123 11119 1126
rect 17953 1123 18019 1126
rect 3049 1050 3115 1053
rect 13169 1050 13235 1053
rect 3049 1048 13235 1050
rect 3049 992 3054 1048
rect 3110 992 13174 1048
rect 13230 992 13235 1048
rect 3049 990 13235 992
rect 3049 987 3115 990
rect 13169 987 13235 990
rect 0 914 480 944
rect 1301 914 1367 917
rect 0 912 1367 914
rect 0 856 1306 912
rect 1362 856 1367 912
rect 0 854 1367 856
rect 0 824 480 854
rect 1301 851 1367 854
rect 8845 914 8911 917
rect 11053 914 11119 917
rect 8845 912 11119 914
rect 8845 856 8850 912
rect 8906 856 11058 912
rect 11114 856 11119 912
rect 8845 854 11119 856
rect 8845 851 8911 854
rect 11053 851 11119 854
rect 26233 914 26299 917
rect 27520 914 28000 944
rect 26233 912 28000 914
rect 26233 856 26238 912
rect 26294 856 28000 912
rect 26233 854 28000 856
rect 26233 851 26299 854
rect 27520 824 28000 854
rect 8753 778 8819 781
rect 18137 778 18203 781
rect 8753 776 18203 778
rect 8753 720 8758 776
rect 8814 720 18142 776
rect 18198 720 18203 776
rect 8753 718 18203 720
rect 8753 715 8819 718
rect 18137 715 18203 718
rect 8017 642 8083 645
rect 18045 642 18111 645
rect 8017 640 18111 642
rect 8017 584 8022 640
rect 8078 584 18050 640
rect 18106 584 18111 640
rect 8017 582 18111 584
rect 8017 579 8083 582
rect 18045 579 18111 582
rect 0 370 480 400
rect 6177 370 6243 373
rect 0 368 6243 370
rect 0 312 6182 368
rect 6238 312 6243 368
rect 0 310 6243 312
rect 0 280 480 310
rect 6177 307 6243 310
rect 10961 370 11027 373
rect 23473 370 23539 373
rect 10961 368 23539 370
rect 10961 312 10966 368
rect 11022 312 23478 368
rect 23534 312 23539 368
rect 10961 310 23539 312
rect 10961 307 11027 310
rect 23473 307 23539 310
rect 26049 370 26115 373
rect 27520 370 28000 400
rect 26049 368 28000 370
rect 26049 312 26054 368
rect 26110 312 28000 368
rect 26049 310 28000 312
rect 26049 307 26115 310
rect 27520 280 28000 310
rect 7005 234 7071 237
rect 8201 234 8267 237
rect 23657 234 23723 237
rect 7005 232 23723 234
rect 7005 176 7010 232
rect 7066 176 8206 232
rect 8262 176 23662 232
rect 23718 176 23723 232
rect 7005 174 23723 176
rect 7005 171 7071 174
rect 8201 171 8267 174
rect 23657 171 23723 174
rect 4429 98 4495 101
rect 22553 98 22619 101
rect 4429 96 22619 98
rect 4429 40 4434 96
rect 4490 40 22558 96
rect 22614 40 22619 96
rect 4429 38 22619 40
rect 4429 35 4495 38
rect 22553 35 22619 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 2820 19076 2884 19140
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 3372 18940 3436 19004
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 24716 17988 24780 18052
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 17908 17172 17972 17236
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 3372 15540 3436 15604
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 5396 14860 5460 14924
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 4660 14588 4724 14652
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 17908 14588 17972 14652
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 19380 14044 19444 14108
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 17908 13092 17972 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 11100 12956 11164 13020
rect 23612 12820 23676 12884
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 4660 12336 4724 12340
rect 4660 12280 4674 12336
rect 4674 12280 4724 12336
rect 4660 12276 4724 12280
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 2820 11732 2884 11796
rect 19380 12276 19444 12340
rect 23428 12276 23492 12340
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 9996 11384 10060 11388
rect 9996 11328 10010 11384
rect 10010 11328 10060 11384
rect 9996 11324 10060 11328
rect 14780 11052 14844 11116
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 23980 9964 24044 10028
rect 18828 9888 18892 9892
rect 18828 9832 18878 9888
rect 18878 9832 18892 9888
rect 18828 9828 18892 9832
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 23980 9420 24044 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 21220 9148 21284 9212
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 4844 8604 4908 8668
rect 12756 8936 12820 8940
rect 12756 8880 12770 8936
rect 12770 8880 12820 8936
rect 12756 8876 12820 8880
rect 23612 9012 23676 9076
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 15884 8468 15948 8532
rect 6868 8332 6932 8396
rect 11652 8196 11716 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 14780 8060 14844 8124
rect 16620 8060 16684 8124
rect 25452 7924 25516 7988
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 5212 7108 5276 7172
rect 14412 7168 14476 7172
rect 14412 7112 14426 7168
rect 14426 7112 14476 7168
rect 14412 7108 14476 7112
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 4844 6972 4908 7036
rect 16988 7032 17052 7036
rect 16988 6976 17038 7032
rect 17038 6976 17052 7032
rect 16988 6972 17052 6976
rect 21220 6896 21284 6900
rect 21220 6840 21270 6896
rect 21270 6840 21284 6896
rect 21220 6836 21284 6840
rect 7972 6564 8036 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 25084 6428 25148 6492
rect 13308 6020 13372 6084
rect 23980 6020 24044 6084
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 4292 5128 4356 5132
rect 4292 5072 4306 5128
rect 4306 5072 4356 5128
rect 4292 5068 4356 5072
rect 17172 5068 17236 5132
rect 15516 4932 15580 4996
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 15332 4660 15396 4724
rect 15332 4388 15396 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 25452 4116 25516 4180
rect 24716 3980 24780 4044
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 980 3300 1044 3364
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 3740 3028 3804 3092
rect 15516 2892 15580 2956
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 6684 2348 6748 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 14596 1804 14660 1868
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 2819 19140 2885 19141
rect 2819 19076 2820 19140
rect 2884 19076 2885 19140
rect 2819 19075 2885 19076
rect 2822 11797 2882 19075
rect 3371 19004 3437 19005
rect 3371 18940 3372 19004
rect 3436 18940 3437 19004
rect 3371 18939 3437 18940
rect 3374 15605 3434 18939
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 3371 15604 3437 15605
rect 3371 15540 3372 15604
rect 3436 15540 3437 15604
rect 3371 15539 3437 15540
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5395 14924 5461 14925
rect 5395 14860 5396 14924
rect 5460 14860 5461 14924
rect 5395 14859 5461 14860
rect 4659 14652 4725 14653
rect 4659 14588 4660 14652
rect 4724 14588 4725 14652
rect 4659 14587 4725 14588
rect 4662 12341 4722 14587
rect 5398 14058 5458 14859
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 4659 12340 4725 12341
rect 4659 12276 4660 12340
rect 4724 12276 4725 12340
rect 4659 12275 4725 12276
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 2819 11796 2885 11797
rect 2819 11732 2820 11796
rect 2884 11732 2885 11796
rect 2819 11731 2885 11732
rect 5610 10912 5931 11936
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 17907 17236 17973 17237
rect 17907 17172 17908 17236
rect 17972 17172 17973 17236
rect 17907 17171 17973 17172
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 17910 14653 17970 17171
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 17907 14652 17973 14653
rect 17907 14588 17908 14652
rect 17972 14588 17973 14652
rect 17907 14587 17973 14588
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 17910 13157 17970 14587
rect 19379 14108 19445 14109
rect 19379 14058 19380 14108
rect 19444 14058 19445 14108
rect 17907 13156 17973 13157
rect 17907 13092 17908 13156
rect 17972 13092 17973 13156
rect 17907 13091 17973 13092
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 11099 13020 11165 13021
rect 11099 12956 11100 13020
rect 11164 12956 11165 13020
rect 11099 12955 11165 12956
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 9995 11388 10061 11389
rect 9995 11324 9996 11388
rect 10060 11324 10061 11388
rect 9995 11323 10061 11324
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 4843 8668 4909 8669
rect 4843 8618 4844 8668
rect 4908 8618 4909 8668
rect 4846 7037 4906 7702
rect 5610 7648 5931 8672
rect 6870 8397 6930 9742
rect 9998 9298 10058 11323
rect 10277 10368 10597 11392
rect 11102 10658 11162 12955
rect 14944 12000 15264 13024
rect 19382 12341 19442 13822
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24715 18052 24781 18053
rect 24715 17988 24716 18052
rect 24780 17988 24781 18052
rect 24715 17987 24781 17988
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 23611 12884 23677 12885
rect 23611 12820 23612 12884
rect 23676 12820 23677 12884
rect 23611 12819 23677 12820
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19379 12340 19445 12341
rect 19379 12276 19380 12340
rect 19444 12276 19445 12340
rect 19379 12275 19445 12276
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14779 11116 14845 11117
rect 14779 11052 14780 11116
rect 14844 11052 14845 11116
rect 14779 11051 14845 11052
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 4843 7036 4909 7037
rect 4843 6972 4844 7036
rect 4908 6972 4909 7036
rect 4843 6971 4909 6972
rect 5610 6560 5931 7584
rect 10277 8192 10597 9216
rect 12755 8940 12821 8941
rect 12755 8876 12756 8940
rect 12820 8876 12821 8940
rect 12755 8875 12821 8876
rect 11651 8260 11717 8261
rect 11651 8196 11652 8260
rect 11716 8196 11717 8260
rect 11651 8195 11717 8196
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 7971 6628 8037 6629
rect 7971 6564 7972 6628
rect 8036 6564 8037 6628
rect 7971 6563 8037 6564
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 7974 5898 8034 6563
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 982 3365 1042 4302
rect 979 3364 1045 3365
rect 979 3300 980 3364
rect 1044 3300 1045 3364
rect 979 3299 1045 3300
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 11654 4538 11714 8195
rect 12758 5898 12818 8875
rect 14782 8125 14842 11051
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 19610 11456 19930 12480
rect 23427 12340 23493 12341
rect 23427 12276 23428 12340
rect 23492 12276 23493 12340
rect 23427 12275 23493 12276
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14779 8124 14845 8125
rect 14779 8060 14780 8124
rect 14844 8060 14845 8124
rect 14779 8059 14845 8060
rect 14944 7648 15264 8672
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 21219 9212 21285 9213
rect 21219 9148 21220 9212
rect 21284 9148 21285 9212
rect 21219 9147 21285 9148
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 16619 8124 16685 8125
rect 16619 8060 16620 8124
rect 16684 8060 16685 8124
rect 16619 8059 16685 8060
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 16622 6578 16682 8059
rect 16990 7037 17050 7702
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 16987 7036 17053 7037
rect 16987 6972 16988 7036
rect 17052 6972 17053 7036
rect 16987 6971 17053 6972
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 13307 6084 13373 6085
rect 13307 6020 13308 6084
rect 13372 6020 13373 6084
rect 13307 6019 13373 6020
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 13310 3178 13370 6019
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 19610 6016 19930 7040
rect 21222 6901 21282 9147
rect 23430 7258 23490 12275
rect 23614 9077 23674 12819
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 23982 10029 24042 10422
rect 23979 10028 24045 10029
rect 23979 9964 23980 10028
rect 24044 9964 24045 10028
rect 23979 9963 24045 9964
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 23979 9484 24045 9485
rect 23979 9420 23980 9484
rect 24044 9420 24045 9484
rect 23979 9419 24045 9420
rect 23982 9298 24042 9419
rect 23611 9076 23677 9077
rect 23611 9012 23612 9076
rect 23676 9012 23677 9076
rect 23611 9011 23677 9012
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 21219 6900 21285 6901
rect 21219 6836 21220 6900
rect 21284 6836 21285 6900
rect 21219 6835 21285 6836
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 23979 6084 24045 6085
rect 23979 6020 23980 6084
rect 24044 6020 24045 6084
rect 23979 6019 24045 6020
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 15515 4996 15581 4997
rect 15515 4932 15516 4996
rect 15580 4932 15581 4996
rect 15515 4931 15581 4932
rect 15331 4724 15397 4725
rect 15331 4660 15332 4724
rect 15396 4660 15397 4724
rect 15331 4659 15397 4660
rect 15334 4453 15394 4659
rect 15331 4452 15397 4453
rect 15331 4388 15332 4452
rect 15396 4388 15397 4452
rect 15331 4387 15397 4388
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2128 10597 2688
rect 14598 1869 14658 2262
rect 14944 2208 15264 3232
rect 15518 2957 15578 4931
rect 19610 4928 19930 5952
rect 23982 5898 24042 6019
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 15515 2956 15581 2957
rect 15515 2892 15516 2956
rect 15580 2892 15581 2956
rect 15515 2891 15581 2892
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24718 4045 24778 17987
rect 25451 7988 25517 7989
rect 25451 7924 25452 7988
rect 25516 7924 25517 7988
rect 25451 7923 25517 7924
rect 25454 4181 25514 7923
rect 25451 4180 25517 4181
rect 25451 4116 25452 4180
rect 25516 4116 25517 4180
rect 25451 4115 25517 4116
rect 24715 4044 24781 4045
rect 24715 3980 24716 4044
rect 24780 3980 24781 4044
rect 24715 3979 24781 3980
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 14595 1868 14661 1869
rect 14595 1804 14596 1868
rect 14660 1804 14661 1868
rect 14595 1803 14661 1804
<< via4 >>
rect 5310 13822 5546 14058
rect 19294 14044 19380 14058
rect 19380 14044 19444 14058
rect 19444 14044 19530 14058
rect 19294 13822 19530 14044
rect 6782 9742 7018 9978
rect 4758 8604 4844 8618
rect 4844 8604 4908 8618
rect 4908 8604 4994 8618
rect 4758 8382 4994 8604
rect 4758 7702 4994 7938
rect 11014 10422 11250 10658
rect 9910 9062 10146 9298
rect 5126 7172 5362 7258
rect 5126 7108 5212 7172
rect 5212 7108 5276 7172
rect 5276 7108 5362 7172
rect 5126 7022 5362 7108
rect 7886 5662 8122 5898
rect 4206 5132 4442 5218
rect 4206 5068 4292 5132
rect 4292 5068 4356 5132
rect 4356 5068 4442 5132
rect 4206 4982 4442 5068
rect 894 4302 1130 4538
rect 3654 3092 3890 3178
rect 3654 3028 3740 3092
rect 3740 3028 3804 3092
rect 3804 3028 3890 3092
rect 3654 2942 3890 3028
rect 18742 9892 18978 9978
rect 18742 9828 18828 9892
rect 18828 9828 18892 9892
rect 18892 9828 18978 9892
rect 18742 9742 18978 9828
rect 15798 8532 16034 8618
rect 15798 8468 15884 8532
rect 15884 8468 15948 8532
rect 15948 8468 16034 8532
rect 15798 8382 16034 8468
rect 14326 7172 14562 7258
rect 14326 7108 14412 7172
rect 14412 7108 14476 7172
rect 14476 7108 14562 7172
rect 14326 7022 14562 7108
rect 16902 7702 17138 7938
rect 12670 5662 12906 5898
rect 11566 4302 11802 4538
rect 16534 6342 16770 6578
rect 23894 10422 24130 10658
rect 23894 9062 24130 9298
rect 23342 7022 23578 7258
rect 17086 5132 17322 5218
rect 17086 5068 17172 5132
rect 17172 5068 17236 5132
rect 17236 5068 17322 5132
rect 17086 4982 17322 5068
rect 13222 2942 13458 3178
rect 6598 2412 6834 2498
rect 6598 2348 6684 2412
rect 6684 2348 6748 2412
rect 6748 2348 6834 2412
rect 6598 2262 6834 2348
rect 14510 2262 14746 2498
rect 23894 5662 24130 5898
rect 24998 6492 25234 6578
rect 24998 6428 25084 6492
rect 25084 6428 25148 6492
rect 25148 6428 25234 6492
rect 24998 6342 25234 6428
<< metal5 >>
rect 5268 14058 19572 14100
rect 5268 13822 5310 14058
rect 5546 13822 19294 14058
rect 19530 13822 19572 14058
rect 5268 13780 19572 13822
rect 10972 10658 24172 10700
rect 10972 10422 11014 10658
rect 11250 10422 23894 10658
rect 24130 10422 24172 10658
rect 10972 10380 24172 10422
rect 6740 9978 19020 10020
rect 6740 9742 6782 9978
rect 7018 9742 18742 9978
rect 18978 9742 19020 9978
rect 6740 9700 19020 9742
rect 9868 9298 24172 9340
rect 9868 9062 9910 9298
rect 10146 9062 23894 9298
rect 24130 9062 24172 9298
rect 9868 9020 24172 9062
rect 4716 8618 16076 8660
rect 4716 8382 4758 8618
rect 4994 8382 15798 8618
rect 16034 8382 16076 8618
rect 4716 8340 16076 8382
rect 4716 7938 17180 7980
rect 4716 7702 4758 7938
rect 4994 7702 16902 7938
rect 17138 7702 17180 7938
rect 4716 7660 17180 7702
rect 5084 7258 23620 7300
rect 5084 7022 5126 7258
rect 5362 7022 14326 7258
rect 14562 7022 23342 7258
rect 23578 7022 23620 7258
rect 5084 6980 23620 7022
rect 16492 6578 25276 6620
rect 16492 6342 16534 6578
rect 16770 6342 24998 6578
rect 25234 6342 25276 6578
rect 16492 6300 25276 6342
rect 7844 5898 24172 5940
rect 7844 5662 7886 5898
rect 8122 5662 12670 5898
rect 12906 5662 23894 5898
rect 24130 5662 24172 5898
rect 7844 5620 24172 5662
rect 4164 5218 17364 5260
rect 4164 4982 4206 5218
rect 4442 4982 17086 5218
rect 17322 4982 17364 5218
rect 4164 4940 17364 4982
rect 852 4538 11844 4580
rect 852 4302 894 4538
rect 1130 4302 11566 4538
rect 11802 4302 11844 4538
rect 852 4260 11844 4302
rect 3612 3178 13500 3220
rect 3612 2942 3654 3178
rect 3890 2942 13222 3178
rect 13458 2942 13500 3178
rect 3612 2900 13500 2942
rect 6556 2498 14788 2540
rect 6556 2262 6598 2498
rect 6834 2262 14510 2498
rect 14746 2262 14788 2498
rect 6556 2220 14788 2262
use sky130_fd_sc_hd__conb_1  _053_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1604681595
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1604681595
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_22
timestamp 1604681595
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 3864 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1604681595
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80
timestamp 1604681595
transform 1 0 8464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1604681595
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1604681595
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1604681595
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1604681595
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12696 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_145
timestamp 1604681595
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_149
timestamp 1604681595
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148
timestamp 1604681595
transform 1 0 14720 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 15180 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_162
timestamp 1604681595
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1604681595
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_174
timestamp 1604681595
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1604681595
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 1604681595
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1604681595
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 17940 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1604681595
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18216 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604681595
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_192
timestamp 1604681595
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_205
timestamp 1604681595
transform 1 0 19964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_228
timestamp 1604681595
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21252 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1604681595
transform 1 0 22632 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_232
timestamp 1604681595
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_240
timestamp 1604681595
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1604681595
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1604681595
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_254
timestamp 1604681595
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_268
timestamp 1604681595
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_272
timestamp 1604681595
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_276
timestamp 1604681595
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_12
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_16
timestamp 1604681595
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1604681595
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1604681595
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_64
timestamp 1604681595
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1604681595
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8924 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1604681595
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_116
timestamp 1604681595
transform 1 0 11776 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1604681595
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1604681595
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1604681595
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1604681595
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1604681595
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1604681595
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18676 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_200
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1604681595
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21620 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24104 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23920 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23552 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_242
timestamp 1604681595
transform 1 0 23368 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_246
timestamp 1604681595
transform 1 0 23736 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_259
timestamp 1604681595
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604681595
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1604681595
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1604681595
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_50
timestamp 1604681595
transform 1 0 5704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_54
timestamp 1604681595
transform 1 0 6072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1604681595
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1604681595
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1604681595
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_96
timestamp 1604681595
transform 1 0 9936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1604681595
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12696 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1604681595
transform 1 0 14444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15456 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_149
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_152
timestamp 1604681595
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1604681595
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1604681595
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_173
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_207
timestamp 1604681595
transform 1 0 20148 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_212
timestamp 1604681595
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_235
timestamp 1604681595
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_239
timestamp 1604681595
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1604681595
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_268
timestamp 1604681595
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_272
timestamp 1604681595
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_12
timestamp 1604681595
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_16
timestamp 1604681595
transform 1 0 2576 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_20
timestamp 1604681595
transform 1 0 2944 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 4232 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_38
timestamp 1604681595
transform 1 0 4600 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5336 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_4_43
timestamp 1604681595
transform 1 0 5060 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_65
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_69
timestamp 1604681595
transform 1 0 7452 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9752 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604681595
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12512 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1604681595
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1604681595
transform 1 0 12236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1604681595
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1604681595
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_162
timestamp 1604681595
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16192 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_183
timestamp 1604681595
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_187
timestamp 1604681595
transform 1 0 18308 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18860 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_228
timestamp 1604681595
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23460 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_241
timestamp 1604681595
transform 1 0 23276 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_245
timestamp 1604681595
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_258
timestamp 1604681595
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_262
timestamp 1604681595
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_266
timestamp 1604681595
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1472 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1604681595
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1604681595
transform 1 0 3864 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_34
timestamp 1604681595
transform 1 0 4232 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_37
timestamp 1604681595
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 6072 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_52
timestamp 1604681595
transform 1 0 5888 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_56
timestamp 1604681595
transform 1 0 6256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_65
timestamp 1604681595
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_69
timestamp 1604681595
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1604681595
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 9384 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1604681595
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_111
timestamp 1604681595
transform 1 0 11316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_115
timestamp 1604681595
transform 1 0 11684 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13892 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1604681595
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1604681595
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1604681595
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1604681595
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_173
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_189
timestamp 1604681595
transform 1 0 18492 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_212
timestamp 1604681595
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1604681595
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_229
timestamp 1604681595
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_233
timestamp 1604681595
transform 1 0 22540 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_237
timestamp 1604681595
transform 1 0 22908 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1604681595
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_268
timestamp 1604681595
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_272
timestamp 1604681595
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_10
timestamp 1604681595
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1604681595
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_37
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_33
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4324 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1604681595
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_54
timestamp 1604681595
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8556 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1604681595
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1604681595
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_80
timestamp 1604681595
transform 1 0 8464 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1604681595
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_98
timestamp 1604681595
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_123
timestamp 1604681595
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_115
timestamp 1604681595
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_127
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1604681595
transform 1 0 13984 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_140
timestamp 1604681595
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14076 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1604681595
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1604681595
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1604681595
transform 1 0 16284 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_160
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15364 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_174
timestamp 1604681595
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1604681595
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_187
timestamp 1604681595
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_178
timestamp 1604681595
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_183
timestamp 1604681595
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_191
timestamp 1604681595
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 1604681595
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_212
timestamp 1604681595
transform 1 0 20608 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_228
timestamp 1604681595
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 21528 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_235
timestamp 1604681595
transform 1 0 22724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_231
timestamp 1604681595
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_238
timestamp 1604681595
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22448 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_242
timestamp 1604681595
transform 1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23184 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23920 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_254
timestamp 1604681595
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_258
timestamp 1604681595
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_261
timestamp 1604681595
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_257
timestamp 1604681595
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1604681595
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_269 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25852 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_265
timestamp 1604681595
transform 1 0 25484 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_272
timestamp 1604681595
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1604681595
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_10
timestamp 1604681595
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5796 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_43
timestamp 1604681595
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1604681595
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_60
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_65
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_77
timestamp 1604681595
transform 1 0 8188 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_83
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10580 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8924 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_99
timestamp 1604681595
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_122
timestamp 1604681595
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1604681595
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_139
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_147
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_158
timestamp 1604681595
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1604681595
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19136 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23368 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23184 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_234
timestamp 1604681595
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_238
timestamp 1604681595
transform 1 0 23000 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_261
timestamp 1604681595
transform 1 0 25116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_265
timestamp 1604681595
transform 1 0 25484 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_269
timestamp 1604681595
transform 1 0 25852 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_14
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1604681595
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_22
timestamp 1604681595
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1604681595
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_90
timestamp 1604681595
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_94
timestamp 1604681595
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_107
timestamp 1604681595
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1604681595
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_115
timestamp 1604681595
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1604681595
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1604681595
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1604681595
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1604681595
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19780 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1604681595
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1604681595
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23092 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_241
timestamp 1604681595
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24564 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_251
timestamp 1604681595
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1604681595
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_268
timestamp 1604681595
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_272
timestamp 1604681595
transform 1 0 26128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604681595
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_6
timestamp 1604681595
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1604681595
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_46
timestamp 1604681595
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_54
timestamp 1604681595
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1604681595
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_71
timestamp 1604681595
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_99
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_103
timestamp 1604681595
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1604681595
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_143
timestamp 1604681595
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 18768 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1604681595
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_204
timestamp 1604681595
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_208
timestamp 1604681595
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1604681595
transform 1 0 21528 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_219
timestamp 1604681595
transform 1 0 21252 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 22540 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22908 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_231
timestamp 1604681595
transform 1 0 22356 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_235
timestamp 1604681595
transform 1 0 22724 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_248
timestamp 1604681595
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24656 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 24472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_252
timestamp 1604681595
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_265
timestamp 1604681595
transform 1 0 25484 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_273
timestamp 1604681595
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_31
timestamp 1604681595
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_44
timestamp 1604681595
transform 1 0 5152 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_50
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_54
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6992 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_11_83
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1604681595
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1604681595
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1604681595
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14352 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_153
timestamp 1604681595
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1604681595
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1604681595
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_165
timestamp 1604681595
transform 1 0 16284 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17664 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18952 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1604681595
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21436 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1604681595
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1604681595
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23092 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_230
timestamp 1604681595
transform 1 0 22264 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_234
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_237
timestamp 1604681595
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_241
timestamp 1604681595
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1604681595
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_268
timestamp 1604681595
transform 1 0 25760 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_6
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1604681595
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 4508 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_40
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1604681595
transform 1 0 6348 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1604681595
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1604681595
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_114
timestamp 1604681595
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13340 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_127
timestamp 1604681595
transform 1 0 12788 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1604681595
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_158
timestamp 1604681595
transform 1 0 15640 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17664 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_172
timestamp 1604681595
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_176
timestamp 1604681595
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1604681595
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1604681595
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22632 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_232
timestamp 1604681595
transform 1 0 22448 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_236
timestamp 1604681595
transform 1 0 22816 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_258
timestamp 1604681595
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_262
timestamp 1604681595
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_266
timestamp 1604681595
transform 1 0 25576 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1604681595
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604681595
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1604681595
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_20
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_40
timestamp 1604681595
transform 1 0 4784 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1604681595
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1604681595
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1604681595
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1604681595
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_68
timestamp 1604681595
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_74
timestamp 1604681595
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7728 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1604681595
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_108
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1604681595
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_116
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_120
timestamp 1604681595
transform 1 0 12144 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_126
timestamp 1604681595
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_127
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1604681595
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_139
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13156 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_14_147
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_151
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1604681595
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1604681595
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 16284 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_13_173
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1604681595
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_192
timestamp 1604681595
transform 1 0 18768 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_193
timestamp 1604681595
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_199
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 19596 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604681595
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604681595
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1604681595
transform 1 0 22080 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_224
timestamp 1604681595
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 21896 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_232
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22632 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_248
timestamp 1604681595
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_243
timestamp 1604681595
transform 1 0 23460 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 24104 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 24380 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_252
timestamp 1604681595
transform 1 0 24288 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_262
timestamp 1604681595
transform 1 0 25208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_266
timestamp 1604681595
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_273
timestamp 1604681595
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604681595
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1656 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_25
timestamp 1604681595
transform 1 0 3404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_29
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1604681595
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_81
timestamp 1604681595
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_85
timestamp 1604681595
transform 1 0 8924 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1604681595
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1604681595
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_111
timestamp 1604681595
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1604681595
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1604681595
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1604681595
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_207
timestamp 1604681595
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1604681595
transform 1 0 21252 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_211
timestamp 1604681595
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_228
timestamp 1604681595
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1604681595
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_239
timestamp 1604681595
transform 1 0 23092 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23828 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_249
timestamp 1604681595
transform 1 0 24012 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24196 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_262
timestamp 1604681595
transform 1 0 25208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_270
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_14
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1604681595
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1604681595
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1604681595
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_38
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4692 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1604681595
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_75
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1604681595
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_118
timestamp 1604681595
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13156 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_126
timestamp 1604681595
transform 1 0 12696 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_140
timestamp 1604681595
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_148
timestamp 1604681595
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1604681595
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_158
timestamp 1604681595
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17940 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_175
timestamp 1604681595
transform 1 0 17204 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_179
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 19504 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_192
timestamp 1604681595
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_196
timestamp 1604681595
transform 1 0 19136 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_204
timestamp 1604681595
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1604681595
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_228
timestamp 1604681595
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22908 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22724 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_232
timestamp 1604681595
transform 1 0 22448 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 25392 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_256
timestamp 1604681595
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_260
timestamp 1604681595
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1604681595
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_38
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_50
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_54
timestamp 1604681595
transform 1 0 6072 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_58
timestamp 1604681595
transform 1 0 6440 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_66
timestamp 1604681595
transform 1 0 7176 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1604681595
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1604681595
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16008 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_146
timestamp 1604681595
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_154
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1604681595
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 19320 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1604681595
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1604681595
transform 1 0 18768 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21896 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_221
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 24104 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23276 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_235
timestamp 1604681595
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_239
timestamp 1604681595
transform 1 0 23092 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_243
timestamp 1604681595
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_273
timestamp 1604681595
transform 1 0 26220 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1604681595
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 5980 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_45
timestamp 1604681595
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10304 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_119
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_127
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17940 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 17756 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1604681595
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_179
timestamp 1604681595
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_207
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1604681595
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_224
timestamp 1604681595
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_228
timestamp 1604681595
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 22816 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22632 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_232
timestamp 1604681595
transform 1 0 22448 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_245
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_249
timestamp 1604681595
transform 1 0 24012 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24380 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_252
timestamp 1604681595
transform 1 0 24288 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_262
timestamp 1604681595
transform 1 0 25208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_266
timestamp 1604681595
transform 1 0 25576 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1604681595
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_17
timestamp 1604681595
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_18
timestamp 1604681595
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_14
timestamp 1604681595
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_25
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1604681595
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_40
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1604681595
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_45
timestamp 1604681595
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 5612 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1604681595
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1604681595
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_64
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_68
timestamp 1604681595
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7728 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_74
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1604681595
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_85
timestamp 1604681595
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9292 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp 1604681595
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_107
timestamp 1604681595
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1604681595
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 1604681595
transform 1 0 12052 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_127
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1604681595
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1604681595
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15180 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16836 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1604681595
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_176
timestamp 1604681595
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_201
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_204
timestamp 1604681595
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1604681595
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 19872 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20332 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_228
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_229
timestamp 1604681595
transform 1 0 22172 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_238
timestamp 1604681595
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_242
timestamp 1604681595
transform 1 0 23368 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_249
timestamp 1604681595
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23552 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23184 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23736 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 24380 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_262
timestamp 1604681595
transform 1 0 25208 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_266
timestamp 1604681595
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_270
timestamp 1604681595
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_265
timestamp 1604681595
transform 1 0 25484 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_274
timestamp 1604681595
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_273
timestamp 1604681595
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2024 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_29
timestamp 1604681595
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_34
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 6900 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1604681595
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_127
timestamp 1604681595
transform 1 0 12788 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_151
timestamp 1604681595
transform 1 0 14996 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_160
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1604681595
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1604681595
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1604681595
transform 1 0 20424 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1604681595
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_254
timestamp 1604681595
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_258
timestamp 1604681595
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_268
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_272
timestamp 1604681595
transform 1 0 26128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_21
timestamp 1604681595
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_25
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5888 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1604681595
transform 1 0 5336 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_61
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1604681595
transform 1 0 7084 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12144 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1604681595
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1604681595
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_139
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_163
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17204 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17020 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_168
timestamp 1604681595
transform 1 0 16560 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_172
timestamp 1604681595
transform 1 0 16928 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1604681595
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1604681595
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_192
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_224
timestamp 1604681595
transform 1 0 21712 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_229
timestamp 1604681595
transform 1 0 22172 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 22724 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_233
timestamp 1604681595
transform 1 0 22540 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 25208 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_254
timestamp 1604681595
transform 1 0 24472 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_258
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 1604681595
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604681595
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_24
timestamp 1604681595
transform 1 0 3312 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1604681595
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604681595
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 1604681595
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_70
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1604681595
transform 1 0 9752 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 14260 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_140
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1604681595
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_166
timestamp 1604681595
transform 1 0 16376 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18216 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_205
timestamp 1604681595
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20700 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1604681595
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_219
timestamp 1604681595
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_223
timestamp 1604681595
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_272
timestamp 1604681595
transform 1 0 26128 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1472 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_13
timestamp 1604681595
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1604681595
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_25
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_21
timestamp 1604681595
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_36
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4508 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_46
timestamp 1604681595
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_50
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_54
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 8372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_100
timestamp 1604681595
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1604681595
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13156 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_127
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_140
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_148
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_160
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_164
timestamp 1604681595
transform 1 0 16192 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17020 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp 1604681595
transform 1 0 16744 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1604681595
transform 1 0 18768 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_196
timestamp 1604681595
transform 1 0 19136 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_199
timestamp 1604681595
transform 1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21160 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_237
timestamp 1604681595
transform 1 0 22908 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_241
timestamp 1604681595
transform 1 0 23276 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_264
timestamp 1604681595
transform 1 0 25392 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_272
timestamp 1604681595
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_12
timestamp 1604681595
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1604681595
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_20
timestamp 1604681595
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1604681595
transform 1 0 4876 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_45
timestamp 1604681595
transform 1 0 5244 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_48
timestamp 1604681595
transform 1 0 5520 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 5612 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_66
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_90 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9384 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_102
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 11040 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_111
timestamp 1604681595
transform 1 0 11316 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13156 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_127
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_140
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_144
timestamp 1604681595
transform 1 0 14352 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_160
timestamp 1604681595
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_164
timestamp 1604681595
transform 1 0 16192 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_170
timestamp 1604681595
transform 1 0 16744 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18124 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19688 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_194
timestamp 1604681595
transform 1 0 18952 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_199
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1604681595
transform 1 0 21804 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_229
timestamp 1604681595
transform 1 0 22172 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1604681595
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_270
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1604681595
transform 1 0 1472 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1604681595
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_13
timestamp 1604681595
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_25
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_38
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1604681595
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_50
timestamp 1604681595
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_42
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1604681595
transform 1 0 6532 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_54
timestamp 1604681595
transform 1 0 6072 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6716 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_47
timestamp 1604681595
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1604681595
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_76
timestamp 1604681595
transform 1 0 8096 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_135
timestamp 1604681595
transform 1 0 13524 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 15824 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16008 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_147
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_164
timestamp 1604681595
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 16928 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_181
timestamp 1604681595
transform 1 0 17756 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_187
timestamp 1604681595
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_168
timestamp 1604681595
transform 1 0 16560 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_190
timestamp 1604681595
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1604681595
transform 1 0 18676 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_200
timestamp 1604681595
transform 1 0 19504 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19320 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19872 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1604681595
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1604681595
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1604681595
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21436 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_234
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_230
timestamp 1604681595
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 22448 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_242
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_247
timestamp 1604681595
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_241
timestamp 1604681595
transform 1 0 23276 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_249
timestamp 1604681595
transform 1 0 24012 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_259
timestamp 1604681595
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_259
timestamp 1604681595
transform 1 0 24932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_255
timestamp 1604681595
transform 1 0 24564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_267
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_263
timestamp 1604681595
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_275
timestamp 1604681595
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1604681595
transform 1 0 1472 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_13
timestamp 1604681595
transform 1 0 2300 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_17
timestamp 1604681595
transform 1 0 2668 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_22
timestamp 1604681595
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604681595
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1604681595
transform 1 0 3496 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1604681595
transform 1 0 4784 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_36
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_48
timestamp 1604681595
transform 1 0 5520 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_60
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 17388 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_174
timestamp 1604681595
transform 1 0 17112 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1604681595
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_192
timestamp 1604681595
transform 1 0 18768 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21804 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604681595
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_223
timestamp 1604681595
transform 1 0 21620 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 22356 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 23460 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_235
timestamp 1604681595
transform 1 0 22724 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_247
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_259
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 1604681595
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3680 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_25
timestamp 1604681595
transform 1 0 3404 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_50
timestamp 1604681595
transform 1 0 5704 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1604681595
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_171
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_176
timestamp 1604681595
transform 1 0 17296 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604681595
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_200
timestamp 1604681595
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_204
timestamp 1604681595
transform 1 0 19872 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 21896 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_216
timestamp 1604681595
transform 1 0 20976 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_224
timestamp 1604681595
transform 1 0 21712 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_228
timestamp 1604681595
transform 1 0 22080 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 22264 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_249
timestamp 1604681595
transform 1 0 24012 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 25392 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 24288 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_256
timestamp 1604681595
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_260
timestamp 1604681595
transform 1 0 25024 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_268
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_272
timestamp 1604681595
transform 1 0 26128 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 2760 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_10
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_14
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_17
timestamp 1604681595
transform 1 0 2668 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_22
timestamp 1604681595
transform 1 0 3128 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1604681595
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_48
timestamp 1604681595
transform 1 0 5520 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_60
timestamp 1604681595
transform 1 0 6624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1604681595
transform 1 0 7728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17112 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1604681595
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_192
timestamp 1604681595
transform 1 0 18768 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 22356 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_235
timestamp 1604681595
transform 1 0 22724 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_247
timestamp 1604681595
transform 1 0 23828 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_259
timestamp 1604681595
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1604681595
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604681595
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_23
timestamp 1604681595
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_35
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1604681595
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 18124 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 1604681595
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1604681595
transform 1 0 19964 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_217
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_229
timestamp 1604681595
transform 1 0 22172 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 22540 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_236
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_259
timestamp 1604681595
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_263
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_275
timestamp 1604681595
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_19
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 23552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_243
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_247
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 24564 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_259
timestamp 1604681595
transform 1 0 24932 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_271
timestamp 1604681595
transform 1 0 26036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_19
timestamp 1604681595
transform 1 0 2852 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_7
timestamp 1604681595
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 4416 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_35
timestamp 1604681595
transform 1 0 4324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_38
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_40
timestamp 1604681595
transform 1 0 4784 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_50
timestamp 1604681595
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_54
timestamp 1604681595
transform 1 0 6072 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_52
timestamp 1604681595
transform 1 0 5888 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_64
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_76
timestamp 1604681595
transform 1 0 8096 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_88
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23828 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_249
timestamp 1604681595
transform 1 0 24012 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 24564 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_259
timestamp 1604681595
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_263
timestamp 1604681595
transform 1 0 25300 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_275
timestamp 1604681595
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1604681595
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_11
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1604681595
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_253
timestamp 1604681595
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_259
timestamp 1604681595
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_263
timestamp 1604681595
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_275
timestamp 1604681595
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604681595
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_12
timestamp 1604681595
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_16
timestamp 1604681595
transform 1 0 2576 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_28
timestamp 1604681595
transform 1 0 3680 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_40
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_52
timestamp 1604681595
transform 1 0 5888 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_60
timestamp 1604681595
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_98
timestamp 1604681595
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1604681595
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19504 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_202
timestamp 1604681595
transform 1 0 19688 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_214
timestamp 1604681595
transform 1 0 20792 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_226
timestamp 1604681595
transform 1 0 21896 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_238
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_7
timestamp 1604681595
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_19
timestamp 1604681595
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1604681595
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1604681595
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_190
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_198
timestamp 1604681595
transform 1 0 19320 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_206
timestamp 1604681595
transform 1 0 20056 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604681595
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1604681595
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_47
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_202
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1604681595
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_253
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604681595
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 27616 480 27736 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 24490 27520 24546 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 27066 0 27122 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_42_
port 4 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_43_
port 5 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_44_
port 6 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_45_
port 7 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_46_
port 8 nsew default input
rlabel metal2 s 3054 0 3110 480 6 bottom_left_grid_pin_47_
port 9 nsew default input
rlabel metal2 s 3606 0 3662 480 6 bottom_left_grid_pin_48_
port 10 nsew default input
rlabel metal2 s 4158 0 4214 480 6 bottom_left_grid_pin_49_
port 11 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 ccff_head
port 12 nsew default input
rlabel metal2 s 17498 27520 17554 28000 6 ccff_tail
port 13 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 chanx_left_in[0]
port 14 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[10]
port 15 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[11]
port 16 nsew default input
rlabel metal3 s 0 11432 480 11552 6 chanx_left_in[12]
port 17 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[13]
port 18 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[14]
port 19 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 20 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 21 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 22 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 23 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 24 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[1]
port 25 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[2]
port 26 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[3]
port 27 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[4]
port 28 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[5]
port 29 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[6]
port 30 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[7]
port 31 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[8]
port 32 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[9]
port 33 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[0]
port 34 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[10]
port 35 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[11]
port 36 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 chanx_left_out[12]
port 37 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[13]
port 38 nsew default tristate
rlabel metal3 s 0 23808 480 23928 6 chanx_left_out[14]
port 39 nsew default tristate
rlabel metal3 s 0 24352 480 24472 6 chanx_left_out[15]
port 40 nsew default tristate
rlabel metal3 s 0 24896 480 25016 6 chanx_left_out[16]
port 41 nsew default tristate
rlabel metal3 s 0 25440 480 25560 6 chanx_left_out[17]
port 42 nsew default tristate
rlabel metal3 s 0 25984 480 26104 6 chanx_left_out[18]
port 43 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[19]
port 44 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[1]
port 45 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[2]
port 46 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 chanx_left_out[3]
port 47 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 chanx_left_out[4]
port 48 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[5]
port 49 nsew default tristate
rlabel metal3 s 0 19320 480 19440 6 chanx_left_out[6]
port 50 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 chanx_left_out[7]
port 51 nsew default tristate
rlabel metal3 s 0 20408 480 20528 6 chanx_left_out[8]
port 52 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[9]
port 53 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[0]
port 54 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[10]
port 55 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[11]
port 56 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[12]
port 57 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_in[13]
port 58 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[14]
port 59 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[15]
port 60 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[16]
port 61 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_in[17]
port 62 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_in[18]
port 63 nsew default input
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_in[19]
port 64 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[1]
port 65 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 66 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[3]
port 67 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[4]
port 68 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[5]
port 69 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[6]
port 70 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[7]
port 71 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[8]
port 72 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[9]
port 73 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_out[0]
port 74 nsew default tristate
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_out[10]
port 75 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[11]
port 76 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[12]
port 77 nsew default tristate
rlabel metal3 s 27520 23672 28000 23792 6 chanx_right_out[13]
port 78 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[14]
port 79 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[15]
port 80 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[16]
port 81 nsew default tristate
rlabel metal3 s 27520 25984 28000 26104 6 chanx_right_out[17]
port 82 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[18]
port 83 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[19]
port 84 nsew default tristate
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_out[1]
port 85 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[2]
port 86 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[3]
port 87 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 88 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 89 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_out[6]
port 90 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 91 nsew default tristate
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_out[8]
port 92 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[9]
port 93 nsew default tristate
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[0]
port 94 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[10]
port 95 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[11]
port 96 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[12]
port 97 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[13]
port 98 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[14]
port 99 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[15]
port 100 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[16]
port 101 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[17]
port 102 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_in[18]
port 103 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[19]
port 104 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[1]
port 105 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[2]
port 106 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[3]
port 107 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[4]
port 108 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[5]
port 109 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[6]
port 110 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[7]
port 111 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[8]
port 112 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[9]
port 113 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[0]
port 114 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[10]
port 115 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 116 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[12]
port 117 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[13]
port 118 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[14]
port 119 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[15]
port 120 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[16]
port 121 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[17]
port 122 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[18]
port 123 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[19]
port 124 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[1]
port 125 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[2]
port 126 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[3]
port 127 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[4]
port 128 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[5]
port 129 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[6]
port 130 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[7]
port 131 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[8]
port 132 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_out[9]
port 133 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 134 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 135 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 136 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 137 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_38_
port 138 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_39_
port 139 nsew default input
rlabel metal3 s 0 3544 480 3664 6 left_bottom_grid_pin_40_
port 140 nsew default input
rlabel metal3 s 0 4088 480 4208 6 left_bottom_grid_pin_41_
port 141 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_1_
port 142 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 prog_clk
port 143 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 144 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 145 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 146 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 147 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_bottom_grid_pin_38_
port 148 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 149 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 150 nsew default input
rlabel metal3 s 27520 4224 28000 4344 6 right_bottom_grid_pin_41_
port 151 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_1_
port 152 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 153 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 154 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
