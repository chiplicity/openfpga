magic
tech sky130A
magscale 1 2
timestamp 1606932241
<< locali >>
rect 8401 19295 8435 19465
rect 4905 18751 4939 18921
rect 6745 18819 6779 18921
rect 8217 18275 8251 18377
rect 12817 18071 12851 18173
rect 4077 17595 4111 17765
rect 17325 17663 17359 17833
rect 3617 16983 3651 17289
rect 14197 16983 14231 17153
rect 4905 16643 4939 16745
rect 11253 16643 11287 16745
rect 19349 16439 19383 16541
rect 1961 15895 1995 15997
rect 6929 15351 6963 15453
rect 4905 14263 4939 14365
rect 6193 12291 6227 12393
rect 4997 12087 5031 12257
rect 9413 12155 9447 12325
rect 19349 12155 19383 12325
rect 6653 11679 6687 11849
rect 10333 10999 10367 11169
rect 12633 11067 12667 11305
rect 7849 10047 7883 10149
rect 16865 9367 16899 9673
rect 17877 9367 17911 9537
rect 18981 9367 19015 9673
rect 9505 8823 9539 9061
rect 10609 8823 10643 9129
rect 13369 8959 13403 9129
rect 11161 8415 11195 8517
rect 7389 7803 7423 8041
rect 12817 7735 12851 7905
rect 20637 6171 20671 6341
rect 16037 5763 16071 5865
rect 22293 5559 22327 5729
rect 13369 5151 13403 5321
rect 13093 3383 13127 3621
rect 15945 3451 15979 3689
<< viali >>
rect 1593 21641 1627 21675
rect 9965 21641 9999 21675
rect 15485 21641 15519 21675
rect 17877 21641 17911 21675
rect 13645 21573 13679 21607
rect 21189 21573 21223 21607
rect 2605 21505 2639 21539
rect 3617 21505 3651 21539
rect 4629 21505 4663 21539
rect 6377 21505 6411 21539
rect 7481 21505 7515 21539
rect 8953 21505 8987 21539
rect 13277 21505 13311 21539
rect 14197 21505 14231 21539
rect 16129 21505 16163 21539
rect 17049 21505 17083 21539
rect 21741 21505 21775 21539
rect 1409 21437 1443 21471
rect 5089 21437 5123 21471
rect 7941 21437 7975 21471
rect 9781 21437 9815 21471
rect 10701 21437 10735 21471
rect 13093 21437 13127 21471
rect 14841 21437 14875 21471
rect 15853 21437 15887 21471
rect 17693 21437 17727 21471
rect 18337 21437 18371 21471
rect 18889 21437 18923 21471
rect 20545 21437 20579 21471
rect 22201 21437 22235 21471
rect 2329 21369 2363 21403
rect 6193 21369 6227 21403
rect 7297 21369 7331 21403
rect 8861 21369 8895 21403
rect 10968 21369 11002 21403
rect 13001 21369 13035 21403
rect 14013 21369 14047 21403
rect 19156 21369 19190 21403
rect 1961 21301 1995 21335
rect 2421 21301 2455 21335
rect 2973 21301 3007 21335
rect 3341 21301 3375 21335
rect 3433 21301 3467 21335
rect 4077 21301 4111 21335
rect 4445 21301 4479 21335
rect 4537 21301 4571 21335
rect 5273 21301 5307 21335
rect 5825 21301 5859 21335
rect 6285 21301 6319 21335
rect 6929 21301 6963 21335
rect 7389 21301 7423 21335
rect 8401 21301 8435 21335
rect 8769 21301 8803 21335
rect 12081 21301 12115 21335
rect 12633 21301 12667 21335
rect 14105 21301 14139 21335
rect 15025 21301 15059 21335
rect 15945 21301 15979 21335
rect 16497 21301 16531 21335
rect 16865 21301 16899 21335
rect 16957 21301 16991 21335
rect 18521 21301 18555 21335
rect 20269 21301 20303 21335
rect 20729 21301 20763 21335
rect 21557 21301 21591 21335
rect 21649 21301 21683 21335
rect 22385 21301 22419 21335
rect 1593 21097 1627 21131
rect 4445 21097 4479 21131
rect 7297 21097 7331 21131
rect 8953 21097 8987 21131
rect 17141 21097 17175 21131
rect 20545 21097 20579 21131
rect 4537 21029 4571 21063
rect 7818 21029 7852 21063
rect 10149 21029 10183 21063
rect 13360 21029 13394 21063
rect 19432 21029 19466 21063
rect 21180 21029 21214 21063
rect 1409 20961 1443 20995
rect 2228 20961 2262 20995
rect 5089 20961 5123 20995
rect 5917 20961 5951 20995
rect 6184 20961 6218 20995
rect 7573 20961 7607 20995
rect 10057 20961 10091 20995
rect 11336 20961 11370 20995
rect 13093 20961 13127 20995
rect 15557 20961 15591 20995
rect 16957 20961 16991 20995
rect 17509 20961 17543 20995
rect 17776 20961 17810 20995
rect 22569 20961 22603 20995
rect 1961 20893 1995 20927
rect 4721 20893 4755 20927
rect 10241 20893 10275 20927
rect 11069 20893 11103 20927
rect 15301 20893 15335 20927
rect 19165 20893 19199 20927
rect 20913 20893 20947 20927
rect 5273 20825 5307 20859
rect 3341 20757 3375 20791
rect 4077 20757 4111 20791
rect 9689 20757 9723 20791
rect 12449 20757 12483 20791
rect 14473 20757 14507 20791
rect 16681 20757 16715 20791
rect 18889 20757 18923 20791
rect 22293 20757 22327 20791
rect 3065 20553 3099 20587
rect 4813 20553 4847 20587
rect 6469 20553 6503 20587
rect 8217 20553 8251 20587
rect 9873 20553 9907 20587
rect 11805 20553 11839 20587
rect 14657 20553 14691 20587
rect 19441 20553 19475 20587
rect 16589 20485 16623 20519
rect 13277 20417 13311 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 20177 20417 20211 20451
rect 20361 20417 20395 20451
rect 1685 20349 1719 20383
rect 3433 20349 3467 20383
rect 3700 20349 3734 20383
rect 5089 20349 5123 20383
rect 5356 20349 5390 20383
rect 6837 20349 6871 20383
rect 7104 20349 7138 20383
rect 8493 20349 8527 20383
rect 8760 20349 8794 20383
rect 10425 20349 10459 20383
rect 10692 20349 10726 20383
rect 12725 20349 12759 20383
rect 13544 20349 13578 20383
rect 14933 20349 14967 20383
rect 15200 20349 15234 20383
rect 18061 20349 18095 20383
rect 20821 20349 20855 20383
rect 21088 20349 21122 20383
rect 22477 20349 22511 20383
rect 1952 20281 1986 20315
rect 16957 20281 16991 20315
rect 18328 20281 18362 20315
rect 20085 20281 20119 20315
rect 12909 20213 12943 20247
rect 16313 20213 16347 20247
rect 19717 20213 19751 20247
rect 22201 20213 22235 20247
rect 22661 20213 22695 20247
rect 3249 20009 3283 20043
rect 6285 20009 6319 20043
rect 6653 20009 6687 20043
rect 11805 20009 11839 20043
rect 13461 20009 13495 20043
rect 14013 20009 14047 20043
rect 19165 20009 19199 20043
rect 19901 20009 19935 20043
rect 4690 19941 4724 19975
rect 6745 19941 6779 19975
rect 8208 19941 8242 19975
rect 9689 19941 9723 19975
rect 12348 19941 12382 19975
rect 13921 19941 13955 19975
rect 15660 19941 15694 19975
rect 17233 19941 17267 19975
rect 19809 19941 19843 19975
rect 1409 19873 1443 19907
rect 1676 19873 1710 19907
rect 3065 19873 3099 19907
rect 7389 19873 7423 19907
rect 9873 19873 9907 19907
rect 10692 19873 10726 19907
rect 12081 19873 12115 19907
rect 14565 19873 14599 19907
rect 14749 19873 14783 19907
rect 17049 19873 17083 19907
rect 18052 19873 18086 19907
rect 21649 19873 21683 19907
rect 22293 19873 22327 19907
rect 22477 19873 22511 19907
rect 4445 19805 4479 19839
rect 6837 19805 6871 19839
rect 7941 19805 7975 19839
rect 10425 19805 10459 19839
rect 14197 19805 14231 19839
rect 15393 19805 15427 19839
rect 17785 19805 17819 19839
rect 20085 19805 20119 19839
rect 21741 19805 21775 19839
rect 21833 19805 21867 19839
rect 5825 19737 5859 19771
rect 16773 19737 16807 19771
rect 21281 19737 21315 19771
rect 2789 19669 2823 19703
rect 7573 19669 7607 19703
rect 9321 19669 9355 19703
rect 10057 19669 10091 19703
rect 13553 19669 13587 19703
rect 17417 19669 17451 19703
rect 19441 19669 19475 19703
rect 22661 19669 22695 19703
rect 2789 19465 2823 19499
rect 4445 19465 4479 19499
rect 8401 19465 8435 19499
rect 14289 19465 14323 19499
rect 19441 19465 19475 19499
rect 7573 19397 7607 19431
rect 5365 19329 5399 19363
rect 6285 19329 6319 19363
rect 8125 19329 8159 19363
rect 15117 19397 15151 19431
rect 10885 19329 10919 19363
rect 11897 19329 11931 19363
rect 13093 19329 13127 19363
rect 14749 19329 14783 19363
rect 14841 19329 14875 19363
rect 15761 19329 15795 19363
rect 16865 19329 16899 19363
rect 20269 19329 20303 19363
rect 1409 19261 1443 19295
rect 3065 19261 3099 19295
rect 3332 19261 3366 19295
rect 5089 19261 5123 19295
rect 7021 19261 7055 19295
rect 7941 19261 7975 19295
rect 8401 19261 8435 19295
rect 8585 19261 8619 19295
rect 12817 19261 12851 19295
rect 13737 19261 13771 19295
rect 15485 19261 15519 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 21005 19261 21039 19295
rect 21272 19261 21306 19295
rect 1676 19193 1710 19227
rect 5181 19193 5215 19227
rect 6101 19193 6135 19227
rect 8830 19193 8864 19227
rect 12909 19193 12943 19227
rect 15577 19193 15611 19227
rect 16773 19193 16807 19227
rect 18328 19193 18362 19227
rect 20085 19193 20119 19227
rect 20177 19193 20211 19227
rect 4721 19125 4755 19159
rect 5733 19125 5767 19159
rect 6193 19125 6227 19159
rect 7205 19125 7239 19159
rect 8033 19125 8067 19159
rect 9965 19125 9999 19159
rect 10333 19125 10367 19159
rect 10701 19125 10735 19159
rect 10793 19125 10827 19159
rect 11345 19125 11379 19159
rect 11713 19125 11747 19159
rect 11805 19125 11839 19159
rect 12449 19125 12483 19159
rect 13921 19125 13955 19159
rect 14657 19125 14691 19159
rect 16129 19125 16163 19159
rect 16313 19125 16347 19159
rect 16681 19125 16715 19159
rect 17601 19125 17635 19159
rect 19717 19125 19751 19159
rect 22385 19125 22419 19159
rect 3709 18921 3743 18955
rect 4445 18921 4479 18955
rect 4905 18921 4939 18955
rect 4537 18853 4571 18887
rect 1777 18785 1811 18819
rect 2329 18785 2363 18819
rect 2596 18785 2630 18819
rect 6745 18921 6779 18955
rect 9321 18921 9355 18955
rect 11621 18921 11655 18955
rect 18797 18921 18831 18955
rect 19533 18921 19567 18955
rect 7297 18853 7331 18887
rect 8208 18853 8242 18887
rect 12142 18853 12176 18887
rect 14013 18853 14047 18887
rect 21548 18853 21582 18887
rect 5457 18785 5491 18819
rect 6285 18785 6319 18819
rect 6745 18785 6779 18819
rect 7205 18785 7239 18819
rect 9689 18785 9723 18819
rect 10508 18785 10542 18819
rect 13921 18785 13955 18819
rect 14657 18785 14691 18819
rect 15393 18785 15427 18819
rect 15660 18785 15694 18819
rect 17417 18785 17451 18819
rect 17684 18785 17718 18819
rect 19441 18785 19475 18819
rect 20085 18785 20119 18819
rect 4721 18717 4755 18751
rect 4905 18717 4939 18751
rect 5549 18717 5583 18751
rect 5733 18717 5767 18751
rect 7481 18717 7515 18751
rect 7941 18717 7975 18751
rect 10241 18717 10275 18751
rect 11897 18717 11931 18751
rect 14105 18717 14139 18751
rect 19717 18717 19751 18751
rect 21281 18717 21315 18751
rect 1961 18649 1995 18683
rect 4077 18649 4111 18683
rect 5089 18581 5123 18615
rect 6469 18581 6503 18615
rect 6837 18581 6871 18615
rect 9873 18581 9907 18615
rect 13277 18581 13311 18615
rect 13553 18581 13587 18615
rect 14841 18581 14875 18615
rect 16773 18581 16807 18615
rect 19073 18581 19107 18615
rect 20269 18581 20303 18615
rect 22661 18581 22695 18615
rect 1961 18377 1995 18411
rect 8217 18377 8251 18411
rect 9965 18377 9999 18411
rect 11621 18377 11655 18411
rect 14381 18377 14415 18411
rect 19441 18377 19475 18411
rect 4261 18309 4295 18343
rect 9689 18309 9723 18343
rect 12633 18309 12667 18343
rect 20637 18309 20671 18343
rect 2329 18241 2363 18275
rect 4629 18241 4663 18275
rect 6837 18241 6871 18275
rect 7941 18241 7975 18275
rect 8217 18241 8251 18275
rect 11897 18241 11931 18275
rect 15209 18241 15243 18275
rect 16221 18241 16255 18275
rect 17325 18241 17359 18275
rect 18061 18241 18095 18275
rect 21189 18241 21223 18275
rect 22477 18241 22511 18275
rect 1777 18173 1811 18207
rect 4077 18173 4111 18207
rect 6285 18173 6319 18207
rect 8309 18173 8343 18207
rect 8576 18173 8610 18207
rect 10149 18173 10183 18207
rect 10241 18173 10275 18207
rect 10508 18173 10542 18207
rect 12449 18173 12483 18207
rect 12817 18173 12851 18207
rect 13001 18173 13035 18207
rect 17049 18173 17083 18207
rect 17877 18173 17911 18207
rect 20085 18173 20119 18207
rect 22293 18173 22327 18207
rect 2596 18105 2630 18139
rect 4874 18105 4908 18139
rect 7757 18105 7791 18139
rect 13268 18105 13302 18139
rect 15025 18105 15059 18139
rect 16129 18105 16163 18139
rect 18328 18105 18362 18139
rect 21097 18105 21131 18139
rect 3709 18037 3743 18071
rect 6009 18037 6043 18071
rect 7297 18037 7331 18071
rect 7665 18037 7699 18071
rect 12817 18037 12851 18071
rect 14657 18037 14691 18071
rect 15117 18037 15151 18071
rect 15669 18037 15703 18071
rect 16037 18037 16071 18071
rect 16681 18037 16715 18071
rect 17141 18037 17175 18071
rect 17693 18037 17727 18071
rect 20269 18037 20303 18071
rect 21005 18037 21039 18071
rect 21833 18037 21867 18071
rect 22201 18037 22235 18071
rect 3617 17833 3651 17867
rect 4445 17833 4479 17867
rect 8125 17833 8159 17867
rect 9873 17833 9907 17867
rect 11713 17833 11747 17867
rect 14289 17833 14323 17867
rect 16957 17833 16991 17867
rect 17325 17833 17359 17867
rect 18797 17833 18831 17867
rect 19533 17833 19567 17867
rect 20453 17833 20487 17867
rect 4077 17765 4111 17799
rect 10600 17765 10634 17799
rect 15546 17765 15580 17799
rect 1685 17697 1719 17731
rect 2237 17697 2271 17731
rect 2493 17697 2527 17731
rect 4261 17697 4295 17731
rect 5080 17697 5114 17731
rect 6725 17697 6759 17731
rect 8493 17697 8527 17731
rect 9689 17697 9723 17731
rect 11989 17697 12023 17731
rect 12909 17697 12943 17731
rect 13176 17697 13210 17731
rect 14657 17697 14691 17731
rect 19441 17765 19475 17799
rect 21640 17765 21674 17799
rect 17684 17697 17718 17731
rect 20269 17697 20303 17731
rect 4813 17629 4847 17663
rect 6469 17629 6503 17663
rect 8585 17629 8619 17663
rect 8677 17629 8711 17663
rect 9137 17629 9171 17663
rect 10333 17629 10367 17663
rect 15301 17629 15335 17663
rect 17325 17629 17359 17663
rect 17417 17629 17451 17663
rect 19717 17629 19751 17663
rect 20913 17629 20947 17663
rect 21373 17629 21407 17663
rect 4077 17561 4111 17595
rect 1869 17493 1903 17527
rect 6193 17493 6227 17527
rect 7849 17493 7883 17527
rect 12173 17493 12207 17527
rect 14841 17493 14875 17527
rect 16681 17493 16715 17527
rect 19073 17493 19107 17527
rect 22753 17493 22787 17527
rect 1777 17289 1811 17323
rect 3525 17289 3559 17323
rect 3617 17289 3651 17323
rect 11713 17289 11747 17323
rect 21649 17289 21683 17323
rect 2145 17153 2179 17187
rect 1593 17085 1627 17119
rect 2412 17017 2446 17051
rect 3801 17221 3835 17255
rect 5917 17221 5951 17255
rect 9873 17221 9907 17255
rect 14013 17221 14047 17255
rect 16497 17221 16531 17255
rect 16773 17221 16807 17255
rect 4353 17153 4387 17187
rect 5365 17153 5399 17187
rect 6837 17153 6871 17187
rect 8493 17153 8527 17187
rect 12633 17153 12667 17187
rect 14197 17153 14231 17187
rect 17325 17153 17359 17187
rect 19257 17153 19291 17187
rect 20269 17153 20303 17187
rect 22477 17153 22511 17187
rect 4169 17085 4203 17119
rect 6101 17085 6135 17119
rect 6193 17085 6227 17119
rect 10333 17085 10367 17119
rect 12900 17085 12934 17119
rect 5181 17017 5215 17051
rect 7104 17017 7138 17051
rect 8760 17017 8794 17051
rect 10600 17017 10634 17051
rect 14473 17085 14507 17119
rect 14565 17085 14599 17119
rect 15117 17085 15151 17119
rect 18061 17085 18095 17119
rect 18981 17085 19015 17119
rect 19717 17085 19751 17119
rect 20536 17085 20570 17119
rect 22293 17085 22327 17119
rect 15384 17017 15418 17051
rect 17233 17017 17267 17051
rect 22385 17017 22419 17051
rect 3617 16949 3651 16983
rect 4261 16949 4295 16983
rect 4813 16949 4847 16983
rect 5273 16949 5307 16983
rect 6377 16949 6411 16983
rect 8217 16949 8251 16983
rect 14197 16949 14231 16983
rect 14289 16949 14323 16983
rect 14749 16949 14783 16983
rect 17141 16949 17175 16983
rect 18245 16949 18279 16983
rect 18613 16949 18647 16983
rect 19073 16949 19107 16983
rect 19901 16949 19935 16983
rect 21925 16949 21959 16983
rect 1593 16745 1627 16779
rect 3341 16745 3375 16779
rect 4077 16745 4111 16779
rect 4445 16745 4479 16779
rect 4905 16745 4939 16779
rect 5089 16745 5123 16779
rect 11069 16745 11103 16779
rect 11253 16745 11287 16779
rect 11345 16745 11379 16779
rect 13369 16745 13403 16779
rect 13829 16745 13863 16779
rect 16681 16745 16715 16779
rect 16957 16745 16991 16779
rect 17417 16745 17451 16779
rect 19165 16745 19199 16779
rect 22569 16745 22603 16779
rect 4537 16677 4571 16711
rect 5549 16677 5583 16711
rect 6552 16677 6586 16711
rect 8208 16677 8242 16711
rect 18052 16677 18086 16711
rect 21180 16677 21214 16711
rect 1409 16609 1443 16643
rect 1961 16609 1995 16643
rect 2228 16609 2262 16643
rect 4905 16609 4939 16643
rect 5457 16609 5491 16643
rect 9945 16609 9979 16643
rect 11253 16609 11287 16643
rect 11529 16609 11563 16643
rect 11713 16609 11747 16643
rect 11980 16609 12014 16643
rect 13737 16609 13771 16643
rect 14657 16609 14691 16643
rect 15301 16609 15335 16643
rect 15568 16609 15602 16643
rect 17141 16609 17175 16643
rect 17233 16609 17267 16643
rect 19809 16609 19843 16643
rect 4629 16541 4663 16575
rect 5641 16541 5675 16575
rect 6285 16541 6319 16575
rect 7941 16541 7975 16575
rect 9689 16541 9723 16575
rect 13921 16541 13955 16575
rect 17785 16541 17819 16575
rect 19349 16541 19383 16575
rect 19901 16541 19935 16575
rect 20085 16541 20119 16575
rect 20913 16541 20947 16575
rect 9321 16473 9355 16507
rect 14841 16473 14875 16507
rect 7665 16405 7699 16439
rect 13093 16405 13127 16439
rect 19349 16405 19383 16439
rect 19441 16405 19475 16439
rect 22293 16405 22327 16439
rect 1685 16201 1719 16235
rect 3433 16201 3467 16235
rect 12633 16201 12667 16235
rect 22753 16201 22787 16235
rect 19441 16133 19475 16167
rect 4540 16065 4574 16099
rect 6837 16065 6871 16099
rect 7343 16065 7377 16099
rect 9276 16065 9310 16099
rect 9459 16065 9493 16099
rect 11621 16065 11655 16099
rect 13369 16065 13403 16099
rect 13692 16065 13726 16099
rect 13832 16065 13866 16099
rect 21373 16065 21407 16099
rect 1501 15997 1535 16031
rect 1961 15997 1995 16031
rect 2053 15997 2087 16031
rect 3985 15997 4019 16031
rect 4077 15997 4111 16031
rect 4813 15997 4847 16031
rect 6193 15997 6227 16031
rect 7573 15997 7607 16031
rect 8953 15997 8987 16031
rect 9689 15997 9723 16031
rect 12449 15997 12483 16031
rect 13277 15997 13311 16031
rect 14105 15997 14139 16031
rect 15577 15997 15611 16031
rect 17233 15997 17267 16031
rect 18061 15997 18095 16031
rect 19717 15997 19751 16031
rect 2320 15929 2354 15963
rect 15822 15929 15856 15963
rect 18328 15929 18362 15963
rect 19984 15929 20018 15963
rect 21618 15929 21652 15963
rect 1961 15861 1995 15895
rect 3801 15861 3835 15895
rect 4543 15861 4577 15895
rect 5917 15861 5951 15895
rect 6377 15861 6411 15895
rect 7303 15861 7337 15895
rect 8677 15861 8711 15895
rect 10793 15861 10827 15895
rect 11069 15861 11103 15895
rect 11437 15861 11471 15895
rect 11529 15861 11563 15895
rect 13093 15861 13127 15895
rect 15209 15861 15243 15895
rect 16957 15861 16991 15895
rect 17417 15861 17451 15895
rect 21097 15861 21131 15895
rect 4629 15657 4663 15691
rect 9229 15657 9263 15691
rect 10149 15657 10183 15691
rect 12909 15657 12943 15691
rect 14841 15657 14875 15691
rect 19349 15657 19383 15691
rect 19809 15657 19843 15691
rect 20177 15589 20211 15623
rect 22569 15589 22603 15623
rect 1501 15521 1535 15555
rect 1768 15521 1802 15555
rect 3157 15521 3191 15555
rect 4445 15521 4479 15555
rect 5320 15521 5354 15555
rect 5733 15521 5767 15555
rect 7113 15521 7147 15555
rect 7380 15521 7414 15555
rect 8953 15521 8987 15555
rect 9045 15521 9079 15555
rect 10057 15521 10091 15555
rect 10977 15521 11011 15555
rect 11069 15521 11103 15555
rect 11392 15521 11426 15555
rect 11805 15521 11839 15555
rect 13441 15521 13475 15555
rect 15025 15521 15059 15555
rect 15301 15521 15335 15555
rect 15624 15521 15658 15555
rect 17417 15521 17451 15555
rect 17969 15521 18003 15555
rect 18225 15521 18259 15555
rect 20269 15521 20303 15555
rect 21169 15521 21203 15555
rect 3341 15453 3375 15487
rect 4997 15453 5031 15487
rect 5503 15453 5537 15487
rect 6929 15453 6963 15487
rect 10333 15453 10367 15487
rect 11532 15453 11566 15487
rect 13185 15453 13219 15487
rect 15764 15453 15798 15487
rect 16037 15453 16071 15487
rect 20453 15453 20487 15487
rect 20913 15453 20947 15487
rect 8769 15385 8803 15419
rect 9689 15385 9723 15419
rect 17601 15385 17635 15419
rect 2881 15317 2915 15351
rect 6837 15317 6871 15351
rect 6929 15317 6963 15351
rect 8493 15317 8527 15351
rect 10793 15317 10827 15351
rect 14565 15317 14599 15351
rect 17141 15317 17175 15351
rect 22293 15317 22327 15351
rect 12081 15113 12115 15147
rect 12449 15113 12483 15147
rect 15025 15113 15059 15147
rect 21189 15113 21223 15147
rect 3801 15045 3835 15079
rect 22661 15045 22695 15079
rect 1869 14977 1903 15011
rect 4675 14977 4709 15011
rect 13001 14977 13035 15011
rect 15853 14977 15887 15011
rect 17417 14977 17451 15011
rect 17601 14977 17635 15011
rect 19855 14977 19889 15011
rect 22017 14977 22051 15011
rect 3617 14909 3651 14943
rect 4169 14909 4203 14943
rect 4905 14909 4939 14943
rect 6837 14909 6871 14943
rect 7104 14909 7138 14943
rect 8953 14909 8987 14943
rect 10701 14909 10735 14943
rect 10957 14909 10991 14943
rect 12909 14909 12943 14943
rect 13461 14909 13495 14943
rect 13717 14909 13751 14943
rect 15209 14909 15243 14943
rect 17325 14909 17359 14943
rect 18245 14909 18279 14943
rect 19349 14909 19383 14943
rect 19672 14909 19706 14943
rect 20085 14909 20119 14943
rect 22477 14909 22511 14943
rect 2136 14841 2170 14875
rect 6285 14841 6319 14875
rect 9220 14841 9254 14875
rect 15761 14841 15795 14875
rect 16313 14841 16347 14875
rect 16497 14841 16531 14875
rect 18889 14841 18923 14875
rect 1409 14773 1443 14807
rect 3249 14773 3283 14807
rect 4635 14773 4669 14807
rect 6009 14773 6043 14807
rect 8217 14773 8251 14807
rect 8493 14773 8527 14807
rect 10333 14773 10367 14807
rect 12817 14773 12851 14807
rect 14841 14773 14875 14807
rect 15301 14773 15335 14807
rect 15669 14773 15703 14807
rect 16957 14773 16991 14807
rect 21465 14773 21499 14807
rect 21833 14773 21867 14807
rect 21925 14773 21959 14807
rect 4445 14569 4479 14603
rect 4537 14569 4571 14603
rect 5089 14569 5123 14603
rect 8309 14569 8343 14603
rect 8677 14569 8711 14603
rect 9321 14569 9355 14603
rect 11529 14569 11563 14603
rect 11897 14569 11931 14603
rect 14381 14569 14415 14603
rect 1952 14501 1986 14535
rect 8769 14501 8803 14535
rect 10140 14501 10174 14535
rect 14289 14501 14323 14535
rect 16589 14501 16623 14535
rect 17325 14501 17359 14535
rect 21434 14501 21468 14535
rect 1685 14433 1719 14467
rect 3433 14433 3467 14467
rect 5457 14433 5491 14467
rect 6101 14433 6135 14467
rect 6909 14433 6943 14467
rect 9505 14433 9539 14467
rect 11989 14433 12023 14467
rect 12449 14433 12483 14467
rect 12716 14433 12750 14467
rect 14749 14433 14783 14467
rect 15669 14433 15703 14467
rect 15761 14433 15795 14467
rect 16497 14433 16531 14467
rect 17417 14433 17451 14467
rect 18052 14433 18086 14467
rect 19809 14433 19843 14467
rect 19901 14433 19935 14467
rect 20637 14433 20671 14467
rect 4629 14365 4663 14399
rect 4905 14365 4939 14399
rect 5549 14365 5583 14399
rect 5641 14365 5675 14399
rect 6653 14365 6687 14399
rect 8861 14365 8895 14399
rect 9873 14365 9907 14399
rect 12173 14365 12207 14399
rect 14473 14365 14507 14399
rect 15853 14365 15887 14399
rect 16681 14365 16715 14399
rect 17601 14365 17635 14399
rect 17785 14365 17819 14399
rect 19993 14365 20027 14399
rect 21189 14365 21223 14399
rect 3065 14297 3099 14331
rect 3617 14297 3651 14331
rect 6285 14297 6319 14331
rect 11253 14297 11287 14331
rect 16957 14297 16991 14331
rect 4077 14229 4111 14263
rect 4905 14229 4939 14263
rect 8033 14229 8067 14263
rect 13829 14229 13863 14263
rect 13921 14229 13955 14263
rect 14933 14229 14967 14263
rect 15301 14229 15335 14263
rect 16129 14229 16163 14263
rect 19165 14229 19199 14263
rect 19441 14229 19475 14263
rect 20453 14229 20487 14263
rect 22569 14229 22603 14263
rect 2881 14025 2915 14059
rect 6285 14025 6319 14059
rect 6837 14025 6871 14059
rect 10149 14025 10183 14059
rect 10701 14025 10735 14059
rect 12633 14025 12667 14059
rect 21557 14025 21591 14059
rect 9689 13957 9723 13991
rect 21833 13957 21867 13991
rect 1501 13889 1535 13923
rect 3709 13889 3743 13923
rect 4905 13889 4939 13923
rect 7389 13889 7423 13923
rect 11345 13889 11379 13923
rect 18061 13889 18095 13923
rect 20040 13889 20074 13923
rect 20223 13889 20257 13923
rect 22477 13889 22511 13923
rect 1768 13821 1802 13855
rect 4445 13821 4479 13855
rect 5172 13821 5206 13855
rect 7297 13821 7331 13855
rect 8309 13821 8343 13855
rect 8576 13821 8610 13855
rect 9965 13821 9999 13855
rect 11161 13821 11195 13855
rect 11713 13821 11747 13855
rect 12081 13821 12115 13855
rect 12449 13821 12483 13855
rect 12817 13821 12851 13855
rect 15853 13821 15887 13855
rect 16313 13821 16347 13855
rect 19717 13821 19751 13855
rect 20453 13821 20487 13855
rect 22293 13821 22327 13855
rect 3525 13753 3559 13787
rect 4261 13753 4295 13787
rect 7205 13753 7239 13787
rect 10425 13753 10459 13787
rect 11897 13753 11931 13787
rect 13084 13753 13118 13787
rect 16037 13753 16071 13787
rect 16580 13753 16614 13787
rect 18306 13753 18340 13787
rect 3157 13685 3191 13719
rect 3617 13685 3651 13719
rect 4629 13685 4663 13719
rect 7849 13685 7883 13719
rect 11069 13685 11103 13719
rect 14197 13685 14231 13719
rect 15301 13685 15335 13719
rect 17693 13685 17727 13719
rect 19441 13685 19475 13719
rect 22201 13685 22235 13719
rect 1869 13481 1903 13515
rect 2697 13481 2731 13515
rect 4077 13481 4111 13515
rect 5917 13481 5951 13515
rect 6377 13481 6411 13515
rect 10149 13481 10183 13515
rect 12081 13481 12115 13515
rect 19717 13481 19751 13515
rect 20913 13481 20947 13515
rect 4804 13413 4838 13447
rect 7012 13413 7046 13447
rect 13890 13413 13924 13447
rect 18512 13413 18546 13447
rect 21640 13413 21674 13447
rect 1685 13345 1719 13379
rect 2605 13345 2639 13379
rect 3433 13345 3467 13379
rect 6193 13345 6227 13379
rect 6745 13345 6779 13379
rect 8769 13345 8803 13379
rect 10057 13345 10091 13379
rect 10968 13345 11002 13379
rect 12173 13345 12207 13379
rect 12429 13345 12463 13379
rect 13645 13345 13679 13379
rect 15301 13345 15335 13379
rect 15557 13345 15591 13379
rect 16773 13345 16807 13379
rect 17029 13345 17063 13379
rect 18245 13345 18279 13379
rect 20085 13345 20119 13379
rect 20177 13345 20211 13379
rect 2789 13277 2823 13311
rect 4537 13277 4571 13311
rect 8861 13277 8895 13311
rect 8953 13277 8987 13311
rect 10333 13277 10367 13311
rect 10701 13277 10735 13311
rect 20269 13277 20303 13311
rect 21373 13277 21407 13311
rect 2237 13209 2271 13243
rect 9689 13209 9723 13243
rect 18153 13209 18187 13243
rect 3617 13141 3651 13175
rect 8125 13141 8159 13175
rect 8401 13141 8435 13175
rect 13553 13141 13587 13175
rect 15025 13141 15059 13175
rect 16681 13141 16715 13175
rect 19625 13141 19659 13175
rect 22753 13141 22787 13175
rect 5365 12937 5399 12971
rect 9505 12937 9539 12971
rect 11805 12937 11839 12971
rect 16589 12937 16623 12971
rect 22385 12937 22419 12971
rect 1685 12869 1719 12903
rect 5089 12869 5123 12903
rect 8493 12869 8527 12903
rect 14013 12869 14047 12903
rect 14197 12869 14231 12903
rect 20545 12869 20579 12903
rect 21189 12869 21223 12903
rect 3709 12801 3743 12835
rect 6009 12801 6043 12835
rect 9045 12801 9079 12835
rect 9965 12801 9999 12835
rect 10057 12801 10091 12835
rect 10425 12801 10459 12835
rect 14841 12801 14875 12835
rect 15209 12801 15243 12835
rect 17417 12801 17451 12835
rect 17601 12801 17635 12835
rect 21649 12801 21683 12835
rect 21833 12801 21867 12835
rect 1501 12733 1535 12767
rect 2053 12733 2087 12767
rect 2320 12733 2354 12767
rect 6837 12733 6871 12767
rect 7104 12733 7138 12767
rect 9873 12733 9907 12767
rect 10692 12733 10726 12767
rect 12265 12733 12299 12767
rect 12633 12733 12667 12767
rect 12900 12733 12934 12767
rect 18061 12733 18095 12767
rect 18245 12733 18279 12767
rect 18705 12733 18739 12767
rect 20361 12733 20395 12767
rect 22201 12733 22235 12767
rect 3976 12665 4010 12699
rect 5733 12665 5767 12699
rect 15476 12665 15510 12699
rect 18972 12665 19006 12699
rect 3433 12597 3467 12631
rect 5825 12597 5859 12631
rect 8217 12597 8251 12631
rect 8861 12597 8895 12631
rect 8953 12597 8987 12631
rect 12081 12597 12115 12631
rect 14565 12597 14599 12631
rect 14657 12597 14691 12631
rect 16957 12597 16991 12631
rect 17325 12597 17359 12631
rect 18429 12597 18463 12631
rect 20085 12597 20119 12631
rect 21557 12597 21591 12631
rect 3617 12393 3651 12427
rect 5089 12393 5123 12427
rect 5365 12393 5399 12427
rect 6193 12393 6227 12427
rect 6561 12393 6595 12427
rect 10057 12393 10091 12427
rect 10609 12393 10643 12427
rect 14933 12393 14967 12427
rect 16497 12393 16531 12427
rect 17049 12393 17083 12427
rect 19165 12393 19199 12427
rect 1860 12325 1894 12359
rect 4445 12325 4479 12359
rect 5733 12325 5767 12359
rect 9413 12325 9447 12359
rect 13185 12325 13219 12359
rect 19349 12325 19383 12359
rect 19901 12325 19935 12359
rect 22569 12325 22603 12359
rect 1593 12257 1627 12291
rect 3433 12257 3467 12291
rect 4997 12257 5031 12291
rect 5273 12257 5307 12291
rect 5825 12257 5859 12291
rect 6193 12257 6227 12291
rect 6377 12257 6411 12291
rect 7021 12257 7055 12291
rect 7288 12257 7322 12291
rect 8861 12257 8895 12291
rect 9045 12257 9079 12291
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 2973 12121 3007 12155
rect 5917 12189 5951 12223
rect 9873 12257 9907 12291
rect 10793 12257 10827 12291
rect 11437 12257 11471 12291
rect 13277 12257 13311 12291
rect 13533 12257 13567 12291
rect 14749 12257 14783 12291
rect 15485 12257 15519 12291
rect 16405 12257 16439 12291
rect 17509 12257 17543 12291
rect 17776 12257 17810 12291
rect 18981 12257 19015 12291
rect 16589 12189 16623 12223
rect 20913 12257 20947 12291
rect 21169 12257 21203 12291
rect 19993 12189 20027 12223
rect 20085 12189 20119 12223
rect 9229 12121 9263 12155
rect 9413 12121 9447 12155
rect 14657 12121 14691 12155
rect 15669 12121 15703 12155
rect 19349 12121 19383 12155
rect 4077 12053 4111 12087
rect 4997 12053 5031 12087
rect 8401 12053 8435 12087
rect 8677 12053 8711 12087
rect 16037 12053 16071 12087
rect 18889 12053 18923 12087
rect 19533 12053 19567 12087
rect 22293 12053 22327 12087
rect 2881 11849 2915 11883
rect 6653 11849 6687 11883
rect 9045 11849 9079 11883
rect 11805 11849 11839 11883
rect 15485 11849 15519 11883
rect 20913 11849 20947 11883
rect 4353 11781 4387 11815
rect 3801 11713 3835 11747
rect 5089 11713 5123 11747
rect 9413 11781 9447 11815
rect 15945 11781 15979 11815
rect 7205 11713 7239 11747
rect 10057 11713 10091 11747
rect 14381 11713 14415 11747
rect 14933 11713 14967 11747
rect 15117 11713 15151 11747
rect 16589 11713 16623 11747
rect 17509 11713 17543 11747
rect 18521 11713 18555 11747
rect 18705 11713 18739 11747
rect 19579 11713 19613 11747
rect 19809 11713 19843 11747
rect 1501 11645 1535 11679
rect 4169 11645 4203 11679
rect 4997 11645 5031 11679
rect 6653 11645 6687 11679
rect 8861 11645 8895 11679
rect 10425 11645 10459 11679
rect 11989 11645 12023 11679
rect 12633 11645 12667 11679
rect 15301 11645 15335 11679
rect 17417 11645 17451 11679
rect 19073 11645 19107 11679
rect 21373 11645 21407 11679
rect 1768 11577 1802 11611
rect 3617 11577 3651 11611
rect 5356 11577 5390 11611
rect 7450 11577 7484 11611
rect 9781 11577 9815 11611
rect 10692 11577 10726 11611
rect 14841 11577 14875 11611
rect 21640 11577 21674 11611
rect 3157 11509 3191 11543
rect 3525 11509 3559 11543
rect 4813 11509 4847 11543
rect 6469 11509 6503 11543
rect 8585 11509 8619 11543
rect 9873 11509 9907 11543
rect 12173 11509 12207 11543
rect 14473 11509 14507 11543
rect 16313 11509 16347 11543
rect 16405 11509 16439 11543
rect 16957 11509 16991 11543
rect 17325 11509 17359 11543
rect 18061 11509 18095 11543
rect 18429 11509 18463 11543
rect 19539 11509 19573 11543
rect 22753 11509 22787 11543
rect 2881 11305 2915 11339
rect 3617 11305 3651 11339
rect 6561 11305 6595 11339
rect 9229 11305 9263 11339
rect 10149 11305 10183 11339
rect 11897 11305 11931 11339
rect 12633 11305 12667 11339
rect 19809 11305 19843 11339
rect 22661 11305 22695 11339
rect 1768 11237 1802 11271
rect 1501 11169 1535 11203
rect 3341 11169 3375 11203
rect 3433 11169 3467 11203
rect 4445 11169 4479 11203
rect 4537 11169 4571 11203
rect 5181 11169 5215 11203
rect 5448 11169 5482 11203
rect 7564 11169 7598 11203
rect 9033 11169 9067 11203
rect 9965 11169 9999 11203
rect 10333 11169 10367 11203
rect 10784 11169 10818 11203
rect 12265 11169 12299 11203
rect 4721 11101 4755 11135
rect 6837 11101 6871 11135
rect 7297 11101 7331 11135
rect 4077 11033 4111 11067
rect 8677 11033 8711 11067
rect 10517 11101 10551 11135
rect 13062 11237 13096 11271
rect 21548 11237 21582 11271
rect 14657 11169 14691 11203
rect 15925 11169 15959 11203
rect 17325 11169 17359 11203
rect 20085 11169 20119 11203
rect 21281 11169 21315 11203
rect 12817 11101 12851 11135
rect 15669 11101 15703 11135
rect 17969 11101 18003 11135
rect 18292 11101 18326 11135
rect 18432 11101 18466 11135
rect 18705 11101 18739 11135
rect 12449 11033 12483 11067
rect 12633 11033 12667 11067
rect 14841 11033 14875 11067
rect 20269 11033 20303 11067
rect 3157 10965 3191 10999
rect 10333 10965 10367 10999
rect 14197 10965 14231 10999
rect 17049 10965 17083 10999
rect 17509 10965 17543 10999
rect 3065 10761 3099 10795
rect 4721 10761 4755 10795
rect 6377 10761 6411 10795
rect 7021 10761 7055 10795
rect 20913 10761 20947 10795
rect 9597 10693 9631 10727
rect 17325 10693 17359 10727
rect 1685 10625 1719 10659
rect 4997 10625 5031 10659
rect 9965 10625 9999 10659
rect 15945 10625 15979 10659
rect 18705 10625 18739 10659
rect 18889 10625 18923 10659
rect 19533 10625 19567 10659
rect 21925 10625 21959 10659
rect 3341 10557 3375 10591
rect 3608 10557 3642 10591
rect 6837 10557 6871 10591
rect 7481 10557 7515 10591
rect 9321 10557 9355 10591
rect 9413 10557 9447 10591
rect 11805 10557 11839 10591
rect 12633 10557 12667 10591
rect 12889 10557 12923 10591
rect 14289 10557 14323 10591
rect 14556 10557 14590 10591
rect 16212 10557 16246 10591
rect 17785 10557 17819 10591
rect 18613 10557 18647 10591
rect 19800 10557 19834 10591
rect 21833 10557 21867 10591
rect 22385 10557 22419 10591
rect 1952 10489 1986 10523
rect 5264 10489 5298 10523
rect 7726 10489 7760 10523
rect 10232 10489 10266 10523
rect 21189 10489 21223 10523
rect 21741 10489 21775 10523
rect 8861 10421 8895 10455
rect 9137 10421 9171 10455
rect 11345 10421 11379 10455
rect 11989 10421 12023 10455
rect 14013 10421 14047 10455
rect 15669 10421 15703 10455
rect 17601 10421 17635 10455
rect 18245 10421 18279 10455
rect 19257 10421 19291 10455
rect 21373 10421 21407 10455
rect 22569 10421 22603 10455
rect 1593 10217 1627 10251
rect 5549 10217 5583 10251
rect 7205 10217 7239 10251
rect 11345 10217 11379 10251
rect 12081 10217 12115 10251
rect 14565 10217 14599 10251
rect 16865 10217 16899 10251
rect 21465 10217 21499 10251
rect 22293 10217 22327 10251
rect 4436 10149 4470 10183
rect 6092 10149 6126 10183
rect 7849 10149 7883 10183
rect 9956 10149 9990 10183
rect 12173 10149 12207 10183
rect 15752 10149 15786 10183
rect 17693 10149 17727 10183
rect 22201 10149 22235 10183
rect 2053 10081 2087 10115
rect 2320 10081 2354 10115
rect 4169 10081 4203 10115
rect 5825 10081 5859 10115
rect 8197 10081 8231 10115
rect 11529 10081 11563 10115
rect 12992 10081 13026 10115
rect 14381 10081 14415 10115
rect 15117 10081 15151 10115
rect 17601 10081 17635 10115
rect 18245 10081 18279 10115
rect 18512 10081 18546 10115
rect 19901 10081 19935 10115
rect 20637 10081 20671 10115
rect 21281 10081 21315 10115
rect 7849 10013 7883 10047
rect 7941 10013 7975 10047
rect 9689 10013 9723 10047
rect 12265 10013 12299 10047
rect 12725 10013 12759 10047
rect 15485 10013 15519 10047
rect 17877 10013 17911 10047
rect 22477 10013 22511 10047
rect 11713 9945 11747 9979
rect 20085 9945 20119 9979
rect 20453 9945 20487 9979
rect 3433 9877 3467 9911
rect 9321 9877 9355 9911
rect 11069 9877 11103 9911
rect 14105 9877 14139 9911
rect 14933 9877 14967 9911
rect 17233 9877 17267 9911
rect 19625 9877 19659 9911
rect 21833 9877 21867 9911
rect 16865 9673 16899 9707
rect 2789 9605 2823 9639
rect 4445 9605 4479 9639
rect 7021 9605 7055 9639
rect 7757 9605 7791 9639
rect 11805 9605 11839 9639
rect 12081 9605 12115 9639
rect 14105 9605 14139 9639
rect 14381 9605 14415 9639
rect 16681 9605 16715 9639
rect 1409 9537 1443 9571
rect 3065 9537 3099 9571
rect 5641 9537 5675 9571
rect 5733 9537 5767 9571
rect 8401 9537 8435 9571
rect 10425 9537 10459 9571
rect 3332 9469 3366 9503
rect 6193 9469 6227 9503
rect 6837 9469 6871 9503
rect 8769 9469 8803 9503
rect 10681 9469 10715 9503
rect 12265 9469 12299 9503
rect 12725 9469 12759 9503
rect 14565 9469 14599 9503
rect 14657 9469 14691 9503
rect 15301 9469 15335 9503
rect 15568 9469 15602 9503
rect 1654 9401 1688 9435
rect 5549 9401 5583 9435
rect 8217 9401 8251 9435
rect 9014 9401 9048 9435
rect 12970 9401 13004 9435
rect 14841 9401 14875 9435
rect 18981 9673 19015 9707
rect 16957 9605 16991 9639
rect 17601 9537 17635 9571
rect 17877 9537 17911 9571
rect 18797 9537 18831 9571
rect 17417 9401 17451 9435
rect 18521 9469 18555 9503
rect 18613 9469 18647 9503
rect 22753 9605 22787 9639
rect 19671 9537 19705 9571
rect 19901 9537 19935 9571
rect 21373 9537 21407 9571
rect 19165 9469 19199 9503
rect 19488 9469 19522 9503
rect 21640 9401 21674 9435
rect 5181 9333 5215 9367
rect 6377 9333 6411 9367
rect 8125 9333 8159 9367
rect 10149 9333 10183 9367
rect 15025 9333 15059 9367
rect 16865 9333 16899 9367
rect 17325 9333 17359 9367
rect 17877 9333 17911 9367
rect 18153 9333 18187 9367
rect 18981 9333 19015 9367
rect 21005 9333 21039 9367
rect 2237 9129 2271 9163
rect 3249 9129 3283 9163
rect 4077 9129 4111 9163
rect 4445 9129 4479 9163
rect 5089 9129 5123 9163
rect 5457 9129 5491 9163
rect 6377 9129 6411 9163
rect 6929 9129 6963 9163
rect 7389 9129 7423 9163
rect 7573 9129 7607 9163
rect 9689 9129 9723 9163
rect 10609 9129 10643 9163
rect 12541 9129 12575 9163
rect 13369 9129 13403 9163
rect 15945 9129 15979 9163
rect 22661 9129 22695 9163
rect 5549 9061 5583 9095
rect 7021 9061 7055 9095
rect 7941 9061 7975 9095
rect 9045 9061 9079 9095
rect 9505 9061 9539 9095
rect 10149 9061 10183 9095
rect 3341 8993 3375 9027
rect 8953 8993 8987 9027
rect 2329 8925 2363 8959
rect 2513 8925 2547 8959
rect 3525 8925 3559 8959
rect 4537 8925 4571 8959
rect 4629 8925 4663 8959
rect 5733 8925 5767 8959
rect 7205 8925 7239 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 9229 8925 9263 8959
rect 2881 8857 2915 8891
rect 10057 8993 10091 9027
rect 10241 8925 10275 8959
rect 1869 8789 1903 8823
rect 6561 8789 6595 8823
rect 8585 8789 8619 8823
rect 9505 8789 9539 8823
rect 11069 9061 11103 9095
rect 12909 9061 12943 9095
rect 11713 8993 11747 9027
rect 12449 8993 12483 9027
rect 13001 8993 13035 9027
rect 21526 9061 21560 9095
rect 13809 8993 13843 9027
rect 15853 8993 15887 9027
rect 16497 8993 16531 9027
rect 16753 8993 16787 9027
rect 20637 8993 20671 9027
rect 21281 8993 21315 9027
rect 11161 8925 11195 8959
rect 11253 8925 11287 8959
rect 13093 8925 13127 8959
rect 13369 8925 13403 8959
rect 13553 8925 13587 8959
rect 16129 8925 16163 8959
rect 18337 8925 18371 8959
rect 18660 8925 18694 8959
rect 18800 8925 18834 8959
rect 19073 8925 19107 8959
rect 10701 8857 10735 8891
rect 20177 8857 20211 8891
rect 10609 8789 10643 8823
rect 11897 8789 11931 8823
rect 12265 8789 12299 8823
rect 14933 8789 14967 8823
rect 15485 8789 15519 8823
rect 17877 8789 17911 8823
rect 20453 8789 20487 8823
rect 2881 8585 2915 8619
rect 4721 8585 4755 8619
rect 15209 8585 15243 8619
rect 18153 8585 18187 8619
rect 20545 8585 20579 8619
rect 22201 8585 22235 8619
rect 5733 8517 5767 8551
rect 7665 8517 7699 8551
rect 8677 8517 8711 8551
rect 11161 8517 11195 8551
rect 11345 8517 11379 8551
rect 13001 8517 13035 8551
rect 14749 8517 14783 8551
rect 22661 8517 22695 8551
rect 3341 8449 3375 8483
rect 3525 8449 3559 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 6377 8449 6411 8483
rect 8125 8449 8159 8483
rect 8217 8449 8251 8483
rect 9321 8449 9355 8483
rect 11897 8449 11931 8483
rect 13369 8449 13403 8483
rect 15577 8449 15611 8483
rect 17509 8449 17543 8483
rect 18797 8449 18831 8483
rect 3249 8381 3283 8415
rect 5089 8381 5123 8415
rect 6101 8381 6135 8415
rect 7113 8381 7147 8415
rect 9045 8381 9079 8415
rect 9689 8381 9723 8415
rect 11161 8381 11195 8415
rect 12817 8381 12851 8415
rect 15025 8381 15059 8415
rect 15833 8381 15867 8415
rect 17233 8381 17267 8415
rect 18613 8381 18647 8415
rect 19165 8381 19199 8415
rect 20821 8381 20855 8415
rect 21077 8381 21111 8415
rect 22477 8381 22511 8415
rect 6193 8313 6227 8347
rect 9137 8313 9171 8347
rect 9956 8313 9990 8347
rect 11713 8313 11747 8347
rect 13636 8313 13670 8347
rect 19410 8313 19444 8347
rect 7297 8245 7331 8279
rect 8033 8245 8067 8279
rect 11069 8245 11103 8279
rect 11805 8245 11839 8279
rect 16957 8245 16991 8279
rect 18521 8245 18555 8279
rect 6561 8041 6595 8075
rect 7021 8041 7055 8075
rect 7389 8041 7423 8075
rect 8585 8041 8619 8075
rect 9045 8041 9079 8075
rect 12725 8041 12759 8075
rect 14381 8041 14415 8075
rect 14841 8041 14875 8075
rect 16405 8041 16439 8075
rect 16957 8041 16991 8075
rect 19349 8041 19383 8075
rect 22201 8041 22235 8075
rect 2513 7905 2547 7939
rect 4721 7905 4755 7939
rect 5825 7905 5859 7939
rect 6469 7905 6503 7939
rect 6929 7905 6963 7939
rect 3157 7837 3191 7871
rect 4905 7837 4939 7871
rect 7205 7837 7239 7871
rect 8953 7973 8987 8007
rect 9956 7973 9990 8007
rect 13268 7973 13302 8007
rect 16313 7973 16347 8007
rect 17325 7973 17359 8007
rect 18214 7973 18248 8007
rect 21281 7973 21315 8007
rect 7941 7905 7975 7939
rect 11601 7905 11635 7939
rect 12817 7905 12851 7939
rect 13001 7905 13035 7939
rect 14657 7905 14691 7939
rect 15393 7905 15427 7939
rect 17969 7905 18003 7939
rect 19993 7905 20027 7939
rect 21005 7905 21039 7939
rect 22109 7905 22143 7939
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 9137 7837 9171 7871
rect 9689 7837 9723 7871
rect 11345 7837 11379 7871
rect 6009 7769 6043 7803
rect 7389 7769 7423 7803
rect 7573 7769 7607 7803
rect 11069 7769 11103 7803
rect 16589 7837 16623 7871
rect 17417 7837 17451 7871
rect 17601 7837 17635 7871
rect 20085 7837 20119 7871
rect 20177 7837 20211 7871
rect 22385 7837 22419 7871
rect 15945 7769 15979 7803
rect 12817 7701 12851 7735
rect 15577 7701 15611 7735
rect 19625 7701 19659 7735
rect 21741 7701 21775 7735
rect 4721 7497 4755 7531
rect 5733 7497 5767 7531
rect 7481 7497 7515 7531
rect 12449 7497 12483 7531
rect 14841 7497 14875 7531
rect 15301 7497 15335 7531
rect 17693 7497 17727 7531
rect 3709 7429 3743 7463
rect 4261 7361 4295 7395
rect 5181 7361 5215 7395
rect 5365 7361 5399 7395
rect 6377 7361 6411 7395
rect 8125 7361 8159 7395
rect 12909 7361 12943 7395
rect 13093 7361 13127 7395
rect 15853 7361 15887 7395
rect 16316 7361 16350 7395
rect 18892 7361 18926 7395
rect 19165 7361 19199 7395
rect 4077 7293 4111 7327
rect 6101 7293 6135 7327
rect 7029 7293 7063 7327
rect 8493 7293 8527 7327
rect 10149 7293 10183 7327
rect 11805 7293 11839 7327
rect 13461 7293 13495 7327
rect 15117 7293 15151 7327
rect 16589 7293 16623 7327
rect 18429 7293 18463 7327
rect 20545 7293 20579 7327
rect 22201 7293 22235 7327
rect 6193 7225 6227 7259
rect 7389 7225 7423 7259
rect 7849 7225 7883 7259
rect 8760 7225 8794 7259
rect 10416 7225 10450 7259
rect 12817 7225 12851 7259
rect 13728 7225 13762 7259
rect 20790 7225 20824 7259
rect 22477 7225 22511 7259
rect 4169 7157 4203 7191
rect 5089 7157 5123 7191
rect 6837 7157 6871 7191
rect 7941 7157 7975 7191
rect 9873 7157 9907 7191
rect 11529 7157 11563 7191
rect 11989 7157 12023 7191
rect 16319 7157 16353 7191
rect 18895 7157 18929 7191
rect 20269 7157 20303 7191
rect 21925 7157 21959 7191
rect 4537 6953 4571 6987
rect 5917 6953 5951 6987
rect 6929 6953 6963 6987
rect 4905 6885 4939 6919
rect 7941 6885 7975 6919
rect 12909 6885 12943 6919
rect 22569 6885 22603 6919
rect 4997 6817 5031 6851
rect 7021 6817 7055 6851
rect 8033 6817 8067 6851
rect 8953 6817 8987 6851
rect 9873 6817 9907 6851
rect 10425 6817 10459 6851
rect 10692 6817 10726 6851
rect 13553 6817 13587 6851
rect 13820 6817 13854 6851
rect 15925 6817 15959 6851
rect 18052 6817 18086 6851
rect 19809 6817 19843 6851
rect 20913 6817 20947 6851
rect 21169 6817 21203 6851
rect 5089 6749 5123 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 7205 6749 7239 6783
rect 8125 6749 8159 6783
rect 9045 6749 9079 6783
rect 9137 6749 9171 6783
rect 12081 6749 12115 6783
rect 13001 6749 13035 6783
rect 13185 6749 13219 6783
rect 15669 6749 15703 6783
rect 17325 6749 17359 6783
rect 17785 6749 17819 6783
rect 19901 6749 19935 6783
rect 19993 6749 20027 6783
rect 5549 6681 5583 6715
rect 6561 6681 6595 6715
rect 8585 6681 8619 6715
rect 7573 6613 7607 6647
rect 10057 6613 10091 6647
rect 11805 6613 11839 6647
rect 12541 6613 12575 6647
rect 14933 6613 14967 6647
rect 17049 6613 17083 6647
rect 19165 6613 19199 6647
rect 19441 6613 19475 6647
rect 22293 6613 22327 6647
rect 5641 6409 5675 6443
rect 7665 6409 7699 6443
rect 9689 6409 9723 6443
rect 17417 6341 17451 6375
rect 18429 6341 18463 6375
rect 20637 6341 20671 6375
rect 6101 6273 6135 6307
rect 6285 6273 6319 6307
rect 8217 6273 8251 6307
rect 9321 6273 9355 6307
rect 10333 6273 10367 6307
rect 10701 6273 10735 6307
rect 12725 6273 12759 6307
rect 16037 6273 16071 6307
rect 6009 6205 6043 6239
rect 8033 6205 8067 6239
rect 8125 6205 8159 6239
rect 9045 6205 9079 6239
rect 10968 6205 11002 6239
rect 14381 6205 14415 6239
rect 16293 6205 16327 6239
rect 17877 6205 17911 6239
rect 18245 6205 18279 6239
rect 18797 6205 18831 6239
rect 19064 6205 19098 6239
rect 21373 6205 21407 6239
rect 9137 6137 9171 6171
rect 12992 6137 13026 6171
rect 14648 6137 14682 6171
rect 20637 6137 20671 6171
rect 20729 6137 20763 6171
rect 20913 6137 20947 6171
rect 21618 6137 21652 6171
rect 8677 6069 8711 6103
rect 10057 6069 10091 6103
rect 10149 6069 10183 6103
rect 12081 6069 12115 6103
rect 14105 6069 14139 6103
rect 15761 6069 15795 6103
rect 17693 6069 17727 6103
rect 20177 6069 20211 6103
rect 21097 6069 21131 6103
rect 22753 6069 22787 6103
rect 5917 5865 5951 5899
rect 6285 5865 6319 5899
rect 6377 5865 6411 5899
rect 8033 5865 8067 5899
rect 8585 5865 8619 5899
rect 9045 5865 9079 5899
rect 13645 5865 13679 5899
rect 14381 5865 14415 5899
rect 14933 5865 14967 5899
rect 16037 5865 16071 5899
rect 18521 5865 18555 5899
rect 19257 5865 19291 5899
rect 21097 5865 21131 5899
rect 21833 5865 21867 5899
rect 8953 5797 8987 5831
rect 7941 5729 7975 5763
rect 10057 5729 10091 5763
rect 10609 5729 10643 5763
rect 10876 5729 10910 5763
rect 12521 5729 12555 5763
rect 14289 5729 14323 5763
rect 15117 5729 15151 5763
rect 15577 5729 15611 5763
rect 16037 5729 16071 5763
rect 16497 5729 16531 5763
rect 16589 5729 16623 5763
rect 17408 5729 17442 5763
rect 19165 5729 19199 5763
rect 20177 5729 20211 5763
rect 20269 5729 20303 5763
rect 20913 5729 20947 5763
rect 21925 5729 21959 5763
rect 22293 5729 22327 5763
rect 22477 5729 22511 5763
rect 6469 5661 6503 5695
rect 8217 5661 8251 5695
rect 9229 5661 9263 5695
rect 12265 5661 12299 5695
rect 14473 5661 14507 5695
rect 16773 5661 16807 5695
rect 17141 5661 17175 5695
rect 19441 5661 19475 5695
rect 20453 5661 20487 5695
rect 22017 5661 22051 5695
rect 7573 5593 7607 5627
rect 11989 5593 12023 5627
rect 15761 5593 15795 5627
rect 19809 5593 19843 5627
rect 22661 5593 22695 5627
rect 10241 5525 10275 5559
rect 13921 5525 13955 5559
rect 16129 5525 16163 5559
rect 18797 5525 18831 5559
rect 21465 5525 21499 5559
rect 22293 5525 22327 5559
rect 7481 5321 7515 5355
rect 11161 5321 11195 5355
rect 12449 5321 12483 5355
rect 13369 5321 13403 5355
rect 14841 5321 14875 5355
rect 19257 5321 19291 5355
rect 19625 5321 19659 5355
rect 22569 5321 22603 5355
rect 8033 5185 8067 5219
rect 9045 5185 9079 5219
rect 10609 5185 10643 5219
rect 10701 5185 10735 5219
rect 11621 5185 11655 5219
rect 11713 5185 11747 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 18061 5253 18095 5287
rect 15209 5185 15243 5219
rect 17417 5185 17451 5219
rect 18613 5185 18647 5219
rect 20085 5185 20119 5219
rect 20177 5185 20211 5219
rect 8861 5117 8895 5151
rect 10517 5117 10551 5151
rect 11529 5117 11563 5151
rect 12817 5117 12851 5151
rect 13369 5117 13403 5151
rect 13461 5117 13495 5151
rect 13728 5117 13762 5151
rect 17325 5117 17359 5151
rect 18521 5117 18555 5151
rect 19073 5117 19107 5151
rect 20637 5117 20671 5151
rect 21189 5117 21223 5151
rect 7849 5049 7883 5083
rect 8953 5049 8987 5083
rect 15454 5049 15488 5083
rect 21456 5049 21490 5083
rect 7941 4981 7975 5015
rect 8493 4981 8527 5015
rect 10149 4981 10183 5015
rect 16589 4981 16623 5015
rect 16865 4981 16899 5015
rect 17233 4981 17267 5015
rect 18429 4981 18463 5015
rect 19993 4981 20027 5015
rect 20821 4981 20855 5015
rect 9873 4777 9907 4811
rect 10333 4777 10367 4811
rect 11345 4777 11379 4811
rect 12265 4777 12299 4811
rect 12909 4777 12943 4811
rect 13277 4777 13311 4811
rect 13921 4777 13955 4811
rect 14381 4777 14415 4811
rect 15301 4777 15335 4811
rect 18153 4777 18187 4811
rect 19165 4777 19199 4811
rect 19809 4777 19843 4811
rect 20177 4777 20211 4811
rect 22477 4777 22511 4811
rect 11253 4709 11287 4743
rect 13369 4709 13403 4743
rect 14289 4709 14323 4743
rect 18245 4709 18279 4743
rect 10241 4641 10275 4675
rect 12357 4641 12391 4675
rect 15761 4641 15795 4675
rect 16017 4641 16051 4675
rect 19257 4641 19291 4675
rect 20269 4641 20303 4675
rect 21364 4641 21398 4675
rect 10517 4573 10551 4607
rect 11529 4573 11563 4607
rect 12449 4573 12483 4607
rect 13461 4573 13495 4607
rect 14473 4573 14507 4607
rect 18337 4573 18371 4607
rect 19349 4573 19383 4607
rect 20361 4573 20395 4607
rect 21097 4573 21131 4607
rect 10885 4505 10919 4539
rect 18797 4505 18831 4539
rect 11897 4437 11931 4471
rect 17141 4437 17175 4471
rect 17785 4437 17819 4471
rect 10333 4165 10367 4199
rect 10977 4097 11011 4131
rect 11897 4097 11931 4131
rect 13277 4097 13311 4131
rect 13553 4097 13587 4131
rect 14289 4097 14323 4131
rect 14657 4097 14691 4131
rect 16313 4097 16347 4131
rect 18613 4097 18647 4131
rect 19073 4097 19107 4131
rect 10701 4029 10735 4063
rect 11805 4029 11839 4063
rect 16569 4029 16603 4063
rect 19533 4029 19567 4063
rect 21373 4029 21407 4063
rect 21640 4029 21674 4063
rect 10793 3961 10827 3995
rect 14013 3961 14047 3995
rect 14924 3961 14958 3995
rect 18521 3961 18555 3995
rect 19778 3961 19812 3995
rect 11345 3893 11379 3927
rect 11713 3893 11747 3927
rect 12633 3893 12667 3927
rect 13001 3893 13035 3927
rect 13093 3893 13127 3927
rect 13645 3893 13679 3927
rect 14105 3893 14139 3927
rect 16037 3893 16071 3927
rect 17693 3893 17727 3927
rect 18061 3893 18095 3927
rect 18429 3893 18463 3927
rect 20913 3893 20947 3927
rect 22753 3893 22787 3927
rect 11161 3689 11195 3723
rect 12541 3689 12575 3723
rect 15945 3689 15979 3723
rect 16129 3689 16163 3723
rect 16497 3689 16531 3723
rect 22753 3689 22787 3723
rect 13093 3621 13127 3655
rect 13553 3621 13587 3655
rect 13645 3621 13679 3655
rect 11529 3553 11563 3587
rect 12633 3553 12667 3587
rect 11621 3485 11655 3519
rect 11805 3485 11839 3519
rect 12817 3485 12851 3519
rect 12173 3417 12207 3451
rect 14565 3553 14599 3587
rect 14657 3553 14691 3587
rect 15577 3553 15611 3587
rect 13737 3485 13771 3519
rect 14749 3485 14783 3519
rect 17408 3621 17442 3655
rect 20913 3621 20947 3655
rect 19248 3553 19282 3587
rect 21373 3553 21407 3587
rect 21640 3553 21674 3587
rect 16589 3485 16623 3519
rect 16681 3485 16715 3519
rect 17141 3485 17175 3519
rect 18981 3485 19015 3519
rect 15945 3417 15979 3451
rect 13093 3349 13127 3383
rect 13185 3349 13219 3383
rect 14197 3349 14231 3383
rect 15761 3349 15795 3383
rect 18521 3349 18555 3383
rect 20361 3349 20395 3383
rect 13277 3145 13311 3179
rect 15301 3145 15335 3179
rect 17693 3145 17727 3179
rect 19625 3145 19659 3179
rect 22109 3145 22143 3179
rect 14289 3077 14323 3111
rect 22569 3077 22603 3111
rect 1961 3009 1995 3043
rect 13921 3009 13955 3043
rect 14749 3009 14783 3043
rect 14933 3009 14967 3043
rect 15945 3009 15979 3043
rect 16313 3009 16347 3043
rect 20729 3009 20763 3043
rect 1777 2941 1811 2975
rect 2519 2941 2553 2975
rect 5089 2941 5123 2975
rect 13645 2941 13679 2975
rect 15669 2941 15703 2975
rect 16580 2941 16614 2975
rect 18245 2941 18279 2975
rect 19993 2941 20027 2975
rect 22385 2941 22419 2975
rect 14657 2873 14691 2907
rect 18512 2873 18546 2907
rect 20269 2873 20303 2907
rect 20974 2873 21008 2907
rect 2697 2805 2731 2839
rect 13737 2805 13771 2839
rect 15761 2805 15795 2839
rect 13369 2601 13403 2635
rect 13829 2601 13863 2635
rect 14841 2601 14875 2635
rect 16221 2601 16255 2635
rect 16681 2601 16715 2635
rect 17601 2601 17635 2635
rect 19717 2601 19751 2635
rect 20085 2601 20119 2635
rect 20545 2601 20579 2635
rect 22569 2601 22603 2635
rect 14749 2533 14783 2567
rect 16589 2533 16623 2567
rect 18604 2533 18638 2567
rect 13737 2465 13771 2499
rect 15669 2465 15703 2499
rect 18337 2465 18371 2499
rect 20453 2465 20487 2499
rect 21189 2465 21223 2499
rect 21445 2465 21479 2499
rect 13921 2397 13955 2431
rect 15025 2397 15059 2431
rect 16865 2397 16899 2431
rect 17693 2397 17727 2431
rect 17785 2397 17819 2431
rect 20637 2397 20671 2431
rect 14381 2261 14415 2295
rect 15853 2261 15887 2295
rect 17233 2261 17267 2295
<< metal1 >>
rect 9950 21904 9956 21956
rect 10008 21944 10014 21956
rect 16942 21944 16948 21956
rect 10008 21916 16948 21944
rect 10008 21904 10014 21916
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 13722 21876 13728 21888
rect 11112 21848 13728 21876
rect 11112 21836 11118 21848
rect 13722 21836 13728 21848
rect 13780 21836 13786 21888
rect 18322 21836 18328 21888
rect 18380 21876 18386 21888
rect 20438 21876 20444 21888
rect 18380 21848 20444 21876
rect 18380 21836 18386 21848
rect 20438 21836 20444 21848
rect 20496 21836 20502 21888
rect 1104 21786 23276 21808
rect 1104 21734 4680 21786
rect 4732 21734 4744 21786
rect 4796 21734 4808 21786
rect 4860 21734 4872 21786
rect 4924 21734 12078 21786
rect 12130 21734 12142 21786
rect 12194 21734 12206 21786
rect 12258 21734 12270 21786
rect 12322 21734 19475 21786
rect 19527 21734 19539 21786
rect 19591 21734 19603 21786
rect 19655 21734 19667 21786
rect 19719 21734 23276 21786
rect 1104 21712 23276 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1544 21644 1593 21672
rect 1544 21632 1550 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 9950 21672 9956 21684
rect 9911 21644 9956 21672
rect 1581 21635 1639 21641
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 15473 21675 15531 21681
rect 15473 21641 15485 21675
rect 15519 21672 15531 21675
rect 16390 21672 16396 21684
rect 15519 21644 16396 21672
rect 15519 21641 15531 21644
rect 15473 21635 15531 21641
rect 16390 21632 16396 21644
rect 16448 21632 16454 21684
rect 17865 21675 17923 21681
rect 17865 21641 17877 21675
rect 17911 21672 17923 21675
rect 19242 21672 19248 21684
rect 17911 21644 19248 21672
rect 17911 21641 17923 21644
rect 17865 21635 17923 21641
rect 19242 21632 19248 21644
rect 19300 21632 19306 21684
rect 13633 21607 13691 21613
rect 13633 21573 13645 21607
rect 13679 21604 13691 21607
rect 16758 21604 16764 21616
rect 13679 21576 16764 21604
rect 13679 21573 13691 21576
rect 13633 21567 13691 21573
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 21177 21607 21235 21613
rect 21177 21573 21189 21607
rect 21223 21604 21235 21607
rect 21818 21604 21824 21616
rect 21223 21576 21824 21604
rect 21223 21573 21235 21576
rect 21177 21567 21235 21573
rect 21818 21564 21824 21576
rect 21876 21564 21882 21616
rect 2590 21536 2596 21548
rect 2551 21508 2596 21536
rect 2590 21496 2596 21508
rect 2648 21496 2654 21548
rect 3605 21539 3663 21545
rect 3605 21505 3617 21539
rect 3651 21536 3663 21539
rect 4617 21539 4675 21545
rect 4617 21536 4629 21539
rect 3651 21508 4629 21536
rect 3651 21505 3663 21508
rect 3605 21499 3663 21505
rect 4617 21505 4629 21508
rect 4663 21536 4675 21539
rect 5534 21536 5540 21548
rect 4663 21508 5540 21536
rect 4663 21505 4675 21508
rect 4617 21499 4675 21505
rect 5534 21496 5540 21508
rect 5592 21536 5598 21548
rect 6365 21539 6423 21545
rect 6365 21536 6377 21539
rect 5592 21508 6377 21536
rect 5592 21496 5598 21508
rect 6365 21505 6377 21508
rect 6411 21536 6423 21539
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 6411 21508 7481 21536
rect 6411 21505 6423 21508
rect 6365 21499 6423 21505
rect 7469 21505 7481 21508
rect 7515 21536 7527 21539
rect 8941 21539 8999 21545
rect 8941 21536 8953 21539
rect 7515 21508 8953 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 8941 21505 8953 21508
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 14182 21536 14188 21548
rect 13311 21508 14188 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 14182 21496 14188 21508
rect 14240 21496 14246 21548
rect 16114 21536 16120 21548
rect 16075 21508 16120 21536
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 16574 21496 16580 21548
rect 16632 21536 16638 21548
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16632 21508 17049 21536
rect 16632 21496 16638 21508
rect 17037 21505 17049 21508
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 21450 21496 21456 21548
rect 21508 21536 21514 21548
rect 21729 21539 21787 21545
rect 21729 21536 21741 21539
rect 21508 21508 21741 21536
rect 21508 21496 21514 21508
rect 21729 21505 21741 21508
rect 21775 21505 21787 21539
rect 21729 21499 21787 21505
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 4154 21428 4160 21480
rect 4212 21468 4218 21480
rect 5074 21468 5080 21480
rect 4212 21440 5080 21468
rect 4212 21428 4218 21440
rect 5074 21428 5080 21440
rect 5132 21428 5138 21480
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 5184 21440 7941 21468
rect 2317 21403 2375 21409
rect 2317 21369 2329 21403
rect 2363 21400 2375 21403
rect 2590 21400 2596 21412
rect 2363 21372 2596 21400
rect 2363 21369 2375 21372
rect 2317 21363 2375 21369
rect 2590 21360 2596 21372
rect 2648 21360 2654 21412
rect 3786 21360 3792 21412
rect 3844 21400 3850 21412
rect 5184 21400 5212 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21468 9827 21471
rect 9950 21468 9956 21480
rect 9815 21440 9956 21468
rect 9815 21437 9827 21440
rect 9769 21431 9827 21437
rect 9950 21428 9956 21440
rect 10008 21428 10014 21480
rect 10410 21428 10416 21480
rect 10468 21468 10474 21480
rect 10689 21471 10747 21477
rect 10689 21468 10701 21471
rect 10468 21440 10701 21468
rect 10468 21428 10474 21440
rect 10689 21437 10701 21440
rect 10735 21437 10747 21471
rect 10689 21431 10747 21437
rect 12158 21428 12164 21480
rect 12216 21468 12222 21480
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12216 21440 13093 21468
rect 12216 21428 12222 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 14826 21468 14832 21480
rect 14787 21440 14832 21468
rect 13081 21431 13139 21437
rect 14826 21428 14832 21440
rect 14884 21428 14890 21480
rect 15470 21428 15476 21480
rect 15528 21468 15534 21480
rect 15841 21471 15899 21477
rect 15841 21468 15853 21471
rect 15528 21440 15853 21468
rect 15528 21428 15534 21440
rect 15841 21437 15853 21440
rect 15887 21437 15899 21471
rect 15841 21431 15899 21437
rect 17681 21471 17739 21477
rect 17681 21437 17693 21471
rect 17727 21468 17739 21471
rect 18230 21468 18236 21480
rect 17727 21440 18236 21468
rect 17727 21437 17739 21440
rect 17681 21431 17739 21437
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 18380 21440 18425 21468
rect 18380 21428 18386 21440
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 18877 21471 18935 21477
rect 18877 21468 18889 21471
rect 18840 21440 18889 21468
rect 18840 21428 18846 21440
rect 18877 21437 18889 21440
rect 18923 21437 18935 21471
rect 19886 21468 19892 21480
rect 18877 21431 18935 21437
rect 18984 21440 19892 21468
rect 3844 21372 5212 21400
rect 6181 21403 6239 21409
rect 3844 21360 3850 21372
rect 6181 21369 6193 21403
rect 6227 21400 6239 21403
rect 6454 21400 6460 21412
rect 6227 21372 6460 21400
rect 6227 21369 6239 21372
rect 6181 21363 6239 21369
rect 6454 21360 6460 21372
rect 6512 21360 6518 21412
rect 7285 21403 7343 21409
rect 7285 21369 7297 21403
rect 7331 21400 7343 21403
rect 7742 21400 7748 21412
rect 7331 21372 7748 21400
rect 7331 21369 7343 21372
rect 7285 21363 7343 21369
rect 7742 21360 7748 21372
rect 7800 21360 7806 21412
rect 8846 21400 8852 21412
rect 8807 21372 8852 21400
rect 8846 21360 8852 21372
rect 8904 21360 8910 21412
rect 10956 21403 11014 21409
rect 10956 21369 10968 21403
rect 11002 21400 11014 21403
rect 11698 21400 11704 21412
rect 11002 21372 11704 21400
rect 11002 21369 11014 21372
rect 10956 21363 11014 21369
rect 11698 21360 11704 21372
rect 11756 21400 11762 21412
rect 12989 21403 13047 21409
rect 12989 21400 13001 21403
rect 11756 21372 13001 21400
rect 11756 21360 11762 21372
rect 12989 21369 13001 21372
rect 13035 21369 13047 21403
rect 12989 21363 13047 21369
rect 14001 21403 14059 21409
rect 14001 21369 14013 21403
rect 14047 21400 14059 21403
rect 14458 21400 14464 21412
rect 14047 21372 14464 21400
rect 14047 21369 14059 21372
rect 14001 21363 14059 21369
rect 14458 21360 14464 21372
rect 14516 21360 14522 21412
rect 18984 21400 19012 21440
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 20530 21468 20536 21480
rect 20491 21440 20536 21468
rect 20530 21428 20536 21440
rect 20588 21428 20594 21480
rect 22189 21471 22247 21477
rect 22189 21437 22201 21471
rect 22235 21468 22247 21471
rect 22278 21468 22284 21480
rect 22235 21440 22284 21468
rect 22235 21437 22247 21440
rect 22189 21431 22247 21437
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 15028 21372 19012 21400
rect 19144 21403 19202 21409
rect 1946 21332 1952 21344
rect 1907 21304 1952 21332
rect 1946 21292 1952 21304
rect 2004 21292 2010 21344
rect 2409 21335 2467 21341
rect 2409 21301 2421 21335
rect 2455 21332 2467 21335
rect 2498 21332 2504 21344
rect 2455 21304 2504 21332
rect 2455 21301 2467 21304
rect 2409 21295 2467 21301
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 2958 21332 2964 21344
rect 2919 21304 2964 21332
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 3326 21332 3332 21344
rect 3287 21304 3332 21332
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 3418 21292 3424 21344
rect 3476 21332 3482 21344
rect 4062 21332 4068 21344
rect 3476 21304 3521 21332
rect 4023 21304 4068 21332
rect 3476 21292 3482 21304
rect 4062 21292 4068 21304
rect 4120 21292 4126 21344
rect 4430 21332 4436 21344
rect 4391 21304 4436 21332
rect 4430 21292 4436 21304
rect 4488 21292 4494 21344
rect 4522 21292 4528 21344
rect 4580 21332 4586 21344
rect 5258 21332 5264 21344
rect 4580 21304 4625 21332
rect 5219 21304 5264 21332
rect 4580 21292 4586 21304
rect 5258 21292 5264 21304
rect 5316 21292 5322 21344
rect 5810 21332 5816 21344
rect 5771 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 5902 21292 5908 21344
rect 5960 21332 5966 21344
rect 6273 21335 6331 21341
rect 6273 21332 6285 21335
rect 5960 21304 6285 21332
rect 5960 21292 5966 21304
rect 6273 21301 6285 21304
rect 6319 21301 6331 21335
rect 6914 21332 6920 21344
rect 6875 21304 6920 21332
rect 6273 21295 6331 21301
rect 6914 21292 6920 21304
rect 6972 21292 6978 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 8389 21335 8447 21341
rect 7432 21304 7477 21332
rect 7432 21292 7438 21304
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 8662 21332 8668 21344
rect 8435 21304 8668 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 8754 21292 8760 21344
rect 8812 21332 8818 21344
rect 12069 21335 12127 21341
rect 8812 21304 8857 21332
rect 8812 21292 8818 21304
rect 12069 21301 12081 21335
rect 12115 21332 12127 21335
rect 12250 21332 12256 21344
rect 12115 21304 12256 21332
rect 12115 21301 12127 21304
rect 12069 21295 12127 21301
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 12621 21335 12679 21341
rect 12621 21301 12633 21335
rect 12667 21332 12679 21335
rect 12894 21332 12900 21344
rect 12667 21304 12900 21332
rect 12667 21301 12679 21304
rect 12621 21295 12679 21301
rect 12894 21292 12900 21304
rect 12952 21292 12958 21344
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 15028 21341 15056 21372
rect 19144 21369 19156 21403
rect 19190 21400 19202 21403
rect 19334 21400 19340 21412
rect 19190 21372 19340 21400
rect 19190 21369 19202 21372
rect 19144 21363 19202 21369
rect 19334 21360 19340 21372
rect 19392 21360 19398 21412
rect 20346 21400 20352 21412
rect 19444 21372 20352 21400
rect 14093 21335 14151 21341
rect 14093 21332 14105 21335
rect 13780 21304 14105 21332
rect 13780 21292 13786 21304
rect 14093 21301 14105 21304
rect 14139 21301 14151 21335
rect 14093 21295 14151 21301
rect 15013 21335 15071 21341
rect 15013 21301 15025 21335
rect 15059 21301 15071 21335
rect 15013 21295 15071 21301
rect 15562 21292 15568 21344
rect 15620 21332 15626 21344
rect 15933 21335 15991 21341
rect 15933 21332 15945 21335
rect 15620 21304 15945 21332
rect 15620 21292 15626 21304
rect 15933 21301 15945 21304
rect 15979 21301 15991 21335
rect 15933 21295 15991 21301
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 16485 21335 16543 21341
rect 16485 21332 16497 21335
rect 16264 21304 16497 21332
rect 16264 21292 16270 21304
rect 16485 21301 16497 21304
rect 16531 21301 16543 21335
rect 16850 21332 16856 21344
rect 16811 21304 16856 21332
rect 16485 21295 16543 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 18509 21335 18567 21341
rect 17000 21304 17045 21332
rect 17000 21292 17006 21304
rect 18509 21301 18521 21335
rect 18555 21332 18567 21335
rect 19444 21332 19472 21372
rect 20346 21360 20352 21372
rect 20404 21360 20410 21412
rect 21910 21400 21916 21412
rect 20732 21372 21916 21400
rect 20254 21332 20260 21344
rect 18555 21304 19472 21332
rect 20215 21304 20260 21332
rect 18555 21301 18567 21304
rect 18509 21295 18567 21301
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 20732 21341 20760 21372
rect 21910 21360 21916 21372
rect 21968 21360 21974 21412
rect 20717 21335 20775 21341
rect 20717 21301 20729 21335
rect 20763 21301 20775 21335
rect 21542 21332 21548 21344
rect 21503 21304 21548 21332
rect 20717 21295 20775 21301
rect 21542 21292 21548 21304
rect 21600 21292 21606 21344
rect 21634 21292 21640 21344
rect 21692 21332 21698 21344
rect 22373 21335 22431 21341
rect 21692 21304 21737 21332
rect 21692 21292 21698 21304
rect 22373 21301 22385 21335
rect 22419 21332 22431 21335
rect 23198 21332 23204 21344
rect 22419 21304 23204 21332
rect 22419 21301 22431 21304
rect 22373 21295 22431 21301
rect 23198 21292 23204 21304
rect 23256 21292 23262 21344
rect 1104 21242 23276 21264
rect 1104 21190 8379 21242
rect 8431 21190 8443 21242
rect 8495 21190 8507 21242
rect 8559 21190 8571 21242
rect 8623 21190 15776 21242
rect 15828 21190 15840 21242
rect 15892 21190 15904 21242
rect 15956 21190 15968 21242
rect 16020 21190 23276 21242
rect 1104 21168 23276 21190
rect 290 21088 296 21140
rect 348 21128 354 21140
rect 1581 21131 1639 21137
rect 1581 21128 1593 21131
rect 348 21100 1593 21128
rect 348 21088 354 21100
rect 1581 21097 1593 21100
rect 1627 21097 1639 21131
rect 1581 21091 1639 21097
rect 4062 21088 4068 21140
rect 4120 21128 4126 21140
rect 4433 21131 4491 21137
rect 4433 21128 4445 21131
rect 4120 21100 4445 21128
rect 4120 21088 4126 21100
rect 4433 21097 4445 21100
rect 4479 21097 4491 21131
rect 4433 21091 4491 21097
rect 7285 21131 7343 21137
rect 7285 21097 7297 21131
rect 7331 21128 7343 21131
rect 7374 21128 7380 21140
rect 7331 21100 7380 21128
rect 7331 21097 7343 21100
rect 7285 21091 7343 21097
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 8941 21131 8999 21137
rect 8941 21128 8953 21131
rect 8904 21100 8953 21128
rect 8904 21088 8910 21100
rect 8941 21097 8953 21100
rect 8987 21097 8999 21131
rect 8941 21091 8999 21097
rect 9030 21088 9036 21140
rect 9088 21128 9094 21140
rect 16482 21128 16488 21140
rect 9088 21100 16488 21128
rect 9088 21088 9094 21100
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 17129 21131 17187 21137
rect 17129 21097 17141 21131
rect 17175 21128 17187 21131
rect 19150 21128 19156 21140
rect 17175 21100 19156 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 19150 21088 19156 21100
rect 19208 21088 19214 21140
rect 20346 21128 20352 21140
rect 19352 21100 20352 21128
rect 2958 21020 2964 21072
rect 3016 21060 3022 21072
rect 4525 21063 4583 21069
rect 4525 21060 4537 21063
rect 3016 21032 4537 21060
rect 3016 21020 3022 21032
rect 4525 21029 4537 21032
rect 4571 21029 4583 21063
rect 5442 21060 5448 21072
rect 4525 21023 4583 21029
rect 4632 21032 5448 21060
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20961 1455 20995
rect 1397 20955 1455 20961
rect 2216 20995 2274 21001
rect 2216 20961 2228 20995
rect 2262 20992 2274 20995
rect 3418 20992 3424 21004
rect 2262 20964 3424 20992
rect 2262 20961 2274 20964
rect 2216 20955 2274 20961
rect 1412 20856 1440 20955
rect 3418 20952 3424 20964
rect 3476 20952 3482 21004
rect 1486 20884 1492 20936
rect 1544 20924 1550 20936
rect 1949 20927 2007 20933
rect 1949 20924 1961 20927
rect 1544 20896 1961 20924
rect 1544 20884 1550 20896
rect 1949 20893 1961 20896
rect 1995 20893 2007 20927
rect 4338 20924 4344 20936
rect 1949 20887 2007 20893
rect 3160 20896 4344 20924
rect 1412 20828 1992 20856
rect 1964 20788 1992 20828
rect 3160 20788 3188 20896
rect 4338 20884 4344 20896
rect 4396 20924 4402 20936
rect 4632 20924 4660 21032
rect 5442 21020 5448 21032
rect 5500 21020 5506 21072
rect 5920 21032 6776 21060
rect 5077 20995 5135 21001
rect 5077 20961 5089 20995
rect 5123 20992 5135 20995
rect 5166 20992 5172 21004
rect 5123 20964 5172 20992
rect 5123 20961 5135 20964
rect 5077 20955 5135 20961
rect 5166 20952 5172 20964
rect 5224 20952 5230 21004
rect 5920 21001 5948 21032
rect 6748 21004 6776 21032
rect 7742 21020 7748 21072
rect 7800 21069 7806 21072
rect 7800 21063 7864 21069
rect 7800 21029 7818 21063
rect 7852 21029 7864 21063
rect 7800 21023 7864 21029
rect 7800 21020 7806 21023
rect 8662 21020 8668 21072
rect 8720 21060 8726 21072
rect 10137 21063 10195 21069
rect 10137 21060 10149 21063
rect 8720 21032 10149 21060
rect 8720 21020 8726 21032
rect 10137 21029 10149 21032
rect 10183 21029 10195 21063
rect 10137 21023 10195 21029
rect 13348 21063 13406 21069
rect 13348 21029 13360 21063
rect 13394 21060 13406 21063
rect 13722 21060 13728 21072
rect 13394 21032 13728 21060
rect 13394 21029 13406 21032
rect 13348 21023 13406 21029
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 18046 21060 18052 21072
rect 17512 21032 18052 21060
rect 5905 20995 5963 21001
rect 5905 20961 5917 20995
rect 5951 20961 5963 20995
rect 5905 20955 5963 20961
rect 6172 20995 6230 21001
rect 6172 20961 6184 20995
rect 6218 20992 6230 20995
rect 6454 20992 6460 21004
rect 6218 20964 6460 20992
rect 6218 20961 6230 20964
rect 6172 20955 6230 20961
rect 6454 20952 6460 20964
rect 6512 20952 6518 21004
rect 6730 20952 6736 21004
rect 6788 20992 6794 21004
rect 7561 20995 7619 21001
rect 7561 20992 7573 20995
rect 6788 20964 7573 20992
rect 6788 20952 6794 20964
rect 7561 20961 7573 20964
rect 7607 20961 7619 20995
rect 10042 20992 10048 21004
rect 10003 20964 10048 20992
rect 7561 20955 7619 20961
rect 10042 20952 10048 20964
rect 10100 20952 10106 21004
rect 11324 20995 11382 21001
rect 11324 20961 11336 20995
rect 11370 20992 11382 20995
rect 12250 20992 12256 21004
rect 11370 20964 12256 20992
rect 11370 20961 11382 20964
rect 11324 20955 11382 20961
rect 12250 20952 12256 20964
rect 12308 20952 12314 21004
rect 13081 20995 13139 21001
rect 13081 20961 13093 20995
rect 13127 20992 13139 20995
rect 13170 20992 13176 21004
rect 13127 20964 13176 20992
rect 13127 20961 13139 20964
rect 13081 20955 13139 20961
rect 13170 20952 13176 20964
rect 13228 20992 13234 21004
rect 13228 20964 14596 20992
rect 13228 20952 13234 20964
rect 4396 20896 4660 20924
rect 4709 20927 4767 20933
rect 4396 20884 4402 20896
rect 4709 20893 4721 20927
rect 4755 20924 4767 20927
rect 10229 20927 10287 20933
rect 4755 20896 5856 20924
rect 4755 20893 4767 20896
rect 4709 20887 4767 20893
rect 3970 20816 3976 20868
rect 4028 20856 4034 20868
rect 5261 20859 5319 20865
rect 5261 20856 5273 20859
rect 4028 20828 5273 20856
rect 4028 20816 4034 20828
rect 5261 20825 5273 20828
rect 5307 20825 5319 20859
rect 5261 20819 5319 20825
rect 3326 20788 3332 20800
rect 1964 20760 3188 20788
rect 3287 20760 3332 20788
rect 3326 20748 3332 20760
rect 3384 20748 3390 20800
rect 4065 20791 4123 20797
rect 4065 20757 4077 20791
rect 4111 20788 4123 20791
rect 4246 20788 4252 20800
rect 4111 20760 4252 20788
rect 4111 20757 4123 20760
rect 4065 20751 4123 20757
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 5828 20788 5856 20896
rect 10229 20893 10241 20927
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 10244 20856 10272 20887
rect 10410 20884 10416 20936
rect 10468 20924 10474 20936
rect 11057 20927 11115 20933
rect 11057 20924 11069 20927
rect 10468 20896 11069 20924
rect 10468 20884 10474 20896
rect 11057 20893 11069 20896
rect 11103 20893 11115 20927
rect 14568 20924 14596 20964
rect 14642 20952 14648 21004
rect 14700 20992 14706 21004
rect 15545 20995 15603 21001
rect 15545 20992 15557 20995
rect 14700 20964 15557 20992
rect 14700 20952 14706 20964
rect 15545 20961 15557 20964
rect 15591 20961 15603 20995
rect 15545 20955 15603 20961
rect 16945 20995 17003 21001
rect 16945 20961 16957 20995
rect 16991 20992 17003 20995
rect 17310 20992 17316 21004
rect 16991 20964 17316 20992
rect 16991 20961 17003 20964
rect 16945 20955 17003 20961
rect 17310 20952 17316 20964
rect 17368 20952 17374 21004
rect 17512 21001 17540 21032
rect 18046 21020 18052 21032
rect 18104 21020 18110 21072
rect 18230 21020 18236 21072
rect 18288 21060 18294 21072
rect 19352 21060 19380 21100
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 20533 21131 20591 21137
rect 20533 21097 20545 21131
rect 20579 21097 20591 21131
rect 20533 21091 20591 21097
rect 18288 21032 19380 21060
rect 19420 21063 19478 21069
rect 18288 21020 18294 21032
rect 19420 21029 19432 21063
rect 19466 21060 19478 21063
rect 20254 21060 20260 21072
rect 19466 21032 20260 21060
rect 19466 21029 19478 21032
rect 19420 21023 19478 21029
rect 20254 21020 20260 21032
rect 20312 21020 20318 21072
rect 20548 21060 20576 21091
rect 21168 21063 21226 21069
rect 21168 21060 21180 21063
rect 20548 21032 21180 21060
rect 21168 21029 21180 21032
rect 21214 21060 21226 21063
rect 21634 21060 21640 21072
rect 21214 21032 21640 21060
rect 21214 21029 21226 21032
rect 21168 21023 21226 21029
rect 21634 21020 21640 21032
rect 21692 21020 21698 21072
rect 17497 20995 17555 21001
rect 17497 20961 17509 20995
rect 17543 20961 17555 20995
rect 17497 20955 17555 20961
rect 17764 20995 17822 21001
rect 17764 20961 17776 20995
rect 17810 20992 17822 20995
rect 19794 20992 19800 21004
rect 17810 20964 19800 20992
rect 17810 20961 17822 20964
rect 17764 20955 17822 20961
rect 19794 20952 19800 20964
rect 19852 20952 19858 21004
rect 20622 20952 20628 21004
rect 20680 20992 20686 21004
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 20680 20964 22569 20992
rect 20680 20952 20686 20964
rect 22557 20961 22569 20964
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 14918 20924 14924 20936
rect 14568 20896 14924 20924
rect 11057 20887 11115 20893
rect 14918 20884 14924 20896
rect 14976 20924 14982 20936
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 14976 20896 15301 20924
rect 14976 20884 14982 20896
rect 15289 20893 15301 20896
rect 15335 20893 15347 20927
rect 15289 20887 15347 20893
rect 18782 20884 18788 20936
rect 18840 20924 18846 20936
rect 19150 20924 19156 20936
rect 18840 20896 19156 20924
rect 18840 20884 18846 20896
rect 19150 20884 19156 20896
rect 19208 20884 19214 20936
rect 20898 20924 20904 20936
rect 20859 20896 20904 20924
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 8496 20828 10272 20856
rect 6822 20788 6828 20800
rect 5828 20760 6828 20788
rect 6822 20748 6828 20760
rect 6880 20788 6886 20800
rect 8496 20788 8524 20828
rect 12250 20816 12256 20868
rect 12308 20856 12314 20868
rect 12308 20828 12664 20856
rect 12308 20816 12314 20828
rect 6880 20760 8524 20788
rect 9677 20791 9735 20797
rect 6880 20748 6886 20760
rect 9677 20757 9689 20791
rect 9723 20788 9735 20791
rect 9766 20788 9772 20800
rect 9723 20760 9772 20788
rect 9723 20757 9735 20760
rect 9677 20751 9735 20757
rect 9766 20748 9772 20760
rect 9824 20748 9830 20800
rect 12437 20791 12495 20797
rect 12437 20757 12449 20791
rect 12483 20788 12495 20791
rect 12526 20788 12532 20800
rect 12483 20760 12532 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 12636 20788 12664 20828
rect 13998 20788 14004 20800
rect 12636 20760 14004 20788
rect 13998 20748 14004 20760
rect 14056 20748 14062 20800
rect 14458 20788 14464 20800
rect 14419 20760 14464 20788
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 16669 20791 16727 20797
rect 16669 20788 16681 20791
rect 15252 20760 16681 20788
rect 15252 20748 15258 20760
rect 16669 20757 16681 20760
rect 16715 20757 16727 20791
rect 16669 20751 16727 20757
rect 18877 20791 18935 20797
rect 18877 20757 18889 20791
rect 18923 20788 18935 20791
rect 19334 20788 19340 20800
rect 18923 20760 19340 20788
rect 18923 20757 18935 20760
rect 18877 20751 18935 20757
rect 19334 20748 19340 20760
rect 19392 20788 19398 20800
rect 20162 20788 20168 20800
rect 19392 20760 20168 20788
rect 19392 20748 19398 20760
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 21542 20748 21548 20800
rect 21600 20788 21606 20800
rect 22281 20791 22339 20797
rect 22281 20788 22293 20791
rect 21600 20760 22293 20788
rect 21600 20748 21606 20760
rect 22281 20757 22293 20760
rect 22327 20757 22339 20791
rect 22281 20751 22339 20757
rect 1104 20698 23276 20720
rect 1104 20646 4680 20698
rect 4732 20646 4744 20698
rect 4796 20646 4808 20698
rect 4860 20646 4872 20698
rect 4924 20646 12078 20698
rect 12130 20646 12142 20698
rect 12194 20646 12206 20698
rect 12258 20646 12270 20698
rect 12322 20646 19475 20698
rect 19527 20646 19539 20698
rect 19591 20646 19603 20698
rect 19655 20646 19667 20698
rect 19719 20646 23276 20698
rect 1104 20624 23276 20646
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 3418 20584 3424 20596
rect 3099 20556 3424 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 3602 20544 3608 20596
rect 3660 20584 3666 20596
rect 3660 20556 4384 20584
rect 3660 20544 3666 20556
rect 4356 20516 4384 20556
rect 4430 20544 4436 20596
rect 4488 20584 4494 20596
rect 4801 20587 4859 20593
rect 4801 20584 4813 20587
rect 4488 20556 4813 20584
rect 4488 20544 4494 20556
rect 4801 20553 4813 20556
rect 4847 20553 4859 20587
rect 6454 20584 6460 20596
rect 4801 20547 4859 20553
rect 4908 20556 6132 20584
rect 6415 20556 6460 20584
rect 4908 20516 4936 20556
rect 4356 20488 4936 20516
rect 6104 20448 6132 20556
rect 6454 20544 6460 20556
rect 6512 20544 6518 20596
rect 7742 20544 7748 20596
rect 7800 20584 7806 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7800 20556 8217 20584
rect 7800 20544 7806 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 8205 20547 8263 20553
rect 8754 20544 8760 20596
rect 8812 20584 8818 20596
rect 9861 20587 9919 20593
rect 9861 20584 9873 20587
rect 8812 20556 9873 20584
rect 8812 20544 8818 20556
rect 9861 20553 9873 20556
rect 9907 20553 9919 20587
rect 9861 20547 9919 20553
rect 11698 20544 11704 20596
rect 11756 20584 11762 20596
rect 11793 20587 11851 20593
rect 11793 20584 11805 20587
rect 11756 20556 11805 20584
rect 11756 20544 11762 20556
rect 11793 20553 11805 20556
rect 11839 20553 11851 20587
rect 14642 20584 14648 20596
rect 14603 20556 14648 20584
rect 11793 20547 11851 20553
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 19242 20584 19248 20596
rect 14936 20556 19248 20584
rect 6104 20420 6960 20448
rect 1394 20340 1400 20392
rect 1452 20380 1458 20392
rect 1673 20383 1731 20389
rect 1673 20380 1685 20383
rect 1452 20352 1685 20380
rect 1452 20340 1458 20352
rect 1673 20349 1685 20352
rect 1719 20380 1731 20383
rect 3050 20380 3056 20392
rect 1719 20352 3056 20380
rect 1719 20349 1731 20352
rect 1673 20343 1731 20349
rect 3050 20340 3056 20352
rect 3108 20380 3114 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3108 20352 3433 20380
rect 3108 20340 3114 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 3688 20383 3746 20389
rect 3688 20349 3700 20383
rect 3734 20380 3746 20383
rect 4522 20380 4528 20392
rect 3734 20352 4528 20380
rect 3734 20349 3746 20352
rect 3688 20343 3746 20349
rect 1940 20315 1998 20321
rect 1940 20281 1952 20315
rect 1986 20312 1998 20315
rect 2314 20312 2320 20324
rect 1986 20284 2320 20312
rect 1986 20281 1998 20284
rect 1940 20275 1998 20281
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 3436 20312 3464 20343
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 5077 20383 5135 20389
rect 5077 20349 5089 20383
rect 5123 20349 5135 20383
rect 5077 20343 5135 20349
rect 5344 20383 5402 20389
rect 5344 20349 5356 20383
rect 5390 20380 5402 20383
rect 5902 20380 5908 20392
rect 5390 20352 5908 20380
rect 5390 20349 5402 20352
rect 5344 20343 5402 20349
rect 5092 20312 5120 20343
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 6730 20340 6736 20392
rect 6788 20380 6794 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6788 20352 6837 20380
rect 6788 20340 6794 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 5626 20312 5632 20324
rect 3436 20284 5632 20312
rect 5626 20272 5632 20284
rect 5684 20312 5690 20324
rect 6362 20312 6368 20324
rect 5684 20284 6368 20312
rect 5684 20272 5690 20284
rect 6362 20272 6368 20284
rect 6420 20312 6426 20324
rect 6748 20312 6776 20340
rect 6420 20284 6776 20312
rect 6932 20312 6960 20420
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 13228 20420 13277 20448
rect 13228 20408 13234 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 14936 20448 14964 20556
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 19794 20584 19800 20596
rect 19475 20556 19800 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 19794 20544 19800 20556
rect 19852 20544 19858 20596
rect 16577 20519 16635 20525
rect 16577 20485 16589 20519
rect 16623 20516 16635 20519
rect 16942 20516 16948 20528
rect 16623 20488 16948 20516
rect 16623 20485 16635 20488
rect 16577 20479 16635 20485
rect 16942 20476 16948 20488
rect 17000 20476 17006 20528
rect 19150 20476 19156 20528
rect 19208 20516 19214 20528
rect 19208 20488 20852 20516
rect 19208 20476 19214 20488
rect 13265 20411 13323 20417
rect 14844 20420 14964 20448
rect 7092 20383 7150 20389
rect 7092 20349 7104 20383
rect 7138 20380 7150 20383
rect 7374 20380 7380 20392
rect 7138 20352 7380 20380
rect 7138 20349 7150 20352
rect 7092 20343 7150 20349
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 7834 20340 7840 20392
rect 7892 20380 7898 20392
rect 8481 20383 8539 20389
rect 8481 20380 8493 20383
rect 7892 20352 8493 20380
rect 7892 20340 7898 20352
rect 8481 20349 8493 20352
rect 8527 20349 8539 20383
rect 8481 20343 8539 20349
rect 8748 20383 8806 20389
rect 8748 20349 8760 20383
rect 8794 20380 8806 20383
rect 9030 20380 9036 20392
rect 8794 20352 9036 20380
rect 8794 20349 8806 20352
rect 8748 20343 8806 20349
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 10226 20340 10232 20392
rect 10284 20380 10290 20392
rect 10410 20380 10416 20392
rect 10284 20352 10416 20380
rect 10284 20340 10290 20352
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10680 20383 10738 20389
rect 10680 20349 10692 20383
rect 10726 20380 10738 20383
rect 11974 20380 11980 20392
rect 10726 20352 11980 20380
rect 10726 20349 10738 20352
rect 10680 20343 10738 20349
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20380 12771 20383
rect 12802 20380 12808 20392
rect 12759 20352 12808 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 13532 20383 13590 20389
rect 13532 20349 13544 20383
rect 13578 20380 13590 20383
rect 14458 20380 14464 20392
rect 13578 20352 14464 20380
rect 13578 20349 13590 20352
rect 13532 20343 13590 20349
rect 14458 20340 14464 20352
rect 14516 20340 14522 20392
rect 10134 20312 10140 20324
rect 6932 20284 10140 20312
rect 6420 20272 6426 20284
rect 10134 20272 10140 20284
rect 10192 20272 10198 20324
rect 11514 20272 11520 20324
rect 11572 20312 11578 20324
rect 12434 20312 12440 20324
rect 11572 20284 12440 20312
rect 11572 20272 11578 20284
rect 12434 20272 12440 20284
rect 12492 20272 12498 20324
rect 14550 20312 14556 20324
rect 12820 20284 14556 20312
rect 842 20204 848 20256
rect 900 20244 906 20256
rect 5258 20244 5264 20256
rect 900 20216 5264 20244
rect 900 20204 906 20216
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 5442 20204 5448 20256
rect 5500 20244 5506 20256
rect 12820 20244 12848 20284
rect 14550 20272 14556 20284
rect 14608 20272 14614 20324
rect 5500 20216 12848 20244
rect 12897 20247 12955 20253
rect 5500 20204 5506 20216
rect 12897 20213 12909 20247
rect 12943 20244 12955 20247
rect 14844 20244 14872 20420
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16816 20420 17049 20448
rect 16816 20408 16822 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 17184 20420 17229 20448
rect 17184 20408 17190 20420
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 19886 20448 19892 20460
rect 19484 20420 19892 20448
rect 19484 20408 19490 20420
rect 19886 20408 19892 20420
rect 19944 20408 19950 20460
rect 20162 20448 20168 20460
rect 20123 20420 20168 20448
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20448 20407 20451
rect 20438 20448 20444 20460
rect 20395 20420 20444 20448
rect 20395 20417 20407 20420
rect 20349 20411 20407 20417
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 14918 20340 14924 20392
rect 14976 20380 14982 20392
rect 15194 20389 15200 20392
rect 15188 20380 15200 20389
rect 14976 20352 15021 20380
rect 15155 20352 15200 20380
rect 14976 20340 14982 20352
rect 15188 20343 15200 20352
rect 15194 20340 15200 20343
rect 15252 20340 15258 20392
rect 16206 20340 16212 20392
rect 16264 20380 16270 20392
rect 18046 20380 18052 20392
rect 16264 20352 17080 20380
rect 18007 20352 18052 20380
rect 16264 20340 16270 20352
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 16945 20315 17003 20321
rect 16945 20312 16957 20315
rect 15344 20284 16957 20312
rect 15344 20272 15350 20284
rect 16945 20281 16957 20284
rect 16991 20281 17003 20315
rect 17052 20312 17080 20352
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 20824 20389 20852 20488
rect 20809 20383 20867 20389
rect 18248 20352 20392 20380
rect 18248 20312 18276 20352
rect 17052 20284 18276 20312
rect 18316 20315 18374 20321
rect 16945 20275 17003 20281
rect 18316 20281 18328 20315
rect 18362 20312 18374 20315
rect 19150 20312 19156 20324
rect 18362 20284 19156 20312
rect 18362 20281 18374 20284
rect 18316 20275 18374 20281
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 19978 20312 19984 20324
rect 19260 20284 19984 20312
rect 16298 20244 16304 20256
rect 12943 20216 14872 20244
rect 16259 20216 16304 20244
rect 12943 20213 12955 20216
rect 12897 20207 12955 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 19260 20244 19288 20284
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 20073 20315 20131 20321
rect 20073 20281 20085 20315
rect 20119 20312 20131 20315
rect 20254 20312 20260 20324
rect 20119 20284 20260 20312
rect 20119 20281 20131 20284
rect 20073 20275 20131 20281
rect 20254 20272 20260 20284
rect 20312 20272 20318 20324
rect 20364 20312 20392 20352
rect 20809 20349 20821 20383
rect 20855 20380 20867 20383
rect 20898 20380 20904 20392
rect 20855 20352 20904 20380
rect 20855 20349 20867 20352
rect 20809 20343 20867 20349
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 21076 20383 21134 20389
rect 21076 20349 21088 20383
rect 21122 20380 21134 20383
rect 21542 20380 21548 20392
rect 21122 20352 21548 20380
rect 21122 20349 21134 20352
rect 21076 20343 21134 20349
rect 21542 20340 21548 20352
rect 21600 20340 21606 20392
rect 22462 20380 22468 20392
rect 22423 20352 22468 20380
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 24026 20312 24032 20324
rect 20364 20284 24032 20312
rect 24026 20272 24032 20284
rect 24084 20272 24090 20324
rect 19702 20244 19708 20256
rect 18012 20216 19288 20244
rect 19663 20216 19708 20244
rect 18012 20204 18018 20216
rect 19702 20204 19708 20216
rect 19760 20204 19766 20256
rect 21726 20204 21732 20256
rect 21784 20244 21790 20256
rect 22189 20247 22247 20253
rect 22189 20244 22201 20247
rect 21784 20216 22201 20244
rect 21784 20204 21790 20216
rect 22189 20213 22201 20216
rect 22235 20213 22247 20247
rect 22189 20207 22247 20213
rect 22649 20247 22707 20253
rect 22649 20213 22661 20247
rect 22695 20244 22707 20247
rect 22922 20244 22928 20256
rect 22695 20216 22928 20244
rect 22695 20213 22707 20216
rect 22649 20207 22707 20213
rect 22922 20204 22928 20216
rect 22980 20204 22986 20256
rect 1104 20154 23276 20176
rect 1104 20102 8379 20154
rect 8431 20102 8443 20154
rect 8495 20102 8507 20154
rect 8559 20102 8571 20154
rect 8623 20102 15776 20154
rect 15828 20102 15840 20154
rect 15892 20102 15904 20154
rect 15956 20102 15968 20154
rect 16020 20102 23276 20154
rect 1104 20080 23276 20102
rect 2130 20000 2136 20052
rect 2188 20040 2194 20052
rect 3237 20043 3295 20049
rect 3237 20040 3249 20043
rect 2188 20012 3249 20040
rect 2188 20000 2194 20012
rect 3237 20009 3249 20012
rect 3283 20009 3295 20043
rect 3237 20003 3295 20009
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 6273 20043 6331 20049
rect 6273 20040 6285 20043
rect 4212 20012 6285 20040
rect 4212 20000 4218 20012
rect 6273 20009 6285 20012
rect 6319 20009 6331 20043
rect 6273 20003 6331 20009
rect 6641 20043 6699 20049
rect 6641 20009 6653 20043
rect 6687 20040 6699 20043
rect 6914 20040 6920 20052
rect 6687 20012 6920 20040
rect 6687 20009 6699 20012
rect 6641 20003 6699 20009
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 9858 20000 9864 20052
rect 9916 20000 9922 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 11606 20040 11612 20052
rect 10192 20012 11612 20040
rect 10192 20000 10198 20012
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 11793 20043 11851 20049
rect 11793 20009 11805 20043
rect 11839 20040 11851 20043
rect 11974 20040 11980 20052
rect 11839 20012 11980 20040
rect 11839 20009 11851 20012
rect 11793 20003 11851 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 13078 20040 13084 20052
rect 12124 20012 13084 20040
rect 12124 20000 12130 20012
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13449 20043 13507 20049
rect 13449 20009 13461 20043
rect 13495 20040 13507 20043
rect 13722 20040 13728 20052
rect 13495 20012 13728 20040
rect 13495 20009 13507 20012
rect 13449 20003 13507 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 13998 20040 14004 20052
rect 13959 20012 14004 20040
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 19150 20040 19156 20052
rect 14608 20012 17356 20040
rect 19111 20012 19156 20040
rect 14608 20000 14614 20012
rect 4430 19932 4436 19984
rect 4488 19972 4494 19984
rect 4678 19975 4736 19981
rect 4678 19972 4690 19975
rect 4488 19944 4690 19972
rect 4488 19932 4494 19944
rect 4678 19941 4690 19944
rect 4724 19941 4736 19975
rect 4678 19935 4736 19941
rect 5074 19932 5080 19984
rect 5132 19972 5138 19984
rect 5132 19944 5764 19972
rect 5132 19932 5138 19944
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 1664 19907 1722 19913
rect 1664 19873 1676 19907
rect 1710 19904 1722 19907
rect 2774 19904 2780 19916
rect 1710 19876 2780 19904
rect 1710 19873 1722 19876
rect 1664 19867 1722 19873
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 3053 19907 3111 19913
rect 3053 19873 3065 19907
rect 3099 19904 3111 19907
rect 3142 19904 3148 19916
rect 3099 19876 3148 19904
rect 3099 19873 3111 19876
rect 3053 19867 3111 19873
rect 3142 19864 3148 19876
rect 3200 19904 3206 19916
rect 3602 19904 3608 19916
rect 3200 19876 3608 19904
rect 3200 19864 3206 19876
rect 3602 19864 3608 19876
rect 3660 19864 3666 19916
rect 5626 19904 5632 19916
rect 4448 19876 5632 19904
rect 4062 19796 4068 19848
rect 4120 19836 4126 19848
rect 4448 19845 4476 19876
rect 5626 19864 5632 19876
rect 5684 19864 5690 19916
rect 4433 19839 4491 19845
rect 4433 19836 4445 19839
rect 4120 19808 4445 19836
rect 4120 19796 4126 19808
rect 4433 19805 4445 19808
rect 4479 19805 4491 19839
rect 5736 19836 5764 19944
rect 5810 19932 5816 19984
rect 5868 19972 5874 19984
rect 6733 19975 6791 19981
rect 6733 19972 6745 19975
rect 5868 19944 6745 19972
rect 5868 19932 5874 19944
rect 6733 19941 6745 19944
rect 6779 19941 6791 19975
rect 6733 19935 6791 19941
rect 8196 19975 8254 19981
rect 8196 19941 8208 19975
rect 8242 19972 8254 19975
rect 8570 19972 8576 19984
rect 8242 19944 8576 19972
rect 8242 19941 8254 19944
rect 8196 19935 8254 19941
rect 8570 19932 8576 19944
rect 8628 19932 8634 19984
rect 9677 19975 9735 19981
rect 9677 19941 9689 19975
rect 9723 19972 9735 19975
rect 9876 19972 9904 20000
rect 12336 19975 12394 19981
rect 9723 19944 9904 19972
rect 10428 19944 12112 19972
rect 9723 19941 9735 19944
rect 9677 19935 9735 19941
rect 7377 19907 7435 19913
rect 7377 19873 7389 19907
rect 7423 19904 7435 19907
rect 9214 19904 9220 19916
rect 7423 19876 9220 19904
rect 7423 19873 7435 19876
rect 7377 19867 7435 19873
rect 9214 19864 9220 19876
rect 9272 19864 9278 19916
rect 9858 19904 9864 19916
rect 9819 19876 9864 19904
rect 9858 19864 9864 19876
rect 9916 19864 9922 19916
rect 6822 19836 6828 19848
rect 5736 19808 6684 19836
rect 6783 19808 6828 19836
rect 4433 19799 4491 19805
rect 3234 19728 3240 19780
rect 3292 19768 3298 19780
rect 3878 19768 3884 19780
rect 3292 19740 3884 19768
rect 3292 19728 3298 19740
rect 3878 19728 3884 19740
rect 3936 19728 3942 19780
rect 5813 19771 5871 19777
rect 5813 19737 5825 19771
rect 5859 19768 5871 19771
rect 5902 19768 5908 19780
rect 5859 19740 5908 19768
rect 5859 19737 5871 19740
rect 5813 19731 5871 19737
rect 5902 19728 5908 19740
rect 5960 19728 5966 19780
rect 6656 19768 6684 19808
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 7834 19796 7840 19848
rect 7892 19836 7898 19848
rect 7929 19839 7987 19845
rect 7929 19836 7941 19839
rect 7892 19808 7941 19836
rect 7892 19796 7898 19808
rect 7929 19805 7941 19808
rect 7975 19805 7987 19839
rect 7929 19799 7987 19805
rect 8938 19796 8944 19848
rect 8996 19836 9002 19848
rect 8996 19808 10180 19836
rect 8996 19796 9002 19808
rect 6656 19740 7972 19768
rect 2314 19660 2320 19712
rect 2372 19700 2378 19712
rect 2777 19703 2835 19709
rect 2777 19700 2789 19703
rect 2372 19672 2789 19700
rect 2372 19660 2378 19672
rect 2777 19669 2789 19672
rect 2823 19700 2835 19703
rect 5074 19700 5080 19712
rect 2823 19672 5080 19700
rect 2823 19669 2835 19672
rect 2777 19663 2835 19669
rect 5074 19660 5080 19672
rect 5132 19660 5138 19712
rect 5442 19660 5448 19712
rect 5500 19700 5506 19712
rect 7282 19700 7288 19712
rect 5500 19672 7288 19700
rect 5500 19660 5506 19672
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7558 19700 7564 19712
rect 7519 19672 7564 19700
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 7944 19700 7972 19740
rect 8202 19700 8208 19712
rect 7944 19672 8208 19700
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 9309 19703 9367 19709
rect 9309 19700 9321 19703
rect 8352 19672 9321 19700
rect 8352 19660 8358 19672
rect 9309 19669 9321 19672
rect 9355 19669 9367 19703
rect 9309 19663 9367 19669
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10045 19703 10103 19709
rect 10045 19700 10057 19703
rect 9732 19672 10057 19700
rect 9732 19660 9738 19672
rect 10045 19669 10057 19672
rect 10091 19669 10103 19703
rect 10152 19700 10180 19808
rect 10226 19796 10232 19848
rect 10284 19836 10290 19848
rect 10428 19845 10456 19944
rect 10686 19913 10692 19916
rect 10680 19904 10692 19913
rect 10647 19876 10692 19904
rect 10680 19867 10692 19876
rect 10686 19864 10692 19867
rect 10744 19864 10750 19916
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11974 19904 11980 19916
rect 11296 19876 11980 19904
rect 11296 19864 11302 19876
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12084 19913 12112 19944
rect 12336 19941 12348 19975
rect 12382 19972 12394 19975
rect 12526 19972 12532 19984
rect 12382 19944 12532 19972
rect 12382 19941 12394 19944
rect 12336 19935 12394 19941
rect 12526 19932 12532 19944
rect 12584 19972 12590 19984
rect 13909 19975 13967 19981
rect 13909 19972 13921 19975
rect 12584 19944 13921 19972
rect 12584 19932 12590 19944
rect 13909 19941 13921 19944
rect 13955 19941 13967 19975
rect 13909 19935 13967 19941
rect 15648 19975 15706 19981
rect 15648 19941 15660 19975
rect 15694 19972 15706 19975
rect 16298 19972 16304 19984
rect 15694 19944 16304 19972
rect 15694 19941 15706 19944
rect 15648 19935 15706 19941
rect 16298 19932 16304 19944
rect 16356 19972 16362 19984
rect 17221 19975 17279 19981
rect 17221 19972 17233 19975
rect 16356 19944 17233 19972
rect 16356 19932 16362 19944
rect 17221 19941 17233 19944
rect 17267 19941 17279 19975
rect 17328 19972 17356 20012
rect 19150 20000 19156 20012
rect 19208 20040 19214 20052
rect 19889 20043 19947 20049
rect 19889 20040 19901 20043
rect 19208 20012 19901 20040
rect 19208 20000 19214 20012
rect 19889 20009 19901 20012
rect 19935 20009 19947 20043
rect 19889 20003 19947 20009
rect 19426 19972 19432 19984
rect 17328 19944 19432 19972
rect 17221 19935 17279 19941
rect 19426 19932 19432 19944
rect 19484 19932 19490 19984
rect 19794 19972 19800 19984
rect 19755 19944 19800 19972
rect 19794 19932 19800 19944
rect 19852 19932 19858 19984
rect 12069 19907 12127 19913
rect 12069 19873 12081 19907
rect 12115 19873 12127 19907
rect 14553 19907 14611 19913
rect 14553 19904 14565 19907
rect 12069 19867 12127 19873
rect 12176 19876 14565 19904
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 10284 19808 10425 19836
rect 10284 19796 10290 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 12176 19836 12204 19876
rect 14553 19873 14565 19876
rect 14599 19904 14611 19907
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14599 19876 14749 19904
rect 14599 19873 14611 19876
rect 14553 19867 14611 19873
rect 14737 19873 14749 19876
rect 14783 19873 14795 19907
rect 14737 19867 14795 19873
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 15068 19876 17049 19904
rect 15068 19864 15074 19876
rect 17037 19873 17049 19876
rect 17083 19873 17095 19907
rect 17037 19867 17095 19873
rect 18040 19907 18098 19913
rect 18040 19873 18052 19907
rect 18086 19904 18098 19907
rect 19334 19904 19340 19916
rect 18086 19876 19340 19904
rect 18086 19873 18098 19876
rect 18040 19867 18098 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 21358 19904 21364 19916
rect 19444 19876 21364 19904
rect 14182 19836 14188 19848
rect 10413 19799 10471 19805
rect 11440 19808 12204 19836
rect 14095 19808 14188 19836
rect 11440 19700 11468 19808
rect 14182 19796 14188 19808
rect 14240 19836 14246 19848
rect 14826 19836 14832 19848
rect 14240 19808 14832 19836
rect 14240 19796 14246 19808
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 14918 19796 14924 19848
rect 14976 19836 14982 19848
rect 15378 19836 15384 19848
rect 14976 19808 15384 19836
rect 14976 19796 14982 19808
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 17552 19808 17785 19836
rect 17552 19796 17558 19808
rect 17773 19805 17785 19808
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 18782 19796 18788 19848
rect 18840 19836 18846 19848
rect 19444 19836 19472 19876
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 21634 19904 21640 19916
rect 21595 19876 21640 19904
rect 21634 19864 21640 19876
rect 21692 19864 21698 19916
rect 22002 19864 22008 19916
rect 22060 19904 22066 19916
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 22060 19876 22293 19904
rect 22060 19864 22066 19876
rect 22281 19873 22293 19876
rect 22327 19873 22339 19907
rect 22281 19867 22339 19873
rect 22465 19907 22523 19913
rect 22465 19873 22477 19907
rect 22511 19904 22523 19907
rect 22646 19904 22652 19916
rect 22511 19876 22652 19904
rect 22511 19873 22523 19876
rect 22465 19867 22523 19873
rect 22646 19864 22652 19876
rect 22704 19864 22710 19916
rect 18840 19808 19472 19836
rect 18840 19796 18846 19808
rect 19886 19796 19892 19848
rect 19944 19836 19950 19848
rect 20073 19839 20131 19845
rect 20073 19836 20085 19839
rect 19944 19808 20085 19836
rect 19944 19796 19950 19808
rect 20073 19805 20085 19808
rect 20119 19836 20131 19839
rect 20438 19836 20444 19848
rect 20119 19808 20444 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 20438 19796 20444 19808
rect 20496 19836 20502 19848
rect 21450 19836 21456 19848
rect 20496 19808 21456 19836
rect 20496 19796 20502 19808
rect 21450 19796 21456 19808
rect 21508 19836 21514 19848
rect 21726 19836 21732 19848
rect 21508 19808 21588 19836
rect 21687 19808 21732 19836
rect 21508 19796 21514 19808
rect 13004 19740 13768 19768
rect 10152 19672 11468 19700
rect 10045 19663 10103 19669
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 12434 19700 12440 19712
rect 11664 19672 12440 19700
rect 11664 19660 11670 19672
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 13004 19700 13032 19740
rect 12768 19672 13032 19700
rect 12768 19660 12774 19672
rect 13078 19660 13084 19712
rect 13136 19700 13142 19712
rect 13541 19703 13599 19709
rect 13541 19700 13553 19703
rect 13136 19672 13553 19700
rect 13136 19660 13142 19672
rect 13541 19669 13553 19672
rect 13587 19669 13599 19703
rect 13740 19700 13768 19740
rect 16482 19728 16488 19780
rect 16540 19768 16546 19780
rect 16761 19771 16819 19777
rect 16761 19768 16773 19771
rect 16540 19740 16773 19768
rect 16540 19728 16546 19740
rect 16761 19737 16773 19740
rect 16807 19737 16819 19771
rect 20806 19768 20812 19780
rect 16761 19731 16819 19737
rect 16868 19740 17540 19768
rect 16868 19700 16896 19740
rect 17402 19700 17408 19712
rect 13740 19672 16896 19700
rect 17363 19672 17408 19700
rect 13541 19663 13599 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 17512 19700 17540 19740
rect 18708 19740 20812 19768
rect 18708 19700 18736 19740
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 21174 19728 21180 19780
rect 21232 19768 21238 19780
rect 21269 19771 21327 19777
rect 21269 19768 21281 19771
rect 21232 19740 21281 19768
rect 21232 19728 21238 19740
rect 21269 19737 21281 19740
rect 21315 19737 21327 19771
rect 21560 19768 21588 19808
rect 21726 19796 21732 19808
rect 21784 19796 21790 19848
rect 21821 19839 21879 19845
rect 21821 19805 21833 19839
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 21836 19768 21864 19799
rect 21560 19740 21864 19768
rect 21269 19731 21327 19737
rect 17512 19672 18736 19700
rect 19429 19703 19487 19709
rect 19429 19669 19441 19703
rect 19475 19700 19487 19703
rect 19886 19700 19892 19712
rect 19475 19672 19892 19700
rect 19475 19669 19487 19672
rect 19429 19663 19487 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 21358 19660 21364 19712
rect 21416 19700 21422 19712
rect 22649 19703 22707 19709
rect 22649 19700 22661 19703
rect 21416 19672 22661 19700
rect 21416 19660 21422 19672
rect 22649 19669 22661 19672
rect 22695 19669 22707 19703
rect 22649 19663 22707 19669
rect 1104 19610 23276 19632
rect 1104 19558 4680 19610
rect 4732 19558 4744 19610
rect 4796 19558 4808 19610
rect 4860 19558 4872 19610
rect 4924 19558 12078 19610
rect 12130 19558 12142 19610
rect 12194 19558 12206 19610
rect 12258 19558 12270 19610
rect 12322 19558 19475 19610
rect 19527 19558 19539 19610
rect 19591 19558 19603 19610
rect 19655 19558 19667 19610
rect 19719 19558 23276 19610
rect 1104 19536 23276 19558
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 4433 19499 4491 19505
rect 2832 19468 4108 19496
rect 2832 19456 2838 19468
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 2406 19292 2412 19304
rect 1443 19264 2412 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 2406 19252 2412 19264
rect 2464 19292 2470 19304
rect 3050 19292 3056 19304
rect 2464 19264 3056 19292
rect 2464 19252 2470 19264
rect 3050 19252 3056 19264
rect 3108 19252 3114 19304
rect 3326 19301 3332 19304
rect 3320 19255 3332 19301
rect 3384 19292 3390 19304
rect 3384 19264 3420 19292
rect 3326 19252 3332 19255
rect 3384 19252 3390 19264
rect 1664 19227 1722 19233
rect 1664 19193 1676 19227
rect 1710 19224 1722 19227
rect 2222 19224 2228 19236
rect 1710 19196 2228 19224
rect 1710 19193 1722 19196
rect 1664 19187 1722 19193
rect 2222 19184 2228 19196
rect 2280 19184 2286 19236
rect 4080 19224 4108 19468
rect 4433 19465 4445 19499
rect 4479 19496 4491 19499
rect 4522 19496 4528 19508
rect 4479 19468 4528 19496
rect 4479 19465 4491 19468
rect 4433 19459 4491 19465
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 6638 19496 6644 19508
rect 4632 19468 6644 19496
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 4396 19332 4476 19360
rect 4396 19320 4402 19332
rect 4448 19304 4476 19332
rect 4522 19320 4528 19372
rect 4580 19360 4586 19372
rect 4632 19360 4660 19468
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 7834 19456 7840 19508
rect 7892 19496 7898 19508
rect 8389 19499 8447 19505
rect 8389 19496 8401 19499
rect 7892 19468 8401 19496
rect 7892 19456 7898 19468
rect 8389 19465 8401 19468
rect 8435 19465 8447 19499
rect 8389 19459 8447 19465
rect 8846 19456 8852 19508
rect 8904 19496 8910 19508
rect 8904 19468 10364 19496
rect 8904 19456 8910 19468
rect 4982 19388 4988 19440
rect 5040 19428 5046 19440
rect 6546 19428 6552 19440
rect 5040 19400 6552 19428
rect 5040 19388 5046 19400
rect 6546 19388 6552 19400
rect 6604 19388 6610 19440
rect 7561 19431 7619 19437
rect 7561 19397 7573 19431
rect 7607 19428 7619 19431
rect 7607 19400 8616 19428
rect 7607 19397 7619 19400
rect 7561 19391 7619 19397
rect 4580 19332 4660 19360
rect 5353 19363 5411 19369
rect 4580 19320 4586 19332
rect 5353 19329 5365 19363
rect 5399 19360 5411 19363
rect 5534 19360 5540 19372
rect 5399 19332 5540 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 5534 19320 5540 19332
rect 5592 19360 5598 19372
rect 6273 19363 6331 19369
rect 6273 19360 6285 19363
rect 5592 19332 6285 19360
rect 5592 19320 5598 19332
rect 6273 19329 6285 19332
rect 6319 19360 6331 19363
rect 6454 19360 6460 19372
rect 6319 19332 6460 19360
rect 6319 19329 6331 19332
rect 6273 19323 6331 19329
rect 6454 19320 6460 19332
rect 6512 19360 6518 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 6512 19332 8125 19360
rect 6512 19320 6518 19332
rect 8113 19329 8125 19332
rect 8159 19329 8171 19363
rect 8588 19360 8616 19400
rect 10336 19360 10364 19468
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 12526 19496 12532 19508
rect 10468 19468 12532 19496
rect 10468 19456 10474 19468
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 14182 19496 14188 19508
rect 12636 19468 14188 19496
rect 10502 19388 10508 19440
rect 10560 19428 10566 19440
rect 11146 19428 11152 19440
rect 10560 19400 11152 19428
rect 10560 19388 10566 19400
rect 11146 19388 11152 19400
rect 11204 19388 11210 19440
rect 10873 19363 10931 19369
rect 10873 19360 10885 19363
rect 8588 19332 8708 19360
rect 10336 19332 10885 19360
rect 8113 19323 8171 19329
rect 4430 19252 4436 19304
rect 4488 19252 4494 19304
rect 5074 19292 5080 19304
rect 5035 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 7009 19295 7067 19301
rect 7009 19261 7021 19295
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 7929 19295 7987 19301
rect 7929 19261 7941 19295
rect 7975 19292 7987 19295
rect 8294 19292 8300 19304
rect 7975 19264 8300 19292
rect 7975 19261 7987 19264
rect 7929 19255 7987 19261
rect 5169 19227 5227 19233
rect 5169 19224 5181 19227
rect 4080 19196 5181 19224
rect 5169 19193 5181 19196
rect 5215 19193 5227 19227
rect 5169 19187 5227 19193
rect 5258 19184 5264 19236
rect 5316 19224 5322 19236
rect 6089 19227 6147 19233
rect 6089 19224 6101 19227
rect 5316 19196 6101 19224
rect 5316 19184 5322 19196
rect 6089 19193 6101 19196
rect 6135 19193 6147 19227
rect 7024 19224 7052 19255
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 8435 19264 8585 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 8573 19261 8585 19264
rect 8619 19261 8631 19295
rect 8680 19292 8708 19332
rect 10873 19329 10885 19332
rect 10919 19360 10931 19363
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 10919 19332 11897 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11885 19329 11897 19332
rect 11931 19360 11943 19363
rect 12636 19360 12664 19468
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19496 14335 19499
rect 15286 19496 15292 19508
rect 14323 19468 15292 19496
rect 14323 19465 14335 19468
rect 14277 19459 14335 19465
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 15396 19468 19012 19496
rect 12820 19400 13860 19428
rect 12820 19360 12848 19400
rect 11931 19332 12664 19360
rect 12728 19332 12848 19360
rect 13081 19363 13139 19369
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 10042 19292 10048 19304
rect 8680 19264 10048 19292
rect 8573 19255 8631 19261
rect 8478 19224 8484 19236
rect 7024 19196 8484 19224
rect 6089 19187 6147 19193
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 8588 19224 8616 19255
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 12728 19292 12756 19332
rect 13081 19329 13093 19363
rect 13127 19360 13139 19363
rect 13630 19360 13636 19372
rect 13127 19332 13636 19360
rect 13127 19329 13139 19332
rect 13081 19323 13139 19329
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 10336 19264 12756 19292
rect 12805 19295 12863 19301
rect 8662 19224 8668 19236
rect 8588 19196 8668 19224
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 8754 19184 8760 19236
rect 8812 19233 8818 19236
rect 8812 19227 8876 19233
rect 8812 19193 8830 19227
rect 8864 19193 8876 19227
rect 8812 19187 8876 19193
rect 8812 19184 8818 19187
rect 4706 19156 4712 19168
rect 4667 19128 4712 19156
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 5718 19156 5724 19168
rect 5679 19128 5724 19156
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 6181 19159 6239 19165
rect 6181 19156 6193 19159
rect 5868 19128 6193 19156
rect 5868 19116 5874 19128
rect 6181 19125 6193 19128
rect 6227 19125 6239 19159
rect 6181 19119 6239 19125
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 6880 19128 7205 19156
rect 6880 19116 6886 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7193 19119 7251 19125
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19156 8079 19159
rect 8110 19156 8116 19168
rect 8067 19128 8116 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 8110 19116 8116 19128
rect 8168 19156 8174 19168
rect 10336 19165 10364 19264
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 12986 19292 12992 19304
rect 12851 19264 12992 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13722 19292 13728 19304
rect 13683 19264 13728 19292
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 13832 19292 13860 19400
rect 14918 19388 14924 19440
rect 14976 19428 14982 19440
rect 15105 19431 15163 19437
rect 15105 19428 15117 19431
rect 14976 19400 15117 19428
rect 14976 19388 14982 19400
rect 15105 19397 15117 19400
rect 15151 19397 15163 19431
rect 15105 19391 15163 19397
rect 14642 19320 14648 19372
rect 14700 19360 14706 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14700 19332 14749 19360
rect 14700 19320 14706 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 14884 19332 14929 19360
rect 14884 19320 14890 19332
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 15396 19360 15424 19468
rect 17126 19428 17132 19440
rect 15764 19400 17132 19428
rect 15764 19372 15792 19400
rect 17126 19388 17132 19400
rect 17184 19388 17190 19440
rect 18984 19428 19012 19468
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 19429 19499 19487 19505
rect 19429 19496 19441 19499
rect 19392 19468 19441 19496
rect 19392 19456 19398 19468
rect 19429 19465 19441 19468
rect 19475 19465 19487 19499
rect 19429 19459 19487 19465
rect 20254 19456 20260 19508
rect 20312 19496 20318 19508
rect 20622 19496 20628 19508
rect 20312 19468 20628 19496
rect 20312 19456 20318 19468
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 20070 19428 20076 19440
rect 18984 19400 20076 19428
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 15746 19360 15752 19372
rect 15068 19332 15424 19360
rect 15659 19332 15752 19360
rect 15068 19320 15074 19332
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16172 19332 16865 19360
rect 16172 19320 16178 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 19794 19320 19800 19372
rect 19852 19360 19858 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 19852 19332 20269 19360
rect 19852 19320 19858 19332
rect 20257 19329 20269 19332
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 15473 19295 15531 19301
rect 15473 19292 15485 19295
rect 13832 19264 15485 19292
rect 15473 19261 15485 19264
rect 15519 19261 15531 19295
rect 15473 19255 15531 19261
rect 17034 19252 17040 19304
rect 17092 19292 17098 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 17092 19264 17417 19292
rect 17092 19252 17098 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 18046 19292 18052 19304
rect 17552 19264 18052 19292
rect 17552 19252 17558 19264
rect 18046 19252 18052 19264
rect 18104 19292 18110 19304
rect 19058 19292 19064 19304
rect 18104 19264 19064 19292
rect 18104 19252 18110 19264
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20956 19264 21005 19292
rect 20956 19252 20962 19264
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21260 19295 21318 19301
rect 21260 19261 21272 19295
rect 21306 19292 21318 19295
rect 21726 19292 21732 19304
rect 21306 19264 21732 19292
rect 21306 19261 21318 19264
rect 21260 19255 21318 19261
rect 12894 19224 12900 19236
rect 11348 19196 12756 19224
rect 12855 19196 12900 19224
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 8168 19128 9965 19156
rect 8168 19116 8174 19128
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 9953 19119 10011 19125
rect 10321 19159 10379 19165
rect 10321 19125 10333 19159
rect 10367 19125 10379 19159
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10321 19119 10379 19125
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 11348 19165 11376 19196
rect 11333 19159 11391 19165
rect 10836 19128 10881 19156
rect 10836 19116 10842 19128
rect 11333 19125 11345 19159
rect 11379 19125 11391 19159
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 11333 19119 11391 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11793 19159 11851 19165
rect 11793 19125 11805 19159
rect 11839 19156 11851 19159
rect 12342 19156 12348 19168
rect 11839 19128 12348 19156
rect 11839 19125 11851 19128
rect 11793 19119 11851 19125
rect 12342 19116 12348 19128
rect 12400 19116 12406 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12728 19156 12756 19196
rect 12894 19184 12900 19196
rect 12952 19184 12958 19236
rect 15565 19227 15623 19233
rect 15565 19224 15577 19227
rect 13004 19196 15577 19224
rect 13004 19156 13032 19196
rect 15565 19193 15577 19196
rect 15611 19193 15623 19227
rect 16761 19227 16819 19233
rect 16761 19224 16773 19227
rect 15565 19187 15623 19193
rect 16132 19196 16773 19224
rect 12492 19128 12537 19156
rect 12728 19128 13032 19156
rect 13909 19159 13967 19165
rect 12492 19116 12498 19128
rect 13909 19125 13921 19159
rect 13955 19156 13967 19159
rect 14458 19156 14464 19168
rect 13955 19128 14464 19156
rect 13955 19125 13967 19128
rect 13909 19119 13967 19125
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 14645 19159 14703 19165
rect 14645 19125 14657 19159
rect 14691 19156 14703 19159
rect 15010 19156 15016 19168
rect 14691 19128 15016 19156
rect 14691 19125 14703 19128
rect 14645 19119 14703 19125
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 16132 19165 16160 19196
rect 16761 19193 16773 19196
rect 16807 19193 16819 19227
rect 16761 19187 16819 19193
rect 18316 19227 18374 19233
rect 18316 19193 18328 19227
rect 18362 19224 18374 19227
rect 18782 19224 18788 19236
rect 18362 19196 18788 19224
rect 18362 19193 18374 19196
rect 18316 19187 18374 19193
rect 18782 19184 18788 19196
rect 18840 19184 18846 19236
rect 20073 19227 20131 19233
rect 20073 19224 20085 19227
rect 18892 19196 20085 19224
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 15344 19128 16129 19156
rect 15344 19116 15350 19128
rect 16117 19125 16129 19128
rect 16163 19125 16175 19159
rect 16298 19156 16304 19168
rect 16259 19128 16304 19156
rect 16117 19119 16175 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16666 19156 16672 19168
rect 16627 19128 16672 19156
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 17589 19159 17647 19165
rect 17589 19125 17601 19159
rect 17635 19156 17647 19159
rect 17678 19156 17684 19168
rect 17635 19128 17684 19156
rect 17635 19125 17647 19128
rect 17589 19119 17647 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 17862 19116 17868 19168
rect 17920 19156 17926 19168
rect 18892 19156 18920 19196
rect 20073 19193 20085 19196
rect 20119 19193 20131 19227
rect 20073 19187 20131 19193
rect 20162 19184 20168 19236
rect 20220 19224 20226 19236
rect 20220 19196 20265 19224
rect 20220 19184 20226 19196
rect 17920 19128 18920 19156
rect 17920 19116 17926 19128
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 19705 19159 19763 19165
rect 19705 19156 19717 19159
rect 19208 19128 19717 19156
rect 19208 19116 19214 19128
rect 19705 19125 19717 19128
rect 19751 19125 19763 19159
rect 21008 19156 21036 19255
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 21266 19156 21272 19168
rect 21008 19128 21272 19156
rect 19705 19119 19763 19125
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21634 19116 21640 19168
rect 21692 19156 21698 19168
rect 22373 19159 22431 19165
rect 22373 19156 22385 19159
rect 21692 19128 22385 19156
rect 21692 19116 21698 19128
rect 22373 19125 22385 19128
rect 22419 19125 22431 19159
rect 22373 19119 22431 19125
rect 1104 19066 23276 19088
rect 1104 19014 8379 19066
rect 8431 19014 8443 19066
rect 8495 19014 8507 19066
rect 8559 19014 8571 19066
rect 8623 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 15904 19066
rect 15956 19014 15968 19066
rect 16020 19014 23276 19066
rect 1104 18992 23276 19014
rect 3697 18955 3755 18961
rect 3697 18921 3709 18955
rect 3743 18952 3755 18955
rect 4433 18955 4491 18961
rect 3743 18924 4200 18952
rect 3743 18921 3755 18924
rect 3697 18915 3755 18921
rect 2222 18844 2228 18896
rect 2280 18884 2286 18896
rect 3712 18884 3740 18915
rect 2280 18856 3740 18884
rect 2280 18844 2286 18856
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2317 18819 2375 18825
rect 2317 18785 2329 18819
rect 2363 18816 2375 18819
rect 2406 18816 2412 18828
rect 2363 18788 2412 18816
rect 2363 18785 2375 18788
rect 2317 18779 2375 18785
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 2584 18819 2642 18825
rect 2584 18785 2596 18819
rect 2630 18816 2642 18819
rect 3694 18816 3700 18828
rect 2630 18788 3700 18816
rect 2630 18785 2642 18788
rect 2584 18779 2642 18785
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 4172 18816 4200 18924
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 4706 18952 4712 18964
rect 4479 18924 4712 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 4893 18955 4951 18961
rect 4893 18921 4905 18955
rect 4939 18952 4951 18955
rect 6638 18952 6644 18964
rect 4939 18924 6644 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 6733 18955 6791 18961
rect 6733 18921 6745 18955
rect 6779 18952 6791 18955
rect 7926 18952 7932 18964
rect 6779 18924 7932 18952
rect 6779 18921 6791 18924
rect 6733 18915 6791 18921
rect 7926 18912 7932 18924
rect 7984 18912 7990 18964
rect 8846 18952 8852 18964
rect 8036 18924 8852 18952
rect 4525 18887 4583 18893
rect 4525 18853 4537 18887
rect 4571 18884 4583 18887
rect 5718 18884 5724 18896
rect 4571 18856 5724 18884
rect 4571 18853 4583 18856
rect 4525 18847 4583 18853
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 7285 18887 7343 18893
rect 7285 18884 7297 18887
rect 5828 18856 7297 18884
rect 5258 18816 5264 18828
rect 4172 18788 5264 18816
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5442 18816 5448 18828
rect 5403 18788 5448 18816
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 5828 18816 5856 18856
rect 7285 18853 7297 18856
rect 7331 18853 7343 18887
rect 7285 18847 7343 18853
rect 7374 18844 7380 18896
rect 7432 18884 7438 18896
rect 8036 18884 8064 18924
rect 8846 18912 8852 18924
rect 8904 18912 8910 18964
rect 9309 18955 9367 18961
rect 9309 18921 9321 18955
rect 9355 18952 9367 18955
rect 9858 18952 9864 18964
rect 9355 18924 9864 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 10744 18924 11621 18952
rect 10744 18912 10750 18924
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 17862 18952 17868 18964
rect 11609 18915 11667 18921
rect 11716 18924 17868 18952
rect 8202 18893 8208 18896
rect 8196 18884 8208 18893
rect 7432 18856 8064 18884
rect 8163 18856 8208 18884
rect 7432 18844 7438 18856
rect 8196 18847 8208 18856
rect 8202 18844 8208 18847
rect 8260 18844 8266 18896
rect 8294 18844 8300 18896
rect 8352 18884 8358 18896
rect 11716 18884 11744 18924
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 18782 18952 18788 18964
rect 18743 18924 18788 18952
rect 18782 18912 18788 18924
rect 18840 18952 18846 18964
rect 19521 18955 19579 18961
rect 19521 18952 19533 18955
rect 18840 18924 19533 18952
rect 18840 18912 18846 18924
rect 19521 18921 19533 18924
rect 19567 18921 19579 18955
rect 19521 18915 19579 18921
rect 8352 18856 11744 18884
rect 8352 18844 8358 18856
rect 11974 18844 11980 18896
rect 12032 18884 12038 18896
rect 12130 18887 12188 18893
rect 12130 18884 12142 18887
rect 12032 18856 12142 18884
rect 12032 18844 12038 18856
rect 12130 18853 12142 18856
rect 12176 18884 12188 18887
rect 14001 18887 14059 18893
rect 14001 18884 14013 18887
rect 12176 18856 14013 18884
rect 12176 18853 12188 18856
rect 12130 18847 12188 18853
rect 14001 18853 14013 18856
rect 14047 18853 14059 18887
rect 21536 18887 21594 18893
rect 14001 18847 14059 18853
rect 14108 18856 20208 18884
rect 5644 18788 5856 18816
rect 6273 18819 6331 18825
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4893 18751 4951 18757
rect 4893 18748 4905 18751
rect 4755 18720 4905 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4893 18717 4905 18720
rect 4939 18717 4951 18751
rect 4893 18711 4951 18717
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 5537 18751 5595 18757
rect 5537 18748 5549 18751
rect 5040 18720 5549 18748
rect 5040 18708 5046 18720
rect 5537 18717 5549 18720
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 1949 18683 2007 18689
rect 1949 18649 1961 18683
rect 1995 18680 2007 18683
rect 2222 18680 2228 18692
rect 1995 18652 2228 18680
rect 1995 18649 2007 18652
rect 1949 18643 2007 18649
rect 2222 18640 2228 18652
rect 2280 18640 2286 18692
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 3252 18652 4077 18680
rect 1762 18572 1768 18624
rect 1820 18612 1826 18624
rect 3252 18612 3280 18652
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4065 18643 4123 18649
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 5644 18680 5672 18788
rect 6273 18785 6285 18819
rect 6319 18816 6331 18819
rect 6733 18819 6791 18825
rect 6733 18816 6745 18819
rect 6319 18788 6745 18816
rect 6319 18785 6331 18788
rect 6273 18779 6331 18785
rect 6733 18785 6745 18788
rect 6779 18785 6791 18819
rect 6733 18779 6791 18785
rect 7193 18819 7251 18825
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 9490 18816 9496 18828
rect 7239 18788 9496 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 9490 18776 9496 18788
rect 9548 18776 9554 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10496 18819 10554 18825
rect 10496 18785 10508 18819
rect 10542 18816 10554 18819
rect 10778 18816 10784 18828
rect 10542 18788 10784 18816
rect 10542 18785 10554 18788
rect 10496 18779 10554 18785
rect 10778 18776 10784 18788
rect 10836 18816 10842 18828
rect 11606 18816 11612 18828
rect 10836 18788 11612 18816
rect 10836 18776 10842 18788
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 12526 18776 12532 18828
rect 12584 18816 12590 18828
rect 12584 18788 12940 18816
rect 12584 18776 12590 18788
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 7558 18748 7564 18760
rect 7515 18720 7564 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 4396 18652 5672 18680
rect 5736 18680 5764 18711
rect 7484 18680 7512 18711
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18717 7987 18751
rect 10226 18748 10232 18760
rect 7929 18711 7987 18717
rect 9600 18720 10232 18748
rect 5736 18652 7512 18680
rect 4396 18640 4402 18652
rect 5074 18612 5080 18624
rect 1820 18584 3280 18612
rect 5035 18584 5080 18612
rect 1820 18572 1826 18584
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 6454 18612 6460 18624
rect 6415 18584 6460 18612
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 6825 18615 6883 18621
rect 6825 18612 6837 18615
rect 6788 18584 6837 18612
rect 6788 18572 6794 18584
rect 6825 18581 6837 18584
rect 6871 18581 6883 18615
rect 7944 18612 7972 18711
rect 9600 18624 9628 18720
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11256 18720 11897 18748
rect 8202 18612 8208 18624
rect 7944 18584 8208 18612
rect 6825 18575 6883 18581
rect 8202 18572 8208 18584
rect 8260 18612 8266 18624
rect 8662 18612 8668 18624
rect 8260 18584 8668 18612
rect 8260 18572 8266 18584
rect 8662 18572 8668 18584
rect 8720 18612 8726 18624
rect 9582 18612 9588 18624
rect 8720 18584 9588 18612
rect 8720 18572 8726 18584
rect 9582 18572 9588 18584
rect 9640 18572 9646 18624
rect 9861 18615 9919 18621
rect 9861 18581 9873 18615
rect 9907 18612 9919 18615
rect 10134 18612 10140 18624
rect 9907 18584 10140 18612
rect 9907 18581 9919 18584
rect 9861 18575 9919 18581
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 10244 18612 10272 18708
rect 11256 18612 11284 18720
rect 11885 18717 11897 18720
rect 11931 18717 11943 18751
rect 12912 18748 12940 18788
rect 13262 18776 13268 18828
rect 13320 18816 13326 18828
rect 13909 18819 13967 18825
rect 13909 18816 13921 18819
rect 13320 18788 13921 18816
rect 13320 18776 13326 18788
rect 13909 18785 13921 18788
rect 13955 18785 13967 18819
rect 14108 18816 14136 18856
rect 13909 18779 13967 18785
rect 14016 18788 14136 18816
rect 14016 18748 14044 18788
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 14645 18819 14703 18825
rect 14645 18816 14657 18819
rect 14240 18788 14657 18816
rect 14240 18776 14246 18788
rect 14645 18785 14657 18788
rect 14691 18785 14703 18819
rect 15378 18816 15384 18828
rect 15339 18788 15384 18816
rect 14645 18779 14703 18785
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 15648 18819 15706 18825
rect 15648 18785 15660 18819
rect 15694 18816 15706 18819
rect 16482 18816 16488 18828
rect 15694 18788 16488 18816
rect 15694 18785 15706 18788
rect 15648 18779 15706 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18816 17463 18819
rect 17494 18816 17500 18828
rect 17451 18788 17500 18816
rect 17451 18785 17463 18788
rect 17405 18779 17463 18785
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 17672 18819 17730 18825
rect 17672 18785 17684 18819
rect 17718 18816 17730 18819
rect 19429 18819 19487 18825
rect 17718 18788 19288 18816
rect 17718 18785 17730 18788
rect 17672 18779 17730 18785
rect 12912 18720 14044 18748
rect 14093 18751 14151 18757
rect 11885 18711 11943 18717
rect 14093 18717 14105 18751
rect 14139 18748 14151 18751
rect 14826 18748 14832 18760
rect 14139 18720 14832 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 14826 18708 14832 18720
rect 14884 18708 14890 18760
rect 19260 18748 19288 18788
rect 19429 18785 19441 18819
rect 19475 18816 19487 18819
rect 19518 18816 19524 18828
rect 19475 18788 19524 18816
rect 19475 18785 19487 18788
rect 19429 18779 19487 18785
rect 19518 18776 19524 18788
rect 19576 18776 19582 18828
rect 20073 18819 20131 18825
rect 20073 18785 20085 18819
rect 20119 18785 20131 18819
rect 20180 18816 20208 18856
rect 21536 18853 21548 18887
rect 21582 18884 21594 18887
rect 21634 18884 21640 18896
rect 21582 18856 21640 18884
rect 21582 18853 21594 18856
rect 21536 18847 21594 18853
rect 21634 18844 21640 18856
rect 21692 18844 21698 18896
rect 22738 18816 22744 18828
rect 20180 18788 22744 18816
rect 20073 18779 20131 18785
rect 19334 18748 19340 18760
rect 19260 18720 19340 18748
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18748 19763 18751
rect 19886 18748 19892 18760
rect 19751 18720 19892 18748
rect 19751 18717 19763 18720
rect 19705 18711 19763 18717
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 18690 18640 18696 18692
rect 18748 18680 18754 18692
rect 20088 18680 20116 18779
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 21266 18748 21272 18760
rect 21227 18720 21272 18748
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 18748 18652 20116 18680
rect 18748 18640 18754 18652
rect 13262 18612 13268 18624
rect 10244 18584 11284 18612
rect 13223 18584 13268 18612
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 13538 18612 13544 18624
rect 13499 18584 13544 18612
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 14829 18615 14887 18621
rect 14829 18612 14841 18615
rect 14792 18584 14841 18612
rect 14792 18572 14798 18584
rect 14829 18581 14841 18584
rect 14875 18581 14887 18615
rect 16758 18612 16764 18624
rect 16719 18584 16764 18612
rect 14829 18575 14887 18581
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 19061 18615 19119 18621
rect 19061 18612 19073 18615
rect 18656 18584 19073 18612
rect 18656 18572 18662 18584
rect 19061 18581 19073 18584
rect 19107 18581 19119 18615
rect 20254 18612 20260 18624
rect 20215 18584 20260 18612
rect 19061 18575 19119 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 22646 18612 22652 18624
rect 22607 18584 22652 18612
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 1104 18522 23276 18544
rect 1104 18470 4680 18522
rect 4732 18470 4744 18522
rect 4796 18470 4808 18522
rect 4860 18470 4872 18522
rect 4924 18470 12078 18522
rect 12130 18470 12142 18522
rect 12194 18470 12206 18522
rect 12258 18470 12270 18522
rect 12322 18470 19475 18522
rect 19527 18470 19539 18522
rect 19591 18470 19603 18522
rect 19655 18470 19667 18522
rect 19719 18470 23276 18522
rect 1104 18448 23276 18470
rect 1949 18411 2007 18417
rect 1949 18377 1961 18411
rect 1995 18408 2007 18411
rect 4982 18408 4988 18420
rect 1995 18380 4988 18408
rect 1995 18377 2007 18380
rect 1949 18371 2007 18377
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 8938 18408 8944 18420
rect 8251 18380 8944 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 9640 18380 9965 18408
rect 9640 18368 9646 18380
rect 9953 18377 9965 18380
rect 9999 18377 10011 18411
rect 11606 18408 11612 18420
rect 11567 18380 11612 18408
rect 9953 18371 10011 18377
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 12434 18368 12440 18420
rect 12492 18408 12498 18420
rect 14369 18411 14427 18417
rect 14369 18408 14381 18411
rect 12492 18380 14381 18408
rect 12492 18368 12498 18380
rect 14369 18377 14381 18380
rect 14415 18377 14427 18411
rect 14369 18371 14427 18377
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 19242 18408 19248 18420
rect 14516 18380 19248 18408
rect 14516 18368 14522 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19429 18411 19487 18417
rect 19429 18408 19441 18411
rect 19392 18380 19441 18408
rect 19392 18368 19398 18380
rect 19429 18377 19441 18380
rect 19475 18377 19487 18411
rect 22002 18408 22008 18420
rect 19429 18371 19487 18377
rect 19536 18380 22008 18408
rect 4062 18300 4068 18352
rect 4120 18300 4126 18352
rect 4249 18343 4307 18349
rect 4249 18309 4261 18343
rect 4295 18340 4307 18343
rect 4338 18340 4344 18352
rect 4295 18312 4344 18340
rect 4295 18309 4307 18312
rect 4249 18303 4307 18309
rect 4338 18300 4344 18312
rect 4396 18300 4402 18352
rect 8294 18340 8300 18352
rect 6840 18312 8300 18340
rect 2314 18272 2320 18284
rect 2275 18244 2320 18272
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 4080 18272 4108 18300
rect 6840 18281 6868 18312
rect 8294 18300 8300 18312
rect 8352 18300 8358 18352
rect 9306 18300 9312 18352
rect 9364 18340 9370 18352
rect 9677 18343 9735 18349
rect 9677 18340 9689 18343
rect 9364 18312 9689 18340
rect 9364 18300 9370 18312
rect 9677 18309 9689 18312
rect 9723 18309 9735 18343
rect 9677 18303 9735 18309
rect 12621 18343 12679 18349
rect 12621 18309 12633 18343
rect 12667 18340 12679 18343
rect 12986 18340 12992 18352
rect 12667 18312 12992 18340
rect 12667 18309 12679 18312
rect 12621 18303 12679 18309
rect 12986 18300 12992 18312
rect 13044 18300 13050 18352
rect 14734 18300 14740 18352
rect 14792 18340 14798 18352
rect 17954 18340 17960 18352
rect 14792 18312 17960 18340
rect 14792 18300 14798 18312
rect 17954 18300 17960 18312
rect 18012 18300 18018 18352
rect 4617 18275 4675 18281
rect 4617 18272 4629 18275
rect 4080 18244 4629 18272
rect 4617 18241 4629 18244
rect 4663 18241 4675 18275
rect 4617 18235 4675 18241
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 7929 18275 7987 18281
rect 7929 18241 7941 18275
rect 7975 18272 7987 18275
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 7975 18244 8217 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 8205 18235 8263 18241
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18272 11943 18275
rect 12894 18272 12900 18284
rect 11931 18244 12900 18272
rect 11931 18241 11943 18244
rect 11885 18235 11943 18241
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 14826 18232 14832 18284
rect 14884 18272 14890 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 14884 18244 15209 18272
rect 14884 18232 14890 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 16206 18272 16212 18284
rect 16167 18244 16212 18272
rect 15197 18235 15255 18241
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 17494 18272 17500 18284
rect 17359 18244 17500 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 18046 18272 18052 18284
rect 18007 18244 18052 18272
rect 18046 18232 18052 18244
rect 18104 18232 18110 18284
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 19426 18272 19432 18284
rect 19208 18244 19432 18272
rect 19208 18232 19214 18244
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2406 18164 2412 18216
rect 2464 18204 2470 18216
rect 4065 18207 4123 18213
rect 2464 18176 4016 18204
rect 2464 18164 2470 18176
rect 2584 18139 2642 18145
rect 2584 18105 2596 18139
rect 2630 18136 2642 18139
rect 3602 18136 3608 18148
rect 2630 18108 3608 18136
rect 2630 18105 2642 18108
rect 2584 18099 2642 18105
rect 3602 18096 3608 18108
rect 3660 18096 3666 18148
rect 3988 18136 4016 18176
rect 4065 18173 4077 18207
rect 4111 18204 4123 18207
rect 4154 18204 4160 18216
rect 4111 18176 4160 18204
rect 4111 18173 4123 18176
rect 4065 18167 4123 18173
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 6273 18207 6331 18213
rect 6273 18204 6285 18207
rect 4724 18176 6285 18204
rect 4724 18136 4752 18176
rect 6273 18173 6285 18176
rect 6319 18173 6331 18207
rect 8294 18204 8300 18216
rect 8255 18176 8300 18204
rect 6273 18167 6331 18173
rect 8294 18164 8300 18176
rect 8352 18164 8358 18216
rect 8564 18207 8622 18213
rect 8564 18173 8576 18207
rect 8610 18204 8622 18207
rect 9858 18204 9864 18216
rect 8610 18176 9864 18204
rect 8610 18173 8622 18176
rect 8564 18167 8622 18173
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10229 18207 10287 18213
rect 10229 18173 10241 18207
rect 10275 18204 10287 18207
rect 10318 18204 10324 18216
rect 10275 18176 10324 18204
rect 10275 18173 10287 18176
rect 10229 18167 10287 18173
rect 3988 18108 4752 18136
rect 4798 18096 4804 18148
rect 4856 18145 4862 18148
rect 4856 18139 4920 18145
rect 4856 18105 4874 18139
rect 4908 18105 4920 18139
rect 4856 18099 4920 18105
rect 7745 18139 7803 18145
rect 7745 18105 7757 18139
rect 7791 18136 7803 18139
rect 10152 18136 10180 18167
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 10496 18207 10554 18213
rect 10496 18173 10508 18207
rect 10542 18204 10554 18207
rect 11698 18204 11704 18216
rect 10542 18176 11704 18204
rect 10542 18173 10554 18176
rect 10496 18167 10554 18173
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 12437 18207 12495 18213
rect 12437 18173 12449 18207
rect 12483 18204 12495 18207
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12483 18176 12817 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 12805 18167 12863 18173
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 13078 18204 13084 18216
rect 13035 18176 13084 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 15930 18164 15936 18216
rect 15988 18204 15994 18216
rect 17037 18207 17095 18213
rect 17037 18204 17049 18207
rect 15988 18176 17049 18204
rect 15988 18164 15994 18176
rect 17037 18173 17049 18176
rect 17083 18173 17095 18207
rect 17037 18167 17095 18173
rect 17678 18164 17684 18216
rect 17736 18204 17742 18216
rect 17865 18207 17923 18213
rect 17865 18204 17877 18207
rect 17736 18176 17877 18204
rect 17736 18164 17742 18176
rect 17865 18173 17877 18176
rect 17911 18173 17923 18207
rect 19536 18204 19564 18380
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 20625 18343 20683 18349
rect 20625 18309 20637 18343
rect 20671 18340 20683 18343
rect 22094 18340 22100 18352
rect 20671 18312 22100 18340
rect 20671 18309 20683 18312
rect 20625 18303 20683 18309
rect 22094 18300 22100 18312
rect 22152 18300 22158 18352
rect 20806 18232 20812 18284
rect 20864 18272 20870 18284
rect 21177 18275 21235 18281
rect 21177 18272 21189 18275
rect 20864 18244 21189 18272
rect 20864 18232 20870 18244
rect 21177 18241 21189 18244
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 22465 18275 22523 18281
rect 22465 18241 22477 18275
rect 22511 18272 22523 18275
rect 22554 18272 22560 18284
rect 22511 18244 22560 18272
rect 22511 18241 22523 18244
rect 22465 18235 22523 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 20070 18204 20076 18216
rect 17865 18167 17923 18173
rect 17972 18176 19564 18204
rect 20031 18176 20076 18204
rect 10962 18136 10968 18148
rect 7791 18108 10088 18136
rect 10152 18108 10968 18136
rect 7791 18105 7803 18108
rect 7745 18099 7803 18105
rect 4856 18096 4862 18099
rect 3694 18068 3700 18080
rect 3607 18040 3700 18068
rect 3694 18028 3700 18040
rect 3752 18068 3758 18080
rect 5810 18068 5816 18080
rect 3752 18040 5816 18068
rect 3752 18028 3758 18040
rect 5810 18028 5816 18040
rect 5868 18028 5874 18080
rect 5994 18068 6000 18080
rect 5955 18040 6000 18068
rect 5994 18028 6000 18040
rect 6052 18028 6058 18080
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 7064 18040 7297 18068
rect 7064 18028 7070 18040
rect 7285 18037 7297 18040
rect 7331 18037 7343 18071
rect 7285 18031 7343 18037
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18068 7711 18071
rect 9582 18068 9588 18080
rect 7699 18040 9588 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10060 18068 10088 18108
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 13256 18139 13314 18145
rect 13256 18105 13268 18139
rect 13302 18136 13314 18139
rect 14274 18136 14280 18148
rect 13302 18108 14280 18136
rect 13302 18105 13314 18108
rect 13256 18099 13314 18105
rect 14274 18096 14280 18108
rect 14332 18136 14338 18148
rect 15013 18139 15071 18145
rect 15013 18136 15025 18139
rect 14332 18108 15025 18136
rect 14332 18096 14338 18108
rect 15013 18105 15025 18108
rect 15059 18105 15071 18139
rect 15013 18099 15071 18105
rect 15746 18096 15752 18148
rect 15804 18136 15810 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15804 18108 16129 18136
rect 15804 18096 15810 18108
rect 16117 18105 16129 18108
rect 16163 18136 16175 18139
rect 16298 18136 16304 18148
rect 16163 18108 16304 18136
rect 16163 18105 16175 18108
rect 16117 18099 16175 18105
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 16758 18136 16764 18148
rect 16671 18108 16764 18136
rect 11606 18068 11612 18080
rect 10060 18040 11612 18068
rect 11606 18028 11612 18040
rect 11664 18028 11670 18080
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 14366 18068 14372 18080
rect 12851 18040 14372 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 14516 18040 14657 18068
rect 14516 18028 14522 18040
rect 14645 18037 14657 18040
rect 14691 18037 14703 18071
rect 15102 18068 15108 18080
rect 15063 18040 15108 18068
rect 14645 18031 14703 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 15436 18040 15669 18068
rect 15436 18028 15442 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 15657 18031 15715 18037
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 16390 18068 16396 18080
rect 16071 18040 16396 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 16684 18077 16712 18108
rect 16758 18096 16764 18108
rect 16816 18136 16822 18148
rect 17972 18136 18000 18176
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 20530 18164 20536 18216
rect 20588 18204 20594 18216
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 20588 18176 22293 18204
rect 20588 18164 20594 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 16816 18108 18000 18136
rect 18316 18139 18374 18145
rect 16816 18096 16822 18108
rect 18316 18105 18328 18139
rect 18362 18136 18374 18139
rect 18782 18136 18788 18148
rect 18362 18108 18788 18136
rect 18362 18105 18374 18108
rect 18316 18099 18374 18105
rect 18782 18096 18788 18108
rect 18840 18096 18846 18148
rect 21085 18139 21143 18145
rect 21085 18136 21097 18139
rect 20272 18108 21097 18136
rect 16669 18071 16727 18077
rect 16669 18037 16681 18071
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 17126 18028 17132 18080
rect 17184 18068 17190 18080
rect 17681 18071 17739 18077
rect 17184 18040 17229 18068
rect 17184 18028 17190 18040
rect 17681 18037 17693 18071
rect 17727 18068 17739 18071
rect 18046 18068 18052 18080
rect 17727 18040 18052 18068
rect 17727 18037 17739 18040
rect 17681 18031 17739 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 20272 18077 20300 18108
rect 21085 18105 21097 18108
rect 21131 18105 21143 18139
rect 21085 18099 21143 18105
rect 20257 18071 20315 18077
rect 20257 18037 20269 18071
rect 20303 18037 20315 18071
rect 20990 18068 20996 18080
rect 20951 18040 20996 18068
rect 20257 18031 20315 18037
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 21726 18028 21732 18080
rect 21784 18068 21790 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 21784 18040 21833 18068
rect 21784 18028 21790 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 22186 18068 22192 18080
rect 22147 18040 22192 18068
rect 21821 18031 21879 18037
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 1104 17978 23276 18000
rect 1104 17926 8379 17978
rect 8431 17926 8443 17978
rect 8495 17926 8507 17978
rect 8559 17926 8571 17978
rect 8623 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 15904 17978
rect 15956 17926 15968 17978
rect 16020 17926 23276 17978
rect 1104 17904 23276 17926
rect 2314 17824 2320 17876
rect 2372 17824 2378 17876
rect 3602 17864 3608 17876
rect 3563 17836 3608 17864
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 5442 17864 5448 17876
rect 4479 17836 5448 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 8113 17867 8171 17873
rect 8113 17864 8125 17867
rect 6972 17836 8125 17864
rect 6972 17824 6978 17836
rect 8113 17833 8125 17836
rect 8159 17833 8171 17867
rect 8113 17827 8171 17833
rect 9490 17824 9496 17876
rect 9548 17864 9554 17876
rect 9861 17867 9919 17873
rect 9861 17864 9873 17867
rect 9548 17836 9873 17864
rect 9548 17824 9554 17836
rect 9861 17833 9873 17836
rect 9907 17833 9919 17867
rect 9861 17827 9919 17833
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 11422 17864 11428 17876
rect 10008 17836 11428 17864
rect 10008 17824 10014 17836
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 11698 17864 11704 17876
rect 11659 17836 11704 17864
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 13630 17864 13636 17876
rect 11940 17836 13636 17864
rect 11940 17824 11946 17836
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 14274 17864 14280 17876
rect 14235 17836 14280 17864
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 14642 17824 14648 17876
rect 14700 17864 14706 17876
rect 15654 17864 15660 17876
rect 14700 17836 15660 17864
rect 14700 17824 14706 17836
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 16850 17824 16856 17876
rect 16908 17864 16914 17876
rect 16945 17867 17003 17873
rect 16945 17864 16957 17867
rect 16908 17836 16957 17864
rect 16908 17824 16914 17836
rect 16945 17833 16957 17836
rect 16991 17833 17003 17867
rect 16945 17827 17003 17833
rect 17313 17867 17371 17873
rect 17313 17833 17325 17867
rect 17359 17864 17371 17867
rect 18046 17864 18052 17876
rect 17359 17836 18052 17864
rect 17359 17833 17371 17836
rect 17313 17827 17371 17833
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 18782 17864 18788 17876
rect 18743 17836 18788 17864
rect 18782 17824 18788 17836
rect 18840 17864 18846 17876
rect 19521 17867 19579 17873
rect 19521 17864 19533 17867
rect 18840 17836 19533 17864
rect 18840 17824 18846 17836
rect 19521 17833 19533 17836
rect 19567 17833 19579 17867
rect 19521 17827 19579 17833
rect 20441 17867 20499 17873
rect 20441 17833 20453 17867
rect 20487 17864 20499 17867
rect 20990 17864 20996 17876
rect 20487 17836 20996 17864
rect 20487 17833 20499 17836
rect 20441 17827 20499 17833
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 2332 17796 2360 17824
rect 2240 17768 2360 17796
rect 4065 17799 4123 17805
rect 1670 17728 1676 17740
rect 1631 17700 1676 17728
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 2130 17688 2136 17740
rect 2188 17728 2194 17740
rect 2240 17737 2268 17768
rect 4065 17765 4077 17799
rect 4111 17796 4123 17799
rect 10410 17796 10416 17808
rect 4111 17768 10416 17796
rect 4111 17765 4123 17768
rect 4065 17759 4123 17765
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 10588 17799 10646 17805
rect 10588 17765 10600 17799
rect 10634 17796 10646 17799
rect 12342 17796 12348 17808
rect 10634 17768 12348 17796
rect 10634 17765 10646 17768
rect 10588 17759 10646 17765
rect 12342 17756 12348 17768
rect 12400 17756 12406 17808
rect 13078 17756 13084 17808
rect 13136 17756 13142 17808
rect 15534 17799 15592 17805
rect 15534 17796 15546 17799
rect 14476 17768 15546 17796
rect 2225 17731 2283 17737
rect 2225 17728 2237 17731
rect 2188 17700 2237 17728
rect 2188 17688 2194 17700
rect 2225 17697 2237 17700
rect 2271 17697 2283 17731
rect 2225 17691 2283 17697
rect 2314 17688 2320 17740
rect 2372 17728 2378 17740
rect 2481 17731 2539 17737
rect 2481 17728 2493 17731
rect 2372 17700 2493 17728
rect 2372 17688 2378 17700
rect 2481 17697 2493 17700
rect 2527 17697 2539 17731
rect 4246 17728 4252 17740
rect 4207 17700 4252 17728
rect 2481 17691 2539 17697
rect 4246 17688 4252 17700
rect 4304 17688 4310 17740
rect 5074 17737 5080 17740
rect 5068 17691 5080 17737
rect 5132 17728 5138 17740
rect 5132 17700 5168 17728
rect 5074 17688 5080 17691
rect 5132 17688 5138 17700
rect 6270 17688 6276 17740
rect 6328 17728 6334 17740
rect 6713 17731 6771 17737
rect 6713 17728 6725 17731
rect 6328 17700 6725 17728
rect 6328 17688 6334 17700
rect 6713 17697 6725 17700
rect 6759 17697 6771 17731
rect 6713 17691 6771 17697
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 9306 17728 9312 17740
rect 8527 17700 9312 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 9306 17688 9312 17700
rect 9364 17688 9370 17740
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 9766 17728 9772 17740
rect 9723 17700 9772 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 11790 17688 11796 17740
rect 11848 17728 11854 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11848 17700 11989 17728
rect 11848 17688 11854 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 12897 17731 12955 17737
rect 12897 17728 12909 17731
rect 12676 17700 12909 17728
rect 12676 17688 12682 17700
rect 12897 17697 12909 17700
rect 12943 17728 12955 17731
rect 13096 17728 13124 17756
rect 12943 17700 13124 17728
rect 13164 17731 13222 17737
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 13164 17697 13176 17731
rect 13210 17728 13222 17731
rect 13998 17728 14004 17740
rect 13210 17700 14004 17728
rect 13210 17697 13222 17700
rect 13164 17691 13222 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 14090 17688 14096 17740
rect 14148 17728 14154 17740
rect 14476 17728 14504 17768
rect 15534 17765 15546 17768
rect 15580 17796 15592 17799
rect 16114 17796 16120 17808
rect 15580 17768 16120 17796
rect 15580 17765 15592 17768
rect 15534 17759 15592 17765
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 17586 17756 17592 17808
rect 17644 17756 17650 17808
rect 19334 17756 19340 17808
rect 19392 17796 19398 17808
rect 19429 17799 19487 17805
rect 19429 17796 19441 17799
rect 19392 17768 19441 17796
rect 19392 17756 19398 17768
rect 19429 17765 19441 17768
rect 19475 17765 19487 17799
rect 19429 17759 19487 17765
rect 21628 17799 21686 17805
rect 21628 17765 21640 17799
rect 21674 17796 21686 17799
rect 22646 17796 22652 17808
rect 21674 17768 22652 17796
rect 21674 17765 21686 17768
rect 21628 17759 21686 17765
rect 22646 17756 22652 17768
rect 22704 17756 22710 17808
rect 14148 17700 14504 17728
rect 14148 17688 14154 17700
rect 14550 17688 14556 17740
rect 14608 17728 14614 17740
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 14608 17700 14657 17728
rect 14608 17688 14614 17700
rect 14645 17697 14657 17700
rect 14691 17697 14703 17731
rect 17604 17728 17632 17756
rect 14645 17691 14703 17697
rect 15212 17700 17632 17728
rect 17672 17731 17730 17737
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 4801 17663 4859 17669
rect 4801 17660 4813 17663
rect 4488 17632 4813 17660
rect 4488 17620 4494 17632
rect 4801 17629 4813 17632
rect 4847 17629 4859 17663
rect 4801 17623 4859 17629
rect 6362 17620 6368 17672
rect 6420 17660 6426 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 6420 17632 6469 17660
rect 6420 17620 6426 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 8665 17663 8723 17669
rect 8665 17629 8677 17663
rect 8711 17660 8723 17663
rect 9125 17663 9183 17669
rect 8711 17632 9076 17660
rect 8711 17629 8723 17632
rect 8665 17623 8723 17629
rect 4065 17595 4123 17601
rect 4065 17592 4077 17595
rect 3620 17564 4077 17592
rect 1857 17527 1915 17533
rect 1857 17493 1869 17527
rect 1903 17524 1915 17527
rect 3620 17524 3648 17564
rect 4065 17561 4077 17564
rect 4111 17561 4123 17595
rect 4065 17555 4123 17561
rect 4154 17552 4160 17604
rect 4212 17592 4218 17604
rect 4522 17592 4528 17604
rect 4212 17564 4528 17592
rect 4212 17552 4218 17564
rect 4522 17552 4528 17564
rect 4580 17552 4586 17604
rect 8588 17592 8616 17623
rect 8754 17592 8760 17604
rect 8588 17564 8760 17592
rect 8754 17552 8760 17564
rect 8812 17552 8818 17604
rect 9048 17592 9076 17632
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 9214 17660 9220 17672
rect 9171 17632 9220 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 10318 17660 10324 17672
rect 10279 17632 10324 17660
rect 10318 17620 10324 17632
rect 10376 17620 10382 17672
rect 10226 17592 10232 17604
rect 9048 17564 10232 17592
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 1903 17496 3648 17524
rect 1903 17493 1915 17496
rect 1857 17487 1915 17493
rect 3694 17484 3700 17536
rect 3752 17524 3758 17536
rect 6086 17524 6092 17536
rect 3752 17496 6092 17524
rect 3752 17484 3758 17496
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 6181 17527 6239 17533
rect 6181 17493 6193 17527
rect 6227 17524 6239 17527
rect 6270 17524 6276 17536
rect 6227 17496 6276 17524
rect 6227 17493 6239 17496
rect 6181 17487 6239 17493
rect 6270 17484 6276 17496
rect 6328 17484 6334 17536
rect 7466 17484 7472 17536
rect 7524 17524 7530 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7524 17496 7849 17524
rect 7524 17484 7530 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 11422 17524 11428 17536
rect 7984 17496 11428 17524
rect 7984 17484 7990 17496
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12161 17527 12219 17533
rect 12161 17524 12173 17527
rect 11756 17496 12173 17524
rect 11756 17484 11762 17496
rect 12161 17493 12173 17496
rect 12207 17493 12219 17527
rect 12161 17487 12219 17493
rect 14829 17527 14887 17533
rect 14829 17493 14841 17527
rect 14875 17524 14887 17527
rect 15212 17524 15240 17700
rect 17672 17697 17684 17731
rect 17718 17728 17730 17731
rect 18966 17728 18972 17740
rect 17718 17700 18972 17728
rect 17718 17697 17730 17700
rect 17672 17691 17730 17697
rect 18966 17688 18972 17700
rect 19024 17688 19030 17740
rect 20070 17688 20076 17740
rect 20128 17728 20134 17740
rect 20257 17731 20315 17737
rect 20257 17728 20269 17731
rect 20128 17700 20269 17728
rect 20128 17688 20134 17700
rect 20257 17697 20269 17700
rect 20303 17697 20315 17731
rect 20257 17691 20315 17697
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 17313 17663 17371 17669
rect 15344 17632 15389 17660
rect 15344 17620 15350 17632
rect 17313 17629 17325 17663
rect 17359 17660 17371 17663
rect 17402 17660 17408 17672
rect 17359 17632 17408 17660
rect 17359 17629 17371 17632
rect 17313 17623 17371 17629
rect 17402 17620 17408 17632
rect 17460 17620 17466 17672
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 19886 17660 19892 17672
rect 19751 17632 19892 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20898 17660 20904 17672
rect 20859 17632 20904 17660
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 20990 17620 20996 17672
rect 21048 17660 21054 17672
rect 21266 17660 21272 17672
rect 21048 17632 21272 17660
rect 21048 17620 21054 17632
rect 21266 17620 21272 17632
rect 21324 17660 21330 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 21324 17632 21373 17660
rect 21324 17620 21330 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 19794 17592 19800 17604
rect 16356 17564 16804 17592
rect 16356 17552 16362 17564
rect 14875 17496 15240 17524
rect 14875 17493 14887 17496
rect 14829 17487 14887 17493
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 16669 17527 16727 17533
rect 16669 17524 16681 17527
rect 15620 17496 16681 17524
rect 15620 17484 15626 17496
rect 16669 17493 16681 17496
rect 16715 17493 16727 17527
rect 16776 17524 16804 17564
rect 18340 17564 19800 17592
rect 18340 17524 18368 17564
rect 19794 17552 19800 17564
rect 19852 17552 19858 17604
rect 19058 17524 19064 17536
rect 16776 17496 18368 17524
rect 19019 17496 19064 17524
rect 16669 17487 16727 17493
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 20806 17484 20812 17536
rect 20864 17524 20870 17536
rect 22741 17527 22799 17533
rect 22741 17524 22753 17527
rect 20864 17496 22753 17524
rect 20864 17484 20870 17496
rect 22741 17493 22753 17496
rect 22787 17493 22799 17527
rect 22741 17487 22799 17493
rect 1104 17434 23276 17456
rect 1104 17382 4680 17434
rect 4732 17382 4744 17434
rect 4796 17382 4808 17434
rect 4860 17382 4872 17434
rect 4924 17382 12078 17434
rect 12130 17382 12142 17434
rect 12194 17382 12206 17434
rect 12258 17382 12270 17434
rect 12322 17382 19475 17434
rect 19527 17382 19539 17434
rect 19591 17382 19603 17434
rect 19655 17382 19667 17434
rect 19719 17382 23276 17434
rect 1104 17360 23276 17382
rect 1765 17323 1823 17329
rect 1765 17289 1777 17323
rect 1811 17320 1823 17323
rect 3513 17323 3571 17329
rect 1811 17292 3470 17320
rect 1811 17289 1823 17292
rect 1765 17283 1823 17289
rect 3442 17252 3470 17292
rect 3513 17289 3525 17323
rect 3559 17320 3571 17323
rect 3605 17323 3663 17329
rect 3605 17320 3617 17323
rect 3559 17292 3617 17320
rect 3559 17289 3571 17292
rect 3513 17283 3571 17289
rect 3605 17289 3617 17292
rect 3651 17320 3663 17323
rect 3651 17292 4660 17320
rect 3651 17289 3663 17292
rect 3605 17283 3663 17289
rect 4632 17264 4660 17292
rect 6086 17280 6092 17332
rect 6144 17320 6150 17332
rect 11701 17323 11759 17329
rect 6144 17292 11284 17320
rect 6144 17280 6150 17292
rect 3694 17252 3700 17264
rect 3442 17224 3700 17252
rect 3694 17212 3700 17224
rect 3752 17212 3758 17264
rect 3789 17255 3847 17261
rect 3789 17221 3801 17255
rect 3835 17252 3847 17255
rect 4522 17252 4528 17264
rect 3835 17224 4528 17252
rect 3835 17221 3847 17224
rect 3789 17215 3847 17221
rect 4522 17212 4528 17224
rect 4580 17212 4586 17264
rect 4614 17212 4620 17264
rect 4672 17212 4678 17264
rect 5905 17255 5963 17261
rect 5905 17221 5917 17255
rect 5951 17252 5963 17255
rect 6362 17252 6368 17264
rect 5951 17224 6368 17252
rect 5951 17221 5963 17224
rect 5905 17215 5963 17221
rect 6362 17212 6368 17224
rect 6420 17252 6426 17264
rect 9861 17255 9919 17261
rect 6420 17224 6868 17252
rect 6420 17212 6426 17224
rect 2130 17184 2136 17196
rect 2091 17156 2136 17184
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 3602 17144 3608 17196
rect 3660 17184 3666 17196
rect 4341 17187 4399 17193
rect 4341 17184 4353 17187
rect 3660 17156 4353 17184
rect 3660 17144 3666 17156
rect 4341 17153 4353 17156
rect 4387 17153 4399 17187
rect 4341 17147 4399 17153
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17085 1639 17119
rect 2774 17116 2780 17128
rect 1581 17079 1639 17085
rect 2240 17088 2780 17116
rect 1596 17048 1624 17079
rect 2240 17048 2268 17088
rect 2774 17076 2780 17088
rect 2832 17076 2838 17128
rect 3694 17116 3700 17128
rect 3068 17088 3700 17116
rect 1596 17020 2268 17048
rect 2400 17051 2458 17057
rect 2400 17017 2412 17051
rect 2446 17048 2458 17051
rect 3068 17048 3096 17088
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 4157 17119 4215 17125
rect 4157 17116 4169 17119
rect 4080 17088 4169 17116
rect 4080 17060 4108 17088
rect 4157 17085 4169 17088
rect 4203 17085 4215 17119
rect 4157 17079 4215 17085
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 5368 17116 5396 17147
rect 5534 17144 5540 17196
rect 5592 17184 5598 17196
rect 6730 17184 6736 17196
rect 5592 17156 6736 17184
rect 5592 17144 5598 17156
rect 6086 17116 6092 17128
rect 4304 17088 5396 17116
rect 6047 17088 6092 17116
rect 4304 17076 4310 17088
rect 6086 17076 6092 17088
rect 6144 17076 6150 17128
rect 6196 17125 6224 17156
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 6840 17193 6868 17224
rect 9861 17221 9873 17255
rect 9907 17221 9919 17255
rect 11256 17252 11284 17292
rect 11701 17289 11713 17323
rect 11747 17320 11759 17323
rect 11974 17320 11980 17332
rect 11747 17292 11980 17320
rect 11747 17289 11759 17292
rect 11701 17283 11759 17289
rect 11974 17280 11980 17292
rect 12032 17280 12038 17332
rect 20990 17320 20996 17332
rect 12268 17292 17356 17320
rect 12268 17264 12296 17292
rect 11882 17252 11888 17264
rect 11256 17224 11888 17252
rect 9861 17215 9919 17221
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 8481 17187 8539 17193
rect 8481 17184 8493 17187
rect 8352 17156 8493 17184
rect 8352 17144 8358 17156
rect 8481 17153 8493 17156
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17085 6239 17119
rect 7834 17116 7840 17128
rect 6181 17079 6239 17085
rect 7024 17088 7840 17116
rect 2446 17020 3096 17048
rect 2446 17017 2458 17020
rect 2400 17011 2458 17017
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 3970 17048 3976 17060
rect 3200 17020 3976 17048
rect 3200 17008 3206 17020
rect 3970 17008 3976 17020
rect 4028 17008 4034 17060
rect 4062 17008 4068 17060
rect 4120 17008 4126 17060
rect 5169 17051 5227 17057
rect 5169 17017 5181 17051
rect 5215 17048 5227 17051
rect 7024 17048 7052 17088
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 9876 17116 9904 17215
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 12250 17212 12256 17264
rect 12308 17212 12314 17264
rect 13998 17252 14004 17264
rect 13911 17224 14004 17252
rect 13998 17212 14004 17224
rect 14056 17252 14062 17264
rect 15102 17252 15108 17264
rect 14056 17224 15108 17252
rect 14056 17212 14062 17224
rect 15102 17212 15108 17224
rect 15160 17212 15166 17264
rect 16485 17255 16543 17261
rect 16485 17221 16497 17255
rect 16531 17252 16543 17255
rect 16574 17252 16580 17264
rect 16531 17224 16580 17252
rect 16531 17221 16543 17224
rect 16485 17215 16543 17221
rect 16574 17212 16580 17224
rect 16632 17212 16638 17264
rect 16761 17255 16819 17261
rect 16761 17221 16773 17255
rect 16807 17252 16819 17255
rect 17126 17252 17132 17264
rect 16807 17224 17132 17252
rect 16807 17221 16819 17224
rect 16761 17215 16819 17221
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 12618 17184 12624 17196
rect 12579 17156 12624 17184
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 17328 17193 17356 17292
rect 20272 17292 20996 17320
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18874 17252 18880 17264
rect 18012 17224 18880 17252
rect 18012 17212 18018 17224
rect 18874 17212 18880 17224
rect 18932 17212 18938 17264
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17184 14243 17187
rect 17313 17187 17371 17193
rect 14231 17156 15148 17184
rect 14231 17153 14243 17156
rect 14185 17147 14243 17153
rect 15120 17128 15148 17156
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17184 19303 17187
rect 19886 17184 19892 17196
rect 19291 17156 19892 17184
rect 19291 17153 19303 17156
rect 19245 17147 19303 17153
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 20272 17193 20300 17292
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 21634 17320 21640 17332
rect 21547 17292 21640 17320
rect 21634 17280 21640 17292
rect 21692 17320 21698 17332
rect 21692 17292 22508 17320
rect 21692 17280 21698 17292
rect 22480 17193 22508 17292
rect 20257 17187 20315 17193
rect 20257 17153 20269 17187
rect 20303 17153 20315 17187
rect 20257 17147 20315 17153
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17153 22523 17187
rect 22465 17147 22523 17153
rect 22738 17144 22744 17196
rect 22796 17184 22802 17196
rect 23382 17184 23388 17196
rect 22796 17156 23388 17184
rect 22796 17144 22802 17156
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 10318 17116 10324 17128
rect 7984 17088 9904 17116
rect 10279 17088 10324 17116
rect 7984 17076 7990 17088
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 12066 17116 12072 17128
rect 11480 17088 12072 17116
rect 11480 17076 11486 17088
rect 12066 17076 12072 17088
rect 12124 17076 12130 17128
rect 12888 17119 12946 17125
rect 12888 17085 12900 17119
rect 12934 17116 12946 17119
rect 13262 17116 13268 17128
rect 12934 17088 13268 17116
rect 12934 17085 12946 17088
rect 12888 17079 12946 17085
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14424 17088 14473 17116
rect 14424 17076 14430 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17116 14611 17119
rect 14826 17116 14832 17128
rect 14599 17088 14832 17116
rect 14599 17085 14611 17088
rect 14553 17079 14611 17085
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 15102 17116 15108 17128
rect 15063 17088 15108 17116
rect 15102 17076 15108 17088
rect 15160 17076 15166 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 15212 17088 18061 17116
rect 5215 17020 7052 17048
rect 7092 17051 7150 17057
rect 5215 17017 5227 17020
rect 5169 17011 5227 17017
rect 7092 17017 7104 17051
rect 7138 17048 7150 17051
rect 7466 17048 7472 17060
rect 7138 17020 7472 17048
rect 7138 17017 7150 17020
rect 7092 17011 7150 17017
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 8748 17051 8806 17057
rect 8748 17048 8760 17051
rect 8220 17020 8760 17048
rect 2314 16940 2320 16992
rect 2372 16980 2378 16992
rect 3605 16983 3663 16989
rect 3605 16980 3617 16983
rect 2372 16952 3617 16980
rect 2372 16940 2378 16952
rect 3605 16949 3617 16952
rect 3651 16949 3663 16983
rect 3605 16943 3663 16949
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4801 16983 4859 16989
rect 4304 16952 4349 16980
rect 4304 16940 4310 16952
rect 4801 16949 4813 16983
rect 4847 16980 4859 16983
rect 4982 16980 4988 16992
rect 4847 16952 4988 16980
rect 4847 16949 4859 16952
rect 4801 16943 4859 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 5258 16940 5264 16992
rect 5316 16980 5322 16992
rect 6365 16983 6423 16989
rect 5316 16952 5361 16980
rect 5316 16940 5322 16952
rect 6365 16949 6377 16983
rect 6411 16980 6423 16983
rect 7650 16980 7656 16992
rect 6411 16952 7656 16980
rect 6411 16949 6423 16952
rect 6365 16943 6423 16949
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 8220 16989 8248 17020
rect 8748 17017 8760 17020
rect 8794 17048 8806 17051
rect 9030 17048 9036 17060
rect 8794 17020 9036 17048
rect 8794 17017 8806 17020
rect 8748 17011 8806 17017
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 9122 17008 9128 17060
rect 9180 17048 9186 17060
rect 10588 17051 10646 17057
rect 9180 17020 9996 17048
rect 9180 17008 9186 17020
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16949 8263 16983
rect 8205 16943 8263 16949
rect 8662 16940 8668 16992
rect 8720 16980 8726 16992
rect 9858 16980 9864 16992
rect 8720 16952 9864 16980
rect 8720 16940 8726 16952
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 9968 16980 9996 17020
rect 10588 17017 10600 17051
rect 10634 17048 10646 17051
rect 11054 17048 11060 17060
rect 10634 17020 11060 17048
rect 10634 17017 10646 17020
rect 10588 17011 10646 17017
rect 11054 17008 11060 17020
rect 11112 17048 11118 17060
rect 11112 17020 12940 17048
rect 11112 17008 11118 17020
rect 11422 16980 11428 16992
rect 9968 16952 11428 16980
rect 11422 16940 11428 16952
rect 11480 16940 11486 16992
rect 12912 16980 12940 17020
rect 12986 17008 12992 17060
rect 13044 17048 13050 17060
rect 15212 17048 15240 17088
rect 18049 17085 18061 17088
rect 18095 17085 18107 17119
rect 18966 17116 18972 17128
rect 18927 17088 18972 17116
rect 18049 17079 18107 17085
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17116 19763 17119
rect 20162 17116 20168 17128
rect 19751 17088 20168 17116
rect 19751 17085 19763 17088
rect 19705 17079 19763 17085
rect 20162 17076 20168 17088
rect 20220 17076 20226 17128
rect 20524 17119 20582 17125
rect 20524 17085 20536 17119
rect 20570 17116 20582 17119
rect 20806 17116 20812 17128
rect 20570 17088 20812 17116
rect 20570 17085 20582 17088
rect 20524 17079 20582 17085
rect 20806 17076 20812 17088
rect 20864 17076 20870 17128
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 20956 17088 22293 17116
rect 20956 17076 20962 17088
rect 22281 17085 22293 17088
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 13044 17020 15240 17048
rect 15372 17051 15430 17057
rect 13044 17008 13050 17020
rect 15372 17017 15384 17051
rect 15418 17048 15430 17051
rect 15562 17048 15568 17060
rect 15418 17020 15568 17048
rect 15418 17017 15430 17020
rect 15372 17011 15430 17017
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 16758 17008 16764 17060
rect 16816 17048 16822 17060
rect 17221 17051 17279 17057
rect 17221 17048 17233 17051
rect 16816 17020 17233 17048
rect 16816 17008 16822 17020
rect 17221 17017 17233 17020
rect 17267 17017 17279 17051
rect 17221 17011 17279 17017
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 21358 17048 21364 17060
rect 19300 17020 21364 17048
rect 19300 17008 19306 17020
rect 21358 17008 21364 17020
rect 21416 17008 21422 17060
rect 22094 17008 22100 17060
rect 22152 17048 22158 17060
rect 22373 17051 22431 17057
rect 22373 17048 22385 17051
rect 22152 17020 22385 17048
rect 22152 17008 22158 17020
rect 22373 17017 22385 17020
rect 22419 17017 22431 17051
rect 22373 17011 22431 17017
rect 14090 16980 14096 16992
rect 12912 16952 14096 16980
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 14185 16983 14243 16989
rect 14185 16949 14197 16983
rect 14231 16980 14243 16983
rect 14277 16983 14335 16989
rect 14277 16980 14289 16983
rect 14231 16952 14289 16980
rect 14231 16949 14243 16952
rect 14185 16943 14243 16949
rect 14277 16949 14289 16952
rect 14323 16949 14335 16983
rect 14277 16943 14335 16949
rect 14737 16983 14795 16989
rect 14737 16949 14749 16983
rect 14783 16980 14795 16983
rect 16206 16980 16212 16992
rect 14783 16952 16212 16980
rect 14783 16949 14795 16952
rect 14737 16943 14795 16949
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 17126 16980 17132 16992
rect 17087 16952 17132 16980
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 18230 16980 18236 16992
rect 18191 16952 18236 16980
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 18601 16983 18659 16989
rect 18601 16980 18613 16983
rect 18564 16952 18613 16980
rect 18564 16940 18570 16952
rect 18601 16949 18613 16952
rect 18647 16949 18659 16983
rect 18601 16943 18659 16949
rect 19061 16983 19119 16989
rect 19061 16949 19073 16983
rect 19107 16980 19119 16983
rect 19794 16980 19800 16992
rect 19107 16952 19800 16980
rect 19107 16949 19119 16952
rect 19061 16943 19119 16949
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 19889 16983 19947 16989
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 19978 16980 19984 16992
rect 19935 16952 19984 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 19978 16940 19984 16952
rect 20036 16940 20042 16992
rect 21913 16983 21971 16989
rect 21913 16949 21925 16983
rect 21959 16980 21971 16983
rect 22002 16980 22008 16992
rect 21959 16952 22008 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 1104 16890 23276 16912
rect 1104 16838 8379 16890
rect 8431 16838 8443 16890
rect 8495 16838 8507 16890
rect 8559 16838 8571 16890
rect 8623 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 15904 16890
rect 15956 16838 15968 16890
rect 16020 16838 23276 16890
rect 1104 16816 23276 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 2774 16776 2780 16788
rect 1627 16748 2780 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 3142 16776 3148 16788
rect 2884 16748 3148 16776
rect 2884 16708 2912 16748
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3329 16779 3387 16785
rect 3329 16745 3341 16779
rect 3375 16776 3387 16779
rect 3602 16776 3608 16788
rect 3375 16748 3608 16776
rect 3375 16745 3387 16748
rect 3329 16739 3387 16745
rect 3602 16736 3608 16748
rect 3660 16736 3666 16788
rect 4065 16779 4123 16785
rect 4065 16745 4077 16779
rect 4111 16776 4123 16779
rect 4246 16776 4252 16788
rect 4111 16748 4252 16776
rect 4111 16745 4123 16748
rect 4065 16739 4123 16745
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 4433 16779 4491 16785
rect 4433 16745 4445 16779
rect 4479 16776 4491 16779
rect 4893 16779 4951 16785
rect 4893 16776 4905 16779
rect 4479 16748 4905 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 4893 16745 4905 16748
rect 4939 16745 4951 16779
rect 4893 16739 4951 16745
rect 5077 16779 5135 16785
rect 5077 16745 5089 16779
rect 5123 16776 5135 16779
rect 5258 16776 5264 16788
rect 5123 16748 5264 16776
rect 5123 16745 5135 16748
rect 5077 16739 5135 16745
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 9122 16776 9128 16788
rect 5368 16748 9128 16776
rect 1412 16680 2912 16708
rect 1412 16649 1440 16680
rect 2958 16668 2964 16720
rect 3016 16708 3022 16720
rect 4525 16711 4583 16717
rect 4525 16708 4537 16711
rect 3016 16680 4016 16708
rect 3016 16668 3022 16680
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16609 1455 16643
rect 1397 16603 1455 16609
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2038 16640 2044 16652
rect 1995 16612 2044 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2216 16643 2274 16649
rect 2216 16609 2228 16643
rect 2262 16640 2274 16643
rect 3418 16640 3424 16652
rect 2262 16612 3424 16640
rect 2262 16609 2274 16612
rect 2216 16603 2274 16609
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 3988 16572 4016 16680
rect 4172 16680 4537 16708
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4172 16640 4200 16680
rect 4525 16677 4537 16680
rect 4571 16677 4583 16711
rect 5368 16708 5396 16748
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9398 16736 9404 16788
rect 9456 16736 9462 16788
rect 11054 16776 11060 16788
rect 11015 16748 11060 16776
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11241 16779 11299 16785
rect 11241 16745 11253 16779
rect 11287 16776 11299 16779
rect 11333 16779 11391 16785
rect 11333 16776 11345 16779
rect 11287 16748 11345 16776
rect 11287 16745 11299 16748
rect 11241 16739 11299 16745
rect 11333 16745 11345 16748
rect 11379 16745 11391 16779
rect 11333 16739 11391 16745
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 11480 16748 11928 16776
rect 11480 16736 11486 16748
rect 4525 16671 4583 16677
rect 4632 16680 5396 16708
rect 5537 16711 5595 16717
rect 4632 16640 4660 16680
rect 5537 16677 5549 16711
rect 5583 16708 5595 16711
rect 5994 16708 6000 16720
rect 5583 16680 6000 16708
rect 5583 16677 5595 16680
rect 5537 16671 5595 16677
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 6540 16711 6598 16717
rect 6540 16677 6552 16711
rect 6586 16708 6598 16711
rect 7742 16708 7748 16720
rect 6586 16680 7748 16708
rect 6586 16677 6598 16680
rect 6540 16671 6598 16677
rect 7742 16668 7748 16680
rect 7800 16708 7806 16720
rect 7926 16708 7932 16720
rect 7800 16680 7932 16708
rect 7800 16668 7806 16680
rect 7926 16668 7932 16680
rect 7984 16668 7990 16720
rect 8196 16711 8254 16717
rect 8196 16677 8208 16711
rect 8242 16708 8254 16711
rect 8846 16708 8852 16720
rect 8242 16680 8852 16708
rect 8242 16677 8254 16680
rect 8196 16671 8254 16677
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 9416 16708 9444 16736
rect 9140 16680 9444 16708
rect 9140 16652 9168 16680
rect 10042 16668 10048 16720
rect 10100 16668 10106 16720
rect 10318 16668 10324 16720
rect 10376 16708 10382 16720
rect 10594 16708 10600 16720
rect 10376 16680 10600 16708
rect 10376 16668 10382 16680
rect 10594 16668 10600 16680
rect 10652 16708 10658 16720
rect 11900 16708 11928 16748
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 12124 16748 13369 16776
rect 12124 16736 12130 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 13357 16739 13415 16745
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 13817 16779 13875 16785
rect 13817 16776 13829 16779
rect 13596 16748 13829 16776
rect 13596 16736 13602 16748
rect 13817 16745 13829 16748
rect 13863 16745 13875 16779
rect 13817 16739 13875 16745
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 16298 16776 16304 16788
rect 14148 16748 16304 16776
rect 14148 16736 14154 16748
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16540 16748 16681 16776
rect 16540 16736 16546 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 16945 16779 17003 16785
rect 16945 16745 16957 16779
rect 16991 16776 17003 16779
rect 17405 16779 17463 16785
rect 16991 16748 17356 16776
rect 16991 16745 17003 16748
rect 16945 16739 17003 16745
rect 10652 16680 11744 16708
rect 11900 16680 14596 16708
rect 10652 16668 10658 16680
rect 4120 16612 4200 16640
rect 4540 16612 4660 16640
rect 4893 16643 4951 16649
rect 4120 16600 4126 16612
rect 4540 16572 4568 16612
rect 4893 16609 4905 16643
rect 4939 16609 4951 16643
rect 4893 16603 4951 16609
rect 3988 16544 4568 16572
rect 4614 16532 4620 16584
rect 4672 16572 4678 16584
rect 4908 16572 4936 16603
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 5445 16643 5503 16649
rect 5445 16640 5457 16643
rect 5040 16612 5457 16640
rect 5040 16600 5046 16612
rect 5445 16609 5457 16612
rect 5491 16609 5503 16643
rect 8662 16640 8668 16652
rect 5445 16603 5503 16609
rect 5552 16612 8668 16640
rect 5552 16572 5580 16612
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9122 16600 9128 16652
rect 9180 16600 9186 16652
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 9933 16643 9991 16649
rect 9933 16640 9945 16643
rect 9456 16612 9945 16640
rect 9456 16600 9462 16612
rect 9933 16609 9945 16612
rect 9979 16609 9991 16643
rect 10060 16640 10088 16668
rect 10060 16612 10712 16640
rect 9933 16603 9991 16609
rect 4672 16544 4717 16572
rect 4908 16544 5580 16572
rect 5629 16575 5687 16581
rect 4672 16532 4678 16544
rect 5629 16541 5641 16575
rect 5675 16541 5687 16575
rect 6270 16572 6276 16584
rect 6231 16544 6276 16572
rect 5629 16535 5687 16541
rect 4246 16464 4252 16516
rect 4304 16504 4310 16516
rect 5166 16504 5172 16516
rect 4304 16476 5172 16504
rect 4304 16464 4310 16476
rect 5166 16464 5172 16476
rect 5224 16464 5230 16516
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 5644 16436 5672 16535
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16541 9735 16575
rect 10684 16572 10712 16612
rect 10962 16600 10968 16652
rect 11020 16640 11026 16652
rect 11716 16649 11744 16680
rect 11974 16649 11980 16652
rect 11241 16643 11299 16649
rect 11241 16640 11253 16643
rect 11020 16612 11253 16640
rect 11020 16600 11026 16612
rect 11241 16609 11253 16612
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16609 11759 16643
rect 11968 16640 11980 16649
rect 11887 16612 11980 16640
rect 11701 16603 11759 16609
rect 11968 16603 11980 16612
rect 12032 16640 12038 16652
rect 12250 16640 12256 16652
rect 12032 16612 12256 16640
rect 11532 16572 11560 16603
rect 11974 16600 11980 16603
rect 12032 16600 12038 16612
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 14458 16640 14464 16652
rect 13771 16612 14464 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 10684 16544 11560 16572
rect 9677 16535 9735 16541
rect 3476 16408 5672 16436
rect 3476 16396 3482 16408
rect 7374 16396 7380 16448
rect 7432 16436 7438 16448
rect 7653 16439 7711 16445
rect 7653 16436 7665 16439
rect 7432 16408 7665 16436
rect 7432 16396 7438 16408
rect 7653 16405 7665 16408
rect 7699 16405 7711 16439
rect 7944 16436 7972 16535
rect 9309 16507 9367 16513
rect 9309 16473 9321 16507
rect 9355 16504 9367 16507
rect 9398 16504 9404 16516
rect 9355 16476 9404 16504
rect 9355 16473 9367 16476
rect 9309 16467 9367 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 9692 16448 9720 16535
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 13909 16575 13967 16581
rect 13909 16572 13921 16575
rect 13688 16544 13921 16572
rect 13688 16532 13694 16544
rect 13909 16541 13921 16544
rect 13955 16541 13967 16575
rect 14568 16572 14596 16680
rect 15010 16668 15016 16720
rect 15068 16708 15074 16720
rect 17328 16708 17356 16748
rect 17405 16745 17417 16779
rect 17451 16776 17463 16779
rect 17586 16776 17592 16788
rect 17451 16748 17592 16776
rect 17451 16745 17463 16748
rect 17405 16739 17463 16745
rect 17586 16736 17592 16748
rect 17644 16736 17650 16788
rect 18966 16736 18972 16788
rect 19024 16776 19030 16788
rect 19153 16779 19211 16785
rect 19153 16776 19165 16779
rect 19024 16748 19165 16776
rect 19024 16736 19030 16748
rect 19153 16745 19165 16748
rect 19199 16745 19211 16779
rect 19153 16739 19211 16745
rect 19794 16736 19800 16788
rect 19852 16736 19858 16788
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 22557 16779 22615 16785
rect 22557 16776 22569 16779
rect 22244 16748 22569 16776
rect 22244 16736 22250 16748
rect 22557 16745 22569 16748
rect 22603 16745 22615 16779
rect 22557 16739 22615 16745
rect 17678 16708 17684 16720
rect 15068 16680 17172 16708
rect 17328 16680 17684 16708
rect 15068 16668 15074 16680
rect 14642 16600 14648 16652
rect 14700 16640 14706 16652
rect 15286 16640 15292 16652
rect 14700 16612 14745 16640
rect 15247 16612 15292 16640
rect 14700 16600 14706 16612
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15556 16643 15614 16649
rect 15556 16609 15568 16643
rect 15602 16640 15614 16643
rect 16574 16640 16580 16652
rect 15602 16612 16580 16640
rect 15602 16609 15614 16612
rect 15556 16603 15614 16609
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 17144 16649 17172 16680
rect 17678 16668 17684 16680
rect 17736 16668 17742 16720
rect 18040 16711 18098 16717
rect 18040 16677 18052 16711
rect 18086 16708 18098 16711
rect 19812 16708 19840 16736
rect 18086 16680 19840 16708
rect 18086 16677 18098 16680
rect 18040 16671 18098 16677
rect 19886 16668 19892 16720
rect 19944 16708 19950 16720
rect 21168 16711 21226 16717
rect 19944 16680 20116 16708
rect 19944 16668 19950 16680
rect 17129 16643 17187 16649
rect 17129 16609 17141 16643
rect 17175 16609 17187 16643
rect 17129 16603 17187 16609
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16640 17279 16643
rect 19242 16640 19248 16652
rect 17267 16612 19248 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19484 16612 19809 16640
rect 19484 16600 19490 16612
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 14568 16544 14872 16572
rect 13909 16535 13967 16541
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 14734 16504 14740 16516
rect 13320 16476 14740 16504
rect 13320 16464 13326 16476
rect 14734 16464 14740 16476
rect 14792 16464 14798 16516
rect 14844 16513 14872 16544
rect 17402 16532 17408 16584
rect 17460 16572 17466 16584
rect 17773 16575 17831 16581
rect 17773 16572 17785 16575
rect 17460 16544 17785 16572
rect 17460 16532 17466 16544
rect 17773 16541 17785 16544
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 19334 16532 19340 16584
rect 19392 16572 19398 16584
rect 20088 16581 20116 16680
rect 21168 16677 21180 16711
rect 21214 16708 21226 16711
rect 21634 16708 21640 16720
rect 21214 16680 21640 16708
rect 21214 16677 21226 16680
rect 21168 16671 21226 16677
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 19889 16575 19947 16581
rect 19392 16544 19437 16572
rect 19392 16532 19398 16544
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16572 20131 16575
rect 20438 16572 20444 16584
rect 20119 16544 20444 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 14829 16507 14887 16513
rect 14829 16473 14841 16507
rect 14875 16473 14887 16507
rect 19904 16504 19932 16535
rect 20438 16532 20444 16544
rect 20496 16532 20502 16584
rect 20898 16572 20904 16584
rect 20859 16544 20904 16572
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 14829 16467 14887 16473
rect 18708 16476 19932 16504
rect 9674 16436 9680 16448
rect 7944 16408 9680 16436
rect 7653 16399 7711 16405
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 9858 16396 9864 16448
rect 9916 16436 9922 16448
rect 13081 16439 13139 16445
rect 13081 16436 13093 16439
rect 9916 16408 13093 16436
rect 9916 16396 9922 16408
rect 13081 16405 13093 16408
rect 13127 16436 13139 16439
rect 17494 16436 17500 16448
rect 13127 16408 17500 16436
rect 13127 16405 13139 16408
rect 13081 16399 13139 16405
rect 17494 16396 17500 16408
rect 17552 16396 17558 16448
rect 18046 16396 18052 16448
rect 18104 16436 18110 16448
rect 18414 16436 18420 16448
rect 18104 16408 18420 16436
rect 18104 16396 18110 16408
rect 18414 16396 18420 16408
rect 18472 16436 18478 16448
rect 18708 16436 18736 16476
rect 18472 16408 18736 16436
rect 18472 16396 18478 16408
rect 18782 16396 18788 16448
rect 18840 16436 18846 16448
rect 19337 16439 19395 16445
rect 19337 16436 19349 16439
rect 18840 16408 19349 16436
rect 18840 16396 18846 16408
rect 19337 16405 19349 16408
rect 19383 16405 19395 16439
rect 19337 16399 19395 16405
rect 19429 16439 19487 16445
rect 19429 16405 19441 16439
rect 19475 16436 19487 16439
rect 19886 16436 19892 16448
rect 19475 16408 19892 16436
rect 19475 16405 19487 16408
rect 19429 16399 19487 16405
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 21542 16396 21548 16448
rect 21600 16436 21606 16448
rect 22281 16439 22339 16445
rect 22281 16436 22293 16439
rect 21600 16408 22293 16436
rect 21600 16396 21606 16408
rect 22281 16405 22293 16408
rect 22327 16405 22339 16439
rect 22281 16399 22339 16405
rect 1104 16346 23276 16368
rect 1104 16294 4680 16346
rect 4732 16294 4744 16346
rect 4796 16294 4808 16346
rect 4860 16294 4872 16346
rect 4924 16294 12078 16346
rect 12130 16294 12142 16346
rect 12194 16294 12206 16346
rect 12258 16294 12270 16346
rect 12322 16294 19475 16346
rect 19527 16294 19539 16346
rect 19591 16294 19603 16346
rect 19655 16294 19667 16346
rect 19719 16294 23276 16346
rect 1104 16272 23276 16294
rect 1673 16235 1731 16241
rect 1673 16201 1685 16235
rect 1719 16232 1731 16235
rect 2774 16232 2780 16244
rect 1719 16204 2780 16232
rect 1719 16201 1731 16204
rect 1673 16195 1731 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 3418 16232 3424 16244
rect 3379 16204 3424 16232
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 3896 16204 12572 16232
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 15997 1547 16031
rect 1489 15991 1547 15997
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1995 16000 2053 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 3896 16028 3924 16204
rect 5626 16124 5632 16176
rect 5684 16164 5690 16176
rect 5684 16136 6868 16164
rect 5684 16124 5690 16136
rect 3988 16068 4384 16096
rect 3988 16037 4016 16068
rect 2041 15991 2099 15997
rect 2148 16000 3924 16028
rect 3973 16031 4031 16037
rect 1504 15960 1532 15991
rect 2148 15960 2176 16000
rect 3973 15997 3985 16031
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4065 16031 4123 16037
rect 4065 15997 4077 16031
rect 4111 15997 4123 16031
rect 4356 16028 4384 16068
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 6086 16096 6092 16108
rect 4580 16068 4625 16096
rect 4724 16068 6092 16096
rect 4580 16056 4586 16068
rect 4724 16028 4752 16068
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 6362 16096 6368 16108
rect 6196 16068 6368 16096
rect 4356 16000 4752 16028
rect 4801 16031 4859 16037
rect 4065 15991 4123 15997
rect 4801 15997 4813 16031
rect 4847 16028 4859 16031
rect 5718 16028 5724 16040
rect 4847 16000 5724 16028
rect 4847 15997 4859 16000
rect 4801 15991 4859 15997
rect 1504 15932 2176 15960
rect 2308 15963 2366 15969
rect 2308 15929 2320 15963
rect 2354 15960 2366 15963
rect 2682 15960 2688 15972
rect 2354 15932 2688 15960
rect 2354 15929 2366 15932
rect 2308 15923 2366 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 3694 15920 3700 15972
rect 3752 15960 3758 15972
rect 4080 15960 4108 15991
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 6196 16037 6224 16068
rect 6362 16056 6368 16068
rect 6420 16056 6426 16108
rect 6840 16105 6868 16136
rect 10318 16124 10324 16176
rect 10376 16164 10382 16176
rect 12544 16164 12572 16204
rect 12618 16192 12624 16244
rect 12676 16232 12682 16244
rect 17126 16232 17132 16244
rect 12676 16204 17132 16232
rect 12676 16192 12682 16204
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 22741 16235 22799 16241
rect 22741 16232 22753 16235
rect 22612 16204 22753 16232
rect 22612 16192 22618 16204
rect 22741 16201 22753 16204
rect 22787 16201 22799 16235
rect 22741 16195 22799 16201
rect 13262 16164 13268 16176
rect 10376 16136 11652 16164
rect 12544 16136 13268 16164
rect 10376 16124 10382 16136
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 7190 16096 7196 16108
rect 6871 16068 7196 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 7331 16099 7389 16105
rect 7331 16065 7343 16099
rect 7377 16096 7389 16099
rect 7650 16096 7656 16108
rect 7377 16068 7656 16096
rect 7377 16065 7389 16068
rect 7331 16059 7389 16065
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 9264 16099 9322 16105
rect 9264 16096 9276 16099
rect 8211 16068 9276 16096
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 15997 6239 16031
rect 6181 15991 6239 15997
rect 6730 15988 6736 16040
rect 6788 16028 6794 16040
rect 7561 16031 7619 16037
rect 7561 16028 7573 16031
rect 6788 16000 7573 16028
rect 6788 15988 6794 16000
rect 7561 15997 7573 16000
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 3752 15932 4108 15960
rect 3752 15920 3758 15932
rect 1854 15852 1860 15904
rect 1912 15892 1918 15904
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1912 15864 1961 15892
rect 1912 15852 1918 15864
rect 1949 15861 1961 15864
rect 1995 15892 2007 15895
rect 3602 15892 3608 15904
rect 1995 15864 3608 15892
rect 1995 15861 2007 15864
rect 1949 15855 2007 15861
rect 3602 15852 3608 15864
rect 3660 15892 3666 15904
rect 3789 15895 3847 15901
rect 3789 15892 3801 15895
rect 3660 15864 3801 15892
rect 3660 15852 3666 15864
rect 3789 15861 3801 15864
rect 3835 15861 3847 15895
rect 3789 15855 3847 15861
rect 4338 15852 4344 15904
rect 4396 15892 4402 15904
rect 4531 15895 4589 15901
rect 4531 15892 4543 15895
rect 4396 15864 4543 15892
rect 4396 15852 4402 15864
rect 4531 15861 4543 15864
rect 4577 15892 4589 15895
rect 4890 15892 4896 15904
rect 4577 15864 4896 15892
rect 4577 15861 4589 15864
rect 4531 15855 4589 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5905 15895 5963 15901
rect 5905 15892 5917 15895
rect 5224 15864 5917 15892
rect 5224 15852 5230 15864
rect 5905 15861 5917 15864
rect 5951 15861 5963 15895
rect 5905 15855 5963 15861
rect 6270 15852 6276 15904
rect 6328 15892 6334 15904
rect 6365 15895 6423 15901
rect 6365 15892 6377 15895
rect 6328 15864 6377 15892
rect 6328 15852 6334 15864
rect 6365 15861 6377 15864
rect 6411 15861 6423 15895
rect 6365 15855 6423 15861
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 7291 15895 7349 15901
rect 7291 15892 7303 15895
rect 7248 15864 7303 15892
rect 7248 15852 7254 15864
rect 7291 15861 7303 15864
rect 7337 15892 7349 15895
rect 7926 15892 7932 15904
rect 7337 15864 7932 15892
rect 7337 15861 7349 15864
rect 7291 15855 7349 15861
rect 7926 15852 7932 15864
rect 7984 15892 7990 15904
rect 8211 15892 8239 16068
rect 9264 16065 9276 16068
rect 9310 16065 9322 16099
rect 9264 16059 9322 16065
rect 9447 16099 9505 16105
rect 9447 16065 9459 16099
rect 9493 16096 9505 16099
rect 11054 16096 11060 16108
rect 9493 16068 11060 16096
rect 9493 16065 9505 16068
rect 9447 16059 9505 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11624 16105 11652 16136
rect 13262 16124 13268 16136
rect 13320 16124 13326 16176
rect 19429 16167 19487 16173
rect 19429 16133 19441 16167
rect 19475 16164 19487 16167
rect 19702 16164 19708 16176
rect 19475 16136 19708 16164
rect 19475 16133 19487 16136
rect 19429 16127 19487 16133
rect 19702 16124 19708 16136
rect 19760 16124 19766 16176
rect 11609 16099 11667 16105
rect 11609 16065 11621 16099
rect 11655 16065 11667 16099
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 11609 16059 11667 16065
rect 11716 16068 13369 16096
rect 8846 15988 8852 16040
rect 8904 16028 8910 16040
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 8904 16000 8953 16028
rect 8904 15988 8910 16000
rect 8941 15997 8953 16000
rect 8987 15997 8999 16031
rect 9677 16031 9735 16037
rect 9677 16028 9689 16031
rect 8941 15991 8999 15997
rect 9048 16000 9689 16028
rect 9048 15960 9076 16000
rect 9677 15997 9689 16000
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 10686 15988 10692 16040
rect 10744 16028 10750 16040
rect 11716 16028 11744 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13630 16056 13636 16108
rect 13688 16105 13694 16108
rect 13688 16099 13738 16105
rect 13688 16065 13692 16099
rect 13726 16065 13738 16099
rect 13814 16096 13820 16108
rect 13778 16068 13820 16096
rect 13688 16059 13738 16065
rect 13688 16056 13694 16059
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 14274 16096 14280 16108
rect 14016 16068 14280 16096
rect 10744 16000 11744 16028
rect 10744 15988 10750 16000
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 13265 16031 13323 16037
rect 12492 16000 12537 16028
rect 12492 15988 12498 16000
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 14016 16028 14044 16068
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14384 16068 15700 16096
rect 13311 16000 14044 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14384 16028 14412 16068
rect 14148 16000 14412 16028
rect 14148 15988 14154 16000
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 15344 16000 15577 16028
rect 15344 15988 15350 16000
rect 15565 15997 15577 16000
rect 15611 15997 15623 16031
rect 15672 16028 15700 16068
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21361 16099 21419 16105
rect 21361 16096 21373 16099
rect 20956 16068 21373 16096
rect 20956 16056 20962 16068
rect 21361 16065 21373 16068
rect 21407 16065 21419 16099
rect 21361 16059 21419 16065
rect 16758 16028 16764 16040
rect 15672 16000 16764 16028
rect 15565 15991 15623 15997
rect 16758 15988 16764 16000
rect 16816 15988 16822 16040
rect 17221 16031 17279 16037
rect 17221 15997 17233 16031
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 12066 15960 12072 15972
rect 8680 15932 9076 15960
rect 10796 15932 12072 15960
rect 8680 15904 8708 15932
rect 8662 15892 8668 15904
rect 7984 15864 8239 15892
rect 8623 15864 8668 15892
rect 7984 15852 7990 15864
rect 8662 15852 8668 15864
rect 8720 15852 8726 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 10410 15892 10416 15904
rect 8904 15864 10416 15892
rect 8904 15852 8910 15864
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 10796 15901 10824 15932
rect 12066 15920 12072 15932
rect 12124 15920 12130 15972
rect 15810 15963 15868 15969
rect 15810 15960 15822 15963
rect 15028 15932 15822 15960
rect 10781 15895 10839 15901
rect 10781 15861 10793 15895
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 11057 15895 11115 15901
rect 11057 15861 11069 15895
rect 11103 15892 11115 15895
rect 11238 15892 11244 15904
rect 11103 15864 11244 15892
rect 11103 15861 11115 15864
rect 11057 15855 11115 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 11422 15892 11428 15904
rect 11383 15864 11428 15892
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 11517 15895 11575 15901
rect 11517 15861 11529 15895
rect 11563 15892 11575 15895
rect 11698 15892 11704 15904
rect 11563 15864 11704 15892
rect 11563 15861 11575 15864
rect 11517 15855 11575 15861
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 13078 15892 13084 15904
rect 13039 15864 13084 15892
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 13170 15852 13176 15904
rect 13228 15892 13234 15904
rect 15028 15892 15056 15932
rect 15810 15929 15822 15932
rect 15856 15960 15868 15963
rect 16482 15960 16488 15972
rect 15856 15932 16488 15960
rect 15856 15929 15868 15932
rect 15810 15923 15868 15929
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 17236 15960 17264 15991
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17920 16000 18061 16028
rect 17920 15988 17926 16000
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 18095 16000 19717 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 19705 15997 19717 16000
rect 19751 16028 19763 16031
rect 20806 16028 20812 16040
rect 19751 16000 20812 16028
rect 19751 15997 19763 16000
rect 19705 15991 19763 15997
rect 20806 15988 20812 16000
rect 20864 15988 20870 16040
rect 18316 15963 18374 15969
rect 17236 15932 18276 15960
rect 15194 15892 15200 15904
rect 13228 15864 15056 15892
rect 15155 15864 15200 15892
rect 13228 15852 13234 15864
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 16945 15895 17003 15901
rect 16945 15892 16957 15895
rect 16816 15864 16957 15892
rect 16816 15852 16822 15864
rect 16945 15861 16957 15864
rect 16991 15861 17003 15895
rect 16945 15855 17003 15861
rect 17405 15895 17463 15901
rect 17405 15861 17417 15895
rect 17451 15892 17463 15895
rect 17494 15892 17500 15904
rect 17451 15864 17500 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 17494 15852 17500 15864
rect 17552 15852 17558 15904
rect 18248 15892 18276 15932
rect 18316 15929 18328 15963
rect 18362 15960 18374 15963
rect 19334 15960 19340 15972
rect 18362 15932 19340 15960
rect 18362 15929 18374 15932
rect 18316 15923 18374 15929
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 19972 15963 20030 15969
rect 19972 15929 19984 15963
rect 20018 15960 20030 15963
rect 20018 15932 21496 15960
rect 20018 15929 20030 15932
rect 19972 15923 20030 15929
rect 19242 15892 19248 15904
rect 18248 15864 19248 15892
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 20990 15852 20996 15904
rect 21048 15892 21054 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 21048 15864 21097 15892
rect 21048 15852 21054 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21468 15892 21496 15932
rect 21542 15920 21548 15972
rect 21600 15969 21606 15972
rect 21600 15963 21664 15969
rect 21600 15929 21618 15963
rect 21652 15929 21664 15963
rect 21600 15923 21664 15929
rect 21600 15920 21606 15923
rect 22554 15892 22560 15904
rect 21468 15864 22560 15892
rect 21085 15855 21143 15861
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 1104 15802 23276 15824
rect 1104 15750 8379 15802
rect 8431 15750 8443 15802
rect 8495 15750 8507 15802
rect 8559 15750 8571 15802
rect 8623 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 15904 15802
rect 15956 15750 15968 15802
rect 16020 15750 23276 15802
rect 1104 15728 23276 15750
rect 3602 15648 3608 15700
rect 3660 15688 3666 15700
rect 4522 15688 4528 15700
rect 3660 15660 4528 15688
rect 3660 15648 3666 15660
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 4617 15691 4675 15697
rect 4617 15657 4629 15691
rect 4663 15688 4675 15691
rect 8846 15688 8852 15700
rect 4663 15660 8852 15688
rect 4663 15657 4675 15660
rect 4617 15651 4675 15657
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 9122 15688 9128 15700
rect 8956 15660 9128 15688
rect 1854 15620 1860 15632
rect 1504 15592 1860 15620
rect 1504 15561 1532 15592
rect 1854 15580 1860 15592
rect 1912 15580 1918 15632
rect 3694 15580 3700 15632
rect 3752 15620 3758 15632
rect 4706 15620 4712 15632
rect 3752 15592 4712 15620
rect 3752 15580 3758 15592
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15521 1547 15555
rect 1489 15515 1547 15521
rect 1756 15555 1814 15561
rect 1756 15521 1768 15555
rect 1802 15552 1814 15555
rect 2958 15552 2964 15564
rect 1802 15524 2964 15552
rect 1802 15521 1814 15524
rect 1756 15515 1814 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15552 3203 15555
rect 4246 15552 4252 15564
rect 3191 15524 4252 15552
rect 3191 15521 3203 15524
rect 3145 15515 3203 15521
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 3326 15484 3332 15496
rect 3287 15456 3332 15484
rect 3326 15444 3332 15456
rect 3384 15444 3390 15496
rect 4246 15376 4252 15428
rect 4304 15416 4310 15428
rect 4356 15416 4384 15592
rect 4706 15580 4712 15592
rect 4764 15580 4770 15632
rect 8956 15620 8984 15660
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9217 15691 9275 15697
rect 9217 15657 9229 15691
rect 9263 15688 9275 15691
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 9263 15660 10149 15688
rect 9263 15657 9275 15660
rect 9217 15651 9275 15657
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 10137 15651 10195 15657
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 10744 15660 11100 15688
rect 10744 15648 10750 15660
rect 10870 15620 10876 15632
rect 7208 15592 8984 15620
rect 9048 15592 10876 15620
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 4304 15388 4384 15416
rect 4304 15376 4310 15388
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 2869 15351 2927 15357
rect 2869 15348 2881 15351
rect 2740 15320 2881 15348
rect 2740 15308 2746 15320
rect 2869 15317 2881 15320
rect 2915 15317 2927 15351
rect 4448 15348 4476 15515
rect 4890 15512 4896 15564
rect 4948 15552 4954 15564
rect 5308 15555 5366 15561
rect 5308 15552 5320 15555
rect 4948 15524 5320 15552
rect 4948 15512 4954 15524
rect 5308 15521 5320 15524
rect 5354 15521 5366 15555
rect 5308 15515 5366 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 5994 15552 6000 15564
rect 5767 15524 6000 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 6822 15552 6828 15564
rect 6420 15524 6828 15552
rect 6420 15512 6426 15524
rect 6822 15512 6828 15524
rect 6880 15552 6886 15564
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 6880 15524 7113 15552
rect 6880 15512 6886 15524
rect 7101 15521 7113 15524
rect 7147 15521 7159 15555
rect 7101 15515 7159 15521
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 4985 15487 5043 15493
rect 4985 15484 4997 15487
rect 4764 15456 4997 15484
rect 4764 15444 4770 15456
rect 4985 15453 4997 15456
rect 5031 15453 5043 15487
rect 4985 15447 5043 15453
rect 5491 15487 5549 15493
rect 5491 15453 5503 15487
rect 5537 15484 5549 15487
rect 5626 15484 5632 15496
rect 5537 15456 5632 15484
rect 5537 15453 5549 15456
rect 5491 15447 5549 15453
rect 5626 15444 5632 15456
rect 5684 15444 5690 15496
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6917 15487 6975 15493
rect 6917 15484 6929 15487
rect 6144 15456 6929 15484
rect 6144 15444 6150 15456
rect 6917 15453 6929 15456
rect 6963 15453 6975 15487
rect 7208 15484 7236 15592
rect 7374 15561 7380 15564
rect 7368 15552 7380 15561
rect 7335 15524 7380 15552
rect 7368 15515 7380 15524
rect 7374 15512 7380 15515
rect 7432 15512 7438 15564
rect 7926 15512 7932 15564
rect 7984 15552 7990 15564
rect 9048 15561 9076 15592
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 11072 15564 11100 15660
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12584 15660 12909 15688
rect 12584 15648 12590 15660
rect 12897 15657 12909 15660
rect 12943 15688 12955 15691
rect 14090 15688 14096 15700
rect 12943 15660 14096 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 14829 15691 14887 15697
rect 14829 15688 14841 15691
rect 14424 15660 14841 15688
rect 14424 15648 14430 15660
rect 14829 15657 14841 15660
rect 14875 15657 14887 15691
rect 19150 15688 19156 15700
rect 14829 15651 14887 15657
rect 15304 15660 19156 15688
rect 8941 15555 8999 15561
rect 7984 15524 8156 15552
rect 7984 15512 7990 15524
rect 6917 15447 6975 15453
rect 7116 15456 7236 15484
rect 8128 15484 8156 15524
rect 8941 15521 8953 15555
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 9033 15555 9091 15561
rect 9033 15521 9045 15555
rect 9079 15521 9091 15555
rect 9858 15552 9864 15564
rect 9033 15515 9091 15521
rect 9140 15524 9864 15552
rect 8956 15484 8984 15515
rect 9140 15496 9168 15524
rect 9858 15512 9864 15524
rect 9916 15512 9922 15564
rect 10042 15552 10048 15564
rect 10003 15524 10048 15552
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10962 15552 10968 15564
rect 10244 15524 10539 15552
rect 10923 15524 10968 15552
rect 9122 15484 9128 15496
rect 8128 15456 8892 15484
rect 8956 15456 9128 15484
rect 7116 15416 7144 15456
rect 8757 15419 8815 15425
rect 8757 15416 8769 15419
rect 6656 15388 7144 15416
rect 8036 15388 8769 15416
rect 6656 15348 6684 15388
rect 4448 15320 6684 15348
rect 2869 15311 2927 15317
rect 6730 15308 6736 15360
rect 6788 15348 6794 15360
rect 6825 15351 6883 15357
rect 6825 15348 6837 15351
rect 6788 15320 6837 15348
rect 6788 15308 6794 15320
rect 6825 15317 6837 15320
rect 6871 15317 6883 15351
rect 6825 15311 6883 15317
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 8036 15348 8064 15388
rect 8757 15385 8769 15388
rect 8803 15385 8815 15419
rect 8864 15416 8892 15456
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 10244 15484 10272 15524
rect 9600 15456 10272 15484
rect 10321 15487 10379 15493
rect 9600 15416 9628 15456
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10410 15484 10416 15496
rect 10367 15456 10416 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 10511 15484 10539 15524
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11380 15555 11438 15561
rect 11112 15524 11205 15552
rect 11112 15512 11118 15524
rect 11380 15521 11392 15555
rect 11426 15552 11438 15555
rect 11606 15552 11612 15564
rect 11426 15524 11612 15552
rect 11426 15521 11438 15524
rect 11380 15515 11438 15521
rect 11395 15484 11423 15515
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 11793 15555 11851 15561
rect 11793 15521 11805 15555
rect 11839 15552 11851 15555
rect 12066 15552 12072 15564
rect 11839 15524 12072 15552
rect 11839 15521 11851 15524
rect 11793 15515 11851 15521
rect 12066 15512 12072 15524
rect 12124 15552 12130 15564
rect 12124 15524 12480 15552
rect 12124 15512 12130 15524
rect 10511 15456 11423 15484
rect 11520 15487 11578 15493
rect 11520 15453 11532 15487
rect 11566 15484 11578 15487
rect 12250 15484 12256 15496
rect 11566 15456 12256 15484
rect 11566 15453 11578 15456
rect 11520 15447 11578 15453
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 12452 15484 12480 15524
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 13429 15555 13487 15561
rect 13429 15552 13441 15555
rect 13320 15524 13441 15552
rect 13320 15512 13326 15524
rect 13429 15521 13441 15524
rect 13475 15552 13487 15555
rect 15010 15552 15016 15564
rect 13475 15524 14872 15552
rect 14971 15524 15016 15552
rect 13475 15521 13487 15524
rect 13429 15515 13487 15521
rect 12452 15456 12848 15484
rect 8864 15388 9628 15416
rect 9677 15419 9735 15425
rect 8757 15379 8815 15385
rect 9677 15385 9689 15419
rect 9723 15416 9735 15419
rect 9723 15388 11100 15416
rect 9723 15385 9735 15388
rect 9677 15379 9735 15385
rect 8478 15348 8484 15360
rect 6963 15320 8064 15348
rect 8439 15320 8484 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 8478 15308 8484 15320
rect 8536 15308 8542 15360
rect 10594 15308 10600 15360
rect 10652 15348 10658 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10652 15320 10793 15348
rect 10652 15308 10658 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 11072 15348 11100 15388
rect 12710 15348 12716 15360
rect 11072 15320 12716 15348
rect 10781 15311 10839 15317
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 12820 15348 12848 15456
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13173 15487 13231 15493
rect 13173 15484 13185 15487
rect 13136 15456 13185 15484
rect 13136 15444 13142 15456
rect 13173 15453 13185 15456
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 13446 15348 13452 15360
rect 12820 15320 13452 15348
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 14550 15348 14556 15360
rect 14511 15320 14556 15348
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 14844 15348 14872 15524
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15304 15561 15332 15660
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19797 15691 19855 15697
rect 19392 15660 19437 15688
rect 19392 15648 19398 15660
rect 19797 15657 19809 15691
rect 19843 15688 19855 15691
rect 20346 15688 20352 15700
rect 19843 15660 20352 15688
rect 19843 15657 19855 15660
rect 19797 15651 19855 15657
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 19702 15620 19708 15632
rect 17420 15592 19708 15620
rect 15654 15561 15660 15564
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15521 15347 15555
rect 15612 15555 15660 15561
rect 15612 15552 15624 15555
rect 15567 15524 15624 15552
rect 15289 15515 15347 15521
rect 15612 15521 15624 15524
rect 15658 15521 15660 15555
rect 15612 15515 15660 15521
rect 15654 15512 15660 15515
rect 15712 15552 15718 15564
rect 17420 15561 17448 15592
rect 19702 15580 19708 15592
rect 19760 15580 19766 15632
rect 20165 15623 20223 15629
rect 20165 15589 20177 15623
rect 20211 15620 20223 15623
rect 22557 15623 22615 15629
rect 22557 15620 22569 15623
rect 20211 15592 22569 15620
rect 20211 15589 20223 15592
rect 20165 15583 20223 15589
rect 22557 15589 22569 15592
rect 22603 15589 22615 15623
rect 22557 15583 22615 15589
rect 17405 15555 17463 15561
rect 15712 15524 16160 15552
rect 15712 15512 15718 15524
rect 15746 15484 15752 15496
rect 15710 15456 15752 15484
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 16022 15484 16028 15496
rect 15983 15456 16028 15484
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 16132 15484 16160 15524
rect 17405 15521 17417 15555
rect 17451 15521 17463 15555
rect 17405 15515 17463 15521
rect 17862 15512 17868 15564
rect 17920 15552 17926 15564
rect 17957 15555 18015 15561
rect 17957 15552 17969 15555
rect 17920 15524 17969 15552
rect 17920 15512 17926 15524
rect 17957 15521 17969 15524
rect 18003 15521 18015 15555
rect 17957 15515 18015 15521
rect 18046 15512 18052 15564
rect 18104 15552 18110 15564
rect 18213 15555 18271 15561
rect 18213 15552 18225 15555
rect 18104 15524 18225 15552
rect 18104 15512 18110 15524
rect 18213 15521 18225 15524
rect 18259 15521 18271 15555
rect 18213 15515 18271 15521
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 18748 15524 20269 15552
rect 18748 15512 18754 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 20990 15512 20996 15564
rect 21048 15552 21054 15564
rect 21157 15555 21215 15561
rect 21157 15552 21169 15555
rect 21048 15524 21169 15552
rect 21048 15512 21054 15524
rect 21157 15521 21169 15524
rect 21203 15521 21215 15555
rect 21157 15515 21215 15521
rect 20441 15487 20499 15493
rect 16132 15456 17715 15484
rect 16850 15376 16856 15428
rect 16908 15416 16914 15428
rect 17589 15419 17647 15425
rect 17589 15416 17601 15419
rect 16908 15388 17601 15416
rect 16908 15376 16914 15388
rect 17589 15385 17601 15388
rect 17635 15385 17647 15419
rect 17589 15379 17647 15385
rect 16758 15348 16764 15360
rect 14844 15320 16764 15348
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 17126 15348 17132 15360
rect 17087 15320 17132 15348
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 17687 15348 17715 15456
rect 20441 15453 20453 15487
rect 20487 15484 20499 15487
rect 20806 15484 20812 15496
rect 20487 15456 20812 15484
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 20898 15444 20904 15496
rect 20956 15484 20962 15496
rect 20956 15456 21001 15484
rect 20956 15444 20962 15456
rect 19794 15348 19800 15360
rect 17687 15320 19800 15348
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 22281 15351 22339 15357
rect 22281 15348 22293 15351
rect 20864 15320 22293 15348
rect 20864 15308 20870 15320
rect 22281 15317 22293 15320
rect 22327 15317 22339 15351
rect 22281 15311 22339 15317
rect 1104 15258 23276 15280
rect 1104 15206 4680 15258
rect 4732 15206 4744 15258
rect 4796 15206 4808 15258
rect 4860 15206 4872 15258
rect 4924 15206 12078 15258
rect 12130 15206 12142 15258
rect 12194 15206 12206 15258
rect 12258 15206 12270 15258
rect 12322 15206 19475 15258
rect 19527 15206 19539 15258
rect 19591 15206 19603 15258
rect 19655 15206 19667 15258
rect 19719 15206 23276 15258
rect 1104 15184 23276 15206
rect 8846 15144 8852 15156
rect 3620 15116 8852 15144
rect 1854 15008 1860 15020
rect 1815 14980 1860 15008
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 3620 14949 3648 15116
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 8938 15104 8944 15156
rect 8996 15144 9002 15156
rect 8996 15116 10712 15144
rect 8996 15104 9002 15116
rect 3789 15079 3847 15085
rect 3789 15045 3801 15079
rect 3835 15045 3847 15079
rect 3789 15039 3847 15045
rect 3804 15008 3832 15039
rect 4663 15011 4721 15017
rect 4663 15008 4675 15011
rect 3804 14980 4675 15008
rect 4663 14977 4675 14980
rect 4709 15008 4721 15011
rect 4982 15008 4988 15020
rect 4709 14980 4988 15008
rect 4709 14977 4721 14980
rect 4663 14971 4721 14977
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 10684 15008 10712 15116
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12069 15147 12127 15153
rect 12069 15144 12081 15147
rect 12032 15116 12081 15144
rect 12032 15104 12038 15116
rect 12069 15113 12081 15116
rect 12115 15113 12127 15147
rect 12069 15107 12127 15113
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 15010 15144 15016 15156
rect 12492 15116 12537 15144
rect 14971 15116 15016 15144
rect 12492 15104 12498 15116
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15470 15144 15476 15156
rect 15344 15116 15476 15144
rect 15344 15104 15350 15116
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 20990 15144 20996 15156
rect 17604 15116 20996 15144
rect 12618 15036 12624 15088
rect 12676 15076 12682 15088
rect 12676 15048 13492 15076
rect 12676 15036 12682 15048
rect 10684 14980 10815 15008
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14940 4215 14943
rect 4246 14940 4252 14952
rect 4203 14912 4252 14940
rect 4203 14909 4215 14912
rect 4157 14903 4215 14909
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4488 14912 4905 14940
rect 4488 14900 4494 14912
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5166 14940 5172 14952
rect 4939 14912 5172 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7092 14943 7150 14949
rect 7092 14909 7104 14943
rect 7138 14940 7150 14943
rect 8478 14940 8484 14952
rect 7138 14912 8484 14940
rect 7138 14909 7150 14912
rect 7092 14903 7150 14909
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14940 8999 14943
rect 10594 14940 10600 14952
rect 8987 14912 10600 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 10594 14900 10600 14912
rect 10652 14940 10658 14952
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 10652 14912 10701 14940
rect 10652 14900 10658 14912
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10787 14940 10815 14980
rect 12250 14968 12256 15020
rect 12308 15008 12314 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12308 14980 13001 15008
rect 12308 14968 12314 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 13464 15008 13492 15048
rect 14458 15036 14464 15088
rect 14516 15076 14522 15088
rect 14516 15048 17448 15076
rect 14516 15036 14522 15048
rect 17420 15020 17448 15048
rect 13464 14980 13564 15008
rect 12989 14971 13047 14977
rect 10962 14949 10968 14952
rect 10945 14943 10968 14949
rect 10945 14940 10957 14943
rect 10787 14912 10957 14940
rect 10689 14903 10747 14909
rect 10945 14909 10957 14912
rect 11020 14940 11026 14952
rect 11020 14912 11093 14940
rect 10945 14903 10968 14909
rect 10962 14900 10968 14903
rect 11020 14900 11026 14912
rect 12342 14900 12348 14952
rect 12400 14940 12406 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12400 14912 12909 14940
rect 12400 14900 12406 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13136 14912 13461 14940
rect 13136 14900 13142 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13536 14940 13564 14980
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15841 15011 15899 15017
rect 15841 15008 15853 15011
rect 14792 14980 15853 15008
rect 14792 14968 14798 14980
rect 15841 14977 15853 14980
rect 15887 14977 15899 15011
rect 17402 15008 17408 15020
rect 17315 14980 17408 15008
rect 15841 14971 15899 14977
rect 17402 14968 17408 14980
rect 17460 14968 17466 15020
rect 17604 15017 17632 15116
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 21174 15144 21180 15156
rect 21135 15116 21180 15144
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 17678 15036 17684 15088
rect 17736 15076 17742 15088
rect 18322 15076 18328 15088
rect 17736 15048 18328 15076
rect 17736 15036 17742 15048
rect 18322 15036 18328 15048
rect 18380 15036 18386 15088
rect 22649 15079 22707 15085
rect 22649 15076 22661 15079
rect 20732 15048 22661 15076
rect 17589 15011 17647 15017
rect 17589 14977 17601 15011
rect 17635 14977 17647 15011
rect 19843 15011 19901 15017
rect 19843 15008 19855 15011
rect 17589 14971 17647 14977
rect 17972 14980 19855 15008
rect 13705 14943 13763 14949
rect 13705 14940 13717 14943
rect 13536 14912 13717 14940
rect 13449 14903 13507 14909
rect 13705 14909 13717 14912
rect 13751 14940 13763 14943
rect 14550 14940 14556 14952
rect 13751 14912 14556 14940
rect 13751 14909 13763 14912
rect 13705 14903 13763 14909
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14940 15255 14943
rect 16206 14940 16212 14952
rect 15243 14912 16212 14940
rect 15243 14909 15255 14912
rect 15197 14903 15255 14909
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 17313 14943 17371 14949
rect 17313 14909 17325 14943
rect 17359 14940 17371 14943
rect 17972 14940 18000 14980
rect 19843 14977 19855 14980
rect 19889 15008 19901 15011
rect 19978 15008 19984 15020
rect 19889 14980 19984 15008
rect 19889 14977 19901 14980
rect 19843 14971 19901 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20438 14968 20444 15020
rect 20496 15008 20502 15020
rect 20732 15008 20760 15048
rect 22649 15045 22661 15048
rect 22695 15045 22707 15079
rect 22649 15039 22707 15045
rect 20496 14980 20760 15008
rect 20496 14968 20502 14980
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 17359 14912 18000 14940
rect 17359 14909 17371 14912
rect 17313 14903 17371 14909
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18233 14943 18291 14949
rect 18233 14940 18245 14943
rect 18196 14912 18245 14940
rect 18196 14900 18202 14912
rect 18233 14909 18245 14912
rect 18279 14940 18291 14943
rect 18782 14940 18788 14952
rect 18279 14912 18788 14940
rect 18279 14909 18291 14912
rect 18233 14903 18291 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 19150 14900 19156 14952
rect 19208 14940 19214 14952
rect 19337 14943 19395 14949
rect 19337 14940 19349 14943
rect 19208 14912 19349 14940
rect 19208 14900 19214 14912
rect 19337 14909 19349 14912
rect 19383 14940 19395 14943
rect 19426 14940 19432 14952
rect 19383 14912 19432 14940
rect 19383 14909 19395 14912
rect 19337 14903 19395 14909
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 19702 14949 19708 14952
rect 19660 14943 19708 14949
rect 19660 14909 19672 14943
rect 19706 14909 19708 14943
rect 19660 14903 19708 14909
rect 19702 14900 19708 14903
rect 19760 14900 19766 14952
rect 20073 14943 20131 14949
rect 20073 14909 20085 14943
rect 20119 14940 20131 14943
rect 20990 14940 20996 14952
rect 20119 14912 20996 14940
rect 20119 14909 20131 14912
rect 20073 14903 20131 14909
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 22462 14940 22468 14952
rect 22423 14912 22468 14940
rect 22462 14900 22468 14912
rect 22520 14900 22526 14952
rect 2124 14875 2182 14881
rect 2124 14841 2136 14875
rect 2170 14872 2182 14875
rect 3050 14872 3056 14884
rect 2170 14844 3056 14872
rect 2170 14841 2182 14844
rect 2124 14835 2182 14841
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 5810 14832 5816 14884
rect 5868 14872 5874 14884
rect 6273 14875 6331 14881
rect 6273 14872 6285 14875
rect 5868 14844 6285 14872
rect 5868 14832 5874 14844
rect 6273 14841 6285 14844
rect 6319 14841 6331 14875
rect 6273 14835 6331 14841
rect 6362 14832 6368 14884
rect 6420 14872 6426 14884
rect 7282 14872 7288 14884
rect 6420 14844 7288 14872
rect 6420 14832 6426 14844
rect 7282 14832 7288 14844
rect 7340 14832 7346 14884
rect 9208 14875 9266 14881
rect 9208 14841 9220 14875
rect 9254 14872 9266 14875
rect 9674 14872 9680 14884
rect 9254 14844 9680 14872
rect 9254 14841 9266 14844
rect 9208 14835 9266 14841
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 15749 14875 15807 14881
rect 15749 14872 15761 14875
rect 12728 14844 15761 14872
rect 1394 14804 1400 14816
rect 1355 14776 1400 14804
rect 1394 14764 1400 14776
rect 1452 14764 1458 14816
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3237 14807 3295 14813
rect 3237 14804 3249 14807
rect 3016 14776 3249 14804
rect 3016 14764 3022 14776
rect 3237 14773 3249 14776
rect 3283 14804 3295 14807
rect 3694 14804 3700 14816
rect 3283 14776 3700 14804
rect 3283 14773 3295 14776
rect 3237 14767 3295 14773
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 4614 14764 4620 14816
rect 4672 14813 4678 14816
rect 4672 14804 4681 14813
rect 5994 14804 6000 14816
rect 4672 14776 4717 14804
rect 5955 14776 6000 14804
rect 4672 14767 4681 14776
rect 4672 14764 4678 14767
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6086 14764 6092 14816
rect 6144 14804 6150 14816
rect 8018 14804 8024 14816
rect 6144 14776 8024 14804
rect 6144 14764 6150 14776
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 10226 14804 10232 14816
rect 8527 14776 10232 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 10318 14764 10324 14816
rect 10376 14804 10382 14816
rect 11514 14804 11520 14816
rect 10376 14776 11520 14804
rect 10376 14764 10382 14776
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12728 14804 12756 14844
rect 15749 14841 15761 14844
rect 15795 14841 15807 14875
rect 16298 14872 16304 14884
rect 16259 14844 16304 14872
rect 15749 14835 15807 14841
rect 16298 14832 16304 14844
rect 16356 14872 16362 14884
rect 16485 14875 16543 14881
rect 16485 14872 16497 14875
rect 16356 14844 16497 14872
rect 16356 14832 16362 14844
rect 16485 14841 16497 14844
rect 16531 14841 16543 14875
rect 18690 14872 18696 14884
rect 16485 14835 16543 14841
rect 16960 14844 18696 14872
rect 12216 14776 12756 14804
rect 12216 14764 12222 14776
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 14826 14804 14832 14816
rect 12860 14776 12905 14804
rect 14787 14776 14832 14804
rect 12860 14764 12866 14776
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15470 14804 15476 14816
rect 15335 14776 15476 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 16960 14813 16988 14844
rect 18690 14832 18696 14844
rect 18748 14832 18754 14884
rect 18874 14872 18880 14884
rect 18835 14844 18880 14872
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 21542 14872 21548 14884
rect 21100 14844 21548 14872
rect 16945 14807 17003 14813
rect 16945 14773 16957 14807
rect 16991 14773 17003 14807
rect 16945 14767 17003 14773
rect 17678 14764 17684 14816
rect 17736 14804 17742 14816
rect 21100 14804 21128 14844
rect 21542 14832 21548 14844
rect 21600 14832 21606 14884
rect 21450 14804 21456 14816
rect 17736 14776 21128 14804
rect 21411 14776 21456 14804
rect 17736 14764 17742 14776
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 21634 14764 21640 14816
rect 21692 14804 21698 14816
rect 21821 14807 21879 14813
rect 21821 14804 21833 14807
rect 21692 14776 21833 14804
rect 21692 14764 21698 14776
rect 21821 14773 21833 14776
rect 21867 14773 21879 14807
rect 21821 14767 21879 14773
rect 21913 14807 21971 14813
rect 21913 14773 21925 14807
rect 21959 14804 21971 14807
rect 22002 14804 22008 14816
rect 21959 14776 22008 14804
rect 21959 14773 21971 14776
rect 21913 14767 21971 14773
rect 22002 14764 22008 14776
rect 22060 14764 22066 14816
rect 1104 14714 23276 14736
rect 1104 14662 8379 14714
rect 8431 14662 8443 14714
rect 8495 14662 8507 14714
rect 8559 14662 8571 14714
rect 8623 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 15904 14714
rect 15956 14662 15968 14714
rect 16020 14662 23276 14714
rect 1104 14640 23276 14662
rect 1394 14560 1400 14612
rect 1452 14600 1458 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 1452 14572 4445 14600
rect 1452 14560 1458 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4433 14563 4491 14569
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 4571 14572 5089 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 8297 14603 8355 14609
rect 8297 14569 8309 14603
rect 8343 14569 8355 14603
rect 8297 14563 8355 14569
rect 8665 14603 8723 14609
rect 8665 14569 8677 14603
rect 8711 14600 8723 14603
rect 8846 14600 8852 14612
rect 8711 14572 8852 14600
rect 8711 14569 8723 14572
rect 8665 14563 8723 14569
rect 1940 14535 1998 14541
rect 1940 14501 1952 14535
rect 1986 14532 1998 14535
rect 2866 14532 2872 14544
rect 1986 14504 2872 14532
rect 1986 14501 1998 14504
rect 1940 14495 1998 14501
rect 2866 14492 2872 14504
rect 2924 14532 2930 14544
rect 8312 14532 8340 14563
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 9180 14572 9321 14600
rect 9180 14560 9186 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 10318 14600 10324 14612
rect 9309 14563 9367 14569
rect 10143 14572 10324 14600
rect 2924 14504 5672 14532
rect 2924 14492 2930 14504
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14464 1731 14467
rect 1762 14464 1768 14476
rect 1719 14436 1768 14464
rect 1719 14433 1731 14436
rect 1673 14427 1731 14433
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 3418 14464 3424 14476
rect 3379 14436 3424 14464
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 3804 14436 5457 14464
rect 3804 14396 3832 14436
rect 5445 14433 5457 14436
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 5644 14405 5672 14504
rect 5736 14504 8340 14532
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 3620 14368 3832 14396
rect 3896 14368 4629 14396
rect 3050 14328 3056 14340
rect 3011 14300 3056 14328
rect 3050 14288 3056 14300
rect 3108 14288 3114 14340
rect 3620 14337 3648 14368
rect 3605 14331 3663 14337
rect 3605 14297 3617 14331
rect 3651 14297 3663 14331
rect 3605 14291 3663 14297
rect 3068 14260 3096 14288
rect 3896 14260 3924 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 4939 14368 5549 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 4338 14288 4344 14340
rect 4396 14328 4402 14340
rect 5736 14328 5764 14504
rect 8570 14492 8576 14544
rect 8628 14532 8634 14544
rect 10143 14541 10171 14572
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 10928 14572 11529 14600
rect 10928 14560 10934 14572
rect 11517 14569 11529 14572
rect 11563 14569 11575 14603
rect 11517 14563 11575 14569
rect 11885 14603 11943 14609
rect 11885 14569 11897 14603
rect 11931 14600 11943 14603
rect 12434 14600 12440 14612
rect 11931 14572 12440 14600
rect 11931 14569 11943 14572
rect 11885 14563 11943 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 12710 14560 12716 14612
rect 12768 14600 12774 14612
rect 14369 14603 14427 14609
rect 14369 14600 14381 14603
rect 12768 14572 14381 14600
rect 12768 14560 12774 14572
rect 14369 14569 14381 14572
rect 14415 14569 14427 14603
rect 19334 14600 19340 14612
rect 14369 14563 14427 14569
rect 14752 14572 19340 14600
rect 8757 14535 8815 14541
rect 8757 14532 8769 14535
rect 8628 14504 8769 14532
rect 8628 14492 8634 14504
rect 8757 14501 8769 14504
rect 8803 14501 8815 14535
rect 8757 14495 8815 14501
rect 10128 14535 10186 14541
rect 10128 14501 10140 14535
rect 10174 14501 10186 14535
rect 10128 14495 10186 14501
rect 10226 14492 10232 14544
rect 10284 14532 10290 14544
rect 14277 14535 14335 14541
rect 14277 14532 14289 14535
rect 10284 14504 14289 14532
rect 10284 14492 10290 14504
rect 14277 14501 14289 14504
rect 14323 14501 14335 14535
rect 14277 14495 14335 14501
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6897 14467 6955 14473
rect 6897 14464 6909 14467
rect 6196 14436 6909 14464
rect 4396 14300 5764 14328
rect 4396 14288 4402 14300
rect 4062 14260 4068 14272
rect 3068 14232 3924 14260
rect 4023 14232 4068 14260
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4893 14263 4951 14269
rect 4893 14260 4905 14263
rect 4304 14232 4905 14260
rect 4304 14220 4310 14232
rect 4893 14229 4905 14232
rect 4939 14229 4951 14263
rect 4893 14223 4951 14229
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 6196 14260 6224 14436
rect 6897 14433 6909 14436
rect 6943 14464 6955 14467
rect 8202 14464 8208 14476
rect 6943 14436 8208 14464
rect 6943 14433 6955 14436
rect 6897 14427 6955 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 9180 14436 9505 14464
rect 9180 14424 9186 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 10008 14436 11989 14464
rect 10008 14424 10014 14436
rect 11977 14433 11989 14436
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12526 14464 12532 14476
rect 12483 14436 12532 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12704 14467 12762 14473
rect 12704 14433 12716 14467
rect 12750 14464 12762 14467
rect 13630 14464 13636 14476
rect 12750 14436 13636 14464
rect 12750 14433 12762 14436
rect 12704 14427 12762 14433
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14752 14473 14780 14572
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 22002 14600 22008 14612
rect 19628 14572 22008 14600
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 16577 14535 16635 14541
rect 16577 14532 16589 14535
rect 15252 14504 16589 14532
rect 15252 14492 15258 14504
rect 16577 14501 16589 14504
rect 16623 14501 16635 14535
rect 16577 14495 16635 14501
rect 17313 14535 17371 14541
rect 17313 14501 17325 14535
rect 17359 14532 17371 14535
rect 17770 14532 17776 14544
rect 17359 14504 17776 14532
rect 17359 14501 17371 14504
rect 17313 14495 17371 14501
rect 17770 14492 17776 14504
rect 17828 14492 17834 14544
rect 17972 14504 18256 14532
rect 14737 14467 14795 14473
rect 13964 14436 14688 14464
rect 13964 14424 13970 14436
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 8846 14396 8852 14408
rect 8807 14368 8852 14396
rect 6641 14359 6699 14365
rect 6273 14331 6331 14337
rect 6273 14297 6285 14331
rect 6319 14328 6331 14331
rect 6362 14328 6368 14340
rect 6319 14300 6368 14328
rect 6319 14297 6331 14300
rect 6273 14291 6331 14297
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 5040 14232 6224 14260
rect 6656 14260 6684 14359
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 6822 14260 6828 14272
rect 6656 14232 6828 14260
rect 5040 14220 5046 14232
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 8018 14260 8024 14272
rect 7979 14232 8024 14260
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 8846 14260 8852 14272
rect 8628 14232 8852 14260
rect 8628 14220 8634 14232
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9876 14260 9904 14359
rect 10962 14288 10968 14340
rect 11020 14328 11026 14340
rect 11241 14331 11299 14337
rect 11241 14328 11253 14331
rect 11020 14300 11253 14328
rect 11020 14288 11026 14300
rect 11241 14297 11253 14300
rect 11287 14297 11299 14331
rect 12176 14328 12204 14359
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14660 14396 14688 14436
rect 14737 14433 14749 14467
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 15672 14396 15700 14427
rect 15746 14424 15752 14476
rect 15804 14464 15810 14476
rect 16482 14464 16488 14476
rect 15804 14436 15849 14464
rect 16443 14436 16488 14464
rect 15804 14424 15810 14436
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 17405 14467 17463 14473
rect 17405 14433 17417 14467
rect 17451 14464 17463 14467
rect 17972 14464 18000 14504
rect 18046 14473 18052 14476
rect 17451 14436 18000 14464
rect 17451 14433 17463 14436
rect 17405 14427 17463 14433
rect 18040 14427 18052 14473
rect 18104 14464 18110 14476
rect 18228 14464 18256 14504
rect 18322 14492 18328 14544
rect 18380 14532 18386 14544
rect 19628 14532 19656 14572
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 18380 14504 19656 14532
rect 19720 14504 20760 14532
rect 18380 14492 18386 14504
rect 19720 14464 19748 14504
rect 18104 14436 18140 14464
rect 18228 14436 19748 14464
rect 19797 14467 19855 14473
rect 18046 14424 18052 14427
rect 18104 14424 18110 14436
rect 19797 14433 19809 14467
rect 19843 14433 19855 14467
rect 19797 14427 19855 14433
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14464 19947 14467
rect 20625 14467 20683 14473
rect 19935 14436 20484 14464
rect 19935 14433 19947 14436
rect 19889 14427 19947 14433
rect 14516 14368 14561 14396
rect 14660 14368 15700 14396
rect 15841 14399 15899 14405
rect 14516 14356 14522 14368
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 12434 14328 12440 14340
rect 12176 14300 12440 14328
rect 11241 14291 11299 14297
rect 12434 14288 12440 14300
rect 12492 14288 12498 14340
rect 15856 14328 15884 14359
rect 16574 14356 16580 14408
rect 16632 14396 16638 14408
rect 16669 14399 16727 14405
rect 16669 14396 16681 14399
rect 16632 14368 16681 14396
rect 16632 14356 16638 14368
rect 16669 14365 16681 14368
rect 16715 14396 16727 14399
rect 16850 14396 16856 14408
rect 16715 14368 16856 14396
rect 16715 14365 16727 14368
rect 16669 14359 16727 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17589 14399 17647 14405
rect 17589 14365 17601 14399
rect 17635 14396 17647 14399
rect 17678 14396 17684 14408
rect 17635 14368 17684 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 17770 14356 17776 14408
rect 17828 14396 17834 14408
rect 17828 14368 17873 14396
rect 17828 14356 17834 14368
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 19812 14396 19840 14427
rect 20456 14408 20484 14436
rect 20625 14433 20637 14467
rect 20671 14433 20683 14467
rect 20732 14464 20760 14504
rect 20806 14492 20812 14544
rect 20864 14532 20870 14544
rect 21422 14535 21480 14541
rect 21422 14532 21434 14535
rect 20864 14504 21434 14532
rect 20864 14492 20870 14504
rect 21422 14501 21434 14504
rect 21468 14501 21480 14535
rect 21422 14495 21480 14501
rect 20990 14464 20996 14476
rect 20732 14436 20996 14464
rect 20625 14427 20683 14433
rect 19208 14368 19840 14396
rect 19981 14399 20039 14405
rect 19208 14356 19214 14368
rect 19981 14365 19993 14399
rect 20027 14365 20039 14399
rect 19981 14359 20039 14365
rect 13372 14300 15884 14328
rect 16945 14331 17003 14337
rect 10594 14260 10600 14272
rect 9876 14232 10600 14260
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 11514 14220 11520 14272
rect 11572 14260 11578 14272
rect 13372 14260 13400 14300
rect 16945 14297 16957 14331
rect 16991 14328 17003 14331
rect 17402 14328 17408 14340
rect 16991 14300 17408 14328
rect 16991 14297 17003 14300
rect 16945 14291 17003 14297
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 19242 14288 19248 14340
rect 19300 14328 19306 14340
rect 19996 14328 20024 14359
rect 20438 14356 20444 14408
rect 20496 14356 20502 14408
rect 20640 14396 20668 14427
rect 20990 14424 20996 14436
rect 21048 14464 21054 14476
rect 21266 14464 21272 14476
rect 21048 14436 21272 14464
rect 21048 14424 21054 14436
rect 21266 14424 21272 14436
rect 21324 14424 21330 14476
rect 20714 14396 20720 14408
rect 20640 14368 20720 14396
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21177 14399 21235 14405
rect 21177 14396 21189 14399
rect 20956 14368 21189 14396
rect 20956 14356 20962 14368
rect 21177 14365 21189 14368
rect 21223 14365 21235 14399
rect 21177 14359 21235 14365
rect 19300 14300 20024 14328
rect 19300 14288 19306 14300
rect 11572 14232 13400 14260
rect 11572 14220 11578 14232
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13817 14263 13875 14269
rect 13817 14260 13829 14263
rect 13504 14232 13829 14260
rect 13504 14220 13510 14232
rect 13817 14229 13829 14232
rect 13863 14229 13875 14263
rect 13817 14223 13875 14229
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 13964 14232 14009 14260
rect 13964 14220 13970 14232
rect 14734 14220 14740 14272
rect 14792 14260 14798 14272
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 14792 14232 14933 14260
rect 14792 14220 14798 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 14921 14223 14979 14229
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 15160 14232 15301 14260
rect 15160 14220 15166 14232
rect 15289 14229 15301 14232
rect 15335 14229 15347 14263
rect 16114 14260 16120 14272
rect 16075 14232 16120 14260
rect 15289 14223 15347 14229
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 19153 14263 19211 14269
rect 19153 14260 19165 14263
rect 18472 14232 19165 14260
rect 18472 14220 18478 14232
rect 19153 14229 19165 14232
rect 19199 14229 19211 14263
rect 19153 14223 19211 14229
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 19392 14232 19441 14260
rect 19392 14220 19398 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 20441 14263 20499 14269
rect 20441 14229 20453 14263
rect 20487 14260 20499 14263
rect 20898 14260 20904 14272
rect 20487 14232 20904 14260
rect 20487 14229 20499 14232
rect 20441 14223 20499 14229
rect 20898 14220 20904 14232
rect 20956 14220 20962 14272
rect 21910 14220 21916 14272
rect 21968 14260 21974 14272
rect 22557 14263 22615 14269
rect 22557 14260 22569 14263
rect 21968 14232 22569 14260
rect 21968 14220 21974 14232
rect 22557 14229 22569 14232
rect 22603 14229 22615 14263
rect 22557 14223 22615 14229
rect 1104 14170 23276 14192
rect 1104 14118 4680 14170
rect 4732 14118 4744 14170
rect 4796 14118 4808 14170
rect 4860 14118 4872 14170
rect 4924 14118 12078 14170
rect 12130 14118 12142 14170
rect 12194 14118 12206 14170
rect 12258 14118 12270 14170
rect 12322 14118 19475 14170
rect 19527 14118 19539 14170
rect 19591 14118 19603 14170
rect 19655 14118 19667 14170
rect 19719 14118 23276 14170
rect 1104 14096 23276 14118
rect 1762 14056 1768 14068
rect 1504 14028 1768 14056
rect 1504 13929 1532 14028
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 4246 14056 4252 14068
rect 3476 14028 4252 14056
rect 3476 14016 3482 14028
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 6273 14059 6331 14065
rect 6273 14056 6285 14059
rect 4540 14028 6285 14056
rect 1489 13923 1547 13929
rect 1489 13889 1501 13923
rect 1535 13889 1547 13923
rect 3694 13920 3700 13932
rect 3655 13892 3700 13920
rect 1489 13883 1547 13889
rect 3694 13880 3700 13892
rect 3752 13880 3758 13932
rect 1756 13855 1814 13861
rect 1756 13821 1768 13855
rect 1802 13852 1814 13855
rect 4433 13855 4491 13861
rect 4433 13852 4445 13855
rect 1802 13824 4445 13852
rect 1802 13821 1814 13824
rect 1756 13815 1814 13821
rect 4433 13821 4445 13824
rect 4479 13852 4491 13855
rect 4540 13852 4568 14028
rect 6273 14025 6285 14028
rect 6319 14025 6331 14059
rect 6273 14019 6331 14025
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 9858 14056 9864 14068
rect 6871 14028 9864 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10042 14016 10048 14068
rect 10100 14056 10106 14068
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 10100 14028 10149 14056
rect 10100 14016 10106 14028
rect 10137 14025 10149 14028
rect 10183 14025 10195 14059
rect 10137 14019 10195 14025
rect 10689 14059 10747 14065
rect 10689 14025 10701 14059
rect 10735 14056 10747 14059
rect 11422 14056 11428 14068
rect 10735 14028 11428 14056
rect 10735 14025 10747 14028
rect 10689 14019 10747 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12492 14028 12633 14056
rect 12492 14016 12498 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 14458 14056 14464 14068
rect 12621 14019 12679 14025
rect 12820 14028 14464 14056
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 6914 13988 6920 14000
rect 6696 13960 6920 13988
rect 6696 13948 6702 13960
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 9674 13988 9680 14000
rect 9587 13960 9680 13988
rect 9674 13948 9680 13960
rect 9732 13988 9738 14000
rect 12820 13988 12848 14028
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 16114 14016 16120 14068
rect 16172 14056 16178 14068
rect 19150 14056 19156 14068
rect 16172 14028 19156 14056
rect 16172 14016 16178 14028
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 21266 14016 21272 14068
rect 21324 14056 21330 14068
rect 21545 14059 21603 14065
rect 21545 14056 21557 14059
rect 21324 14028 21557 14056
rect 21324 14016 21330 14028
rect 21545 14025 21557 14028
rect 21591 14025 21603 14059
rect 21545 14019 21603 14025
rect 9732 13960 12848 13988
rect 9732 13948 9738 13960
rect 15562 13948 15568 14000
rect 15620 13988 15626 14000
rect 16022 13988 16028 14000
rect 15620 13960 16028 13988
rect 15620 13948 15626 13960
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 21821 13991 21879 13997
rect 21821 13957 21833 13991
rect 21867 13957 21879 13991
rect 21821 13951 21879 13957
rect 4614 13880 4620 13932
rect 4672 13920 4678 13932
rect 4890 13920 4896 13932
rect 4672 13892 4896 13920
rect 4672 13880 4678 13892
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 6420 13892 7389 13920
rect 6420 13880 6426 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 10410 13920 10416 13932
rect 7377 13883 7435 13889
rect 9784 13892 10416 13920
rect 4479 13824 4568 13852
rect 5160 13855 5218 13861
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 5160 13821 5172 13855
rect 5206 13852 5218 13855
rect 5206 13824 5948 13852
rect 5206 13821 5218 13824
rect 5160 13815 5218 13821
rect 5920 13796 5948 13824
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6144 13824 7297 13852
rect 6144 13812 6150 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 8564 13855 8622 13861
rect 8564 13821 8576 13855
rect 8610 13852 8622 13855
rect 9784 13852 9812 13892
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 11333 13923 11391 13929
rect 11333 13889 11345 13923
rect 11379 13889 11391 13923
rect 11333 13883 11391 13889
rect 9950 13852 9956 13864
rect 8610 13824 9812 13852
rect 9911 13824 9956 13852
rect 8610 13821 8622 13824
rect 8564 13815 8622 13821
rect 3513 13787 3571 13793
rect 3513 13753 3525 13787
rect 3559 13784 3571 13787
rect 4062 13784 4068 13796
rect 3559 13756 4068 13784
rect 3559 13753 3571 13756
rect 3513 13747 3571 13753
rect 4062 13744 4068 13756
rect 4120 13744 4126 13796
rect 4246 13784 4252 13796
rect 4207 13756 4252 13784
rect 4246 13744 4252 13756
rect 4304 13744 4310 13796
rect 5902 13744 5908 13796
rect 5960 13784 5966 13796
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 5960 13756 7205 13784
rect 5960 13744 5966 13756
rect 7193 13753 7205 13756
rect 7239 13753 7251 13787
rect 8312 13784 8340 13815
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10134 13812 10140 13864
rect 10192 13852 10198 13864
rect 10318 13852 10324 13864
rect 10192 13824 10324 13852
rect 10192 13812 10198 13824
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 10744 13824 11161 13852
rect 10744 13812 10750 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11348 13852 11376 13883
rect 11422 13880 11428 13932
rect 11480 13920 11486 13932
rect 11882 13920 11888 13932
rect 11480 13892 11888 13920
rect 11480 13880 11486 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12584 13892 12756 13920
rect 12584 13880 12590 13892
rect 12728 13864 12756 13892
rect 17862 13880 17868 13932
rect 17920 13920 17926 13932
rect 18049 13923 18107 13929
rect 18049 13920 18061 13923
rect 17920 13892 18061 13920
rect 17920 13880 17926 13892
rect 18049 13889 18061 13892
rect 18095 13889 18107 13923
rect 18049 13883 18107 13889
rect 11514 13852 11520 13864
rect 11348 13824 11520 13852
rect 11149 13815 11207 13821
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11664 13824 11713 13852
rect 11664 13812 11670 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 12069 13855 12127 13861
rect 12069 13821 12081 13855
rect 12115 13852 12127 13855
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12115 13824 12449 13852
rect 12115 13821 12127 13824
rect 12069 13815 12127 13821
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12768 13824 12817 13852
rect 12768 13812 12774 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 15102 13812 15108 13864
rect 15160 13852 15166 13864
rect 15841 13855 15899 13861
rect 15841 13852 15853 13855
rect 15160 13824 15853 13852
rect 15160 13812 15166 13824
rect 15841 13821 15853 13824
rect 15887 13852 15899 13855
rect 16301 13855 16359 13861
rect 15887 13824 15956 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 7193 13747 7251 13753
rect 7291 13756 8340 13784
rect 3142 13716 3148 13728
rect 3103 13688 3148 13716
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 3605 13719 3663 13725
rect 3605 13685 3617 13719
rect 3651 13716 3663 13719
rect 4430 13716 4436 13728
rect 3651 13688 4436 13716
rect 3651 13685 3663 13688
rect 3605 13679 3663 13685
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 4614 13716 4620 13728
rect 4575 13688 4620 13716
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 7291 13716 7319 13756
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10413 13787 10471 13793
rect 10413 13784 10425 13787
rect 9824 13756 10425 13784
rect 9824 13744 9830 13756
rect 10413 13753 10425 13756
rect 10459 13753 10471 13787
rect 10413 13747 10471 13753
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 11882 13784 11888 13796
rect 10652 13756 11192 13784
rect 11843 13756 11888 13784
rect 10652 13744 10658 13756
rect 7834 13716 7840 13728
rect 6880 13688 7319 13716
rect 7795 13688 7840 13716
rect 6880 13676 6886 13688
rect 7834 13676 7840 13688
rect 7892 13676 7898 13728
rect 8202 13676 8208 13728
rect 8260 13716 8266 13728
rect 10042 13716 10048 13728
rect 8260 13688 10048 13716
rect 8260 13676 8266 13688
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 11054 13716 11060 13728
rect 11015 13688 11060 13716
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 11164 13716 11192 13756
rect 11882 13744 11888 13756
rect 11940 13744 11946 13796
rect 13072 13787 13130 13793
rect 13072 13753 13084 13787
rect 13118 13753 13130 13787
rect 15928 13784 15956 13824
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 18064 13852 18092 13883
rect 19978 13880 19984 13932
rect 20036 13929 20042 13932
rect 20036 13923 20086 13929
rect 20036 13889 20040 13923
rect 20074 13889 20086 13923
rect 20036 13883 20086 13889
rect 20211 13923 20269 13929
rect 20211 13889 20223 13923
rect 20257 13920 20269 13923
rect 21836 13920 21864 13951
rect 20257 13892 21864 13920
rect 22465 13923 22523 13929
rect 20257 13889 20269 13892
rect 20211 13883 20269 13889
rect 22465 13889 22477 13923
rect 22511 13920 22523 13923
rect 22830 13920 22836 13932
rect 22511 13892 22836 13920
rect 22511 13889 22523 13892
rect 22465 13883 22523 13889
rect 20036 13880 20042 13883
rect 22830 13880 22836 13892
rect 22888 13880 22894 13932
rect 18690 13852 18696 13864
rect 16347 13824 18696 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19208 13824 19717 13852
rect 19208 13812 19214 13824
rect 19705 13821 19717 13824
rect 19751 13852 19763 13855
rect 19794 13852 19800 13864
rect 19751 13824 19800 13852
rect 19751 13821 19763 13824
rect 19705 13815 19763 13821
rect 19794 13812 19800 13824
rect 19852 13812 19858 13864
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13852 20499 13855
rect 20487 13824 21404 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 16025 13787 16083 13793
rect 16025 13784 16037 13787
rect 15928 13756 16037 13784
rect 13072 13747 13130 13753
rect 16025 13753 16037 13756
rect 16071 13753 16083 13787
rect 16025 13747 16083 13753
rect 16568 13787 16626 13793
rect 16568 13753 16580 13787
rect 16614 13784 16626 13787
rect 17862 13784 17868 13796
rect 16614 13756 17868 13784
rect 16614 13753 16626 13756
rect 16568 13747 16626 13753
rect 12158 13716 12164 13728
rect 11164 13688 12164 13716
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 12977 13676 12983 13728
rect 13035 13716 13041 13728
rect 13087 13716 13115 13747
rect 17862 13744 17868 13756
rect 17920 13744 17926 13796
rect 18322 13793 18328 13796
rect 18294 13787 18328 13793
rect 18294 13784 18306 13787
rect 17972 13756 18306 13784
rect 13035 13688 13115 13716
rect 13035 13676 13041 13688
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14185 13719 14243 13725
rect 14185 13716 14197 13719
rect 13872 13688 14197 13716
rect 13872 13676 13878 13688
rect 14185 13685 14197 13688
rect 14231 13685 14243 13719
rect 14185 13679 14243 13685
rect 15289 13719 15347 13725
rect 15289 13685 15301 13719
rect 15335 13716 15347 13719
rect 16758 13716 16764 13728
rect 15335 13688 16764 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 17681 13719 17739 13725
rect 17681 13685 17693 13719
rect 17727 13716 17739 13719
rect 17972 13716 18000 13756
rect 18294 13753 18306 13756
rect 18380 13784 18386 13796
rect 21376 13784 21404 13824
rect 21450 13812 21456 13864
rect 21508 13852 21514 13864
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 21508 13824 22293 13852
rect 21508 13812 21514 13824
rect 22281 13821 22293 13824
rect 22327 13821 22339 13855
rect 22281 13815 22339 13821
rect 21634 13784 21640 13796
rect 18380 13756 18442 13784
rect 21376 13756 21640 13784
rect 18294 13747 18328 13753
rect 18322 13744 18328 13747
rect 18380 13744 18386 13756
rect 21634 13744 21640 13756
rect 21692 13744 21698 13796
rect 17727 13688 18000 13716
rect 17727 13685 17739 13688
rect 17681 13679 17739 13685
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18966 13716 18972 13728
rect 18104 13688 18972 13716
rect 18104 13676 18110 13688
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 19429 13719 19487 13725
rect 19429 13685 19441 13719
rect 19475 13716 19487 13719
rect 19702 13716 19708 13728
rect 19475 13688 19708 13716
rect 19475 13685 19487 13688
rect 19429 13679 19487 13685
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20530 13716 20536 13728
rect 20036 13688 20536 13716
rect 20036 13676 20042 13688
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 22186 13716 22192 13728
rect 22147 13688 22192 13716
rect 22186 13676 22192 13688
rect 22244 13676 22250 13728
rect 1104 13626 23276 13648
rect 1104 13574 8379 13626
rect 8431 13574 8443 13626
rect 8495 13574 8507 13626
rect 8559 13574 8571 13626
rect 8623 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 15904 13626
rect 15956 13574 15968 13626
rect 16020 13574 23276 13626
rect 1104 13552 23276 13574
rect 1854 13512 1860 13524
rect 1815 13484 1860 13512
rect 1854 13472 1860 13484
rect 1912 13472 1918 13524
rect 2685 13515 2743 13521
rect 2685 13481 2697 13515
rect 2731 13512 2743 13515
rect 3142 13512 3148 13524
rect 2731 13484 3148 13512
rect 2731 13481 2743 13484
rect 2685 13475 2743 13481
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 4065 13515 4123 13521
rect 4065 13481 4077 13515
rect 4111 13512 4123 13515
rect 4154 13512 4160 13524
rect 4111 13484 4160 13512
rect 4111 13481 4123 13484
rect 4065 13475 4123 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 5902 13512 5908 13524
rect 5863 13484 5908 13512
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 6411 13484 10149 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 10137 13481 10149 13484
rect 10183 13481 10195 13515
rect 10137 13475 10195 13481
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10468 13484 11192 13512
rect 10468 13472 10474 13484
rect 4614 13444 4620 13456
rect 1688 13416 4620 13444
rect 1688 13385 1716 13416
rect 4614 13404 4620 13416
rect 4672 13404 4678 13456
rect 4792 13447 4850 13453
rect 4792 13413 4804 13447
rect 4838 13444 4850 13447
rect 5534 13444 5540 13456
rect 4838 13416 5540 13444
rect 4838 13413 4850 13416
rect 4792 13407 4850 13413
rect 5534 13404 5540 13416
rect 5592 13444 5598 13456
rect 6086 13444 6092 13456
rect 5592 13416 6092 13444
rect 5592 13404 5598 13416
rect 6086 13404 6092 13416
rect 6144 13404 6150 13456
rect 6638 13444 6644 13456
rect 6196 13416 6644 13444
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13345 1731 13379
rect 2590 13376 2596 13388
rect 2551 13348 2596 13376
rect 1673 13339 1731 13345
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 6196 13385 6224 13416
rect 6638 13404 6644 13416
rect 6696 13404 6702 13456
rect 6894 13444 6900 13456
rect 6748 13416 6900 13444
rect 6748 13385 6776 13416
rect 6894 13404 6900 13416
rect 6952 13404 6958 13456
rect 7000 13447 7058 13453
rect 7000 13413 7012 13447
rect 7046 13444 7058 13447
rect 7558 13444 7564 13456
rect 7046 13416 7564 13444
rect 7046 13413 7058 13416
rect 7000 13407 7058 13413
rect 7558 13404 7564 13416
rect 7616 13444 7622 13456
rect 8018 13444 8024 13456
rect 7616 13416 8024 13444
rect 7616 13404 7622 13416
rect 8018 13404 8024 13416
rect 8076 13404 8082 13456
rect 8110 13404 8116 13456
rect 8168 13444 8174 13456
rect 8570 13444 8576 13456
rect 8168 13416 8576 13444
rect 8168 13404 8174 13416
rect 8570 13404 8576 13416
rect 8628 13444 8634 13456
rect 8628 13416 8892 13444
rect 8628 13404 8634 13416
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13376 3479 13379
rect 6181 13379 6239 13385
rect 3467 13348 6132 13376
rect 3467 13345 3479 13348
rect 3421 13339 3479 13345
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 2740 13280 2789 13308
rect 2740 13268 2746 13280
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 3970 13308 3976 13320
rect 2777 13271 2835 13277
rect 3160 13280 3976 13308
rect 2225 13243 2283 13249
rect 2225 13209 2237 13243
rect 2271 13240 2283 13243
rect 3160 13240 3188 13280
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 4522 13308 4528 13320
rect 4483 13280 4528 13308
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 6104 13308 6132 13348
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 6840 13348 7880 13376
rect 6840 13308 6868 13348
rect 6104 13280 6868 13308
rect 2271 13212 3188 13240
rect 2271 13209 2283 13212
rect 2225 13203 2283 13209
rect 3234 13200 3240 13252
rect 3292 13240 3298 13252
rect 3510 13240 3516 13252
rect 3292 13212 3516 13240
rect 3292 13200 3298 13212
rect 3510 13200 3516 13212
rect 3568 13200 3574 13252
rect 7852 13240 7880 13348
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8757 13379 8815 13385
rect 8757 13376 8769 13379
rect 7984 13348 8769 13376
rect 7984 13336 7990 13348
rect 8757 13345 8769 13348
rect 8803 13345 8815 13379
rect 8864 13376 8892 13416
rect 11054 13404 11060 13456
rect 11112 13404 11118 13456
rect 11164 13444 11192 13484
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11940 13484 12081 13512
rect 11940 13472 11946 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 16574 13512 16580 13524
rect 12069 13475 12127 13481
rect 15212 13484 16580 13512
rect 12084 13444 12112 13475
rect 11164 13416 12020 13444
rect 12084 13416 12296 13444
rect 10042 13376 10048 13388
rect 8864 13348 8984 13376
rect 10003 13348 10048 13376
rect 8757 13339 8815 13345
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8956 13317 8984 13348
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 10956 13379 11014 13385
rect 10956 13345 10968 13379
rect 11002 13376 11014 13379
rect 11072 13376 11100 13404
rect 11790 13376 11796 13388
rect 11002 13348 11796 13376
rect 11002 13345 11014 13348
rect 10956 13339 11014 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 8849 13311 8907 13317
rect 8849 13308 8861 13311
rect 8076 13280 8861 13308
rect 8076 13268 8082 13280
rect 8849 13277 8861 13280
rect 8895 13277 8907 13311
rect 8849 13271 8907 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 9490 13240 9496 13252
rect 7852 13212 9496 13240
rect 9490 13200 9496 13212
rect 9548 13200 9554 13252
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 9950 13240 9956 13252
rect 9723 13212 9956 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 3605 13175 3663 13181
rect 3605 13141 3617 13175
rect 3651 13172 3663 13175
rect 7926 13172 7932 13184
rect 3651 13144 7932 13172
rect 3651 13141 3663 13144
rect 3605 13135 3663 13141
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 8110 13172 8116 13184
rect 8071 13144 8116 13172
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8389 13175 8447 13181
rect 8389 13141 8401 13175
rect 8435 13172 8447 13175
rect 8938 13172 8944 13184
rect 8435 13144 8944 13172
rect 8435 13141 8447 13144
rect 8389 13135 8447 13141
rect 8938 13132 8944 13144
rect 8996 13132 9002 13184
rect 10336 13172 10364 13271
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 10468 13280 10701 13308
rect 10468 13268 10474 13280
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 11422 13172 11428 13184
rect 10336 13144 11428 13172
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11992 13172 12020 13416
rect 12158 13376 12164 13388
rect 12119 13348 12164 13376
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 12268 13376 12296 13416
rect 12710 13404 12716 13456
rect 12768 13444 12774 13456
rect 13078 13444 13084 13456
rect 12768 13416 13084 13444
rect 12768 13404 12774 13416
rect 13078 13404 13084 13416
rect 13136 13444 13142 13456
rect 13136 13416 13676 13444
rect 13136 13404 13142 13416
rect 13648 13385 13676 13416
rect 13814 13404 13820 13456
rect 13872 13453 13878 13456
rect 13872 13447 13936 13453
rect 13872 13413 13890 13447
rect 13924 13413 13936 13447
rect 13872 13407 13936 13413
rect 13872 13404 13878 13407
rect 14918 13404 14924 13456
rect 14976 13444 14982 13456
rect 15212 13444 15240 13484
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 19705 13515 19763 13521
rect 19705 13512 19717 13515
rect 17460 13484 19717 13512
rect 17460 13472 17466 13484
rect 19705 13481 19717 13484
rect 19751 13481 19763 13515
rect 19705 13475 19763 13481
rect 19978 13472 19984 13524
rect 20036 13512 20042 13524
rect 20346 13512 20352 13524
rect 20036 13484 20352 13512
rect 20036 13472 20042 13484
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 20901 13515 20959 13521
rect 20901 13481 20913 13515
rect 20947 13512 20959 13515
rect 22186 13512 22192 13524
rect 20947 13484 22192 13512
rect 20947 13481 20959 13484
rect 20901 13475 20959 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 18500 13447 18558 13453
rect 14976 13416 15240 13444
rect 15304 13416 16804 13444
rect 14976 13404 14982 13416
rect 12417 13379 12475 13385
rect 12417 13376 12429 13379
rect 12268 13348 12429 13376
rect 12417 13345 12429 13348
rect 12463 13345 12475 13379
rect 12417 13339 12475 13345
rect 13633 13379 13691 13385
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 15102 13376 15108 13388
rect 13679 13348 15108 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 15102 13336 15108 13348
rect 15160 13376 15166 13388
rect 15304 13385 15332 13416
rect 16776 13385 16804 13416
rect 18500 13413 18512 13447
rect 18546 13444 18558 13447
rect 21628 13447 21686 13453
rect 18546 13416 19748 13444
rect 18546 13413 18558 13416
rect 18500 13407 18558 13413
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 15160 13348 15301 13376
rect 15160 13336 15166 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15545 13379 15603 13385
rect 15545 13376 15557 13379
rect 15289 13339 15347 13345
rect 15387 13348 15557 13376
rect 15387 13308 15415 13348
rect 15545 13345 15557 13348
rect 15591 13345 15603 13379
rect 15545 13339 15603 13345
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13345 16819 13379
rect 16761 13339 16819 13345
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 17017 13379 17075 13385
rect 17017 13376 17029 13379
rect 16908 13348 17029 13376
rect 16908 13336 16914 13348
rect 17017 13345 17029 13348
rect 17063 13345 17075 13379
rect 17017 13339 17075 13345
rect 17770 13336 17776 13388
rect 17828 13376 17834 13388
rect 18233 13379 18291 13385
rect 18233 13376 18245 13379
rect 17828 13348 18245 13376
rect 17828 13336 17834 13348
rect 18233 13345 18245 13348
rect 18279 13345 18291 13379
rect 18233 13339 18291 13345
rect 18966 13336 18972 13388
rect 19024 13376 19030 13388
rect 19024 13348 19656 13376
rect 19024 13336 19030 13348
rect 15028 13280 15415 13308
rect 15028 13184 15056 13280
rect 17770 13200 17776 13252
rect 17828 13240 17834 13252
rect 18141 13243 18199 13249
rect 18141 13240 18153 13243
rect 17828 13212 18153 13240
rect 17828 13200 17834 13212
rect 18141 13209 18153 13212
rect 18187 13209 18199 13243
rect 18141 13203 18199 13209
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 11992 13144 13553 13172
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 15010 13172 15016 13184
rect 14971 13144 15016 13172
rect 13541 13135 13599 13141
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 16669 13175 16727 13181
rect 16669 13172 16681 13175
rect 15620 13144 16681 13172
rect 15620 13132 15626 13144
rect 16669 13141 16681 13144
rect 16715 13141 16727 13175
rect 16669 13135 16727 13141
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 18874 13172 18880 13184
rect 16816 13144 18880 13172
rect 16816 13132 16822 13144
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19628 13181 19656 13348
rect 19720 13320 19748 13416
rect 21628 13413 21640 13447
rect 21674 13444 21686 13447
rect 21910 13444 21916 13456
rect 21674 13416 21916 13444
rect 21674 13413 21686 13416
rect 21628 13407 21686 13413
rect 21910 13404 21916 13416
rect 21968 13404 21974 13456
rect 19794 13336 19800 13388
rect 19852 13376 19858 13388
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 19852 13348 20085 13376
rect 19852 13336 19858 13348
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 20165 13379 20223 13385
rect 20165 13345 20177 13379
rect 20211 13376 20223 13379
rect 20346 13376 20352 13388
rect 20211 13348 20352 13376
rect 20211 13345 20223 13348
rect 20165 13339 20223 13345
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 19702 13268 19708 13320
rect 19760 13308 19766 13320
rect 20257 13311 20315 13317
rect 20257 13308 20269 13311
rect 19760 13280 20269 13308
rect 19760 13268 19766 13280
rect 20257 13277 20269 13280
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 20898 13268 20904 13320
rect 20956 13308 20962 13320
rect 21361 13311 21419 13317
rect 21361 13308 21373 13311
rect 20956 13280 21373 13308
rect 20956 13268 20962 13280
rect 21361 13277 21373 13280
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 19613 13175 19671 13181
rect 19613 13141 19625 13175
rect 19659 13141 19671 13175
rect 19613 13135 19671 13141
rect 22741 13175 22799 13181
rect 22741 13141 22753 13175
rect 22787 13172 22799 13175
rect 22830 13172 22836 13184
rect 22787 13144 22836 13172
rect 22787 13141 22799 13144
rect 22741 13135 22799 13141
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 1104 13082 23276 13104
rect 1104 13030 4680 13082
rect 4732 13030 4744 13082
rect 4796 13030 4808 13082
rect 4860 13030 4872 13082
rect 4924 13030 12078 13082
rect 12130 13030 12142 13082
rect 12194 13030 12206 13082
rect 12258 13030 12270 13082
rect 12322 13030 19475 13082
rect 19527 13030 19539 13082
rect 19591 13030 19603 13082
rect 19655 13030 19667 13082
rect 19719 13030 23276 13082
rect 1104 13008 23276 13030
rect 5353 12971 5411 12977
rect 2056 12940 3648 12968
rect 1670 12900 1676 12912
rect 1631 12872 1676 12900
rect 1670 12860 1676 12872
rect 1728 12860 1734 12912
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12733 1547 12767
rect 1489 12727 1547 12733
rect 1504 12696 1532 12727
rect 1578 12724 1584 12776
rect 1636 12764 1642 12776
rect 2056 12773 2084 12940
rect 3620 12832 3648 12940
rect 5353 12937 5365 12971
rect 5399 12968 5411 12971
rect 9490 12968 9496 12980
rect 5399 12940 9168 12968
rect 9451 12940 9496 12968
rect 5399 12937 5411 12940
rect 5353 12931 5411 12937
rect 5077 12903 5135 12909
rect 5077 12869 5089 12903
rect 5123 12900 5135 12903
rect 5534 12900 5540 12912
rect 5123 12872 5540 12900
rect 5123 12869 5135 12872
rect 5077 12863 5135 12869
rect 5534 12860 5540 12872
rect 5592 12860 5598 12912
rect 8481 12903 8539 12909
rect 8481 12869 8493 12903
rect 8527 12900 8539 12903
rect 8846 12900 8852 12912
rect 8527 12872 8852 12900
rect 8527 12869 8539 12872
rect 8481 12863 8539 12869
rect 8846 12860 8852 12872
rect 8904 12860 8910 12912
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3620 12804 3709 12832
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 2041 12767 2099 12773
rect 2041 12764 2053 12767
rect 1636 12736 2053 12764
rect 1636 12724 1642 12736
rect 2041 12733 2053 12736
rect 2087 12733 2099 12767
rect 2041 12727 2099 12733
rect 2308 12767 2366 12773
rect 2308 12733 2320 12767
rect 2354 12764 2366 12767
rect 2682 12764 2688 12776
rect 2354 12736 2688 12764
rect 2354 12733 2366 12736
rect 2308 12727 2366 12733
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 3712 12764 3740 12795
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 5997 12835 6055 12841
rect 5997 12832 6009 12835
rect 5776 12804 6009 12832
rect 5776 12792 5782 12804
rect 5997 12801 6009 12804
rect 6043 12832 6055 12835
rect 6362 12832 6368 12844
rect 6043 12804 6368 12832
rect 6043 12801 6055 12804
rect 5997 12795 6055 12801
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 7892 12804 8248 12832
rect 7892 12792 7898 12804
rect 4890 12764 4896 12776
rect 3712 12736 4896 12764
rect 4890 12724 4896 12736
rect 4948 12764 4954 12776
rect 6822 12764 6828 12776
rect 4948 12736 6828 12764
rect 4948 12724 4954 12736
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7092 12767 7150 12773
rect 7092 12733 7104 12767
rect 7138 12764 7150 12767
rect 8110 12764 8116 12776
rect 7138 12736 8116 12764
rect 7138 12733 7150 12736
rect 7092 12727 7150 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8220 12764 8248 12804
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8628 12804 9045 12832
rect 8628 12792 8634 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9140 12832 9168 12940
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13262 12968 13268 12980
rect 12636 12940 13268 12968
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 9140 12804 9965 12832
rect 9033 12795 9091 12801
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 10045 12795 10103 12801
rect 8220 12736 8708 12764
rect 2866 12696 2872 12708
rect 1504 12668 2872 12696
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 3964 12699 4022 12705
rect 3964 12696 3976 12699
rect 3436 12668 3976 12696
rect 3436 12637 3464 12668
rect 3964 12665 3976 12668
rect 4010 12696 4022 12699
rect 5721 12699 5779 12705
rect 5721 12696 5733 12699
rect 4010 12668 5733 12696
rect 4010 12665 4022 12668
rect 3964 12659 4022 12665
rect 5721 12665 5733 12668
rect 5767 12665 5779 12699
rect 8680 12696 8708 12736
rect 9214 12724 9220 12776
rect 9272 12764 9278 12776
rect 9490 12764 9496 12776
rect 9272 12736 9496 12764
rect 9272 12724 9278 12736
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 9858 12764 9864 12776
rect 9819 12736 9864 12764
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 10060 12696 10088 12795
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 12636 12832 12664 12940
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 16577 12971 16635 12977
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 16850 12968 16856 12980
rect 16623 12940 16856 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 18966 12968 18972 12980
rect 17604 12940 18972 12968
rect 13630 12860 13636 12912
rect 13688 12900 13694 12912
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 13688 12872 14013 12900
rect 13688 12860 13694 12872
rect 14001 12869 14013 12872
rect 14047 12869 14059 12903
rect 14001 12863 14059 12869
rect 14185 12903 14243 12909
rect 14185 12869 14197 12903
rect 14231 12900 14243 12903
rect 14458 12900 14464 12912
rect 14231 12872 14464 12900
rect 14231 12869 14243 12872
rect 14185 12863 14243 12869
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 11664 12804 12664 12832
rect 14829 12835 14887 12841
rect 11664 12792 11670 12804
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 14918 12832 14924 12844
rect 14875 12804 14924 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 15102 12792 15108 12844
rect 15160 12832 15166 12844
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 15160 12804 15209 12832
rect 15160 12792 15166 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 17402 12832 17408 12844
rect 17363 12804 17408 12832
rect 15197 12795 15255 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 17604 12841 17632 12940
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 20622 12928 20628 12980
rect 20680 12968 20686 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 20680 12940 22385 12968
rect 20680 12928 20686 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22373 12931 22431 12937
rect 19702 12860 19708 12912
rect 19760 12900 19766 12912
rect 20533 12903 20591 12909
rect 20533 12900 20545 12903
rect 19760 12872 20545 12900
rect 19760 12860 19766 12872
rect 20533 12869 20545 12872
rect 20579 12869 20591 12903
rect 20533 12863 20591 12869
rect 21177 12903 21235 12909
rect 21177 12869 21189 12903
rect 21223 12900 21235 12903
rect 22278 12900 22284 12912
rect 21223 12872 22284 12900
rect 21223 12869 21235 12872
rect 21177 12863 21235 12869
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 21634 12832 21640 12844
rect 17589 12795 17647 12801
rect 17687 12804 18828 12832
rect 21595 12804 21640 12832
rect 10686 12773 10692 12776
rect 10680 12764 10692 12773
rect 10647 12736 10692 12764
rect 10680 12727 10692 12736
rect 10686 12724 10692 12727
rect 10744 12724 10750 12776
rect 12253 12767 12311 12773
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12764 12679 12767
rect 12710 12764 12716 12776
rect 12667 12736 12716 12764
rect 12667 12733 12679 12736
rect 12621 12727 12679 12733
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 12888 12767 12946 12773
rect 12888 12733 12900 12767
rect 12934 12764 12946 12767
rect 13446 12764 13452 12776
rect 12934 12736 13452 12764
rect 12934 12733 12946 12736
rect 12888 12727 12946 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 17687 12764 17715 12804
rect 18046 12764 18052 12776
rect 13556 12736 17715 12764
rect 18007 12736 18052 12764
rect 8680 12668 10088 12696
rect 5721 12659 5779 12665
rect 10318 12656 10324 12708
rect 10376 12696 10382 12708
rect 11238 12696 11244 12708
rect 10376 12668 11244 12696
rect 10376 12656 10382 12668
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 11422 12656 11428 12708
rect 11480 12696 11486 12708
rect 13556 12696 13584 12736
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12764 18291 12767
rect 18322 12764 18328 12776
rect 18279 12736 18328 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 18322 12724 18328 12736
rect 18380 12724 18386 12776
rect 18690 12764 18696 12776
rect 18651 12736 18696 12764
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 18800 12764 18828 12804
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12832 21879 12835
rect 22094 12832 22100 12844
rect 21867 12804 22100 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 20349 12767 20407 12773
rect 20349 12764 20361 12767
rect 18800 12736 20361 12764
rect 20349 12733 20361 12736
rect 20395 12733 20407 12767
rect 20349 12727 20407 12733
rect 21726 12724 21732 12776
rect 21784 12764 21790 12776
rect 21910 12764 21916 12776
rect 21784 12736 21916 12764
rect 21784 12724 21790 12736
rect 21910 12724 21916 12736
rect 21968 12724 21974 12776
rect 22189 12767 22247 12773
rect 22189 12733 22201 12767
rect 22235 12764 22247 12767
rect 22370 12764 22376 12776
rect 22235 12736 22376 12764
rect 22235 12733 22247 12736
rect 22189 12727 22247 12733
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 11480 12668 13584 12696
rect 15464 12699 15522 12705
rect 11480 12656 11486 12668
rect 15464 12665 15476 12699
rect 15510 12696 15522 12699
rect 15562 12696 15568 12708
rect 15510 12668 15568 12696
rect 15510 12665 15522 12668
rect 15464 12659 15522 12665
rect 15562 12656 15568 12668
rect 15620 12656 15626 12708
rect 17770 12696 17776 12708
rect 16960 12668 17776 12696
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12597 3479 12631
rect 3421 12591 3479 12597
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 5813 12631 5871 12637
rect 5813 12628 5825 12631
rect 4120 12600 5825 12628
rect 4120 12588 4126 12600
rect 5813 12597 5825 12600
rect 5859 12597 5871 12631
rect 5813 12591 5871 12597
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 8076 12600 8217 12628
rect 8076 12588 8082 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8205 12591 8263 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 8996 12600 9041 12628
rect 8996 12588 9002 12600
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 11112 12600 12081 12628
rect 11112 12588 11118 12600
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 12069 12591 12127 12597
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 13630 12628 13636 12640
rect 13320 12600 13636 12628
rect 13320 12588 13326 12600
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 14550 12628 14556 12640
rect 14511 12600 14556 12628
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 14645 12631 14703 12637
rect 14645 12597 14657 12631
rect 14691 12628 14703 12631
rect 16758 12628 16764 12640
rect 14691 12600 16764 12628
rect 14691 12597 14703 12600
rect 14645 12591 14703 12597
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 16960 12637 16988 12668
rect 17770 12656 17776 12668
rect 17828 12656 17834 12708
rect 18966 12705 18972 12708
rect 18960 12696 18972 12705
rect 18927 12668 18972 12696
rect 18960 12659 18972 12668
rect 18966 12656 18972 12659
rect 19024 12656 19030 12708
rect 20806 12696 20812 12708
rect 19076 12668 20812 12696
rect 16945 12631 17003 12637
rect 16945 12597 16957 12631
rect 16991 12597 17003 12631
rect 16945 12591 17003 12597
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 17276 12600 17325 12628
rect 17276 12588 17282 12600
rect 17313 12597 17325 12600
rect 17359 12597 17371 12631
rect 18414 12628 18420 12640
rect 18375 12600 18420 12628
rect 17313 12591 17371 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 19076 12628 19104 12668
rect 20806 12656 20812 12668
rect 20864 12656 20870 12708
rect 18932 12600 19104 12628
rect 18932 12588 18938 12600
rect 19702 12588 19708 12640
rect 19760 12628 19766 12640
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 19760 12600 20085 12628
rect 19760 12588 19766 12600
rect 20073 12597 20085 12600
rect 20119 12597 20131 12631
rect 21542 12628 21548 12640
rect 21503 12600 21548 12628
rect 20073 12591 20131 12597
rect 21542 12588 21548 12600
rect 21600 12588 21606 12640
rect 1104 12538 23276 12560
rect 1104 12486 8379 12538
rect 8431 12486 8443 12538
rect 8495 12486 8507 12538
rect 8559 12486 8571 12538
rect 8623 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 15904 12538
rect 15956 12486 15968 12538
rect 16020 12486 23276 12538
rect 1104 12464 23276 12486
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 3660 12396 3705 12424
rect 3660 12384 3666 12396
rect 4890 12384 4896 12436
rect 4948 12424 4954 12436
rect 5077 12427 5135 12433
rect 5077 12424 5089 12427
rect 4948 12396 5089 12424
rect 4948 12384 4954 12396
rect 5077 12393 5089 12396
rect 5123 12393 5135 12427
rect 5077 12387 5135 12393
rect 5258 12384 5264 12436
rect 5316 12424 5322 12436
rect 5353 12427 5411 12433
rect 5353 12424 5365 12427
rect 5316 12396 5365 12424
rect 5316 12384 5322 12396
rect 5353 12393 5365 12396
rect 5399 12393 5411 12427
rect 5353 12387 5411 12393
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 6181 12427 6239 12433
rect 6181 12424 6193 12427
rect 5500 12396 6193 12424
rect 5500 12384 5506 12396
rect 6181 12393 6193 12396
rect 6227 12393 6239 12427
rect 6181 12387 6239 12393
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 8846 12424 8852 12436
rect 6595 12396 8852 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 10045 12427 10103 12433
rect 10045 12424 10057 12427
rect 10008 12396 10057 12424
rect 10008 12384 10014 12396
rect 10045 12393 10057 12396
rect 10091 12393 10103 12427
rect 10045 12387 10103 12393
rect 10597 12427 10655 12433
rect 10597 12393 10609 12427
rect 10643 12424 10655 12427
rect 10962 12424 10968 12436
rect 10643 12396 10968 12424
rect 10643 12393 10655 12396
rect 10597 12387 10655 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 12802 12424 12808 12436
rect 11348 12396 12808 12424
rect 1848 12359 1906 12365
rect 1848 12325 1860 12359
rect 1894 12356 1906 12359
rect 2774 12356 2780 12368
rect 1894 12328 2780 12356
rect 1894 12325 1906 12328
rect 1848 12319 1906 12325
rect 2774 12316 2780 12328
rect 2832 12356 2838 12368
rect 4433 12359 4491 12365
rect 4433 12356 4445 12359
rect 2832 12328 4445 12356
rect 2832 12316 2838 12328
rect 4433 12325 4445 12328
rect 4479 12325 4491 12359
rect 4433 12319 4491 12325
rect 5721 12359 5779 12365
rect 5721 12325 5733 12359
rect 5767 12356 5779 12359
rect 5767 12328 6592 12356
rect 5767 12325 5779 12328
rect 5721 12319 5779 12325
rect 6564 12300 6592 12328
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 7558 12356 7564 12368
rect 7248 12328 7564 12356
rect 7248 12316 7254 12328
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 8202 12356 8208 12368
rect 7984 12328 8208 12356
rect 7984 12316 7990 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 9401 12359 9459 12365
rect 9401 12325 9413 12359
rect 9447 12356 9459 12359
rect 11348 12356 11376 12396
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 14921 12427 14979 12433
rect 13065 12396 13952 12424
rect 9447 12328 11376 12356
rect 9447 12325 9459 12328
rect 9401 12319 9459 12325
rect 12618 12316 12624 12368
rect 12676 12356 12682 12368
rect 13065 12356 13093 12396
rect 13170 12356 13176 12368
rect 12676 12328 13093 12356
rect 13131 12328 13176 12356
rect 12676 12316 12682 12328
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 13924 12356 13952 12396
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15194 12424 15200 12436
rect 14967 12396 15200 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 16485 12427 16543 12433
rect 16485 12424 16497 12427
rect 15304 12396 16497 12424
rect 15304 12356 15332 12396
rect 16485 12393 16497 12396
rect 16531 12393 16543 12427
rect 16485 12387 16543 12393
rect 17037 12427 17095 12433
rect 17037 12393 17049 12427
rect 17083 12424 17095 12427
rect 18322 12424 18328 12436
rect 17083 12396 18328 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 13924 12328 15332 12356
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 15562 12356 15568 12368
rect 15436 12328 15568 12356
rect 15436 12316 15442 12328
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 16500 12356 16528 12387
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 19153 12427 19211 12433
rect 19153 12393 19165 12427
rect 19199 12424 19211 12427
rect 19242 12424 19248 12436
rect 19199 12396 19248 12424
rect 19199 12393 19211 12396
rect 19153 12387 19211 12393
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 19978 12384 19984 12436
rect 20036 12424 20042 12436
rect 20036 12396 20116 12424
rect 20036 12384 20042 12396
rect 17402 12356 17408 12368
rect 16500 12328 17408 12356
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 17862 12356 17868 12368
rect 17512 12328 17868 12356
rect 1578 12288 1584 12300
rect 1539 12260 1584 12288
rect 1578 12248 1584 12260
rect 1636 12248 1642 12300
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 4338 12288 4344 12300
rect 3467 12260 4344 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12288 5043 12291
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 5031 12260 5273 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 5813 12291 5871 12297
rect 5813 12257 5825 12291
rect 5859 12288 5871 12291
rect 6181 12291 6239 12297
rect 5859 12260 6132 12288
rect 5859 12257 5871 12260
rect 5813 12251 5871 12257
rect 3050 12180 3056 12232
rect 3108 12220 3114 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 3108 12192 4537 12220
rect 3108 12180 3114 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4672 12192 4721 12220
rect 4672 12180 4678 12192
rect 4709 12189 4721 12192
rect 4755 12220 4767 12223
rect 5718 12220 5724 12232
rect 4755 12192 5724 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 5718 12180 5724 12192
rect 5776 12220 5782 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5776 12192 5917 12220
rect 5776 12180 5782 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 2682 12112 2688 12164
rect 2740 12152 2746 12164
rect 2961 12155 3019 12161
rect 2961 12152 2973 12155
rect 2740 12124 2973 12152
rect 2740 12112 2746 12124
rect 2961 12121 2973 12124
rect 3007 12152 3019 12155
rect 3970 12152 3976 12164
rect 3007 12124 3976 12152
rect 3007 12121 3019 12124
rect 2961 12115 3019 12121
rect 3970 12112 3976 12124
rect 4028 12112 4034 12164
rect 4890 12112 4896 12164
rect 4948 12152 4954 12164
rect 4948 12124 5304 12152
rect 4948 12112 4954 12124
rect 5276 12096 5304 12124
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3292 12056 4077 12084
rect 3292 12044 3298 12056
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 4065 12047 4123 12053
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 4985 12087 5043 12093
rect 4985 12084 4997 12087
rect 4488 12056 4997 12084
rect 4488 12044 4494 12056
rect 4985 12053 4997 12056
rect 5031 12053 5043 12087
rect 4985 12047 5043 12053
rect 5258 12044 5264 12096
rect 5316 12044 5322 12096
rect 6104 12084 6132 12260
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 6227 12260 6377 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6546 12248 6552 12300
rect 6604 12248 6610 12300
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 7282 12297 7288 12300
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6880 12260 7021 12288
rect 6880 12248 6886 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7276 12288 7288 12297
rect 7243 12260 7288 12288
rect 7009 12251 7067 12257
rect 7276 12251 7288 12260
rect 7340 12288 7346 12300
rect 8018 12288 8024 12300
rect 7340 12260 8024 12288
rect 7282 12248 7288 12251
rect 7340 12248 7346 12260
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 8846 12288 8852 12300
rect 8807 12260 8852 12288
rect 8846 12248 8852 12260
rect 8904 12248 8910 12300
rect 9033 12291 9091 12297
rect 9033 12257 9045 12291
rect 9079 12288 9091 12291
rect 9079 12260 9812 12288
rect 9079 12257 9091 12260
rect 9033 12251 9091 12257
rect 9784 12220 9812 12260
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10781 12291 10839 12297
rect 9916 12260 9961 12288
rect 9916 12248 9922 12260
rect 10781 12257 10793 12291
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 10318 12220 10324 12232
rect 9784 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10796 12220 10824 12251
rect 10962 12248 10968 12300
rect 11020 12288 11026 12300
rect 11425 12291 11483 12297
rect 11425 12288 11437 12291
rect 11020 12260 11437 12288
rect 11020 12248 11026 12260
rect 11425 12257 11437 12260
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 13136 12260 13277 12288
rect 13136 12248 13142 12260
rect 13265 12257 13277 12260
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13354 12248 13360 12300
rect 13412 12288 13418 12300
rect 13521 12291 13579 12297
rect 13521 12288 13533 12291
rect 13412 12260 13533 12288
rect 13412 12248 13418 12260
rect 13521 12257 13533 12260
rect 13567 12257 13579 12291
rect 13521 12251 13579 12257
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 14148 12260 14749 12288
rect 14148 12248 14154 12260
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 14737 12251 14795 12257
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 17512 12297 17540 12328
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 18414 12316 18420 12368
rect 18472 12356 18478 12368
rect 19337 12359 19395 12365
rect 18472 12328 19012 12356
rect 18472 12316 18478 12328
rect 16393 12291 16451 12297
rect 16393 12288 16405 12291
rect 15804 12260 16405 12288
rect 15804 12248 15810 12260
rect 16393 12257 16405 12260
rect 16439 12257 16451 12291
rect 16393 12251 16451 12257
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 17764 12291 17822 12297
rect 17764 12257 17776 12291
rect 17810 12288 17822 12291
rect 18690 12288 18696 12300
rect 17810 12260 18696 12288
rect 17810 12257 17822 12260
rect 17764 12251 17822 12257
rect 18690 12248 18696 12260
rect 18748 12248 18754 12300
rect 18984 12297 19012 12328
rect 19337 12325 19349 12359
rect 19383 12356 19395 12359
rect 19889 12359 19947 12365
rect 19889 12356 19901 12359
rect 19383 12328 19901 12356
rect 19383 12325 19395 12328
rect 19337 12319 19395 12325
rect 19889 12325 19901 12328
rect 19935 12325 19947 12359
rect 19889 12319 19947 12325
rect 18969 12291 19027 12297
rect 18969 12257 18981 12291
rect 19015 12257 19027 12291
rect 20088 12288 20116 12396
rect 20714 12316 20720 12368
rect 20772 12356 20778 12368
rect 22557 12359 22615 12365
rect 22557 12356 22569 12359
rect 20772 12328 22569 12356
rect 20772 12316 20778 12328
rect 22557 12325 22569 12328
rect 22603 12325 22615 12359
rect 22557 12319 22615 12325
rect 20346 12288 20352 12300
rect 20088 12260 20352 12288
rect 18969 12251 19027 12257
rect 20346 12248 20352 12260
rect 20404 12248 20410 12300
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 20990 12248 20996 12300
rect 21048 12288 21054 12300
rect 21157 12291 21215 12297
rect 21157 12288 21169 12291
rect 21048 12260 21169 12288
rect 21048 12248 21054 12260
rect 21157 12257 21169 12260
rect 21203 12257 21215 12291
rect 21157 12251 21215 12257
rect 10796 12192 13308 12220
rect 8846 12112 8852 12164
rect 8904 12112 8910 12164
rect 9217 12155 9275 12161
rect 9217 12121 9229 12155
rect 9263 12152 9275 12155
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 9263 12124 9413 12152
rect 9263 12121 9275 12124
rect 9217 12115 9275 12121
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 11882 12152 11888 12164
rect 9732 12124 11888 12152
rect 9732 12112 9738 12124
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 6270 12084 6276 12096
rect 6104 12056 6276 12084
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8076 12056 8401 12084
rect 8076 12044 8082 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8389 12047 8447 12053
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 8665 12087 8723 12093
rect 8665 12084 8677 12087
rect 8628 12056 8677 12084
rect 8628 12044 8634 12056
rect 8665 12053 8677 12056
rect 8711 12053 8723 12087
rect 8864 12084 8892 12112
rect 11330 12084 11336 12096
rect 8864 12056 11336 12084
rect 8665 12047 8723 12053
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 12434 12044 12440 12096
rect 12492 12084 12498 12096
rect 13078 12084 13084 12096
rect 12492 12056 13084 12084
rect 12492 12044 12498 12056
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13280 12084 13308 12192
rect 15378 12180 15384 12232
rect 15436 12220 15442 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 15436 12192 16589 12220
rect 15436 12180 15442 12192
rect 16577 12189 16589 12192
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 19794 12180 19800 12232
rect 19852 12220 19858 12232
rect 19981 12223 20039 12229
rect 19981 12220 19993 12223
rect 19852 12192 19993 12220
rect 19852 12180 19858 12192
rect 19981 12189 19993 12192
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 20070 12180 20076 12232
rect 20128 12220 20134 12232
rect 20128 12192 20173 12220
rect 20128 12180 20134 12192
rect 14274 12112 14280 12164
rect 14332 12152 14338 12164
rect 14645 12155 14703 12161
rect 14645 12152 14657 12155
rect 14332 12124 14657 12152
rect 14332 12112 14338 12124
rect 14645 12121 14657 12124
rect 14691 12121 14703 12155
rect 14645 12115 14703 12121
rect 15657 12155 15715 12161
rect 15657 12121 15669 12155
rect 15703 12152 15715 12155
rect 16482 12152 16488 12164
rect 15703 12124 16488 12152
rect 15703 12121 15715 12124
rect 15657 12115 15715 12121
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 18506 12112 18512 12164
rect 18564 12152 18570 12164
rect 19337 12155 19395 12161
rect 19337 12152 19349 12155
rect 18564 12124 19349 12152
rect 18564 12112 18570 12124
rect 19337 12121 19349 12124
rect 19383 12121 19395 12155
rect 19337 12115 19395 12121
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 20088 12152 20116 12180
rect 19760 12124 20116 12152
rect 19760 12112 19766 12124
rect 14458 12084 14464 12096
rect 13280 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15528 12056 16037 12084
rect 15528 12044 15534 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18782 12084 18788 12096
rect 18196 12056 18788 12084
rect 18196 12044 18202 12056
rect 18782 12044 18788 12056
rect 18840 12084 18846 12096
rect 18877 12087 18935 12093
rect 18877 12084 18889 12087
rect 18840 12056 18889 12084
rect 18840 12044 18846 12056
rect 18877 12053 18889 12056
rect 18923 12053 18935 12087
rect 18877 12047 18935 12053
rect 19521 12087 19579 12093
rect 19521 12053 19533 12087
rect 19567 12084 19579 12087
rect 20622 12084 20628 12096
rect 19567 12056 20628 12084
rect 19567 12053 19579 12056
rect 19521 12047 19579 12053
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 22244 12056 22293 12084
rect 22244 12044 22250 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22281 12047 22339 12053
rect 1104 11994 23276 12016
rect 1104 11942 4680 11994
rect 4732 11942 4744 11994
rect 4796 11942 4808 11994
rect 4860 11942 4872 11994
rect 4924 11942 12078 11994
rect 12130 11942 12142 11994
rect 12194 11942 12206 11994
rect 12258 11942 12270 11994
rect 12322 11942 19475 11994
rect 19527 11942 19539 11994
rect 19591 11942 19603 11994
rect 19655 11942 19667 11994
rect 19719 11942 23276 11994
rect 1104 11920 23276 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2832 11852 2881 11880
rect 2832 11840 2838 11852
rect 2869 11849 2881 11852
rect 2915 11849 2927 11883
rect 5258 11880 5264 11892
rect 2869 11843 2927 11849
rect 5092 11852 5264 11880
rect 4341 11815 4399 11821
rect 4341 11781 4353 11815
rect 4387 11812 4399 11815
rect 4798 11812 4804 11824
rect 4387 11784 4804 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 3970 11744 3976 11756
rect 3835 11716 3976 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 3970 11704 3976 11716
rect 4028 11744 4034 11756
rect 4522 11744 4528 11756
rect 4028 11716 4528 11744
rect 4028 11704 4034 11716
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5092 11753 5120 11852
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 8570 11880 8576 11892
rect 6687 11852 8576 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 8570 11840 8576 11852
rect 8628 11880 8634 11892
rect 8938 11880 8944 11892
rect 8628 11852 8944 11880
rect 8628 11840 8634 11852
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9033 11883 9091 11889
rect 9033 11849 9045 11883
rect 9079 11880 9091 11883
rect 10042 11880 10048 11892
rect 9079 11852 10048 11880
rect 9079 11849 9091 11852
rect 9033 11843 9091 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 10744 11852 11805 11880
rect 10744 11840 10750 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 15473 11883 15531 11889
rect 15473 11880 15485 11883
rect 14608 11852 15485 11880
rect 14608 11840 14614 11852
rect 15473 11849 15485 11852
rect 15519 11849 15531 11883
rect 15473 11843 15531 11849
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 19334 11880 19340 11892
rect 15712 11852 19340 11880
rect 15712 11840 15718 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 20162 11840 20168 11892
rect 20220 11880 20226 11892
rect 20714 11880 20720 11892
rect 20220 11852 20720 11880
rect 20220 11840 20226 11852
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 21634 11880 21640 11892
rect 20947 11852 21640 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 9401 11815 9459 11821
rect 9401 11781 9413 11815
rect 9447 11812 9459 11815
rect 9950 11812 9956 11824
rect 9447 11784 9956 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10410 11772 10416 11824
rect 10468 11772 10474 11824
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 15838 11812 15844 11824
rect 12584 11784 15844 11812
rect 12584 11772 12590 11784
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 15933 11815 15991 11821
rect 15933 11781 15945 11815
rect 15979 11781 15991 11815
rect 15933 11775 15991 11781
rect 5077 11747 5135 11753
rect 5077 11744 5089 11747
rect 4948 11716 5089 11744
rect 4948 11704 4954 11716
rect 5077 11713 5089 11716
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 6880 11716 7205 11744
rect 6880 11704 6886 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 10042 11744 10048 11756
rect 10003 11716 10048 11744
rect 7193 11707 7251 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 1486 11676 1492 11688
rect 1447 11648 1492 11676
rect 1486 11636 1492 11648
rect 1544 11636 1550 11688
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 4120 11648 4169 11676
rect 4120 11636 4126 11648
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4985 11679 5043 11685
rect 4985 11645 4997 11679
rect 5031 11676 5043 11679
rect 6641 11679 6699 11685
rect 6641 11676 6653 11679
rect 5031 11648 6653 11676
rect 5031 11645 5043 11648
rect 4985 11639 5043 11645
rect 6641 11645 6653 11648
rect 6687 11645 6699 11679
rect 6641 11639 6699 11645
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 10428 11685 10456 11772
rect 14182 11744 14188 11756
rect 12636 11716 14188 11744
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 7800 11648 8861 11676
rect 7800 11636 7806 11648
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 12636 11685 12664 11716
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11744 14427 11747
rect 14458 11744 14464 11756
rect 14415 11716 14464 11744
rect 14415 11713 14427 11716
rect 14369 11707 14427 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14568 11716 14933 11744
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11204 11648 11989 11676
rect 11204 11636 11210 11648
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 13078 11636 13084 11688
rect 13136 11676 13142 11688
rect 14568 11676 14596 11716
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 15102 11744 15108 11756
rect 15063 11716 15108 11744
rect 14921 11707 14979 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15948 11744 15976 11775
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 16080 11784 16620 11812
rect 16080 11772 16086 11784
rect 16390 11744 16396 11756
rect 15948 11716 16396 11744
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 16592 11753 16620 11784
rect 18874 11772 18880 11824
rect 18932 11812 18938 11824
rect 19058 11812 19064 11824
rect 18932 11784 19064 11812
rect 18932 11772 18938 11784
rect 19058 11772 19064 11784
rect 19116 11772 19122 11824
rect 16577 11747 16635 11753
rect 16577 11713 16589 11747
rect 16623 11744 16635 11747
rect 17494 11744 17500 11756
rect 16623 11716 17500 11744
rect 16623 11713 16635 11716
rect 16577 11707 16635 11713
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 17770 11704 17776 11756
rect 17828 11744 17834 11756
rect 18506 11744 18512 11756
rect 17828 11716 18512 11744
rect 17828 11704 17834 11716
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 18690 11744 18696 11756
rect 18603 11716 18696 11744
rect 18690 11704 18696 11716
rect 18748 11744 18754 11756
rect 19610 11753 19616 11756
rect 19567 11747 19616 11753
rect 18748 11716 19472 11744
rect 18748 11704 18754 11716
rect 13136 11648 14596 11676
rect 13136 11636 13142 11648
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 15289 11679 15347 11685
rect 15289 11676 15301 11679
rect 15252 11648 15301 11676
rect 15252 11636 15258 11648
rect 15289 11645 15301 11648
rect 15335 11645 15347 11679
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 15289 11639 15347 11645
rect 15387 11648 17417 11676
rect 1756 11611 1814 11617
rect 1756 11577 1768 11611
rect 1802 11608 1814 11611
rect 3050 11608 3056 11620
rect 1802 11580 3056 11608
rect 1802 11577 1814 11580
rect 1756 11571 1814 11577
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 3605 11611 3663 11617
rect 3605 11608 3617 11611
rect 3476 11580 3617 11608
rect 3476 11568 3482 11580
rect 3605 11577 3617 11580
rect 3651 11608 3663 11611
rect 5344 11611 5402 11617
rect 3651 11580 4936 11608
rect 3651 11577 3663 11580
rect 3605 11571 3663 11577
rect 3142 11540 3148 11552
rect 3103 11512 3148 11540
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 4798 11540 4804 11552
rect 4488 11512 4804 11540
rect 4488 11500 4494 11512
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 4908 11540 4936 11580
rect 5344 11577 5356 11611
rect 5390 11608 5402 11611
rect 6546 11608 6552 11620
rect 5390 11580 6552 11608
rect 5390 11577 5402 11580
rect 5344 11571 5402 11577
rect 6546 11568 6552 11580
rect 6604 11608 6610 11620
rect 6914 11608 6920 11620
rect 6604 11580 6920 11608
rect 6604 11568 6610 11580
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7098 11568 7104 11620
rect 7156 11608 7162 11620
rect 7438 11611 7496 11617
rect 7438 11608 7450 11611
rect 7156 11580 7450 11608
rect 7156 11568 7162 11580
rect 7438 11577 7450 11580
rect 7484 11608 7496 11611
rect 8018 11608 8024 11620
rect 7484 11580 8024 11608
rect 7484 11577 7496 11580
rect 7438 11571 7496 11577
rect 8018 11568 8024 11580
rect 8076 11568 8082 11620
rect 9769 11611 9827 11617
rect 9769 11577 9781 11611
rect 9815 11608 9827 11611
rect 10680 11611 10738 11617
rect 10680 11608 10692 11611
rect 9815 11580 10692 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 10680 11577 10692 11580
rect 10726 11608 10738 11611
rect 11882 11608 11888 11620
rect 10726 11580 11888 11608
rect 10726 11577 10738 11580
rect 10680 11571 10738 11577
rect 11882 11568 11888 11580
rect 11940 11568 11946 11620
rect 14642 11608 14648 11620
rect 13556 11580 14648 11608
rect 6457 11543 6515 11549
rect 6457 11540 6469 11543
rect 4908 11512 6469 11540
rect 6457 11509 6469 11512
rect 6503 11509 6515 11543
rect 6457 11503 6515 11509
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 7616 11512 8585 11540
rect 7616 11500 7622 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 9858 11540 9864 11552
rect 9819 11512 9864 11540
rect 8573 11503 8631 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 11514 11540 11520 11552
rect 10100 11512 11520 11540
rect 10100 11500 10106 11512
rect 11514 11500 11520 11512
rect 11572 11540 11578 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11572 11512 12173 11540
rect 11572 11500 11578 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 13556 11540 13584 11580
rect 14642 11568 14648 11580
rect 14700 11568 14706 11620
rect 14829 11611 14887 11617
rect 14829 11577 14841 11611
rect 14875 11608 14887 11611
rect 15010 11608 15016 11620
rect 14875 11580 15016 11608
rect 14875 11577 14887 11580
rect 14829 11571 14887 11577
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 12308 11512 13584 11540
rect 12308 11500 12314 11512
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 14274 11540 14280 11552
rect 13964 11512 14280 11540
rect 13964 11500 13970 11512
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14461 11543 14519 11549
rect 14461 11509 14473 11543
rect 14507 11540 14519 11543
rect 14550 11540 14556 11552
rect 14507 11512 14556 11540
rect 14507 11509 14519 11512
rect 14461 11503 14519 11509
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 15387 11540 15415 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 17920 11648 19073 11676
rect 17920 11636 17926 11648
rect 19061 11645 19073 11648
rect 19107 11676 19119 11679
rect 19150 11676 19156 11688
rect 19107 11648 19156 11676
rect 19107 11645 19119 11648
rect 19061 11639 19119 11645
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 19444 11676 19472 11716
rect 19567 11713 19579 11747
rect 19613 11713 19616 11747
rect 19567 11707 19616 11713
rect 19610 11704 19616 11707
rect 19668 11704 19674 11756
rect 19794 11744 19800 11756
rect 19755 11716 19800 11744
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 19444 11648 20484 11676
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 18564 11580 18828 11608
rect 18564 11568 18570 11580
rect 14976 11512 15415 11540
rect 14976 11500 14982 11512
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16264 11512 16313 11540
rect 16264 11500 16270 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 16448 11512 16493 11540
rect 16448 11500 16454 11512
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16816 11512 16957 11540
rect 16816 11500 16822 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17313 11543 17371 11549
rect 17313 11540 17325 11543
rect 17184 11512 17325 11540
rect 17184 11500 17190 11512
rect 17313 11509 17325 11512
rect 17359 11509 17371 11543
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 17313 11503 17371 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18417 11543 18475 11549
rect 18417 11509 18429 11543
rect 18463 11540 18475 11543
rect 18690 11540 18696 11552
rect 18463 11512 18696 11540
rect 18463 11509 18475 11512
rect 18417 11503 18475 11509
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 18800 11540 18828 11580
rect 19527 11543 19585 11549
rect 19527 11540 19539 11543
rect 18800 11512 19539 11540
rect 19527 11509 19539 11512
rect 19573 11540 19585 11543
rect 20254 11540 20260 11552
rect 19573 11512 20260 11540
rect 19573 11509 19585 11512
rect 19527 11503 19585 11509
rect 20254 11500 20260 11512
rect 20312 11500 20318 11552
rect 20456 11540 20484 11648
rect 21266 11636 21272 11688
rect 21324 11676 21330 11688
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 21324 11648 21373 11676
rect 21324 11636 21330 11648
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 21628 11611 21686 11617
rect 21628 11577 21640 11611
rect 21674 11608 21686 11611
rect 22646 11608 22652 11620
rect 21674 11580 22652 11608
rect 21674 11577 21686 11580
rect 21628 11571 21686 11577
rect 22646 11568 22652 11580
rect 22704 11568 22710 11620
rect 22741 11543 22799 11549
rect 22741 11540 22753 11543
rect 20456 11512 22753 11540
rect 22741 11509 22753 11512
rect 22787 11509 22799 11543
rect 22741 11503 22799 11509
rect 1104 11450 23276 11472
rect 1104 11398 8379 11450
rect 8431 11398 8443 11450
rect 8495 11398 8507 11450
rect 8559 11398 8571 11450
rect 8623 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 15904 11450
rect 15956 11398 15968 11450
rect 16020 11398 23276 11450
rect 1104 11376 23276 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3050 11336 3056 11348
rect 2915 11308 3056 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 3605 11339 3663 11345
rect 3605 11305 3617 11339
rect 3651 11336 3663 11339
rect 3694 11336 3700 11348
rect 3651 11308 3700 11336
rect 3651 11305 3663 11308
rect 3605 11299 3663 11305
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 5258 11296 5264 11348
rect 5316 11336 5322 11348
rect 5442 11336 5448 11348
rect 5316 11308 5448 11336
rect 5316 11296 5322 11308
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 6328 11308 6561 11336
rect 6328 11296 6334 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 8846 11296 8852 11348
rect 8904 11296 8910 11348
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 9674 11336 9680 11348
rect 9263 11308 9680 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11882 11336 11888 11348
rect 11843 11308 11888 11336
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 12621 11339 12679 11345
rect 12621 11305 12633 11339
rect 12667 11336 12679 11339
rect 13538 11336 13544 11348
rect 12667 11308 13544 11336
rect 12667 11305 12679 11308
rect 12621 11299 12679 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 15620 11308 17356 11336
rect 15620 11296 15626 11308
rect 1756 11271 1814 11277
rect 1756 11237 1768 11271
rect 1802 11268 1814 11271
rect 4798 11268 4804 11280
rect 1802 11240 2728 11268
rect 1802 11237 1814 11240
rect 1756 11231 1814 11237
rect 1486 11200 1492 11212
rect 1447 11172 1492 11200
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 2700 11132 2728 11240
rect 3344 11240 4804 11268
rect 3344 11209 3372 11240
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11200 3479 11203
rect 4430 11200 4436 11212
rect 3467 11172 4016 11200
rect 4391 11172 4436 11200
rect 3467 11169 3479 11172
rect 3421 11163 3479 11169
rect 3510 11132 3516 11144
rect 2700 11104 3516 11132
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 3145 10999 3203 11005
rect 3145 10965 3157 10999
rect 3191 10996 3203 10999
rect 3326 10996 3332 11008
rect 3191 10968 3332 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 3988 10996 4016 11172
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 4540 11132 4568 11163
rect 4890 11160 4896 11212
rect 4948 11200 4954 11212
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 4948 11172 5181 11200
rect 4948 11160 4954 11172
rect 5169 11169 5181 11172
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5436 11203 5494 11209
rect 5436 11169 5448 11203
rect 5482 11200 5494 11203
rect 5718 11200 5724 11212
rect 5482 11172 5724 11200
rect 5482 11169 5494 11172
rect 5436 11163 5494 11169
rect 5718 11160 5724 11172
rect 5776 11200 5782 11212
rect 6362 11200 6368 11212
rect 5776 11172 6368 11200
rect 5776 11160 5782 11172
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7558 11209 7564 11212
rect 7552 11200 7564 11209
rect 7519 11172 7564 11200
rect 7552 11163 7564 11172
rect 7558 11160 7564 11163
rect 7616 11160 7622 11212
rect 8864 11200 8892 11296
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 12434 11268 12440 11280
rect 9180 11240 12440 11268
rect 9180 11228 9186 11240
rect 12434 11228 12440 11240
rect 12492 11228 12498 11280
rect 12986 11228 12992 11280
rect 13044 11277 13050 11280
rect 13044 11271 13108 11277
rect 13044 11237 13062 11271
rect 13096 11237 13108 11271
rect 16298 11268 16304 11280
rect 13044 11231 13108 11237
rect 14660 11240 16304 11268
rect 13044 11228 13050 11231
rect 9021 11203 9079 11209
rect 9021 11200 9033 11203
rect 8864 11172 9033 11200
rect 9021 11169 9033 11172
rect 9067 11169 9079 11203
rect 9021 11163 9079 11169
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10772 11203 10830 11209
rect 10772 11200 10784 11203
rect 10367 11172 10784 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 10772 11169 10784 11172
rect 10818 11200 10830 11203
rect 11790 11200 11796 11212
rect 10818 11172 11796 11200
rect 10818 11169 10830 11172
rect 10772 11163 10830 11169
rect 4706 11132 4712 11144
rect 4448 11104 4568 11132
rect 4667 11104 4712 11132
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4338 11064 4344 11076
rect 4111 11036 4344 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 4448 11064 4476 11104
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 6822 11132 6828 11144
rect 6783 11104 6828 11132
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 4522 11064 4528 11076
rect 4448 11036 4528 11064
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 7300 11064 7328 11095
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 9968 11132 9996 11163
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 12250 11200 12256 11212
rect 12211 11172 12256 11200
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13354 11200 13360 11212
rect 12952 11172 13360 11200
rect 12952 11160 12958 11172
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 14660 11209 14688 11240
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 16574 11228 16580 11280
rect 16632 11268 16638 11280
rect 17034 11268 17040 11280
rect 16632 11240 17040 11268
rect 16632 11228 16638 11240
rect 17034 11228 17040 11240
rect 17092 11228 17098 11280
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 15913 11203 15971 11209
rect 15913 11200 15925 11203
rect 15620 11172 15925 11200
rect 15620 11160 15626 11172
rect 15913 11169 15925 11172
rect 15959 11200 15971 11203
rect 16482 11200 16488 11212
rect 15959 11172 16488 11200
rect 15959 11169 15971 11172
rect 15913 11163 15971 11169
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 17328 11209 17356 11308
rect 17402 11296 17408 11348
rect 17460 11336 17466 11348
rect 19794 11336 19800 11348
rect 17460 11308 19380 11336
rect 19755 11308 19800 11336
rect 17460 11296 17466 11308
rect 17313 11203 17371 11209
rect 17313 11169 17325 11203
rect 17359 11169 17371 11203
rect 19352 11200 19380 11308
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 22646 11336 22652 11348
rect 22607 11308 22652 11336
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 21536 11271 21594 11277
rect 21536 11237 21548 11271
rect 21582 11268 21594 11271
rect 22186 11268 22192 11280
rect 21582 11240 22192 11268
rect 21582 11237 21594 11240
rect 21536 11231 21594 11237
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 20073 11203 20131 11209
rect 20073 11200 20085 11203
rect 17313 11163 17371 11169
rect 17420 11172 18828 11200
rect 19352 11172 20085 11200
rect 8812 11104 9996 11132
rect 8812 11092 8818 11104
rect 10410 11092 10416 11144
rect 10468 11132 10474 11144
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 10468 11104 10517 11132
rect 10468 11092 10474 11104
rect 10505 11101 10517 11104
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12768 11104 12817 11132
rect 12768 11092 12774 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 8665 11067 8723 11073
rect 8665 11064 8677 11067
rect 6604 11036 7328 11064
rect 8220 11036 8677 11064
rect 6604 11024 6610 11036
rect 7006 10996 7012 11008
rect 3988 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8220 10996 8248 11036
rect 8665 11033 8677 11036
rect 8711 11033 8723 11067
rect 8665 11027 8723 11033
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10428 11064 10456 11092
rect 10008 11036 10456 11064
rect 12437 11067 12495 11073
rect 10008 11024 10014 11036
rect 12437 11033 12449 11067
rect 12483 11064 12495 11067
rect 12621 11067 12679 11073
rect 12621 11064 12633 11067
rect 12483 11036 12633 11064
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 12621 11033 12633 11036
rect 12667 11033 12679 11067
rect 12621 11027 12679 11033
rect 14642 11024 14648 11076
rect 14700 11064 14706 11076
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 14700 11036 14841 11064
rect 14700 11024 14706 11036
rect 14829 11033 14841 11036
rect 14875 11033 14887 11067
rect 14829 11027 14887 11033
rect 15010 11024 15016 11076
rect 15068 11064 15074 11076
rect 15194 11064 15200 11076
rect 15068 11036 15200 11064
rect 15068 11024 15074 11036
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 8076 10968 8248 10996
rect 8076 10956 8082 10968
rect 9858 10956 9864 11008
rect 9916 10996 9922 11008
rect 10321 10999 10379 11005
rect 10321 10996 10333 10999
rect 9916 10968 10333 10996
rect 9916 10956 9922 10968
rect 10321 10965 10333 10968
rect 10367 10965 10379 10999
rect 10321 10959 10379 10965
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13722 10996 13728 11008
rect 12860 10968 13728 10996
rect 12860 10956 12866 10968
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 13906 10956 13912 11008
rect 13964 10996 13970 11008
rect 14185 10999 14243 11005
rect 14185 10996 14197 10999
rect 13964 10968 14197 10996
rect 13964 10956 13970 10968
rect 14185 10965 14197 10968
rect 14231 10965 14243 10999
rect 15672 10996 15700 11095
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 17420 11132 17448 11172
rect 16724 11104 17448 11132
rect 16724 11092 16730 11104
rect 17862 11092 17868 11144
rect 17920 11132 17926 11144
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 17920 11104 17969 11132
rect 17920 11092 17926 11104
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 18230 11092 18236 11144
rect 18288 11141 18294 11144
rect 18288 11135 18338 11141
rect 18288 11101 18292 11135
rect 18326 11101 18338 11135
rect 18288 11095 18338 11101
rect 18288 11092 18294 11095
rect 18414 11092 18420 11144
rect 18472 11132 18478 11144
rect 18690 11132 18696 11144
rect 18472 11104 18517 11132
rect 18651 11104 18696 11132
rect 18472 11092 18478 11104
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 18800 11132 18828 11172
rect 20073 11169 20085 11172
rect 20119 11169 20131 11203
rect 21266 11200 21272 11212
rect 21227 11172 21272 11200
rect 20073 11163 20131 11169
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 18800 11104 20300 11132
rect 20272 11073 20300 11104
rect 20257 11067 20315 11073
rect 20257 11033 20269 11067
rect 20303 11033 20315 11067
rect 20257 11027 20315 11033
rect 15930 10996 15936 11008
rect 15672 10968 15936 10996
rect 14185 10959 14243 10965
rect 15930 10956 15936 10968
rect 15988 10956 15994 11008
rect 17034 10996 17040 11008
rect 16995 10968 17040 10996
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 17494 10996 17500 11008
rect 17455 10968 17500 10996
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 18506 10996 18512 11008
rect 18288 10968 18512 10996
rect 18288 10956 18294 10968
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 18598 10956 18604 11008
rect 18656 10996 18662 11008
rect 19150 10996 19156 11008
rect 18656 10968 19156 10996
rect 18656 10956 18662 10968
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 1104 10906 23276 10928
rect 1104 10854 4680 10906
rect 4732 10854 4744 10906
rect 4796 10854 4808 10906
rect 4860 10854 4872 10906
rect 4924 10854 12078 10906
rect 12130 10854 12142 10906
rect 12194 10854 12206 10906
rect 12258 10854 12270 10906
rect 12322 10854 19475 10906
rect 19527 10854 19539 10906
rect 19591 10854 19603 10906
rect 19655 10854 19667 10906
rect 19719 10854 23276 10906
rect 1104 10832 23276 10854
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 3510 10792 3516 10804
rect 3099 10764 3516 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3510 10752 3516 10764
rect 3568 10752 3574 10804
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 4488 10764 4721 10792
rect 4488 10752 4494 10764
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 6362 10792 6368 10804
rect 6323 10764 6368 10792
rect 4709 10755 4767 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 7009 10795 7067 10801
rect 7009 10761 7021 10795
rect 7055 10792 7067 10795
rect 7466 10792 7472 10804
rect 7055 10764 7472 10792
rect 7055 10761 7067 10764
rect 7009 10755 7067 10761
rect 1486 10616 1492 10668
rect 1544 10656 1550 10668
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1544 10628 1685 10656
rect 1544 10616 1550 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 4890 10616 4896 10668
rect 4948 10656 4954 10668
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4948 10628 4997 10656
rect 4948 10616 4954 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 3326 10588 3332 10600
rect 3287 10560 3332 10588
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 3596 10591 3654 10597
rect 3596 10557 3608 10591
rect 3642 10588 3654 10591
rect 4522 10588 4528 10600
rect 3642 10560 4528 10588
rect 3642 10557 3654 10560
rect 3596 10551 3654 10557
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6236 10560 6837 10588
rect 6236 10548 6242 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 1940 10523 1998 10529
rect 1940 10489 1952 10523
rect 1986 10489 1998 10523
rect 1940 10483 1998 10489
rect 5252 10523 5310 10529
rect 5252 10489 5264 10523
rect 5298 10520 5310 10523
rect 5534 10520 5540 10532
rect 5298 10492 5540 10520
rect 5298 10489 5310 10492
rect 5252 10483 5310 10489
rect 1955 10452 1983 10483
rect 5534 10480 5540 10492
rect 5592 10480 5598 10532
rect 3418 10452 3424 10464
rect 1955 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 7024 10452 7052 10755
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 17034 10792 17040 10804
rect 13639 10764 17040 10792
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 9674 10724 9680 10736
rect 9631 10696 9680 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 9950 10656 9956 10668
rect 8579 10628 9956 10656
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 8579 10588 8607 10628
rect 9692 10600 9720 10628
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 11572 10628 12747 10656
rect 11572 10616 11578 10628
rect 7515 10560 8607 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8996 10560 9321 10588
rect 8996 10548 9002 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 7374 10480 7380 10532
rect 7432 10520 7438 10532
rect 7714 10523 7772 10529
rect 7714 10520 7726 10523
rect 7432 10492 7726 10520
rect 7432 10480 7438 10492
rect 7714 10489 7726 10492
rect 7760 10520 7772 10523
rect 8018 10520 8024 10532
rect 7760 10492 8024 10520
rect 7760 10489 7772 10492
rect 7714 10483 7772 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 9416 10520 9444 10551
rect 9674 10548 9680 10600
rect 9732 10548 9738 10600
rect 10778 10588 10784 10600
rect 10152 10560 10784 10588
rect 10152 10520 10180 10560
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 11793 10591 11851 10597
rect 11793 10557 11805 10591
rect 11839 10588 11851 10591
rect 12434 10588 12440 10600
rect 11839 10560 12440 10588
rect 11839 10557 11851 10560
rect 11793 10551 11851 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12621 10591 12679 10597
rect 12621 10557 12633 10591
rect 12667 10557 12679 10591
rect 12719 10588 12747 10628
rect 12877 10591 12935 10597
rect 12877 10588 12889 10591
rect 12719 10560 12889 10588
rect 12621 10551 12679 10557
rect 12877 10557 12889 10560
rect 12923 10588 12935 10591
rect 13639 10588 13667 10764
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 17402 10752 17408 10804
rect 17460 10792 17466 10804
rect 20254 10792 20260 10804
rect 17460 10764 20260 10792
rect 17460 10752 17466 10764
rect 20254 10752 20260 10764
rect 20312 10752 20318 10804
rect 20901 10795 20959 10801
rect 20901 10761 20913 10795
rect 20947 10792 20959 10795
rect 20990 10792 20996 10804
rect 20947 10764 20996 10792
rect 20947 10761 20959 10764
rect 20901 10755 20959 10761
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 17313 10727 17371 10733
rect 17313 10693 17325 10727
rect 17359 10693 17371 10727
rect 17313 10687 17371 10693
rect 15930 10656 15936 10668
rect 15891 10628 15936 10656
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 17034 10616 17040 10668
rect 17092 10656 17098 10668
rect 17218 10656 17224 10668
rect 17092 10628 17224 10656
rect 17092 10616 17098 10628
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 12923 10560 13667 10588
rect 12923 10557 12935 10560
rect 12877 10551 12935 10557
rect 9416 10492 10180 10520
rect 10220 10523 10278 10529
rect 10220 10489 10232 10523
rect 10266 10489 10278 10523
rect 12526 10520 12532 10532
rect 10220 10483 10278 10489
rect 10796 10492 12532 10520
rect 6236 10424 7052 10452
rect 6236 10412 6242 10424
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8849 10455 8907 10461
rect 8849 10452 8861 10455
rect 8260 10424 8861 10452
rect 8260 10412 8266 10424
rect 8849 10421 8861 10424
rect 8895 10421 8907 10455
rect 8849 10415 8907 10421
rect 8938 10412 8944 10464
rect 8996 10452 9002 10464
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 8996 10424 9137 10452
rect 8996 10412 9002 10424
rect 9125 10421 9137 10424
rect 9171 10421 9183 10455
rect 9125 10415 9183 10421
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 9582 10452 9588 10464
rect 9364 10424 9588 10452
rect 9364 10412 9370 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10244 10452 10272 10483
rect 10796 10464 10824 10492
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12636 10520 12664 10551
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14240 10560 14289 10588
rect 14240 10548 14246 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14544 10591 14602 10597
rect 14544 10557 14556 10591
rect 14590 10588 14602 10591
rect 14918 10588 14924 10600
rect 14590 10560 14924 10588
rect 14590 10557 14602 10560
rect 14544 10551 14602 10557
rect 12710 10520 12716 10532
rect 12636 10492 12716 10520
rect 12710 10480 12716 10492
rect 12768 10480 12774 10532
rect 10008 10424 10272 10452
rect 10008 10412 10014 10424
rect 10778 10412 10784 10464
rect 10836 10412 10842 10464
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 11333 10455 11391 10461
rect 11333 10452 11345 10455
rect 11020 10424 11345 10452
rect 11020 10412 11026 10424
rect 11333 10421 11345 10424
rect 11379 10421 11391 10455
rect 11333 10415 11391 10421
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 11977 10455 12035 10461
rect 11977 10452 11989 10455
rect 11940 10424 11989 10452
rect 11940 10412 11946 10424
rect 11977 10421 11989 10424
rect 12023 10421 12035 10455
rect 11977 10415 12035 10421
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14559 10452 14587 10551
rect 14918 10548 14924 10560
rect 14976 10548 14982 10600
rect 16206 10597 16212 10600
rect 16200 10588 16212 10597
rect 16167 10560 16212 10588
rect 16200 10551 16212 10560
rect 16206 10548 16212 10551
rect 16264 10548 16270 10600
rect 16482 10548 16488 10600
rect 16540 10588 16546 10600
rect 17328 10588 17356 10687
rect 18230 10684 18236 10736
rect 18288 10724 18294 10736
rect 19058 10724 19064 10736
rect 18288 10696 19064 10724
rect 18288 10684 18294 10696
rect 19058 10684 19064 10696
rect 19116 10724 19122 10736
rect 19242 10724 19248 10736
rect 19116 10696 19248 10724
rect 19116 10684 19122 10696
rect 19242 10684 19248 10696
rect 19300 10724 19306 10736
rect 19300 10696 19564 10724
rect 19300 10684 19306 10696
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 19536 10665 19564 10696
rect 18693 10659 18751 10665
rect 18693 10656 18705 10659
rect 18104 10628 18705 10656
rect 18104 10616 18110 10628
rect 18693 10625 18705 10628
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10625 18935 10659
rect 18877 10619 18935 10625
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10625 19579 10659
rect 21008 10656 21036 10752
rect 21913 10659 21971 10665
rect 21913 10656 21925 10659
rect 21008 10628 21925 10656
rect 19521 10619 19579 10625
rect 21913 10625 21925 10628
rect 21959 10625 21971 10659
rect 21913 10619 21971 10625
rect 16540 10560 17356 10588
rect 16540 10548 16546 10560
rect 17494 10548 17500 10600
rect 17552 10588 17558 10600
rect 17773 10591 17831 10597
rect 17773 10588 17785 10591
rect 17552 10560 17785 10588
rect 17552 10548 17558 10560
rect 17773 10557 17785 10560
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 18322 10548 18328 10600
rect 18380 10588 18386 10600
rect 18601 10591 18659 10597
rect 18601 10588 18613 10591
rect 18380 10560 18613 10588
rect 18380 10548 18386 10560
rect 18601 10557 18613 10560
rect 18647 10557 18659 10591
rect 18601 10551 18659 10557
rect 18782 10548 18788 10600
rect 18840 10588 18846 10600
rect 18892 10588 18920 10619
rect 18840 10560 18920 10588
rect 19788 10591 19846 10597
rect 18840 10548 18846 10560
rect 19788 10557 19800 10591
rect 19834 10588 19846 10591
rect 20070 10588 20076 10600
rect 19834 10560 20076 10588
rect 19834 10557 19846 10560
rect 19788 10551 19846 10557
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 21821 10591 21879 10597
rect 21821 10588 21833 10591
rect 20680 10560 21833 10588
rect 20680 10548 20686 10560
rect 21821 10557 21833 10560
rect 21867 10557 21879 10591
rect 21821 10551 21879 10557
rect 22002 10548 22008 10600
rect 22060 10588 22066 10600
rect 22373 10591 22431 10597
rect 22373 10588 22385 10591
rect 22060 10560 22385 10588
rect 22060 10548 22066 10560
rect 22373 10557 22385 10560
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 15010 10480 15016 10532
rect 15068 10520 15074 10532
rect 19334 10520 19340 10532
rect 15068 10492 19340 10520
rect 15068 10480 15074 10492
rect 19334 10480 19340 10492
rect 19392 10480 19398 10532
rect 21174 10520 21180 10532
rect 21135 10492 21180 10520
rect 21174 10480 21180 10492
rect 21232 10520 21238 10532
rect 21729 10523 21787 10529
rect 21729 10520 21741 10523
rect 21232 10492 21741 10520
rect 21232 10480 21238 10492
rect 21729 10489 21741 10492
rect 21775 10489 21787 10523
rect 21729 10483 21787 10489
rect 14047 10424 14587 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14642 10412 14648 10464
rect 14700 10452 14706 10464
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 14700 10424 15669 10452
rect 14700 10412 14706 10424
rect 15657 10421 15669 10424
rect 15703 10452 15715 10455
rect 17126 10452 17132 10464
rect 15703 10424 17132 10452
rect 15703 10421 15715 10424
rect 15657 10415 15715 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17589 10455 17647 10461
rect 17589 10452 17601 10455
rect 17276 10424 17601 10452
rect 17276 10412 17282 10424
rect 17589 10421 17601 10424
rect 17635 10421 17647 10455
rect 17589 10415 17647 10421
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 18104 10424 18245 10452
rect 18104 10412 18110 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 18233 10415 18291 10421
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 18380 10424 19257 10452
rect 18380 10412 18386 10424
rect 19245 10421 19257 10424
rect 19291 10421 19303 10455
rect 19245 10415 19303 10421
rect 19610 10412 19616 10464
rect 19668 10452 19674 10464
rect 19886 10452 19892 10464
rect 19668 10424 19892 10452
rect 19668 10412 19674 10424
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 21361 10455 21419 10461
rect 21361 10452 21373 10455
rect 20312 10424 21373 10452
rect 20312 10412 20318 10424
rect 21361 10421 21373 10424
rect 21407 10421 21419 10455
rect 21361 10415 21419 10421
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 22557 10455 22615 10461
rect 22557 10452 22569 10455
rect 21600 10424 22569 10452
rect 21600 10412 21606 10424
rect 22557 10421 22569 10424
rect 22603 10421 22615 10455
rect 22557 10415 22615 10421
rect 1104 10362 23276 10384
rect 1104 10310 8379 10362
rect 8431 10310 8443 10362
rect 8495 10310 8507 10362
rect 8559 10310 8571 10362
rect 8623 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 15904 10362
rect 15956 10310 15968 10362
rect 16020 10310 23276 10362
rect 1104 10288 23276 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2590 10248 2596 10260
rect 1627 10220 2596 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 5534 10248 5540 10260
rect 5495 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 6972 10220 7205 10248
rect 6972 10208 6978 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 8938 10248 8944 10260
rect 7193 10211 7251 10217
rect 7760 10220 8944 10248
rect 4430 10189 4436 10192
rect 4424 10180 4436 10189
rect 2056 10152 2912 10180
rect 4391 10152 4436 10180
rect 1486 10072 1492 10124
rect 1544 10112 1550 10124
rect 2056 10121 2084 10152
rect 2041 10115 2099 10121
rect 2041 10112 2053 10115
rect 1544 10084 2053 10112
rect 1544 10072 1550 10084
rect 2041 10081 2053 10084
rect 2087 10081 2099 10115
rect 2041 10075 2099 10081
rect 2308 10115 2366 10121
rect 2308 10081 2320 10115
rect 2354 10112 2366 10115
rect 2774 10112 2780 10124
rect 2354 10084 2780 10112
rect 2354 10081 2366 10084
rect 2308 10075 2366 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 2884 10112 2912 10152
rect 4424 10143 4436 10152
rect 4430 10140 4436 10143
rect 4488 10140 4494 10192
rect 6080 10183 6138 10189
rect 6080 10149 6092 10183
rect 6126 10180 6138 10183
rect 6270 10180 6276 10192
rect 6126 10152 6276 10180
rect 6126 10149 6138 10152
rect 6080 10143 6138 10149
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 7760 10180 7788 10220
rect 8938 10208 8944 10220
rect 8996 10248 9002 10260
rect 8996 10220 10364 10248
rect 8996 10208 9002 10220
rect 7064 10152 7788 10180
rect 7837 10183 7895 10189
rect 7064 10140 7070 10152
rect 7837 10149 7849 10183
rect 7883 10180 7895 10183
rect 9674 10180 9680 10192
rect 7883 10152 9680 10180
rect 7883 10149 7895 10152
rect 7837 10143 7895 10149
rect 9674 10140 9680 10152
rect 9732 10140 9738 10192
rect 9944 10183 10002 10189
rect 9944 10149 9956 10183
rect 9990 10180 10002 10183
rect 10134 10180 10140 10192
rect 9990 10152 10140 10180
rect 9990 10149 10002 10152
rect 9944 10143 10002 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 10336 10180 10364 10220
rect 10410 10208 10416 10260
rect 10468 10248 10474 10260
rect 11333 10251 11391 10257
rect 11333 10248 11345 10251
rect 10468 10220 11345 10248
rect 10468 10208 10474 10220
rect 11333 10217 11345 10220
rect 11379 10217 11391 10251
rect 11333 10211 11391 10217
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 13446 10248 13452 10260
rect 12115 10220 13452 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 14553 10251 14611 10257
rect 14553 10217 14565 10251
rect 14599 10248 14611 10251
rect 15286 10248 15292 10260
rect 14599 10220 15292 10248
rect 14599 10217 14611 10220
rect 14553 10211 14611 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 16264 10220 16865 10248
rect 16264 10208 16270 10220
rect 16853 10217 16865 10220
rect 16899 10217 16911 10251
rect 21453 10251 21511 10257
rect 21453 10248 21465 10251
rect 16853 10211 16911 10217
rect 16960 10220 21465 10248
rect 12161 10183 12219 10189
rect 10336 10152 11560 10180
rect 3050 10112 3056 10124
rect 2884 10084 3056 10112
rect 3050 10072 3056 10084
rect 3108 10112 3114 10124
rect 3326 10112 3332 10124
rect 3108 10084 3332 10112
rect 3108 10072 3114 10084
rect 3326 10072 3332 10084
rect 3384 10112 3390 10124
rect 4157 10115 4215 10121
rect 4157 10112 4169 10115
rect 3384 10084 4169 10112
rect 3384 10072 3390 10084
rect 4157 10081 4169 10084
rect 4203 10112 4215 10115
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 4203 10084 5825 10112
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 5813 10081 5825 10084
rect 5859 10112 5871 10115
rect 6546 10112 6552 10124
rect 5859 10084 6552 10112
rect 5859 10081 5871 10084
rect 5813 10075 5871 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 8202 10121 8208 10124
rect 8185 10115 8208 10121
rect 8185 10112 8197 10115
rect 6972 10084 8197 10112
rect 6972 10072 6978 10084
rect 8185 10081 8197 10084
rect 8260 10112 8266 10124
rect 8260 10084 8333 10112
rect 8185 10075 8208 10081
rect 8202 10072 8208 10075
rect 8260 10072 8266 10084
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 11532 10121 11560 10152
rect 12161 10149 12173 10183
rect 12207 10180 12219 10183
rect 13722 10180 13728 10192
rect 12207 10152 13728 10180
rect 12207 10149 12219 10152
rect 12161 10143 12219 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 14642 10180 14648 10192
rect 14200 10152 14648 10180
rect 11517 10115 11575 10121
rect 10468 10084 10712 10112
rect 10468 10072 10474 10084
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 7883 10016 7941 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 7929 10013 7941 10016
rect 7975 10013 7987 10047
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 7929 10007 7987 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10684 10044 10712 10084
rect 11517 10081 11529 10115
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 12980 10115 13038 10121
rect 12980 10081 12992 10115
rect 13026 10112 13038 10115
rect 14200 10112 14228 10152
rect 14642 10140 14648 10152
rect 14700 10140 14706 10192
rect 15740 10183 15798 10189
rect 15740 10149 15752 10183
rect 15786 10180 15798 10183
rect 16390 10180 16396 10192
rect 15786 10152 16396 10180
rect 15786 10149 15798 10152
rect 15740 10143 15798 10149
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 16960 10180 16988 10220
rect 21453 10217 21465 10220
rect 21499 10217 21511 10251
rect 22278 10248 22284 10260
rect 22239 10220 22284 10248
rect 21453 10211 21511 10217
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 16632 10152 16988 10180
rect 17681 10183 17739 10189
rect 16632 10140 16638 10152
rect 17681 10149 17693 10183
rect 17727 10180 17739 10183
rect 19794 10180 19800 10192
rect 17727 10152 19800 10180
rect 17727 10149 17739 10152
rect 17681 10143 17739 10149
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 20806 10140 20812 10192
rect 20864 10180 20870 10192
rect 22189 10183 22247 10189
rect 22189 10180 22201 10183
rect 20864 10152 22201 10180
rect 20864 10140 20870 10152
rect 22189 10149 22201 10152
rect 22235 10149 22247 10183
rect 22189 10143 22247 10149
rect 13026 10084 14228 10112
rect 14369 10115 14427 10121
rect 13026 10081 13038 10084
rect 12980 10075 13038 10081
rect 14369 10081 14381 10115
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 12253 10047 12311 10053
rect 10684 10016 11744 10044
rect 11716 9985 11744 10016
rect 12253 10013 12265 10047
rect 12299 10013 12311 10047
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12253 10007 12311 10013
rect 11701 9979 11759 9985
rect 11701 9945 11713 9979
rect 11747 9945 11759 9979
rect 11701 9939 11759 9945
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 12268 9976 12296 10007
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 14384 10044 14412 10075
rect 14458 10072 14464 10124
rect 14516 10112 14522 10124
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 14516 10084 15117 10112
rect 14516 10072 14522 10084
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 16942 10112 16948 10124
rect 15105 10075 15163 10081
rect 15396 10084 16948 10112
rect 15396 10044 15424 10084
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10112 17647 10115
rect 17770 10112 17776 10124
rect 17635 10084 17776 10112
rect 17635 10081 17647 10084
rect 17589 10075 17647 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 18230 10112 18236 10124
rect 18191 10084 18236 10112
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 18500 10115 18558 10121
rect 18500 10081 18512 10115
rect 18546 10112 18558 10115
rect 18782 10112 18788 10124
rect 18546 10084 18788 10112
rect 18546 10081 18558 10084
rect 18500 10075 18558 10081
rect 18782 10072 18788 10084
rect 18840 10112 18846 10124
rect 19610 10112 19616 10124
rect 18840 10084 19616 10112
rect 18840 10072 18846 10084
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10112 19947 10115
rect 20438 10112 20444 10124
rect 19935 10084 20444 10112
rect 19935 10081 19947 10084
rect 19889 10075 19947 10081
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 20625 10115 20683 10121
rect 20625 10081 20637 10115
rect 20671 10112 20683 10115
rect 20990 10112 20996 10124
rect 20671 10084 20996 10112
rect 20671 10081 20683 10084
rect 20625 10075 20683 10081
rect 20990 10072 20996 10084
rect 21048 10072 21054 10124
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10112 21327 10115
rect 21450 10112 21456 10124
rect 21315 10084 21456 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 14384 10016 15424 10044
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10013 15531 10047
rect 17494 10044 17500 10056
rect 15473 10007 15531 10013
rect 16960 10016 17500 10044
rect 11940 9948 12296 9976
rect 11940 9936 11946 9948
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 15286 9976 15292 9988
rect 14240 9948 15292 9976
rect 14240 9936 14246 9948
rect 15286 9936 15292 9948
rect 15344 9976 15350 9988
rect 15488 9976 15516 10007
rect 15344 9948 15516 9976
rect 15344 9936 15350 9948
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3421 9911 3479 9917
rect 3421 9908 3433 9911
rect 3384 9880 3433 9908
rect 3384 9868 3390 9880
rect 3421 9877 3433 9880
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 8904 9880 9321 9908
rect 8904 9868 8910 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 11057 9911 11115 9917
rect 11057 9908 11069 9911
rect 10008 9880 11069 9908
rect 10008 9868 10014 9880
rect 11057 9877 11069 9880
rect 11103 9877 11115 9911
rect 11057 9871 11115 9877
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12986 9908 12992 9920
rect 12492 9880 12992 9908
rect 12492 9868 12498 9880
rect 12986 9868 12992 9880
rect 13044 9908 13050 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13044 9880 14105 9908
rect 13044 9868 13050 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14918 9908 14924 9920
rect 14879 9880 14924 9908
rect 14093 9871 14151 9877
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 15102 9868 15108 9920
rect 15160 9908 15166 9920
rect 16206 9908 16212 9920
rect 15160 9880 16212 9908
rect 15160 9868 15166 9880
rect 16206 9868 16212 9880
rect 16264 9908 16270 9920
rect 16960 9908 16988 10016
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17865 10047 17923 10053
rect 17865 10013 17877 10047
rect 17911 10044 17923 10047
rect 18046 10044 18052 10056
rect 17911 10016 18052 10044
rect 17911 10013 17923 10016
rect 17865 10007 17923 10013
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 19242 10004 19248 10056
rect 19300 10044 19306 10056
rect 22465 10047 22523 10053
rect 19300 10016 20760 10044
rect 19300 10004 19306 10016
rect 20456 9985 20484 10016
rect 20732 9988 20760 10016
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 22646 10044 22652 10056
rect 22511 10016 22652 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 20073 9979 20131 9985
rect 20073 9976 20085 9979
rect 19168 9948 20085 9976
rect 17218 9908 17224 9920
rect 16264 9880 16988 9908
rect 17179 9880 17224 9908
rect 16264 9868 16270 9880
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 18230 9868 18236 9920
rect 18288 9908 18294 9920
rect 19168 9908 19196 9948
rect 20073 9945 20085 9948
rect 20119 9945 20131 9979
rect 20073 9939 20131 9945
rect 20441 9979 20499 9985
rect 20441 9945 20453 9979
rect 20487 9945 20499 9979
rect 20441 9939 20499 9945
rect 20714 9936 20720 9988
rect 20772 9976 20778 9988
rect 21266 9976 21272 9988
rect 20772 9948 21272 9976
rect 20772 9936 20778 9948
rect 21266 9936 21272 9948
rect 21324 9936 21330 9988
rect 18288 9880 19196 9908
rect 18288 9868 18294 9880
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19392 9880 19625 9908
rect 19392 9868 19398 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 21821 9911 21879 9917
rect 21821 9908 21833 9911
rect 19944 9880 21833 9908
rect 19944 9868 19950 9880
rect 21821 9877 21833 9880
rect 21867 9877 21879 9911
rect 21821 9871 21879 9877
rect 1104 9818 23276 9840
rect 1104 9766 4680 9818
rect 4732 9766 4744 9818
rect 4796 9766 4808 9818
rect 4860 9766 4872 9818
rect 4924 9766 12078 9818
rect 12130 9766 12142 9818
rect 12194 9766 12206 9818
rect 12258 9766 12270 9818
rect 12322 9766 19475 9818
rect 19527 9766 19539 9818
rect 19591 9766 19603 9818
rect 19655 9766 19667 9818
rect 19719 9766 23276 9818
rect 1104 9744 23276 9766
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 4028 9676 5351 9704
rect 4028 9664 4034 9676
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 4433 9639 4491 9645
rect 2832 9608 2877 9636
rect 2832 9596 2838 9608
rect 4433 9605 4445 9639
rect 4479 9636 4491 9639
rect 4522 9636 4528 9648
rect 4479 9608 4528 9636
rect 4479 9605 4491 9608
rect 4433 9599 4491 9605
rect 4522 9596 4528 9608
rect 4580 9596 4586 9648
rect 5323 9636 5351 9676
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 7190 9704 7196 9716
rect 6328 9676 7196 9704
rect 6328 9664 6334 9676
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 15010 9704 15016 9716
rect 9732 9676 15016 9704
rect 9732 9664 9738 9676
rect 15010 9664 15016 9676
rect 15068 9704 15074 9716
rect 16574 9704 16580 9716
rect 15068 9676 16580 9704
rect 15068 9664 15074 9676
rect 16574 9664 16580 9676
rect 16632 9664 16638 9716
rect 16853 9707 16911 9713
rect 16853 9673 16865 9707
rect 16899 9704 16911 9707
rect 18138 9704 18144 9716
rect 16899 9676 18144 9704
rect 16899 9673 16911 9676
rect 16853 9667 16911 9673
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 18690 9664 18696 9716
rect 18748 9704 18754 9716
rect 18969 9707 19027 9713
rect 18969 9704 18981 9707
rect 18748 9676 18981 9704
rect 18748 9664 18754 9676
rect 18969 9673 18981 9676
rect 19015 9673 19027 9707
rect 18969 9667 19027 9673
rect 20622 9664 20628 9716
rect 20680 9704 20686 9716
rect 20990 9704 20996 9716
rect 20680 9676 20996 9704
rect 20680 9664 20686 9676
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 7009 9639 7067 9645
rect 7009 9636 7021 9639
rect 5323 9608 7021 9636
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 3050 9568 3056 9580
rect 3011 9540 3056 9568
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 5736 9577 5764 9608
rect 7009 9605 7021 9608
rect 7055 9605 7067 9639
rect 7009 9599 7067 9605
rect 7745 9639 7803 9645
rect 7745 9605 7757 9639
rect 7791 9636 7803 9639
rect 8754 9636 8760 9648
rect 7791 9608 8760 9636
rect 7791 9605 7803 9608
rect 7745 9599 7803 9605
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 11790 9636 11796 9648
rect 11751 9608 11796 9636
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 12069 9639 12127 9645
rect 12069 9605 12081 9639
rect 12115 9636 12127 9639
rect 12710 9636 12716 9648
rect 12115 9608 12716 9636
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 12710 9596 12716 9608
rect 12768 9596 12774 9648
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 13780 9608 14105 9636
rect 13780 9596 13786 9608
rect 14093 9605 14105 9608
rect 14139 9605 14151 9639
rect 14093 9599 14151 9605
rect 14369 9639 14427 9645
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 15102 9636 15108 9648
rect 14415 9608 15108 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 15102 9596 15108 9608
rect 15160 9596 15166 9648
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 16448 9608 16681 9636
rect 16448 9596 16454 9608
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 16942 9636 16948 9648
rect 16903 9608 16948 9636
rect 16669 9599 16727 9605
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 18230 9636 18236 9648
rect 17052 9608 18236 9636
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5592 9540 5641 9568
rect 5592 9528 5598 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9568 5779 9571
rect 5767 9540 5801 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 5902 9528 5908 9580
rect 5960 9568 5966 9580
rect 5960 9540 6868 9568
rect 5960 9528 5966 9540
rect 3326 9509 3332 9512
rect 3320 9500 3332 9509
rect 3287 9472 3332 9500
rect 3320 9463 3332 9472
rect 3326 9460 3332 9463
rect 3384 9460 3390 9512
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 5258 9500 5264 9512
rect 4948 9472 5264 9500
rect 4948 9460 4954 9472
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 6840 9509 6868 9540
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7650 9568 7656 9580
rect 7248 9540 7656 9568
rect 7248 9528 7254 9540
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8386 9568 8392 9580
rect 8260 9540 8392 9568
rect 8260 9528 8266 9540
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 10226 9568 10232 9580
rect 9784 9540 10232 9568
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9469 6239 9503
rect 6181 9463 6239 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 1486 9392 1492 9444
rect 1544 9432 1550 9444
rect 1642 9435 1700 9441
rect 1642 9432 1654 9435
rect 1544 9404 1654 9432
rect 1544 9392 1550 9404
rect 1642 9401 1654 9404
rect 1688 9401 1700 9435
rect 1642 9395 1700 9401
rect 3694 9392 3700 9444
rect 3752 9432 3758 9444
rect 5537 9435 5595 9441
rect 3752 9404 5396 9432
rect 3752 9392 3758 9404
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5368 9364 5396 9404
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 5718 9432 5724 9444
rect 5583 9404 5724 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 6196 9432 6224 9463
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8110 9500 8116 9512
rect 7984 9472 8116 9500
rect 7984 9460 7990 9472
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9784 9500 9812 9540
rect 10226 9528 10232 9540
rect 10284 9568 10290 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 10284 9540 10425 9568
rect 10284 9528 10290 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 17052 9568 17080 9608
rect 18230 9596 18236 9608
rect 18288 9596 18294 9648
rect 19150 9596 19156 9648
rect 19208 9596 19214 9648
rect 22741 9639 22799 9645
rect 22741 9605 22753 9639
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 16356 9540 17080 9568
rect 17589 9571 17647 9577
rect 16356 9528 16362 9540
rect 17589 9537 17601 9571
rect 17635 9568 17647 9571
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17635 9540 17877 9568
rect 17635 9537 17647 9540
rect 17589 9531 17647 9537
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 18785 9571 18843 9577
rect 17865 9531 17923 9537
rect 17972 9540 18552 9568
rect 8803 9472 9812 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 10669 9503 10727 9509
rect 10669 9500 10681 9503
rect 9916 9472 10681 9500
rect 9916 9460 9922 9472
rect 10669 9469 10681 9472
rect 10715 9500 10727 9503
rect 10962 9500 10968 9512
rect 10715 9472 10968 9500
rect 10715 9469 10727 9472
rect 10669 9463 10727 9469
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12618 9500 12624 9512
rect 12299 9472 12624 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12710 9460 12716 9512
rect 12768 9500 12774 9512
rect 13354 9500 13360 9512
rect 12768 9472 13360 9500
rect 12768 9460 12774 9472
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 13872 9472 14565 9500
rect 13872 9460 13878 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 14645 9503 14703 9509
rect 14645 9469 14657 9503
rect 14691 9500 14703 9503
rect 14691 9472 15240 9500
rect 14691 9469 14703 9472
rect 14645 9463 14703 9469
rect 6196 9404 6868 9432
rect 6840 9376 6868 9404
rect 7650 9392 7656 9444
rect 7708 9432 7714 9444
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 7708 9404 8217 9432
rect 7708 9392 7714 9404
rect 8205 9401 8217 9404
rect 8251 9401 8263 9435
rect 8205 9395 8263 9401
rect 8846 9392 8852 9444
rect 8904 9432 8910 9444
rect 9002 9435 9060 9441
rect 9002 9432 9014 9435
rect 8904 9404 9014 9432
rect 8904 9392 8910 9404
rect 9002 9401 9014 9404
rect 9048 9401 9060 9435
rect 9002 9395 9060 9401
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 9674 9432 9680 9444
rect 9548 9404 9680 9432
rect 9548 9392 9554 9404
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 9824 9404 10456 9432
rect 9824 9392 9830 9404
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 5368 9336 6377 9364
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 6822 9324 6828 9376
rect 6880 9324 6886 9376
rect 8110 9364 8116 9376
rect 8071 9336 8116 9364
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10428 9364 10456 9404
rect 10502 9392 10508 9444
rect 10560 9432 10566 9444
rect 11146 9432 11152 9444
rect 10560 9404 11152 9432
rect 10560 9392 10566 9404
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 12342 9392 12348 9444
rect 12400 9432 12406 9444
rect 12958 9435 13016 9441
rect 12958 9432 12970 9435
rect 12400 9404 12970 9432
rect 12400 9392 12406 9404
rect 12958 9401 12970 9404
rect 13004 9401 13016 9435
rect 12958 9395 13016 9401
rect 14829 9435 14887 9441
rect 14829 9401 14841 9435
rect 14875 9432 14887 9435
rect 15102 9432 15108 9444
rect 14875 9404 15108 9432
rect 14875 9401 14887 9404
rect 14829 9395 14887 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 10686 9364 10692 9376
rect 10428 9336 10692 9364
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14366 9364 14372 9376
rect 13964 9336 14372 9364
rect 13964 9324 13970 9336
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 15010 9364 15016 9376
rect 14971 9336 15016 9364
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 15212 9364 15240 9472
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15556 9503 15614 9509
rect 15344 9472 15437 9500
rect 15344 9460 15350 9472
rect 15556 9469 15568 9503
rect 15602 9500 15614 9503
rect 16942 9500 16948 9512
rect 15602 9472 16948 9500
rect 15602 9469 15614 9472
rect 15556 9463 15614 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17972 9500 18000 9540
rect 18524 9509 18552 9540
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 19168 9568 19196 9596
rect 19334 9568 19340 9580
rect 18831 9540 19340 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19702 9577 19708 9580
rect 19659 9571 19708 9577
rect 19659 9537 19671 9571
rect 19705 9537 19708 9571
rect 19659 9531 19708 9537
rect 19702 9528 19708 9531
rect 19760 9528 19766 9580
rect 19794 9528 19800 9580
rect 19852 9568 19858 9580
rect 19889 9571 19947 9577
rect 19889 9568 19901 9571
rect 19852 9540 19901 9568
rect 19852 9528 19858 9540
rect 19889 9537 19901 9540
rect 19935 9537 19947 9571
rect 19889 9531 19947 9537
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 21266 9568 21272 9580
rect 20772 9540 21272 9568
rect 20772 9528 20778 9540
rect 21266 9528 21272 9540
rect 21324 9568 21330 9580
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 21324 9540 21373 9568
rect 21324 9528 21330 9540
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 17052 9472 18000 9500
rect 18509 9503 18567 9509
rect 15304 9432 15332 9460
rect 16390 9432 16396 9444
rect 15304 9404 16396 9432
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 16574 9392 16580 9444
rect 16632 9432 16638 9444
rect 17052 9432 17080 9472
rect 18509 9469 18521 9503
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 19153 9503 19211 9509
rect 18656 9472 18701 9500
rect 18656 9460 18662 9472
rect 19153 9469 19165 9503
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 16632 9404 17080 9432
rect 17405 9435 17463 9441
rect 16632 9392 16638 9404
rect 17405 9401 17417 9435
rect 17451 9432 17463 9435
rect 17451 9404 18368 9432
rect 17451 9401 17463 9404
rect 17405 9395 17463 9401
rect 16853 9367 16911 9373
rect 16853 9364 16865 9367
rect 15212 9336 16865 9364
rect 16853 9333 16865 9336
rect 16899 9333 16911 9367
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 16853 9327 16911 9333
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17862 9364 17868 9376
rect 17823 9336 17868 9364
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18138 9364 18144 9376
rect 18099 9336 18144 9364
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 18340 9364 18368 9404
rect 18414 9392 18420 9444
rect 18472 9432 18478 9444
rect 19168 9432 19196 9463
rect 19426 9460 19432 9512
rect 19484 9509 19490 9512
rect 19484 9503 19534 9509
rect 19484 9469 19488 9503
rect 19522 9469 19534 9503
rect 19484 9463 19534 9469
rect 19484 9460 19490 9463
rect 19978 9460 19984 9512
rect 20036 9500 20042 9512
rect 22756 9500 22784 9599
rect 20036 9472 22784 9500
rect 20036 9460 20042 9472
rect 18472 9404 19196 9432
rect 21628 9435 21686 9441
rect 18472 9392 18478 9404
rect 21628 9401 21640 9435
rect 21674 9432 21686 9435
rect 22646 9432 22652 9444
rect 21674 9404 22652 9432
rect 21674 9401 21686 9404
rect 21628 9395 21686 9401
rect 22646 9392 22652 9404
rect 22704 9392 22710 9444
rect 18969 9367 19027 9373
rect 18969 9364 18981 9367
rect 18340 9336 18981 9364
rect 18969 9333 18981 9336
rect 19015 9364 19027 9367
rect 20993 9367 21051 9373
rect 20993 9364 21005 9367
rect 19015 9336 21005 9364
rect 19015 9333 19027 9336
rect 18969 9327 19027 9333
rect 20993 9333 21005 9336
rect 21039 9333 21051 9367
rect 20993 9327 21051 9333
rect 1104 9274 23276 9296
rect 1104 9222 8379 9274
rect 8431 9222 8443 9274
rect 8495 9222 8507 9274
rect 8559 9222 8571 9274
rect 8623 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 15904 9274
rect 15956 9222 15968 9274
rect 16020 9222 23276 9274
rect 1104 9200 23276 9222
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9160 2283 9163
rect 2406 9160 2412 9172
rect 2271 9132 2412 9160
rect 2271 9129 2283 9132
rect 2225 9123 2283 9129
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3326 9160 3332 9172
rect 3283 9132 3332 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 4062 9160 4068 9172
rect 4023 9132 4068 9160
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4396 9132 4445 9160
rect 4396 9120 4402 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 5077 9163 5135 9169
rect 5077 9160 5089 9163
rect 4948 9132 5089 9160
rect 4948 9120 4954 9132
rect 5077 9129 5089 9132
rect 5123 9129 5135 9163
rect 5077 9123 5135 9129
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 5408 9132 5457 9160
rect 5408 9120 5414 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6365 9163 6423 9169
rect 6365 9160 6377 9163
rect 6144 9132 6377 9160
rect 6144 9120 6150 9132
rect 6365 9129 6377 9132
rect 6411 9160 6423 9163
rect 6917 9163 6975 9169
rect 6917 9160 6929 9163
rect 6411 9132 6929 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 6917 9129 6929 9132
rect 6963 9160 6975 9163
rect 7377 9163 7435 9169
rect 7377 9160 7389 9163
rect 6963 9132 7389 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7377 9129 7389 9132
rect 7423 9129 7435 9163
rect 7377 9123 7435 9129
rect 7561 9163 7619 9169
rect 7561 9129 7573 9163
rect 7607 9160 7619 9163
rect 7742 9160 7748 9172
rect 7607 9132 7748 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 9306 9160 9312 9172
rect 8036 9132 9312 9160
rect 1946 9052 1952 9104
rect 2004 9092 2010 9104
rect 2004 9064 4936 9092
rect 2004 9052 2010 9064
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3329 9027 3387 9033
rect 3329 9024 3341 9027
rect 2832 8996 3341 9024
rect 2832 8984 2838 8996
rect 3329 8993 3341 8996
rect 3375 8993 3387 9027
rect 4908 9024 4936 9064
rect 5258 9052 5264 9104
rect 5316 9092 5322 9104
rect 5537 9095 5595 9101
rect 5537 9092 5549 9095
rect 5316 9064 5549 9092
rect 5316 9052 5322 9064
rect 5537 9061 5549 9064
rect 5583 9061 5595 9095
rect 7009 9095 7067 9101
rect 7009 9092 7021 9095
rect 5537 9055 5595 9061
rect 5644 9064 7021 9092
rect 5644 9024 5672 9064
rect 7009 9061 7021 9064
rect 7055 9061 7067 9095
rect 7929 9095 7987 9101
rect 7929 9092 7941 9095
rect 7009 9055 7067 9061
rect 7116 9064 7941 9092
rect 4908 8996 5672 9024
rect 3329 8987 3387 8993
rect 6178 8984 6184 9036
rect 6236 8984 6242 9036
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2958 8956 2964 8968
rect 2547 8928 2964 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 3970 8956 3976 8968
rect 3559 8928 3976 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 4663 8928 5733 8956
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 5721 8925 5733 8928
rect 5767 8956 5779 8959
rect 6196 8956 6224 8984
rect 5767 8928 6224 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 4540 8888 4568 8919
rect 2915 8860 4568 8888
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8820 1915 8823
rect 3602 8820 3608 8832
rect 1903 8792 3608 8820
rect 1903 8789 1915 8792
rect 1857 8783 1915 8789
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 4632 8820 4660 8919
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7116 8956 7144 9064
rect 7929 9061 7941 9064
rect 7975 9061 7987 9095
rect 7929 9055 7987 9061
rect 8036 9024 8064 9132
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9766 9160 9772 9172
rect 9723 9132 9772 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10410 9160 10416 9172
rect 10060 9132 10416 9160
rect 9033 9095 9091 9101
rect 9033 9061 9045 9095
rect 9079 9092 9091 9095
rect 9493 9095 9551 9101
rect 9493 9092 9505 9095
rect 9079 9064 9505 9092
rect 9079 9061 9091 9064
rect 9033 9055 9091 9061
rect 9493 9061 9505 9064
rect 9539 9061 9551 9095
rect 10060 9092 10088 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 12529 9163 12587 9169
rect 12529 9160 12541 9163
rect 10643 9132 12541 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 12529 9129 12541 9132
rect 12575 9129 12587 9163
rect 13354 9160 13360 9172
rect 13267 9132 13360 9160
rect 12529 9123 12587 9129
rect 13354 9120 13360 9132
rect 13412 9160 13418 9172
rect 14182 9160 14188 9172
rect 13412 9132 14188 9160
rect 13412 9120 13418 9132
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 17218 9160 17224 9172
rect 15979 9132 17224 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 22646 9160 22652 9172
rect 17920 9132 20392 9160
rect 22607 9132 22652 9160
rect 17920 9120 17926 9132
rect 9493 9055 9551 9061
rect 9600 9064 10088 9092
rect 10137 9095 10195 9101
rect 7944 8996 8064 9024
rect 8941 9027 8999 9033
rect 6880 8928 7144 8956
rect 7193 8959 7251 8965
rect 6880 8916 6886 8928
rect 7193 8925 7205 8959
rect 7239 8956 7251 8959
rect 7944 8956 7972 8996
rect 8941 8993 8953 9027
rect 8987 9024 8999 9027
rect 9600 9024 9628 9064
rect 10137 9061 10149 9095
rect 10183 9092 10195 9095
rect 11057 9095 11115 9101
rect 10183 9064 10640 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 8987 8996 9628 9024
rect 10045 9027 10103 9033
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10091 8996 10447 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 7239 8928 7972 8956
rect 8021 8959 8079 8965
rect 7239 8925 7251 8928
rect 7193 8919 7251 8925
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8202 8956 8208 8968
rect 8163 8928 8208 8956
rect 8021 8919 8079 8925
rect 6178 8848 6184 8900
rect 6236 8848 6242 8900
rect 8036 8888 8064 8919
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 9030 8956 9036 8968
rect 8628 8928 9036 8956
rect 8628 8916 8634 8928
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9263 8928 10171 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 10042 8888 10048 8900
rect 6380 8860 8064 8888
rect 8220 8860 10048 8888
rect 3752 8792 4660 8820
rect 6196 8820 6224 8848
rect 6380 8820 6408 8860
rect 8220 8832 8248 8860
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 10143 8888 10171 8928
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 10284 8928 10329 8956
rect 10284 8916 10290 8928
rect 10244 8888 10272 8916
rect 10143 8860 10272 8888
rect 10419 8888 10447 8996
rect 10612 8956 10640 9064
rect 11057 9061 11069 9095
rect 11103 9092 11115 9095
rect 11146 9092 11152 9104
rect 11103 9064 11152 9092
rect 11103 9061 11115 9064
rect 11057 9055 11115 9061
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 12342 9052 12348 9104
rect 12400 9092 12406 9104
rect 12897 9095 12955 9101
rect 12897 9092 12909 9095
rect 12400 9064 12909 9092
rect 12400 9052 12406 9064
rect 12897 9061 12909 9064
rect 12943 9092 12955 9095
rect 14366 9092 14372 9104
rect 12943 9064 14372 9092
rect 12943 9061 12955 9064
rect 12897 9055 12955 9061
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 14458 9052 14464 9104
rect 14516 9092 14522 9104
rect 16298 9092 16304 9104
rect 14516 9064 16304 9092
rect 14516 9052 14522 9064
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 20364 9092 20392 9132
rect 22646 9120 22652 9132
rect 22704 9120 22710 9172
rect 21514 9095 21572 9101
rect 21514 9092 21526 9095
rect 20364 9064 21526 9092
rect 21514 9061 21526 9064
rect 21560 9092 21572 9095
rect 22186 9092 22192 9104
rect 21560 9064 22192 9092
rect 21560 9061 21572 9064
rect 21514 9055 21572 9061
rect 22186 9052 22192 9064
rect 22244 9052 22250 9104
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 10744 8996 11713 9024
rect 10744 8984 10750 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 12437 9027 12495 9033
rect 12437 8993 12449 9027
rect 12483 9024 12495 9027
rect 12989 9027 13047 9033
rect 12483 8996 12940 9024
rect 12483 8993 12495 8996
rect 12437 8987 12495 8993
rect 12912 8968 12940 8996
rect 12989 8993 13001 9027
rect 13035 9024 13047 9027
rect 13262 9024 13268 9036
rect 13035 8996 13268 9024
rect 13035 8993 13047 8996
rect 12989 8987 13047 8993
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13446 8984 13452 9036
rect 13504 9024 13510 9036
rect 13797 9027 13855 9033
rect 13797 9024 13809 9027
rect 13504 8996 13809 9024
rect 13504 8984 13510 8996
rect 13797 8993 13809 8996
rect 13843 8993 13855 9027
rect 15838 9024 15844 9036
rect 15799 8996 15844 9024
rect 13797 8987 13855 8993
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16448 8996 16497 9024
rect 16448 8984 16454 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16741 9027 16799 9033
rect 16741 9024 16753 9027
rect 16632 8996 16753 9024
rect 16632 8984 16638 8996
rect 16741 8993 16753 8996
rect 16787 8993 16799 9027
rect 16741 8987 16799 8993
rect 17310 8984 17316 9036
rect 17368 9024 17374 9036
rect 17368 8996 18000 9024
rect 17368 8984 17374 8996
rect 11146 8956 11152 8968
rect 10612 8928 11008 8956
rect 11107 8928 11152 8956
rect 10689 8891 10747 8897
rect 10689 8888 10701 8891
rect 10419 8860 10701 8888
rect 10689 8857 10701 8860
rect 10735 8857 10747 8891
rect 10980 8888 11008 8928
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11882 8956 11888 8968
rect 11287 8928 11888 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11882 8916 11888 8928
rect 11940 8956 11946 8968
rect 11940 8928 12848 8956
rect 11940 8916 11946 8928
rect 11330 8888 11336 8900
rect 10980 8860 11336 8888
rect 10689 8851 10747 8857
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 12820 8888 12848 8928
rect 12894 8916 12900 8968
rect 12952 8916 12958 8968
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 13403 8928 13553 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8956 16175 8959
rect 16298 8956 16304 8968
rect 16163 8928 16304 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 13096 8888 13124 8919
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 12820 8860 13124 8888
rect 14844 8860 16528 8888
rect 6546 8820 6552 8832
rect 6196 8792 6408 8820
rect 6507 8792 6552 8820
rect 3752 8780 3758 8792
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8018 8820 8024 8832
rect 7800 8792 8024 8820
rect 7800 8780 7806 8792
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8202 8780 8208 8832
rect 8260 8780 8266 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 9030 8820 9036 8832
rect 8619 8792 9036 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 9539 8792 10609 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10597 8783 10655 8789
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11848 8792 11897 8820
rect 11848 8780 11854 8792
rect 11885 8789 11897 8792
rect 11931 8789 11943 8823
rect 11885 8783 11943 8789
rect 12253 8823 12311 8829
rect 12253 8789 12265 8823
rect 12299 8820 12311 8823
rect 12710 8820 12716 8832
rect 12299 8792 12716 8820
rect 12299 8789 12311 8792
rect 12253 8783 12311 8789
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 14844 8820 14872 8860
rect 12952 8792 14872 8820
rect 14921 8823 14979 8829
rect 12952 8780 12958 8792
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15102 8820 15108 8832
rect 14967 8792 15108 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15102 8780 15108 8792
rect 15160 8820 15166 8832
rect 15286 8820 15292 8832
rect 15160 8792 15292 8820
rect 15160 8780 15166 8792
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15473 8823 15531 8829
rect 15473 8789 15485 8823
rect 15519 8820 15531 8823
rect 15562 8820 15568 8832
rect 15519 8792 15568 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 15562 8780 15568 8792
rect 15620 8820 15626 8832
rect 16390 8820 16396 8832
rect 15620 8792 16396 8820
rect 15620 8780 15626 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 16500 8820 16528 8860
rect 17126 8820 17132 8832
rect 16500 8792 17132 8820
rect 17126 8780 17132 8792
rect 17184 8780 17190 8832
rect 17862 8820 17868 8832
rect 17823 8792 17868 8820
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 17972 8820 18000 8996
rect 18138 8984 18144 9036
rect 18196 9024 18202 9036
rect 18196 8996 18831 9024
rect 18196 8984 18202 8996
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18288 8928 18337 8956
rect 18288 8916 18294 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 18803 8965 18831 8996
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 20625 9027 20683 9033
rect 20625 9024 20637 9027
rect 19392 8996 20637 9024
rect 19392 8984 19398 8996
rect 20625 8993 20637 8996
rect 20671 8993 20683 9027
rect 21266 9024 21272 9036
rect 21227 8996 21272 9024
rect 20625 8987 20683 8993
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 18648 8959 18706 8965
rect 18648 8956 18660 8959
rect 18564 8928 18660 8956
rect 18564 8916 18570 8928
rect 18648 8925 18660 8928
rect 18694 8925 18706 8959
rect 18648 8919 18706 8925
rect 18788 8959 18846 8965
rect 18788 8925 18800 8959
rect 18834 8925 18846 8959
rect 18788 8919 18846 8925
rect 19061 8959 19119 8965
rect 19061 8925 19073 8959
rect 19107 8956 19119 8959
rect 20070 8956 20076 8968
rect 19107 8928 20076 8956
rect 19107 8925 19119 8928
rect 19061 8919 19119 8925
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 19702 8848 19708 8900
rect 19760 8848 19766 8900
rect 19794 8848 19800 8900
rect 19852 8888 19858 8900
rect 20165 8891 20223 8897
rect 20165 8888 20177 8891
rect 19852 8860 20177 8888
rect 19852 8848 19858 8860
rect 20165 8857 20177 8860
rect 20211 8857 20223 8891
rect 20165 8851 20223 8857
rect 19720 8820 19748 8848
rect 17972 8792 19748 8820
rect 19978 8780 19984 8832
rect 20036 8820 20042 8832
rect 20441 8823 20499 8829
rect 20441 8820 20453 8823
rect 20036 8792 20453 8820
rect 20036 8780 20042 8792
rect 20441 8789 20453 8792
rect 20487 8820 20499 8823
rect 20622 8820 20628 8832
rect 20487 8792 20628 8820
rect 20487 8789 20499 8792
rect 20441 8783 20499 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 22370 8780 22376 8832
rect 22428 8820 22434 8832
rect 23014 8820 23020 8832
rect 22428 8792 23020 8820
rect 22428 8780 22434 8792
rect 23014 8780 23020 8792
rect 23072 8780 23078 8832
rect 1104 8730 23276 8752
rect 1104 8678 4680 8730
rect 4732 8678 4744 8730
rect 4796 8678 4808 8730
rect 4860 8678 4872 8730
rect 4924 8678 12078 8730
rect 12130 8678 12142 8730
rect 12194 8678 12206 8730
rect 12258 8678 12270 8730
rect 12322 8678 19475 8730
rect 19527 8678 19539 8730
rect 19591 8678 19603 8730
rect 19655 8678 19667 8730
rect 19719 8678 23276 8730
rect 1104 8656 23276 8678
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 5074 8616 5080 8628
rect 4755 8588 5080 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 5074 8576 5080 8588
rect 5132 8576 5138 8628
rect 8570 8616 8576 8628
rect 7576 8588 8576 8616
rect 2314 8508 2320 8560
rect 2372 8548 2378 8560
rect 5721 8551 5779 8557
rect 2372 8520 5488 8548
rect 2372 8508 2378 8520
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 3200 8452 3341 8480
rect 3200 8440 3206 8452
rect 3329 8449 3341 8452
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 3694 8480 3700 8492
rect 3559 8452 3700 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 5166 8480 5172 8492
rect 5127 8452 5172 8480
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5350 8480 5356 8492
rect 5311 8452 5356 8480
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 5460 8480 5488 8520
rect 5721 8517 5733 8551
rect 5767 8548 5779 8551
rect 7006 8548 7012 8560
rect 5767 8520 7012 8548
rect 5767 8517 5779 8520
rect 5721 8511 5779 8517
rect 7006 8508 7012 8520
rect 7064 8508 7070 8560
rect 6365 8483 6423 8489
rect 5460 8452 5764 8480
rect 5736 8424 5764 8452
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 7576 8480 7604 8588
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 15102 8616 15108 8628
rect 9088 8588 15108 8616
rect 9088 8576 9094 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15378 8616 15384 8628
rect 15243 8588 15384 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 18141 8619 18199 8625
rect 15896 8588 18092 8616
rect 15896 8576 15902 8588
rect 7653 8551 7711 8557
rect 7653 8517 7665 8551
rect 7699 8548 7711 8551
rect 8478 8548 8484 8560
rect 7699 8520 8484 8548
rect 7699 8517 7711 8520
rect 7653 8511 7711 8517
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 8665 8551 8723 8557
rect 8665 8517 8677 8551
rect 8711 8548 8723 8551
rect 9122 8548 9128 8560
rect 8711 8520 9128 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 9674 8548 9680 8560
rect 9600 8520 9680 8548
rect 6411 8452 7604 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 8113 8483 8171 8489
rect 8113 8480 8125 8483
rect 8076 8452 8125 8480
rect 8076 8440 8082 8452
rect 8113 8449 8125 8452
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8202 8440 8208 8492
rect 8260 8480 8266 8492
rect 8260 8452 8305 8480
rect 8260 8440 8266 8452
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9490 8480 9496 8492
rect 9355 8452 9496 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 3234 8412 3240 8424
rect 3195 8384 3240 8412
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 5077 8415 5135 8421
rect 5077 8381 5089 8415
rect 5123 8412 5135 8415
rect 5534 8412 5540 8424
rect 5123 8384 5540 8412
rect 5123 8381 5135 8384
rect 5077 8375 5135 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5718 8372 5724 8424
rect 5776 8372 5782 8424
rect 6086 8412 6092 8424
rect 6047 8384 6092 8412
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 8404 8412 8432 8440
rect 7147 8384 8432 8412
rect 9033 8415 9091 8421
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9600 8412 9628 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 11149 8551 11207 8557
rect 11149 8548 11161 8551
rect 10695 8520 11161 8548
rect 9079 8384 9628 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10695 8412 10723 8520
rect 11149 8517 11161 8520
rect 11195 8517 11207 8551
rect 11330 8548 11336 8560
rect 11291 8520 11336 8548
rect 11149 8511 11207 8517
rect 11330 8508 11336 8520
rect 11388 8508 11394 8560
rect 12989 8551 13047 8557
rect 12989 8517 13001 8551
rect 13035 8548 13047 8551
rect 13078 8548 13084 8560
rect 13035 8520 13084 8548
rect 13035 8517 13047 8520
rect 12989 8511 13047 8517
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 14737 8551 14795 8557
rect 14737 8548 14749 8551
rect 14384 8520 14749 8548
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11238 8480 11244 8492
rect 10836 8452 11244 8480
rect 10836 8440 10842 8452
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11882 8480 11888 8492
rect 11843 8452 11888 8480
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 13354 8480 13360 8492
rect 13315 8452 13360 8480
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 9732 8384 9777 8412
rect 9876 8384 10723 8412
rect 11149 8415 11207 8421
rect 9732 8372 9738 8384
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 6104 8316 6193 8344
rect 6104 8288 6132 8316
rect 6181 8313 6193 8316
rect 6227 8344 6239 8347
rect 6546 8344 6552 8356
rect 6227 8316 6552 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 8294 8344 8300 8356
rect 7300 8316 8300 8344
rect 6086 8236 6092 8288
rect 6144 8236 6150 8288
rect 7300 8285 7328 8316
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 9125 8347 9183 8353
rect 9125 8313 9137 8347
rect 9171 8344 9183 8347
rect 9876 8344 9904 8384
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 11790 8412 11796 8424
rect 11195 8384 11796 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12802 8412 12808 8424
rect 12763 8384 12808 8412
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 13446 8372 13452 8424
rect 13504 8412 13510 8424
rect 14384 8412 14412 8520
rect 14737 8517 14749 8520
rect 14783 8517 14795 8551
rect 14737 8511 14795 8517
rect 15562 8480 15568 8492
rect 15523 8452 15568 8480
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8480 17555 8483
rect 17954 8480 17960 8492
rect 17543 8452 17960 8480
rect 17543 8449 17555 8452
rect 17497 8443 17555 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18064 8480 18092 8588
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18598 8616 18604 8628
rect 18187 8588 18604 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 18708 8588 20545 8616
rect 18414 8508 18420 8560
rect 18472 8548 18478 8560
rect 18708 8548 18736 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 22186 8616 22192 8628
rect 22147 8588 22192 8616
rect 20533 8579 20591 8585
rect 18472 8520 18736 8548
rect 18472 8508 18478 8520
rect 18064 8452 18736 8480
rect 15010 8412 15016 8424
rect 13504 8384 14412 8412
rect 14971 8384 15016 8412
rect 13504 8372 13510 8384
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 15286 8372 15292 8424
rect 15344 8412 15350 8424
rect 15821 8415 15879 8421
rect 15821 8412 15833 8415
rect 15344 8384 15833 8412
rect 15344 8372 15350 8384
rect 15821 8381 15833 8384
rect 15867 8381 15879 8415
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 15821 8375 15879 8381
rect 16868 8384 17233 8412
rect 9171 8316 9904 8344
rect 9944 8347 10002 8353
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 9944 8313 9956 8347
rect 9990 8344 10002 8347
rect 11701 8347 11759 8353
rect 11701 8344 11713 8347
rect 9990 8316 11713 8344
rect 9990 8313 10002 8316
rect 9944 8307 10002 8313
rect 11701 8313 11713 8316
rect 11747 8344 11759 8347
rect 12618 8344 12624 8356
rect 11747 8316 12624 8344
rect 11747 8313 11759 8316
rect 11701 8307 11759 8313
rect 12618 8304 12624 8316
rect 12676 8304 12682 8356
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 13624 8347 13682 8353
rect 12768 8316 13584 8344
rect 12768 8304 12774 8316
rect 7285 8279 7343 8285
rect 7285 8245 7297 8279
rect 7331 8245 7343 8279
rect 7285 8239 7343 8245
rect 8021 8279 8079 8285
rect 8021 8245 8033 8279
rect 8067 8276 8079 8279
rect 10042 8276 10048 8288
rect 8067 8248 10048 8276
rect 8067 8245 8079 8248
rect 8021 8239 8079 8245
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 10226 8236 10232 8288
rect 10284 8276 10290 8288
rect 10962 8276 10968 8288
rect 10284 8248 10968 8276
rect 10284 8236 10290 8248
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 11057 8279 11115 8285
rect 11057 8245 11069 8279
rect 11103 8276 11115 8279
rect 11146 8276 11152 8288
rect 11103 8248 11152 8276
rect 11103 8245 11115 8248
rect 11057 8239 11115 8245
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 11793 8279 11851 8285
rect 11793 8276 11805 8279
rect 11296 8248 11805 8276
rect 11296 8236 11302 8248
rect 11793 8245 11805 8248
rect 11839 8245 11851 8279
rect 11793 8239 11851 8245
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13078 8276 13084 8288
rect 12952 8248 13084 8276
rect 12952 8236 12958 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 13556 8276 13584 8316
rect 13624 8313 13636 8347
rect 13670 8344 13682 8347
rect 13814 8344 13820 8356
rect 13670 8316 13820 8344
rect 13670 8313 13682 8316
rect 13624 8307 13682 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 14550 8344 14556 8356
rect 13924 8316 14556 8344
rect 13924 8276 13952 8316
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 13556 8248 13952 8276
rect 14182 8236 14188 8288
rect 14240 8276 14246 8288
rect 16868 8276 16896 8384
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 17236 8344 17264 8375
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 17770 8412 17776 8424
rect 17460 8384 17776 8412
rect 17460 8372 17466 8384
rect 17770 8372 17776 8384
rect 17828 8412 17834 8424
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 17828 8384 18613 8412
rect 17828 8372 17834 8384
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18708 8412 18736 8452
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 20548 8480 20576 8579
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 22370 8508 22376 8560
rect 22428 8548 22434 8560
rect 22649 8551 22707 8557
rect 22649 8548 22661 8551
rect 22428 8520 22661 8548
rect 22428 8508 22434 8520
rect 22649 8517 22661 8520
rect 22695 8517 22707 8551
rect 22649 8511 22707 8517
rect 18840 8452 18885 8480
rect 18984 8452 19279 8480
rect 20548 8452 20944 8480
rect 18840 8440 18846 8452
rect 18984 8412 19012 8452
rect 18708 8384 19012 8412
rect 18601 8375 18659 8381
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 19116 8384 19165 8412
rect 19116 8372 19122 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19251 8412 19279 8452
rect 20162 8412 20168 8424
rect 19251 8384 20168 8412
rect 19153 8375 19211 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 20809 8415 20867 8421
rect 20809 8412 20821 8415
rect 20772 8384 20821 8412
rect 20772 8372 20778 8384
rect 20809 8381 20821 8384
rect 20855 8381 20867 8415
rect 20916 8412 20944 8452
rect 21065 8415 21123 8421
rect 21065 8412 21077 8415
rect 20916 8384 21077 8412
rect 20809 8375 20867 8381
rect 21065 8381 21077 8384
rect 21111 8381 21123 8415
rect 21065 8375 21123 8381
rect 22278 8372 22284 8424
rect 22336 8412 22342 8424
rect 22465 8415 22523 8421
rect 22465 8412 22477 8415
rect 22336 8384 22477 8412
rect 22336 8372 22342 8384
rect 22465 8381 22477 8384
rect 22511 8381 22523 8415
rect 22465 8375 22523 8381
rect 17494 8344 17500 8356
rect 17236 8316 17500 8344
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 18046 8304 18052 8356
rect 18104 8344 18110 8356
rect 19242 8344 19248 8356
rect 18104 8316 19248 8344
rect 18104 8304 18110 8316
rect 19242 8304 19248 8316
rect 19300 8344 19306 8356
rect 19398 8347 19456 8353
rect 19398 8344 19410 8347
rect 19300 8316 19410 8344
rect 19300 8304 19306 8316
rect 19398 8313 19410 8316
rect 19444 8313 19456 8347
rect 19398 8307 19456 8313
rect 20346 8304 20352 8356
rect 20404 8344 20410 8356
rect 20622 8344 20628 8356
rect 20404 8316 20628 8344
rect 20404 8304 20410 8316
rect 20622 8304 20628 8316
rect 20680 8304 20686 8356
rect 14240 8248 16896 8276
rect 16945 8279 17003 8285
rect 14240 8236 14246 8248
rect 16945 8245 16957 8279
rect 16991 8276 17003 8279
rect 17126 8276 17132 8288
rect 16991 8248 17132 8276
rect 16991 8245 17003 8248
rect 16945 8239 17003 8245
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 18509 8279 18567 8285
rect 18509 8245 18521 8279
rect 18555 8276 18567 8279
rect 20070 8276 20076 8288
rect 18555 8248 20076 8276
rect 18555 8245 18567 8248
rect 18509 8239 18567 8245
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 1104 8186 23276 8208
rect 1104 8134 8379 8186
rect 8431 8134 8443 8186
rect 8495 8134 8507 8186
rect 8559 8134 8571 8186
rect 8623 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 15904 8186
rect 15956 8134 15968 8186
rect 16020 8134 23276 8186
rect 1104 8112 23276 8134
rect 5442 8032 5448 8084
rect 5500 8072 5506 8084
rect 5994 8072 6000 8084
rect 5500 8044 6000 8072
rect 5500 8032 5506 8044
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 6546 8072 6552 8084
rect 6507 8044 6552 8072
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 7006 8072 7012 8084
rect 6967 8044 7012 8072
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7377 8075 7435 8081
rect 7377 8041 7389 8075
rect 7423 8072 7435 8075
rect 7742 8072 7748 8084
rect 7423 8044 7748 8072
rect 7423 8041 7435 8044
rect 7377 8035 7435 8041
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8754 8072 8760 8084
rect 8619 8044 8760 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9030 8072 9036 8084
rect 8991 8044 9036 8072
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9876 8044 12572 8072
rect 8018 7964 8024 8016
rect 8076 8004 8082 8016
rect 8076 7976 8156 8004
rect 8076 7964 8082 7976
rect 2498 7936 2504 7948
rect 2459 7908 2504 7936
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7936 4767 7939
rect 5074 7936 5080 7948
rect 4755 7908 5080 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7936 5871 7939
rect 5902 7936 5908 7948
rect 5859 7908 5908 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6503 7908 6929 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 3160 7732 3188 7831
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4212 7840 4905 7868
rect 4212 7828 4218 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 6932 7868 6960 7899
rect 7006 7896 7012 7948
rect 7064 7936 7070 7948
rect 7558 7936 7564 7948
rect 7064 7908 7564 7936
rect 7064 7896 7070 7908
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 7742 7896 7748 7948
rect 7800 7936 7806 7948
rect 7929 7939 7987 7945
rect 7929 7936 7941 7939
rect 7800 7908 7941 7936
rect 7800 7896 7806 7908
rect 7929 7905 7941 7908
rect 7975 7905 7987 7939
rect 8128 7936 8156 7976
rect 8662 7964 8668 8016
rect 8720 8004 8726 8016
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 8720 7976 8953 8004
rect 8720 7964 8726 7976
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 8941 7967 8999 7973
rect 9876 7936 9904 8044
rect 9944 8007 10002 8013
rect 9944 7973 9956 8007
rect 9990 8004 10002 8007
rect 11146 8004 11152 8016
rect 9990 7976 11152 8004
rect 9990 7973 10002 7976
rect 9944 7967 10002 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 8128 7908 9904 7936
rect 7929 7899 7987 7905
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11589 7939 11647 7945
rect 11589 7936 11601 7939
rect 11296 7908 11601 7936
rect 11296 7896 11302 7908
rect 11589 7905 11601 7908
rect 11635 7905 11647 7939
rect 11589 7899 11647 7905
rect 7193 7871 7251 7877
rect 6932 7840 7052 7868
rect 4893 7831 4951 7837
rect 5997 7803 6055 7809
rect 5997 7769 6009 7803
rect 6043 7800 6055 7803
rect 6638 7800 6644 7812
rect 6043 7772 6644 7800
rect 6043 7769 6055 7772
rect 5997 7763 6055 7769
rect 6638 7760 6644 7772
rect 6696 7760 6702 7812
rect 7024 7800 7052 7840
rect 7193 7837 7205 7871
rect 7239 7868 7251 7871
rect 8018 7868 8024 7880
rect 7239 7840 7880 7868
rect 7979 7840 8024 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 7024 7772 7389 7800
rect 7377 7769 7389 7772
rect 7423 7769 7435 7803
rect 7558 7800 7564 7812
rect 7519 7772 7564 7800
rect 7377 7763 7435 7769
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 7852 7800 7880 7840
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8202 7868 8208 7880
rect 8163 7840 8208 7868
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9140 7800 9168 7831
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 11333 7871 11391 7877
rect 9732 7840 9777 7868
rect 9732 7828 9738 7840
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 12544 7868 12572 8044
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12713 8075 12771 8081
rect 12713 8072 12725 8075
rect 12676 8044 12725 8072
rect 12676 8032 12682 8044
rect 12713 8041 12725 8044
rect 12759 8041 12771 8075
rect 13354 8072 13360 8084
rect 12713 8035 12771 8041
rect 13004 8044 13360 8072
rect 13004 7945 13032 8044
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 14366 8072 14372 8084
rect 14327 8044 14372 8072
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14829 8075 14887 8081
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 14875 8044 16405 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 16393 8041 16405 8044
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17402 8072 17408 8084
rect 16991 8044 17408 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 18322 8072 18328 8084
rect 17788 8044 18328 8072
rect 13262 8013 13268 8016
rect 13256 7967 13268 8013
rect 13320 8004 13326 8016
rect 15470 8004 15476 8016
rect 13320 7976 13356 8004
rect 14660 7976 15476 8004
rect 13262 7964 13268 7967
rect 13320 7964 13326 7976
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7936 12863 7939
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12851 7908 13001 7936
rect 12851 7905 12863 7908
rect 12805 7899 12863 7905
rect 12989 7905 13001 7908
rect 13035 7905 13047 7939
rect 14182 7936 14188 7948
rect 12989 7899 13047 7905
rect 13096 7908 14188 7936
rect 13096 7868 13124 7908
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 14660 7945 14688 7976
rect 15470 7964 15476 7976
rect 15528 7964 15534 8016
rect 16301 8007 16359 8013
rect 16301 7973 16313 8007
rect 16347 8004 16359 8007
rect 16482 8004 16488 8016
rect 16347 7976 16488 8004
rect 16347 7973 16359 7976
rect 16301 7967 16359 7973
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 17313 8007 17371 8013
rect 17313 7973 17325 8007
rect 17359 8004 17371 8007
rect 17788 8004 17816 8044
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 19242 8032 19248 8084
rect 19300 8072 19306 8084
rect 19337 8075 19395 8081
rect 19337 8072 19349 8075
rect 19300 8044 19349 8072
rect 19300 8032 19306 8044
rect 19337 8041 19349 8044
rect 19383 8041 19395 8075
rect 22189 8075 22247 8081
rect 22189 8072 22201 8075
rect 19337 8035 19395 8041
rect 19536 8044 22201 8072
rect 17359 7976 17816 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 18202 8007 18260 8013
rect 18202 8004 18214 8007
rect 17920 7976 18214 8004
rect 17920 7964 17926 7976
rect 18202 7973 18214 7976
rect 18248 7973 18260 8007
rect 19058 8004 19064 8016
rect 18202 7967 18260 7973
rect 18892 7976 19064 8004
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 15381 7939 15439 7945
rect 15381 7905 15393 7939
rect 15427 7936 15439 7939
rect 15654 7936 15660 7948
rect 15427 7908 15660 7936
rect 15427 7905 15439 7908
rect 15381 7899 15439 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 16408 7908 17540 7936
rect 16408 7868 16436 7908
rect 16574 7868 16580 7880
rect 12544 7840 13124 7868
rect 15488 7840 16436 7868
rect 16487 7840 16580 7868
rect 11333 7831 11391 7837
rect 9398 7800 9404 7812
rect 7852 7772 9076 7800
rect 9140 7772 9404 7800
rect 8478 7732 8484 7744
rect 3160 7704 8484 7732
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 9048 7732 9076 7772
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 11054 7800 11060 7812
rect 11015 7772 11060 7800
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 10962 7732 10968 7744
rect 9048 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11348 7732 11376 7831
rect 12805 7735 12863 7741
rect 12805 7732 12817 7735
rect 11348 7704 12817 7732
rect 12805 7701 12817 7704
rect 12851 7701 12863 7735
rect 12805 7695 12863 7701
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 15488 7732 15516 7840
rect 16574 7828 16580 7840
rect 16632 7868 16638 7880
rect 17126 7868 17132 7880
rect 16632 7840 17132 7868
rect 16632 7828 16638 7840
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7800 15991 7803
rect 17420 7800 17448 7831
rect 15979 7772 17448 7800
rect 15979 7769 15991 7772
rect 15933 7763 15991 7769
rect 12952 7704 15516 7732
rect 15565 7735 15623 7741
rect 12952 7692 12958 7704
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 17218 7732 17224 7744
rect 15611 7704 17224 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 17512 7732 17540 7908
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 17880 7868 17908 7964
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7936 18015 7939
rect 18892 7936 18920 7976
rect 19058 7964 19064 7976
rect 19116 7964 19122 8016
rect 19150 7964 19156 8016
rect 19208 8004 19214 8016
rect 19536 8004 19564 8044
rect 22189 8041 22201 8044
rect 22235 8041 22247 8075
rect 22189 8035 22247 8041
rect 21266 8004 21272 8016
rect 19208 7976 19564 8004
rect 21227 7976 21272 8004
rect 19208 7964 19214 7976
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 19981 7939 20039 7945
rect 19981 7936 19993 7939
rect 18003 7908 18920 7936
rect 18984 7908 19993 7936
rect 18003 7905 18015 7908
rect 17957 7899 18015 7905
rect 17635 7840 17908 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17954 7732 17960 7744
rect 17512 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7732 18018 7744
rect 18984 7732 19012 7908
rect 19981 7905 19993 7908
rect 20027 7905 20039 7939
rect 20990 7936 20996 7948
rect 20951 7908 20996 7936
rect 19981 7899 20039 7905
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 21174 7896 21180 7948
rect 21232 7936 21238 7948
rect 22097 7939 22155 7945
rect 22097 7936 22109 7939
rect 21232 7908 22109 7936
rect 21232 7896 21238 7908
rect 22097 7905 22109 7908
rect 22143 7905 22155 7939
rect 22097 7899 22155 7905
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19208 7840 20085 7868
rect 19208 7828 19214 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 22373 7871 22431 7877
rect 22373 7837 22385 7871
rect 22419 7868 22431 7871
rect 22646 7868 22652 7880
rect 22419 7840 22652 7868
rect 22419 7837 22431 7840
rect 22373 7831 22431 7837
rect 19426 7760 19432 7812
rect 19484 7800 19490 7812
rect 20180 7800 20208 7831
rect 22646 7828 22652 7840
rect 22704 7828 22710 7880
rect 19484 7772 20208 7800
rect 19484 7760 19490 7772
rect 18012 7704 19012 7732
rect 19613 7735 19671 7741
rect 18012 7692 18018 7704
rect 19613 7701 19625 7735
rect 19659 7732 19671 7735
rect 19794 7732 19800 7744
rect 19659 7704 19800 7732
rect 19659 7701 19671 7704
rect 19613 7695 19671 7701
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 19886 7692 19892 7744
rect 19944 7732 19950 7744
rect 21729 7735 21787 7741
rect 21729 7732 21741 7735
rect 19944 7704 21741 7732
rect 19944 7692 19950 7704
rect 21729 7701 21741 7704
rect 21775 7732 21787 7735
rect 22186 7732 22192 7744
rect 21775 7704 22192 7732
rect 21775 7701 21787 7704
rect 21729 7695 21787 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 1104 7642 23276 7664
rect 1104 7590 4680 7642
rect 4732 7590 4744 7642
rect 4796 7590 4808 7642
rect 4860 7590 4872 7642
rect 4924 7590 12078 7642
rect 12130 7590 12142 7642
rect 12194 7590 12206 7642
rect 12258 7590 12270 7642
rect 12322 7590 19475 7642
rect 19527 7590 19539 7642
rect 19591 7590 19603 7642
rect 19655 7590 19667 7642
rect 19719 7590 23276 7642
rect 1104 7568 23276 7590
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 5534 7528 5540 7540
rect 4755 7500 5540 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 5721 7531 5779 7537
rect 5721 7497 5733 7531
rect 5767 7528 5779 7531
rect 6178 7528 6184 7540
rect 5767 7500 6184 7528
rect 5767 7497 5779 7500
rect 5721 7491 5779 7497
rect 6178 7488 6184 7500
rect 6236 7488 6242 7540
rect 7469 7531 7527 7537
rect 6748 7500 7135 7528
rect 3697 7463 3755 7469
rect 3697 7429 3709 7463
rect 3743 7460 3755 7463
rect 6086 7460 6092 7472
rect 3743 7432 6092 7460
rect 3743 7429 3755 7432
rect 3697 7423 3755 7429
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 3936 7364 4261 7392
rect 3936 7352 3942 7364
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 5040 7364 5181 7392
rect 5040 7352 5046 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 5399 7364 6377 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 6365 7361 6377 7364
rect 6411 7392 6423 7395
rect 6748 7392 6776 7500
rect 7006 7460 7012 7472
rect 6932 7432 7012 7460
rect 6932 7392 6960 7432
rect 7006 7420 7012 7432
rect 7064 7420 7070 7472
rect 7107 7460 7135 7500
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 7558 7528 7564 7540
rect 7515 7500 7564 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 8018 7488 8024 7540
rect 8076 7528 8082 7540
rect 12437 7531 12495 7537
rect 8076 7500 11100 7528
rect 8076 7488 8082 7500
rect 8478 7460 8484 7472
rect 7107 7432 7604 7460
rect 7576 7404 7604 7432
rect 8128 7432 8484 7460
rect 6411 7364 6776 7392
rect 6840 7364 6960 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 3844 7296 4077 7324
rect 3844 7284 3850 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 4065 7287 4123 7293
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7324 6147 7327
rect 6840 7324 6868 7364
rect 7558 7352 7564 7404
rect 7616 7352 7622 7404
rect 8128 7401 8156 7432
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 11072 7460 11100 7500
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 12483 7500 13216 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 12710 7460 12716 7472
rect 11072 7432 12716 7460
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 9824 7364 10272 7392
rect 9824 7352 9830 7364
rect 7006 7324 7012 7336
rect 7064 7333 7070 7336
rect 6135 7296 6868 7324
rect 6975 7296 7012 7324
rect 6135 7293 6147 7296
rect 6089 7287 6147 7293
rect 7006 7284 7012 7296
rect 7064 7287 7075 7333
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 7300 7296 8493 7324
rect 7064 7284 7070 7287
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 7098 7256 7104 7268
rect 6227 7228 7104 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 4522 7188 4528 7200
rect 4203 7160 4528 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 6270 7188 6276 7200
rect 5123 7160 6276 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 7300 7188 7328 7296
rect 8481 7293 8493 7296
rect 8527 7324 8539 7327
rect 9674 7324 9680 7336
rect 8527 7296 9680 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 9674 7284 9680 7296
rect 9732 7324 9738 7336
rect 10042 7324 10048 7336
rect 9732 7296 10048 7324
rect 9732 7284 9738 7296
rect 10042 7284 10048 7296
rect 10100 7324 10106 7336
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 10100 7296 10149 7324
rect 10100 7284 10106 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10244 7324 10272 7364
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 12526 7392 12532 7404
rect 11204 7364 12532 7392
rect 11204 7352 11210 7364
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13188 7392 13216 7500
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 14829 7531 14887 7537
rect 14829 7528 14841 7531
rect 13320 7500 14841 7528
rect 13320 7488 13326 7500
rect 14829 7497 14841 7500
rect 14875 7497 14887 7531
rect 14829 7491 14887 7497
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15252 7500 15301 7528
rect 15252 7488 15258 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 16942 7528 16948 7540
rect 15289 7491 15347 7497
rect 15396 7500 16948 7528
rect 14458 7420 14464 7472
rect 14516 7460 14522 7472
rect 15396 7460 15424 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17681 7531 17739 7537
rect 17681 7497 17693 7531
rect 17727 7528 17739 7531
rect 19150 7528 19156 7540
rect 17727 7500 19156 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 14516 7432 15424 7460
rect 14516 7420 14522 7432
rect 18414 7420 18420 7472
rect 18472 7420 18478 7472
rect 13188 7364 13584 7392
rect 13081 7355 13139 7361
rect 10244 7296 11192 7324
rect 10137 7287 10195 7293
rect 7377 7259 7435 7265
rect 7377 7225 7389 7259
rect 7423 7256 7435 7259
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7423 7228 7849 7256
rect 7423 7225 7435 7228
rect 7377 7219 7435 7225
rect 7837 7225 7849 7228
rect 7883 7256 7895 7259
rect 8018 7256 8024 7268
rect 7883 7228 8024 7256
rect 7883 7225 7895 7228
rect 7837 7219 7895 7225
rect 8018 7216 8024 7228
rect 8076 7216 8082 7268
rect 8748 7259 8806 7265
rect 8748 7225 8760 7259
rect 8794 7256 8806 7259
rect 10226 7256 10232 7268
rect 8794 7228 10232 7256
rect 8794 7225 8806 7228
rect 8748 7219 8806 7225
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 10404 7259 10462 7265
rect 10404 7225 10416 7259
rect 10450 7256 10462 7259
rect 11054 7256 11060 7268
rect 10450 7228 11060 7256
rect 10450 7225 10462 7228
rect 10404 7219 10462 7225
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11164 7256 11192 7296
rect 11330 7284 11336 7336
rect 11388 7324 11394 7336
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11388 7296 11805 7324
rect 11388 7284 11394 7296
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 11793 7287 11851 7293
rect 12805 7259 12863 7265
rect 11164 7228 12020 7256
rect 6871 7160 7328 7188
rect 7929 7191 7987 7197
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 7929 7157 7941 7191
rect 7975 7188 7987 7191
rect 9122 7188 9128 7200
rect 7975 7160 9128 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 9861 7191 9919 7197
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 11238 7188 11244 7200
rect 9907 7160 11244 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11606 7188 11612 7200
rect 11563 7160 11612 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11992 7197 12020 7228
rect 12805 7225 12817 7259
rect 12851 7256 12863 7259
rect 12894 7256 12900 7268
rect 12851 7228 12900 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7157 12035 7191
rect 13096 7188 13124 7355
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 13412 7296 13461 7324
rect 13412 7284 13418 7296
rect 13449 7293 13461 7296
rect 13495 7293 13507 7327
rect 13556 7324 13584 7364
rect 14918 7352 14924 7404
rect 14976 7392 14982 7404
rect 15841 7395 15899 7401
rect 15841 7392 15853 7395
rect 14976 7364 15853 7392
rect 14976 7352 14982 7364
rect 15841 7361 15853 7364
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 16114 7352 16120 7404
rect 16172 7392 16178 7404
rect 16304 7395 16362 7401
rect 16304 7392 16316 7395
rect 16172 7364 16316 7392
rect 16172 7352 16178 7364
rect 16304 7361 16316 7364
rect 16350 7361 16362 7395
rect 18432 7392 18460 7420
rect 18880 7395 18938 7401
rect 18880 7392 18892 7395
rect 18432 7364 18892 7392
rect 16304 7355 16362 7361
rect 18880 7361 18892 7364
rect 18926 7361 18938 7395
rect 19150 7392 19156 7404
rect 19111 7364 19156 7392
rect 18880 7355 18938 7361
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 14734 7324 14740 7336
rect 13556 7296 14740 7324
rect 13449 7287 13507 7293
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 15102 7324 15108 7336
rect 15063 7296 15108 7324
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 16577 7327 16635 7333
rect 16577 7293 16589 7327
rect 16623 7324 16635 7327
rect 16942 7324 16948 7336
rect 16623 7296 16948 7324
rect 16623 7293 16635 7296
rect 16577 7287 16635 7293
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18288 7296 18429 7324
rect 18288 7284 18294 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 18690 7284 18696 7336
rect 18748 7324 18754 7336
rect 19058 7324 19064 7336
rect 18748 7296 19064 7324
rect 18748 7284 18754 7296
rect 19058 7284 19064 7296
rect 19116 7324 19122 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 19116 7296 20545 7324
rect 19116 7284 19122 7296
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 22189 7327 22247 7333
rect 22189 7293 22201 7327
rect 22235 7324 22247 7327
rect 22738 7324 22744 7336
rect 22235 7296 22744 7324
rect 22235 7293 22247 7296
rect 22189 7287 22247 7293
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 13716 7259 13774 7265
rect 13716 7225 13728 7259
rect 13762 7256 13774 7259
rect 14918 7256 14924 7268
rect 13762 7228 14924 7256
rect 13762 7225 13774 7228
rect 13716 7219 13774 7225
rect 14918 7216 14924 7228
rect 14976 7216 14982 7268
rect 20714 7216 20720 7268
rect 20772 7265 20778 7268
rect 20772 7259 20836 7265
rect 20772 7225 20790 7259
rect 20824 7225 20836 7259
rect 22462 7256 22468 7268
rect 22423 7228 22468 7256
rect 20772 7219 20836 7225
rect 20772 7216 20778 7219
rect 22462 7216 22468 7228
rect 22520 7216 22526 7268
rect 15102 7188 15108 7200
rect 13096 7160 15108 7188
rect 11977 7151 12035 7157
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 16307 7191 16365 7197
rect 16307 7157 16319 7191
rect 16353 7188 16365 7191
rect 18506 7188 18512 7200
rect 16353 7160 18512 7188
rect 16353 7157 16365 7160
rect 16307 7151 16365 7157
rect 18506 7148 18512 7160
rect 18564 7188 18570 7200
rect 18883 7191 18941 7197
rect 18883 7188 18895 7191
rect 18564 7160 18895 7188
rect 18564 7148 18570 7160
rect 18883 7157 18895 7160
rect 18929 7157 18941 7191
rect 18883 7151 18941 7157
rect 20070 7148 20076 7200
rect 20128 7188 20134 7200
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 20128 7160 20269 7188
rect 20128 7148 20134 7160
rect 20257 7157 20269 7160
rect 20303 7188 20315 7191
rect 20438 7188 20444 7200
rect 20303 7160 20444 7188
rect 20303 7157 20315 7160
rect 20257 7151 20315 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20990 7148 20996 7200
rect 21048 7188 21054 7200
rect 21913 7191 21971 7197
rect 21913 7188 21925 7191
rect 21048 7160 21925 7188
rect 21048 7148 21054 7160
rect 21913 7157 21925 7160
rect 21959 7157 21971 7191
rect 21913 7151 21971 7157
rect 1104 7098 23276 7120
rect 1104 7046 8379 7098
rect 8431 7046 8443 7098
rect 8495 7046 8507 7098
rect 8559 7046 8571 7098
rect 8623 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 15904 7098
rect 15956 7046 15968 7098
rect 16020 7046 23276 7098
rect 1104 7024 23276 7046
rect 4522 6984 4528 6996
rect 4483 6956 4528 6984
rect 4522 6944 4528 6956
rect 4580 6944 4586 6996
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 5905 6987 5963 6993
rect 5905 6984 5917 6987
rect 5868 6956 5917 6984
rect 5868 6944 5874 6956
rect 5905 6953 5917 6956
rect 5951 6953 5963 6987
rect 6914 6984 6920 6996
rect 6875 6956 6920 6984
rect 5905 6947 5963 6953
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 9858 6984 9864 6996
rect 7024 6956 9864 6984
rect 4430 6876 4436 6928
rect 4488 6916 4494 6928
rect 4893 6919 4951 6925
rect 4893 6916 4905 6919
rect 4488 6888 4905 6916
rect 4488 6876 4494 6888
rect 4893 6885 4905 6888
rect 4939 6885 4951 6919
rect 4893 6879 4951 6885
rect 5074 6876 5080 6928
rect 5132 6916 5138 6928
rect 7024 6916 7052 6956
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 10870 6984 10876 6996
rect 9968 6956 10876 6984
rect 5132 6888 7052 6916
rect 7929 6919 7987 6925
rect 5132 6876 5138 6888
rect 7929 6885 7941 6919
rect 7975 6916 7987 6919
rect 9582 6916 9588 6928
rect 7975 6888 9588 6916
rect 7975 6885 7987 6888
rect 7929 6879 7987 6885
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6848 5043 6851
rect 6362 6848 6368 6860
rect 5031 6820 6368 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 7374 6848 7380 6860
rect 7055 6820 7380 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8076 6820 8121 6848
rect 8076 6808 8082 6820
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8754 6848 8760 6860
rect 8352 6820 8760 6848
rect 8352 6808 8358 6820
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9674 6848 9680 6860
rect 8987 6820 9680 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 9858 6848 9864 6860
rect 9819 6820 9864 6848
rect 9858 6808 9864 6820
rect 9916 6808 9922 6860
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4304 6752 5089 6780
rect 4304 6740 4310 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5684 6752 6009 6780
rect 5684 6740 5690 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 7193 6783 7251 6789
rect 6227 6752 7144 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 5534 6712 5540 6724
rect 5495 6684 5540 6712
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 6549 6715 6607 6721
rect 6549 6681 6561 6715
rect 6595 6712 6607 6715
rect 6822 6712 6828 6724
rect 6595 6684 6828 6712
rect 6595 6681 6607 6684
rect 6549 6675 6607 6681
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 7116 6712 7144 6752
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 7558 6780 7564 6792
rect 7239 6752 7564 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7558 6740 7564 6752
rect 7616 6780 7622 6792
rect 7742 6780 7748 6792
rect 7616 6752 7748 6780
rect 7616 6740 7622 6752
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8159 6752 8340 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8202 6712 8208 6724
rect 7116 6684 8208 6712
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 7558 6644 7564 6656
rect 7519 6616 7564 6644
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 8312 6644 8340 6752
rect 8496 6752 9045 6780
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 8496 6712 8524 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9398 6780 9404 6792
rect 9171 6752 9404 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9968 6780 9996 6956
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 10962 6944 10968 6996
rect 11020 6984 11026 6996
rect 22738 6984 22744 6996
rect 11020 6956 22744 6984
rect 11020 6944 11026 6956
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 10226 6876 10232 6928
rect 10284 6916 10290 6928
rect 12897 6919 12955 6925
rect 10284 6888 12664 6916
rect 10284 6876 10290 6888
rect 10042 6808 10048 6860
rect 10100 6808 10106 6860
rect 10410 6848 10416 6860
rect 10323 6820 10416 6848
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10680 6851 10738 6857
rect 10680 6817 10692 6851
rect 10726 6848 10738 6851
rect 11606 6848 11612 6860
rect 10726 6820 11612 6848
rect 10726 6817 10738 6820
rect 10680 6811 10738 6817
rect 11606 6808 11612 6820
rect 11664 6808 11670 6860
rect 9600 6752 9996 6780
rect 8444 6684 8524 6712
rect 8573 6715 8631 6721
rect 8444 6672 8450 6684
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 9600 6712 9628 6752
rect 8619 6684 9628 6712
rect 10060 6712 10088 6808
rect 10419 6712 10447 6808
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 12032 6752 12081 6780
rect 12032 6740 12038 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12636 6780 12664 6888
rect 12897 6885 12909 6919
rect 12943 6916 12955 6919
rect 22557 6919 22615 6925
rect 22557 6916 22569 6919
rect 12943 6888 22569 6916
rect 12943 6885 12955 6888
rect 12897 6879 12955 6885
rect 22557 6885 22569 6888
rect 22603 6885 22615 6919
rect 22557 6879 22615 6885
rect 12710 6808 12716 6860
rect 12768 6848 12774 6860
rect 13354 6848 13360 6860
rect 12768 6820 13360 6848
rect 12768 6808 12774 6820
rect 13354 6808 13360 6820
rect 13412 6848 13418 6860
rect 13541 6851 13599 6857
rect 13541 6848 13553 6851
rect 13412 6820 13553 6848
rect 13412 6808 13418 6820
rect 13541 6817 13553 6820
rect 13587 6817 13599 6851
rect 13541 6811 13599 6817
rect 13808 6851 13866 6857
rect 13808 6817 13820 6851
rect 13854 6848 13866 6851
rect 14826 6848 14832 6860
rect 13854 6820 14832 6848
rect 13854 6817 13866 6820
rect 13808 6811 13866 6817
rect 14826 6808 14832 6820
rect 14884 6808 14890 6860
rect 15102 6808 15108 6860
rect 15160 6848 15166 6860
rect 15913 6851 15971 6857
rect 15913 6848 15925 6851
rect 15160 6820 15925 6848
rect 15160 6808 15166 6820
rect 15913 6817 15925 6820
rect 15959 6848 15971 6851
rect 17402 6848 17408 6860
rect 15959 6820 17408 6848
rect 15959 6817 15971 6820
rect 15913 6811 15971 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 18040 6851 18098 6857
rect 18040 6817 18052 6851
rect 18086 6848 18098 6851
rect 18506 6848 18512 6860
rect 18086 6820 18512 6848
rect 18086 6817 18098 6820
rect 18040 6811 18098 6817
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 19794 6848 19800 6860
rect 19755 6820 19800 6848
rect 19794 6808 19800 6820
rect 19852 6808 19858 6860
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20864 6820 20913 6848
rect 20864 6808 20870 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21157 6851 21215 6857
rect 21157 6848 21169 6851
rect 21048 6820 21169 6848
rect 21048 6808 21054 6820
rect 21157 6817 21169 6820
rect 21203 6817 21215 6851
rect 21157 6811 21215 6817
rect 12894 6780 12900 6792
rect 12636 6752 12900 6780
rect 12069 6743 12127 6749
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 13262 6780 13268 6792
rect 13219 6752 13268 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 12618 6712 12624 6724
rect 10060 6684 10447 6712
rect 11624 6684 12624 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 9674 6644 9680 6656
rect 8312 6616 9680 6644
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 11624 6644 11652 6684
rect 12618 6672 12624 6684
rect 12676 6672 12682 6724
rect 11790 6644 11796 6656
rect 10091 6616 11652 6644
rect 11751 6616 11796 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 12526 6644 12532 6656
rect 12487 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 13004 6644 13032 6743
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 15654 6780 15660 6792
rect 15615 6752 15660 6780
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 17276 6752 17325 6780
rect 17276 6740 17282 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 17552 6752 17785 6780
rect 17552 6740 17558 6752
rect 17773 6749 17785 6752
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 19702 6780 19708 6792
rect 18840 6752 19708 6780
rect 18840 6740 18846 6752
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 19886 6780 19892 6792
rect 19847 6752 19892 6780
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 19058 6672 19064 6724
rect 19116 6712 19122 6724
rect 19996 6712 20024 6743
rect 19116 6684 20024 6712
rect 19116 6672 19122 6684
rect 13814 6644 13820 6656
rect 13004 6616 13820 6644
rect 13814 6604 13820 6616
rect 13872 6604 13878 6656
rect 14918 6644 14924 6656
rect 14879 6616 14924 6644
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 17000 6616 17049 6644
rect 17000 6604 17006 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 19153 6647 19211 6653
rect 19153 6613 19165 6647
rect 19199 6644 19211 6647
rect 19334 6644 19340 6656
rect 19199 6616 19340 6644
rect 19199 6613 19211 6616
rect 19153 6607 19211 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 20898 6644 20904 6656
rect 19475 6616 20904 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 21082 6604 21088 6656
rect 21140 6644 21146 6656
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 21140 6616 22293 6644
rect 21140 6604 21146 6616
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 1104 6554 23276 6576
rect 1104 6502 4680 6554
rect 4732 6502 4744 6554
rect 4796 6502 4808 6554
rect 4860 6502 4872 6554
rect 4924 6502 12078 6554
rect 12130 6502 12142 6554
rect 12194 6502 12206 6554
rect 12258 6502 12270 6554
rect 12322 6502 19475 6554
rect 19527 6502 19539 6554
rect 19591 6502 19603 6554
rect 19655 6502 19667 6554
rect 19719 6502 23276 6554
rect 1104 6480 23276 6502
rect 5626 6440 5632 6452
rect 5587 6412 5632 6440
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 7650 6440 7656 6452
rect 7611 6412 7656 6440
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 8202 6440 8208 6452
rect 7800 6412 8208 6440
rect 7800 6400 7806 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9306 6440 9312 6452
rect 8812 6412 9312 6440
rect 8812 6400 8818 6412
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 11330 6440 11336 6452
rect 9723 6412 11336 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 23014 6440 23020 6452
rect 12584 6412 23020 6440
rect 12584 6400 12590 6412
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 10134 6372 10140 6384
rect 8036 6344 10140 6372
rect 6086 6304 6092 6316
rect 6047 6276 6092 6304
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 7466 6304 7472 6316
rect 6319 6276 7472 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 8036 6245 8064 6344
rect 10134 6332 10140 6344
rect 10192 6332 10198 6384
rect 10594 6372 10600 6384
rect 10244 6344 10600 6372
rect 8202 6304 8208 6316
rect 8163 6276 8208 6304
rect 8202 6264 8208 6276
rect 8260 6264 8266 6316
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9398 6304 9404 6316
rect 9355 6276 9404 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9398 6264 9404 6276
rect 9456 6264 9462 6316
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5500 6208 6009 6236
rect 5500 6196 5506 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6236 8171 6239
rect 8294 6236 8300 6248
rect 8159 6208 8300 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 9030 6236 9036 6248
rect 8991 6208 9036 6236
rect 9030 6196 9036 6208
rect 9088 6196 9094 6248
rect 10244 6236 10272 6344
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 17402 6372 17408 6384
rect 17363 6344 17408 6372
rect 17402 6332 17408 6344
rect 17460 6332 17466 6384
rect 18414 6372 18420 6384
rect 18375 6344 18420 6372
rect 18414 6332 18420 6344
rect 18472 6332 18478 6384
rect 18782 6332 18788 6384
rect 18840 6332 18846 6384
rect 20625 6375 20683 6381
rect 20625 6341 20637 6375
rect 20671 6372 20683 6375
rect 20714 6372 20720 6384
rect 20671 6344 20720 6372
rect 20671 6341 20683 6344
rect 20625 6335 20683 6341
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 9876 6208 10272 6236
rect 10336 6236 10364 6267
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10468 6276 10701 6304
rect 10468 6264 10474 6276
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12710 6304 12716 6316
rect 12308 6276 12716 6304
rect 12308 6264 12314 6276
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 15712 6276 16037 6304
rect 15712 6264 15718 6276
rect 16025 6273 16037 6276
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 18800 6304 18828 6332
rect 17092 6276 18828 6304
rect 17092 6264 17098 6276
rect 20070 6264 20076 6316
rect 20128 6304 20134 6316
rect 20128 6276 21476 6304
rect 20128 6264 20134 6276
rect 10778 6236 10784 6248
rect 10336 6208 10784 6236
rect 9122 6168 9128 6180
rect 9083 6140 9128 6168
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 9876 6100 9904 6208
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 10956 6239 11014 6245
rect 10956 6205 10968 6239
rect 11002 6236 11014 6239
rect 11790 6236 11796 6248
rect 11002 6208 11796 6236
rect 11002 6205 11014 6208
rect 10956 6199 11014 6205
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 14366 6236 14372 6248
rect 13320 6208 14228 6236
rect 14327 6208 14372 6236
rect 13320 6196 13326 6208
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 12980 6171 13038 6177
rect 10652 6140 12204 6168
rect 10652 6128 10658 6140
rect 10042 6100 10048 6112
rect 8711 6072 9904 6100
rect 10003 6072 10048 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 11146 6100 11152 6112
rect 10183 6072 11152 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 12032 6072 12081 6100
rect 12032 6060 12038 6072
rect 12069 6069 12081 6072
rect 12115 6069 12127 6103
rect 12176 6100 12204 6140
rect 12980 6137 12992 6171
rect 13026 6168 13038 6171
rect 13630 6168 13636 6180
rect 13026 6140 13636 6168
rect 13026 6137 13038 6140
rect 12980 6131 13038 6137
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 14200 6168 14228 6208
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 16281 6239 16339 6245
rect 16281 6236 16293 6239
rect 14568 6208 16293 6236
rect 14568 6168 14596 6208
rect 16281 6205 16293 6208
rect 16327 6236 16339 6239
rect 17865 6239 17923 6245
rect 16327 6208 17816 6236
rect 16327 6205 16339 6208
rect 16281 6199 16339 6205
rect 14642 6177 14648 6180
rect 14200 6140 14596 6168
rect 14636 6131 14648 6177
rect 14700 6168 14706 6180
rect 14700 6140 14736 6168
rect 14642 6128 14648 6131
rect 14700 6128 14706 6140
rect 13170 6100 13176 6112
rect 12176 6072 13176 6100
rect 12069 6063 12127 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14274 6100 14280 6112
rect 14139 6072 14280 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 15528 6072 15761 6100
rect 15528 6060 15534 6072
rect 15749 6069 15761 6072
rect 15795 6069 15807 6103
rect 15749 6063 15807 6069
rect 17126 6060 17132 6112
rect 17184 6100 17190 6112
rect 17494 6100 17500 6112
rect 17184 6072 17500 6100
rect 17184 6060 17190 6072
rect 17494 6060 17500 6072
rect 17552 6100 17558 6112
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 17552 6072 17693 6100
rect 17552 6060 17558 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17788 6100 17816 6208
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 18138 6236 18144 6248
rect 17911 6208 18144 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 18248 6168 18276 6199
rect 18690 6196 18696 6248
rect 18748 6236 18754 6248
rect 18785 6239 18843 6245
rect 18785 6236 18797 6239
rect 18748 6208 18797 6236
rect 18748 6196 18754 6208
rect 18785 6205 18797 6208
rect 18831 6205 18843 6239
rect 18785 6199 18843 6205
rect 19052 6239 19110 6245
rect 19052 6205 19064 6239
rect 19098 6236 19110 6239
rect 19334 6236 19340 6248
rect 19098 6208 19340 6236
rect 19098 6205 19110 6208
rect 19052 6199 19110 6205
rect 19334 6196 19340 6208
rect 19392 6196 19398 6248
rect 21082 6236 21088 6248
rect 19904 6208 21088 6236
rect 19794 6168 19800 6180
rect 18248 6140 19800 6168
rect 19794 6128 19800 6140
rect 19852 6128 19858 6180
rect 19904 6100 19932 6208
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 21266 6196 21272 6248
rect 21324 6236 21330 6248
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 21324 6208 21373 6236
rect 21324 6196 21330 6208
rect 21361 6205 21373 6208
rect 21407 6205 21419 6239
rect 21448 6236 21476 6276
rect 22370 6236 22376 6248
rect 21448 6208 22376 6236
rect 21361 6199 21419 6205
rect 22370 6196 22376 6208
rect 22428 6196 22434 6248
rect 20625 6171 20683 6177
rect 20625 6168 20637 6171
rect 20180 6140 20637 6168
rect 17788 6072 19932 6100
rect 17681 6063 17739 6069
rect 19978 6060 19984 6112
rect 20036 6100 20042 6112
rect 20180 6109 20208 6140
rect 20625 6137 20637 6140
rect 20671 6137 20683 6171
rect 20625 6131 20683 6137
rect 20717 6171 20775 6177
rect 20717 6137 20729 6171
rect 20763 6168 20775 6171
rect 20806 6168 20812 6180
rect 20763 6140 20812 6168
rect 20763 6137 20775 6140
rect 20717 6131 20775 6137
rect 20806 6128 20812 6140
rect 20864 6128 20870 6180
rect 20901 6171 20959 6177
rect 20901 6137 20913 6171
rect 20947 6168 20959 6171
rect 21606 6171 21664 6177
rect 21606 6168 21618 6171
rect 20947 6140 21618 6168
rect 20947 6137 20959 6140
rect 20901 6131 20959 6137
rect 21606 6137 21618 6140
rect 21652 6168 21664 6171
rect 22554 6168 22560 6180
rect 21652 6140 22560 6168
rect 21652 6137 21664 6140
rect 21606 6131 21664 6137
rect 22554 6128 22560 6140
rect 22612 6128 22618 6180
rect 20165 6103 20223 6109
rect 20165 6100 20177 6103
rect 20036 6072 20177 6100
rect 20036 6060 20042 6072
rect 20165 6069 20177 6072
rect 20211 6069 20223 6103
rect 21082 6100 21088 6112
rect 21043 6072 21088 6100
rect 20165 6063 20223 6069
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 22738 6100 22744 6112
rect 22699 6072 22744 6100
rect 22738 6060 22744 6072
rect 22796 6060 22802 6112
rect 1104 6010 23276 6032
rect 1104 5958 8379 6010
rect 8431 5958 8443 6010
rect 8495 5958 8507 6010
rect 8559 5958 8571 6010
rect 8623 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 15904 6010
rect 15956 5958 15968 6010
rect 16020 5958 23276 6010
rect 1104 5936 23276 5958
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 5905 5899 5963 5905
rect 5905 5896 5917 5899
rect 5776 5868 5917 5896
rect 5776 5856 5782 5868
rect 5905 5865 5917 5868
rect 5951 5865 5963 5899
rect 5905 5859 5963 5865
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 6144 5868 6285 5896
rect 6144 5856 6150 5868
rect 6273 5865 6285 5868
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 6365 5899 6423 5905
rect 6365 5865 6377 5899
rect 6411 5896 6423 5899
rect 6730 5896 6736 5908
rect 6411 5868 6736 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7984 5868 8033 5896
rect 7984 5856 7990 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 8168 5868 8585 5896
rect 8168 5856 8174 5868
rect 8573 5865 8585 5868
rect 8619 5865 8631 5899
rect 8573 5859 8631 5865
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9950 5896 9956 5908
rect 9079 5868 9956 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 11238 5896 11244 5908
rect 10100 5868 11244 5896
rect 10100 5856 10106 5868
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 12986 5896 12992 5908
rect 11388 5868 12992 5896
rect 11388 5856 11394 5868
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13630 5896 13636 5908
rect 13591 5868 13636 5896
rect 13630 5856 13636 5868
rect 13688 5896 13694 5908
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 13688 5868 14381 5896
rect 13688 5856 13694 5868
rect 14369 5865 14381 5868
rect 14415 5865 14427 5899
rect 14369 5859 14427 5865
rect 14458 5856 14464 5908
rect 14516 5896 14522 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 14516 5868 14933 5896
rect 14516 5856 14522 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 14921 5859 14979 5865
rect 16025 5899 16083 5905
rect 16025 5865 16037 5899
rect 16071 5896 16083 5899
rect 18046 5896 18052 5908
rect 16071 5868 18052 5896
rect 16071 5865 16083 5868
rect 16025 5859 16083 5865
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18506 5896 18512 5908
rect 18467 5868 18512 5896
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19245 5899 19303 5905
rect 19245 5865 19257 5899
rect 19291 5896 19303 5899
rect 21085 5899 21143 5905
rect 21085 5896 21097 5899
rect 19291 5868 21097 5896
rect 19291 5865 19303 5868
rect 19245 5859 19303 5865
rect 21085 5865 21097 5868
rect 21131 5865 21143 5899
rect 21085 5859 21143 5865
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 21821 5899 21879 5905
rect 21821 5896 21833 5899
rect 21692 5868 21833 5896
rect 21692 5856 21698 5868
rect 21821 5865 21833 5868
rect 21867 5865 21879 5899
rect 21821 5859 21879 5865
rect 8941 5831 8999 5837
rect 8941 5797 8953 5831
rect 8987 5828 8999 5831
rect 9766 5828 9772 5840
rect 8987 5800 9772 5828
rect 8987 5797 8999 5800
rect 8941 5791 8999 5797
rect 9766 5788 9772 5800
rect 9824 5788 9830 5840
rect 9858 5788 9864 5840
rect 9916 5828 9922 5840
rect 9916 5800 21128 5828
rect 9916 5788 9922 5800
rect 21100 5772 21128 5800
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7929 5763 7987 5769
rect 7929 5760 7941 5763
rect 7340 5732 7941 5760
rect 7340 5720 7346 5732
rect 7929 5729 7941 5732
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10226 5760 10232 5772
rect 10091 5732 10232 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 10597 5763 10655 5769
rect 10597 5760 10609 5763
rect 10468 5732 10609 5760
rect 10468 5720 10474 5732
rect 10597 5729 10609 5732
rect 10643 5729 10655 5763
rect 10597 5723 10655 5729
rect 10864 5763 10922 5769
rect 10864 5729 10876 5763
rect 10910 5760 10922 5763
rect 11974 5760 11980 5772
rect 10910 5732 11980 5760
rect 10910 5729 10922 5732
rect 10864 5723 10922 5729
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12509 5763 12567 5769
rect 12509 5760 12521 5763
rect 12084 5732 12521 5760
rect 6454 5692 6460 5704
rect 6415 5664 6460 5692
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 8202 5692 8208 5704
rect 8115 5664 8208 5692
rect 8202 5652 8208 5664
rect 8260 5692 8266 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8260 5664 9229 5692
rect 8260 5652 8266 5664
rect 9217 5661 9229 5664
rect 9263 5692 9275 5695
rect 9306 5692 9312 5704
rect 9263 5664 9312 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 7561 5627 7619 5633
rect 7561 5593 7573 5627
rect 7607 5624 7619 5627
rect 8754 5624 8760 5636
rect 7607 5596 8760 5624
rect 7607 5593 7619 5596
rect 7561 5587 7619 5593
rect 8754 5584 8760 5596
rect 8812 5584 8818 5636
rect 11977 5627 12035 5633
rect 11977 5593 11989 5627
rect 12023 5624 12035 5627
rect 12084 5624 12112 5732
rect 12509 5729 12521 5732
rect 12555 5760 12567 5763
rect 12986 5760 12992 5772
rect 12555 5732 12992 5760
rect 12555 5729 12567 5732
rect 12509 5723 12567 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 14274 5760 14280 5772
rect 14235 5732 14280 5760
rect 14274 5720 14280 5732
rect 14332 5720 14338 5772
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 15105 5763 15163 5769
rect 15105 5760 15117 5763
rect 14608 5732 15117 5760
rect 14608 5720 14614 5732
rect 15105 5729 15117 5732
rect 15151 5729 15163 5763
rect 15105 5723 15163 5729
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5760 15623 5763
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 15611 5732 16037 5760
rect 15611 5729 15623 5732
rect 15565 5723 15623 5729
rect 16025 5729 16037 5732
rect 16071 5729 16083 5763
rect 16482 5760 16488 5772
rect 16443 5732 16488 5760
rect 16025 5723 16083 5729
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5760 16635 5763
rect 17034 5760 17040 5772
rect 16623 5732 17040 5760
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 17034 5720 17040 5732
rect 17092 5720 17098 5772
rect 17396 5763 17454 5769
rect 17396 5729 17408 5763
rect 17442 5760 17454 5763
rect 19150 5760 19156 5772
rect 17442 5732 19012 5760
rect 19111 5732 19156 5760
rect 17442 5729 17454 5732
rect 17396 5723 17454 5729
rect 12250 5692 12256 5704
rect 12211 5664 12256 5692
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 14458 5692 14464 5704
rect 14419 5664 14464 5692
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 16666 5692 16672 5704
rect 15672 5664 16672 5692
rect 15672 5624 15700 5664
rect 16666 5652 16672 5664
rect 16724 5652 16730 5704
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5692 16819 5695
rect 16942 5692 16948 5704
rect 16807 5664 16948 5692
rect 16807 5661 16819 5664
rect 16761 5655 16819 5661
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 17126 5692 17132 5704
rect 17087 5664 17132 5692
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 18984 5692 19012 5732
rect 19150 5720 19156 5732
rect 19208 5720 19214 5772
rect 20070 5720 20076 5772
rect 20128 5760 20134 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 20128 5732 20177 5760
rect 20128 5720 20134 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 20257 5763 20315 5769
rect 20257 5729 20269 5763
rect 20303 5760 20315 5763
rect 20898 5760 20904 5772
rect 20303 5732 20760 5760
rect 20859 5732 20904 5760
rect 20303 5729 20315 5732
rect 20257 5723 20315 5729
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 18984 5664 19441 5692
rect 19429 5661 19441 5664
rect 19475 5692 19487 5695
rect 19610 5692 19616 5704
rect 19475 5664 19616 5692
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5661 20499 5695
rect 20441 5655 20499 5661
rect 12023 5596 12112 5624
rect 13740 5596 15700 5624
rect 15749 5627 15807 5633
rect 12023 5593 12035 5596
rect 11977 5587 12035 5593
rect 10229 5559 10287 5565
rect 10229 5525 10241 5559
rect 10275 5556 10287 5559
rect 13740 5556 13768 5596
rect 15749 5593 15761 5627
rect 15795 5624 15807 5627
rect 15795 5596 16988 5624
rect 15795 5593 15807 5596
rect 15749 5587 15807 5593
rect 10275 5528 13768 5556
rect 10275 5525 10287 5528
rect 10229 5519 10287 5525
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 13909 5559 13967 5565
rect 13909 5556 13921 5559
rect 13872 5528 13921 5556
rect 13872 5516 13878 5528
rect 13909 5525 13921 5528
rect 13955 5525 13967 5559
rect 13909 5519 13967 5525
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 16117 5559 16175 5565
rect 16117 5556 16129 5559
rect 15620 5528 16129 5556
rect 15620 5516 15626 5528
rect 16117 5525 16129 5528
rect 16163 5556 16175 5559
rect 16758 5556 16764 5568
rect 16163 5528 16764 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 16960 5556 16988 5596
rect 18414 5584 18420 5636
rect 18472 5624 18478 5636
rect 19242 5624 19248 5636
rect 18472 5596 19248 5624
rect 18472 5584 18478 5596
rect 19242 5584 19248 5596
rect 19300 5584 19306 5636
rect 19794 5624 19800 5636
rect 19755 5596 19800 5624
rect 19794 5584 19800 5596
rect 19852 5584 19858 5636
rect 18138 5556 18144 5568
rect 16960 5528 18144 5556
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 18782 5556 18788 5568
rect 18743 5528 18788 5556
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 18966 5516 18972 5568
rect 19024 5556 19030 5568
rect 20456 5556 20484 5655
rect 20732 5624 20760 5732
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21082 5720 21088 5772
rect 21140 5720 21146 5772
rect 21910 5760 21916 5772
rect 21871 5732 21916 5760
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 22281 5763 22339 5769
rect 22281 5729 22293 5763
rect 22327 5760 22339 5763
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 22327 5732 22477 5760
rect 22327 5729 22339 5732
rect 22281 5723 22339 5729
rect 22465 5729 22477 5732
rect 22511 5729 22523 5763
rect 22465 5723 22523 5729
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 21542 5692 21548 5704
rect 20864 5664 21548 5692
rect 20864 5652 20870 5664
rect 21542 5652 21548 5664
rect 21600 5692 21606 5704
rect 22005 5695 22063 5701
rect 22005 5692 22017 5695
rect 21600 5664 22017 5692
rect 21600 5652 21606 5664
rect 22005 5661 22017 5664
rect 22051 5661 22063 5695
rect 22005 5655 22063 5661
rect 22649 5627 22707 5633
rect 22649 5624 22661 5627
rect 20732 5596 22661 5624
rect 22649 5593 22661 5596
rect 22695 5593 22707 5627
rect 22649 5587 22707 5593
rect 19024 5528 20484 5556
rect 19024 5516 19030 5528
rect 20714 5516 20720 5568
rect 20772 5556 20778 5568
rect 21453 5559 21511 5565
rect 21453 5556 21465 5559
rect 20772 5528 21465 5556
rect 20772 5516 20778 5528
rect 21453 5525 21465 5528
rect 21499 5525 21511 5559
rect 21453 5519 21511 5525
rect 21542 5516 21548 5568
rect 21600 5556 21606 5568
rect 22281 5559 22339 5565
rect 22281 5556 22293 5559
rect 21600 5528 22293 5556
rect 21600 5516 21606 5528
rect 22281 5525 22293 5528
rect 22327 5525 22339 5559
rect 22281 5519 22339 5525
rect 1104 5466 23276 5488
rect 1104 5414 4680 5466
rect 4732 5414 4744 5466
rect 4796 5414 4808 5466
rect 4860 5414 4872 5466
rect 4924 5414 12078 5466
rect 12130 5414 12142 5466
rect 12194 5414 12206 5466
rect 12258 5414 12270 5466
rect 12322 5414 19475 5466
rect 19527 5414 19539 5466
rect 19591 5414 19603 5466
rect 19655 5414 19667 5466
rect 19719 5414 23276 5466
rect 1104 5392 23276 5414
rect 7466 5352 7472 5364
rect 7427 5324 7472 5352
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 10778 5312 10784 5364
rect 10836 5312 10842 5364
rect 11146 5352 11152 5364
rect 11107 5324 11152 5352
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 12437 5355 12495 5361
rect 12437 5352 12449 5355
rect 11296 5324 12449 5352
rect 11296 5312 11302 5324
rect 12437 5321 12449 5324
rect 12483 5321 12495 5355
rect 12437 5315 12495 5321
rect 13357 5355 13415 5361
rect 13357 5321 13369 5355
rect 13403 5352 13415 5355
rect 14366 5352 14372 5364
rect 13403 5324 14372 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 14826 5352 14832 5364
rect 14787 5324 14832 5352
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 17310 5352 17316 5364
rect 16816 5324 17316 5352
rect 16816 5312 16822 5324
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 19245 5355 19303 5361
rect 19245 5352 19257 5355
rect 19208 5324 19257 5352
rect 19208 5312 19214 5324
rect 19245 5321 19257 5324
rect 19291 5321 19303 5355
rect 19245 5315 19303 5321
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 21542 5352 21548 5364
rect 19659 5324 21548 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 21542 5312 21548 5324
rect 21600 5312 21606 5364
rect 22554 5352 22560 5364
rect 22515 5324 22560 5352
rect 22554 5312 22560 5324
rect 22612 5312 22618 5364
rect 8846 5244 8852 5296
rect 8904 5244 8910 5296
rect 10796 5284 10824 5312
rect 13446 5284 13452 5296
rect 10796 5256 13452 5284
rect 13446 5244 13452 5256
rect 13504 5244 13510 5296
rect 14384 5284 14412 5312
rect 14384 5256 15240 5284
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 7892 5188 8033 5216
rect 7892 5176 7898 5188
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8864 5216 8892 5244
rect 9033 5219 9091 5225
rect 9033 5216 9045 5219
rect 8864 5188 9045 5216
rect 8021 5179 8079 5185
rect 9033 5185 9045 5188
rect 9079 5185 9091 5219
rect 10594 5216 10600 5228
rect 10555 5188 10600 5216
rect 9033 5179 9091 5185
rect 10594 5176 10600 5188
rect 10652 5176 10658 5228
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10744 5188 10789 5216
rect 10744 5176 10750 5188
rect 11330 5176 11336 5228
rect 11388 5176 11394 5228
rect 11606 5216 11612 5228
rect 11567 5188 11612 5216
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 11882 5216 11888 5228
rect 11747 5188 11888 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 11974 5176 11980 5228
rect 12032 5216 12038 5228
rect 15212 5225 15240 5256
rect 17954 5244 17960 5296
rect 18012 5284 18018 5296
rect 18049 5287 18107 5293
rect 18049 5284 18061 5287
rect 18012 5256 18061 5284
rect 18012 5244 18018 5256
rect 18049 5253 18061 5256
rect 18095 5253 18107 5287
rect 18049 5247 18107 5253
rect 18506 5244 18512 5296
rect 18564 5284 18570 5296
rect 18564 5256 18644 5284
rect 18564 5244 18570 5256
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12032 5188 12909 5216
rect 12032 5176 12038 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 15197 5219 15255 5225
rect 13127 5188 13216 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 7248 5120 8861 5148
rect 7248 5108 7254 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5148 10563 5151
rect 11348 5148 11376 5176
rect 10551 5120 11376 5148
rect 11517 5151 11575 5157
rect 10551 5117 10563 5120
rect 10505 5111 10563 5117
rect 11517 5117 11529 5151
rect 11563 5148 11575 5151
rect 11790 5148 11796 5160
rect 11563 5120 11796 5148
rect 11563 5117 11575 5120
rect 11517 5111 11575 5117
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 11900 5148 11928 5176
rect 12805 5151 12863 5157
rect 11900 5120 12664 5148
rect 7837 5083 7895 5089
rect 7837 5049 7849 5083
rect 7883 5080 7895 5083
rect 7883 5052 8616 5080
rect 7883 5049 7895 5052
rect 7837 5043 7895 5049
rect 7929 5015 7987 5021
rect 7929 4981 7941 5015
rect 7975 5012 7987 5015
rect 8481 5015 8539 5021
rect 8481 5012 8493 5015
rect 7975 4984 8493 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8481 4981 8493 4984
rect 8527 4981 8539 5015
rect 8588 5012 8616 5052
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 8941 5083 8999 5089
rect 8941 5080 8953 5083
rect 8720 5052 8953 5080
rect 8720 5040 8726 5052
rect 8941 5049 8953 5052
rect 8987 5049 8999 5083
rect 8941 5043 8999 5049
rect 11330 5040 11336 5092
rect 11388 5080 11394 5092
rect 12636 5080 12664 5120
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 12986 5148 12992 5160
rect 12851 5120 12992 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13188 5080 13216 5188
rect 15197 5185 15209 5219
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 17402 5216 17408 5228
rect 16816 5188 17408 5216
rect 16816 5176 16822 5188
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 18616 5225 18644 5256
rect 19058 5244 19064 5296
rect 19116 5284 19122 5296
rect 19116 5256 20208 5284
rect 19116 5244 19122 5256
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 20180 5225 20208 5256
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 18748 5188 20085 5216
rect 18748 5176 18754 5188
rect 20073 5185 20085 5188
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 13403 5120 13461 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 13716 5151 13774 5157
rect 13716 5117 13728 5151
rect 13762 5148 13774 5151
rect 14274 5148 14280 5160
rect 13762 5120 14280 5148
rect 13762 5117 13774 5120
rect 13716 5111 13774 5117
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 15580 5120 17325 5148
rect 15580 5092 15608 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5148 18567 5151
rect 18782 5148 18788 5160
rect 18555 5120 18788 5148
rect 18555 5117 18567 5120
rect 18509 5111 18567 5117
rect 18782 5108 18788 5120
rect 18840 5108 18846 5160
rect 19061 5151 19119 5157
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 19334 5148 19340 5160
rect 19107 5120 19340 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 19334 5108 19340 5120
rect 19392 5148 19398 5160
rect 19978 5148 19984 5160
rect 19392 5120 19984 5148
rect 19392 5108 19398 5120
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 20625 5151 20683 5157
rect 20625 5117 20637 5151
rect 20671 5117 20683 5151
rect 20625 5111 20683 5117
rect 14458 5080 14464 5092
rect 11388 5052 12572 5080
rect 12636 5052 14464 5080
rect 11388 5040 11394 5052
rect 9490 5012 9496 5024
rect 8588 4984 9496 5012
rect 8481 4975 8539 4981
rect 9490 4972 9496 4984
rect 9548 4972 9554 5024
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 12250 5012 12256 5024
rect 10183 4984 12256 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 12544 5012 12572 5052
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 15470 5089 15476 5092
rect 15442 5083 15476 5089
rect 15442 5080 15454 5083
rect 14568 5052 15454 5080
rect 14568 5012 14596 5052
rect 15442 5049 15454 5052
rect 15442 5043 15476 5049
rect 15470 5040 15476 5043
rect 15528 5040 15534 5092
rect 15562 5040 15568 5092
rect 15620 5040 15626 5092
rect 20640 5080 20668 5111
rect 21082 5108 21088 5160
rect 21140 5148 21146 5160
rect 21177 5151 21235 5157
rect 21177 5148 21189 5151
rect 21140 5120 21189 5148
rect 21140 5108 21146 5120
rect 21177 5117 21189 5120
rect 21223 5148 21235 5151
rect 21266 5148 21272 5160
rect 21223 5120 21272 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 21266 5108 21272 5120
rect 21324 5108 21330 5160
rect 16868 5052 20668 5080
rect 21444 5083 21502 5089
rect 12544 4984 14596 5012
rect 15010 4972 15016 5024
rect 15068 5012 15074 5024
rect 16868 5021 16896 5052
rect 21444 5049 21456 5083
rect 21490 5080 21502 5083
rect 22094 5080 22100 5092
rect 21490 5052 22100 5080
rect 21490 5049 21502 5052
rect 21444 5043 21502 5049
rect 22094 5040 22100 5052
rect 22152 5040 22158 5092
rect 16577 5015 16635 5021
rect 16577 5012 16589 5015
rect 15068 4984 16589 5012
rect 15068 4972 15074 4984
rect 16577 4981 16589 4984
rect 16623 4981 16635 5015
rect 16577 4975 16635 4981
rect 16853 5015 16911 5021
rect 16853 4981 16865 5015
rect 16899 4981 16911 5015
rect 16853 4975 16911 4981
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17221 5015 17279 5021
rect 17221 5012 17233 5015
rect 17184 4984 17233 5012
rect 17184 4972 17190 4984
rect 17221 4981 17233 4984
rect 17267 4981 17279 5015
rect 17221 4975 17279 4981
rect 18417 5015 18475 5021
rect 18417 4981 18429 5015
rect 18463 5012 18475 5015
rect 19058 5012 19064 5024
rect 18463 4984 19064 5012
rect 18463 4981 18475 4984
rect 18417 4975 18475 4981
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20806 5012 20812 5024
rect 20767 4984 20812 5012
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 1104 4922 23276 4944
rect 1104 4870 8379 4922
rect 8431 4870 8443 4922
rect 8495 4870 8507 4922
rect 8559 4870 8571 4922
rect 8623 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 15904 4922
rect 15956 4870 15968 4922
rect 16020 4870 23276 4922
rect 1104 4848 23276 4870
rect 9858 4808 9864 4820
rect 9819 4780 9864 4808
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10318 4808 10324 4820
rect 10279 4780 10324 4808
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 11330 4808 11336 4820
rect 11291 4780 11336 4808
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 12526 4808 12532 4820
rect 12299 4780 12532 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12860 4780 12909 4808
rect 12860 4768 12866 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 12897 4771 12955 4777
rect 13265 4811 13323 4817
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 13909 4811 13967 4817
rect 13909 4808 13921 4811
rect 13311 4780 13921 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13909 4777 13921 4780
rect 13955 4777 13967 4811
rect 13909 4771 13967 4777
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 14826 4808 14832 4820
rect 14415 4780 14832 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 16206 4808 16212 4820
rect 15335 4780 16212 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 16942 4808 16948 4820
rect 16316 4780 16948 4808
rect 11241 4743 11299 4749
rect 11241 4709 11253 4743
rect 11287 4740 11299 4743
rect 13357 4743 13415 4749
rect 11287 4712 13308 4740
rect 11287 4709 11299 4712
rect 11241 4703 11299 4709
rect 10226 4672 10232 4684
rect 10187 4644 10232 4672
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 12342 4672 12348 4684
rect 11756 4644 12020 4672
rect 12303 4644 12348 4672
rect 11756 4632 11762 4644
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4604 11575 4607
rect 11882 4604 11888 4616
rect 11563 4576 11888 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 11992 4604 12020 4644
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 13280 4672 13308 4712
rect 13357 4709 13369 4743
rect 13403 4740 13415 4743
rect 13814 4740 13820 4752
rect 13403 4712 13820 4740
rect 13403 4709 13415 4712
rect 13357 4703 13415 4709
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 14277 4743 14335 4749
rect 14277 4709 14289 4743
rect 14323 4740 14335 4743
rect 14918 4740 14924 4752
rect 14323 4712 14924 4740
rect 14323 4709 14335 4712
rect 14277 4703 14335 4709
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 16316 4740 16344 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 19153 4811 19211 4817
rect 19153 4777 19165 4811
rect 19199 4808 19211 4811
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19199 4780 19809 4808
rect 19199 4777 19211 4780
rect 19153 4771 19211 4777
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 20165 4811 20223 4817
rect 20165 4777 20177 4811
rect 20211 4808 20223 4811
rect 22094 4808 22100 4820
rect 20211 4780 22100 4808
rect 20211 4777 20223 4780
rect 20165 4771 20223 4777
rect 22094 4768 22100 4780
rect 22152 4808 22158 4820
rect 22465 4811 22523 4817
rect 22465 4808 22477 4811
rect 22152 4780 22477 4808
rect 22152 4768 22158 4780
rect 22465 4777 22477 4780
rect 22511 4777 22523 4811
rect 22465 4771 22523 4777
rect 15212 4712 16344 4740
rect 13280 4644 14964 4672
rect 14936 4616 14964 4644
rect 15212 4616 15240 4712
rect 16666 4700 16672 4752
rect 16724 4700 16730 4752
rect 18233 4743 18291 4749
rect 18233 4709 18245 4743
rect 18279 4740 18291 4743
rect 20806 4740 20812 4752
rect 18279 4712 20812 4740
rect 18279 4709 18291 4712
rect 18233 4703 18291 4709
rect 20806 4700 20812 4712
rect 20864 4700 20870 4752
rect 15654 4632 15660 4684
rect 15712 4672 15718 4684
rect 15749 4675 15807 4681
rect 15749 4672 15761 4675
rect 15712 4644 15761 4672
rect 15712 4632 15718 4644
rect 15749 4641 15761 4644
rect 15795 4641 15807 4675
rect 15749 4635 15807 4641
rect 15838 4632 15844 4684
rect 15896 4672 15902 4684
rect 16005 4675 16063 4681
rect 16005 4672 16017 4675
rect 15896 4644 16017 4672
rect 15896 4632 15902 4644
rect 16005 4641 16017 4644
rect 16051 4641 16063 4675
rect 16684 4672 16712 4700
rect 18966 4672 18972 4684
rect 16684 4644 18972 4672
rect 16005 4635 16063 4641
rect 12437 4607 12495 4613
rect 12437 4604 12449 4607
rect 11992 4576 12449 4604
rect 12437 4573 12449 4576
rect 12483 4573 12495 4607
rect 13446 4604 13452 4616
rect 13407 4576 13452 4604
rect 12437 4567 12495 4573
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 14458 4604 14464 4616
rect 14419 4576 14464 4604
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 14918 4564 14924 4616
rect 14976 4564 14982 4616
rect 15194 4564 15200 4616
rect 15252 4564 15258 4616
rect 18340 4613 18368 4644
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19245 4675 19303 4681
rect 19245 4641 19257 4675
rect 19291 4672 19303 4675
rect 19886 4672 19892 4684
rect 19291 4644 19892 4672
rect 19291 4641 19303 4644
rect 19245 4635 19303 4641
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 21358 4681 21364 4684
rect 20257 4675 20315 4681
rect 20257 4641 20269 4675
rect 20303 4672 20315 4675
rect 21352 4672 21364 4681
rect 20303 4644 21364 4672
rect 20303 4641 20315 4644
rect 20257 4635 20315 4641
rect 21352 4635 21364 4644
rect 21358 4632 21364 4635
rect 21416 4632 21422 4684
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 18506 4564 18512 4616
rect 18564 4604 18570 4616
rect 19150 4604 19156 4616
rect 18564 4576 19156 4604
rect 18564 4564 18570 4576
rect 19150 4564 19156 4576
rect 19208 4604 19214 4616
rect 19337 4607 19395 4613
rect 19337 4604 19349 4607
rect 19208 4576 19349 4604
rect 19208 4564 19214 4576
rect 19337 4573 19349 4576
rect 19383 4573 19395 4607
rect 19337 4567 19395 4573
rect 19794 4564 19800 4616
rect 19852 4604 19858 4616
rect 20349 4607 20407 4613
rect 20349 4604 20361 4607
rect 19852 4576 20361 4604
rect 19852 4564 19858 4576
rect 20349 4573 20361 4576
rect 20395 4604 20407 4607
rect 20395 4576 20668 4604
rect 20395 4573 20407 4576
rect 20349 4567 20407 4573
rect 10873 4539 10931 4545
rect 10873 4505 10885 4539
rect 10919 4536 10931 4539
rect 15562 4536 15568 4548
rect 10919 4508 15568 4536
rect 10919 4505 10931 4508
rect 10873 4499 10931 4505
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 18785 4539 18843 4545
rect 18785 4505 18797 4539
rect 18831 4536 18843 4539
rect 20640 4536 20668 4576
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21082 4604 21088 4616
rect 20772 4576 21088 4604
rect 20772 4564 20778 4576
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 20898 4536 20904 4548
rect 18831 4508 20484 4536
rect 20640 4508 20904 4536
rect 18831 4505 18843 4508
rect 18785 4499 18843 4505
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 14090 4468 14096 4480
rect 11931 4440 14096 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 14274 4428 14280 4480
rect 14332 4468 14338 4480
rect 14550 4468 14556 4480
rect 14332 4440 14556 4468
rect 14332 4428 14338 4440
rect 14550 4428 14556 4440
rect 14608 4468 14614 4480
rect 15286 4468 15292 4480
rect 14608 4440 15292 4468
rect 14608 4428 14614 4440
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 15746 4428 15752 4480
rect 15804 4468 15810 4480
rect 16666 4468 16672 4480
rect 15804 4440 16672 4468
rect 15804 4428 15810 4440
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 16942 4428 16948 4480
rect 17000 4468 17006 4480
rect 17129 4471 17187 4477
rect 17129 4468 17141 4471
rect 17000 4440 17141 4468
rect 17000 4428 17006 4440
rect 17129 4437 17141 4440
rect 17175 4437 17187 4471
rect 17129 4431 17187 4437
rect 17773 4471 17831 4477
rect 17773 4437 17785 4471
rect 17819 4468 17831 4471
rect 19334 4468 19340 4480
rect 17819 4440 19340 4468
rect 17819 4437 17831 4440
rect 17773 4431 17831 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 20456 4468 20484 4508
rect 20898 4496 20904 4508
rect 20956 4496 20962 4548
rect 22278 4468 22284 4480
rect 20456 4440 22284 4468
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 1104 4378 23276 4400
rect 1104 4326 4680 4378
rect 4732 4326 4744 4378
rect 4796 4326 4808 4378
rect 4860 4326 4872 4378
rect 4924 4326 12078 4378
rect 12130 4326 12142 4378
rect 12194 4326 12206 4378
rect 12258 4326 12270 4378
rect 12322 4326 19475 4378
rect 19527 4326 19539 4378
rect 19591 4326 19603 4378
rect 19655 4326 19667 4378
rect 19719 4326 23276 4378
rect 1104 4304 23276 4326
rect 10226 4224 10232 4276
rect 10284 4264 10290 4276
rect 13998 4264 14004 4276
rect 10284 4236 14004 4264
rect 10284 4224 10290 4236
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 14274 4264 14280 4276
rect 14108 4236 14280 4264
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 10321 4199 10379 4205
rect 10321 4196 10333 4199
rect 9640 4168 10333 4196
rect 9640 4156 9646 4168
rect 10321 4165 10333 4168
rect 10367 4165 10379 4199
rect 10321 4159 10379 4165
rect 10502 4156 10508 4208
rect 10560 4196 10566 4208
rect 11790 4196 11796 4208
rect 10560 4168 11796 4196
rect 10560 4156 10566 4168
rect 10980 4137 11008 4168
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 12618 4156 12624 4208
rect 12676 4196 12682 4208
rect 14108 4196 14136 4236
rect 14274 4224 14280 4236
rect 14332 4224 14338 4276
rect 16206 4264 16212 4276
rect 14384 4236 16212 4264
rect 14384 4196 14412 4236
rect 16206 4224 16212 4236
rect 16264 4264 16270 4276
rect 23198 4264 23204 4276
rect 16264 4236 23204 4264
rect 16264 4224 16270 4236
rect 23198 4224 23204 4236
rect 23256 4224 23262 4276
rect 12676 4168 14136 4196
rect 14292 4168 14412 4196
rect 12676 4156 12682 4168
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 13280 4137 13308 4168
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11756 4100 11897 4128
rect 11756 4088 11762 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13998 4128 14004 4140
rect 13587 4100 14004 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 14292 4137 14320 4168
rect 17770 4156 17776 4208
rect 17828 4196 17834 4208
rect 19518 4196 19524 4208
rect 17828 4168 19524 4196
rect 17828 4156 17834 4168
rect 19518 4156 19524 4168
rect 19576 4156 19582 4208
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14424 4100 14657 4128
rect 14424 4088 14430 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 15654 4088 15660 4140
rect 15712 4128 15718 4140
rect 16298 4128 16304 4140
rect 15712 4100 16304 4128
rect 15712 4088 15718 4100
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 18506 4128 18512 4140
rect 17460 4100 18512 4128
rect 17460 4088 17466 4100
rect 18506 4088 18512 4100
rect 18564 4128 18570 4140
rect 18601 4131 18659 4137
rect 18601 4128 18613 4131
rect 18564 4100 18613 4128
rect 18564 4088 18570 4100
rect 18601 4097 18613 4100
rect 18647 4097 18659 4131
rect 19058 4128 19064 4140
rect 19019 4100 19064 4128
rect 18601 4091 18659 4097
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4060 10747 4063
rect 11054 4060 11060 4072
rect 10735 4032 11060 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 15194 4060 15200 4072
rect 11839 4032 15200 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15286 4020 15292 4072
rect 15344 4060 15350 4072
rect 16557 4063 16615 4069
rect 16557 4060 16569 4063
rect 15344 4032 16569 4060
rect 15344 4020 15350 4032
rect 16557 4029 16569 4032
rect 16603 4060 16615 4063
rect 16942 4060 16948 4072
rect 16603 4032 16948 4060
rect 16603 4029 16615 4032
rect 16557 4023 16615 4029
rect 16942 4020 16948 4032
rect 17000 4020 17006 4072
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 19521 4063 19579 4069
rect 19521 4060 19533 4063
rect 19024 4032 19533 4060
rect 19024 4020 19030 4032
rect 19521 4029 19533 4032
rect 19567 4060 19579 4063
rect 20714 4060 20720 4072
rect 19567 4032 20720 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 20714 4020 20720 4032
rect 20772 4060 20778 4072
rect 21634 4069 21640 4072
rect 21361 4063 21419 4069
rect 21361 4060 21373 4063
rect 20772 4032 21373 4060
rect 20772 4020 20778 4032
rect 21361 4029 21373 4032
rect 21407 4029 21419 4063
rect 21628 4060 21640 4069
rect 21595 4032 21640 4060
rect 21361 4023 21419 4029
rect 21628 4023 21640 4032
rect 21634 4020 21640 4023
rect 21692 4020 21698 4072
rect 10781 3995 10839 4001
rect 10781 3961 10793 3995
rect 10827 3992 10839 3995
rect 12434 3992 12440 4004
rect 10827 3964 12440 3992
rect 10827 3961 10839 3964
rect 10781 3955 10839 3961
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 13814 3992 13820 4004
rect 12636 3964 13820 3992
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 11422 3924 11428 3936
rect 11379 3896 11428 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 11514 3884 11520 3936
rect 11572 3924 11578 3936
rect 12636 3933 12664 3964
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 14918 4001 14924 4004
rect 14001 3995 14059 4001
rect 14001 3961 14013 3995
rect 14047 3992 14059 3995
rect 14047 3964 14872 3992
rect 14047 3961 14059 3964
rect 14001 3955 14059 3961
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11572 3896 11713 3924
rect 11572 3884 11578 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3893 12679 3927
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12621 3887 12679 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13136 3896 13181 3924
rect 13136 3884 13142 3896
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 13633 3927 13691 3933
rect 13633 3924 13645 3927
rect 13320 3896 13645 3924
rect 13320 3884 13326 3896
rect 13633 3893 13645 3896
rect 13679 3893 13691 3927
rect 13633 3887 13691 3893
rect 14093 3927 14151 3933
rect 14093 3893 14105 3927
rect 14139 3924 14151 3927
rect 14642 3924 14648 3936
rect 14139 3896 14648 3924
rect 14139 3893 14151 3896
rect 14093 3887 14151 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 14844 3924 14872 3964
rect 14912 3955 14924 4001
rect 14976 3992 14982 4004
rect 14976 3964 15012 3992
rect 14918 3952 14924 3955
rect 14976 3952 14982 3964
rect 15102 3952 15108 4004
rect 15160 3992 15166 4004
rect 18509 3995 18567 4001
rect 18509 3992 18521 3995
rect 15160 3964 18521 3992
rect 15160 3952 15166 3964
rect 18509 3961 18521 3964
rect 18555 3961 18567 3995
rect 18509 3955 18567 3961
rect 19150 3952 19156 4004
rect 19208 3992 19214 4004
rect 19766 3995 19824 4001
rect 19766 3992 19778 3995
rect 19208 3964 19778 3992
rect 19208 3952 19214 3964
rect 19766 3961 19778 3964
rect 19812 3961 19824 3995
rect 19766 3955 19824 3961
rect 15562 3924 15568 3936
rect 14844 3896 15568 3924
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 16025 3927 16083 3933
rect 16025 3924 16037 3927
rect 15712 3896 16037 3924
rect 15712 3884 15718 3896
rect 16025 3893 16037 3896
rect 16071 3893 16083 3927
rect 16025 3887 16083 3893
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 17681 3927 17739 3933
rect 17681 3924 17693 3927
rect 16632 3896 17693 3924
rect 16632 3884 16638 3896
rect 17681 3893 17693 3896
rect 17727 3893 17739 3927
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 17681 3887 17739 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18414 3924 18420 3936
rect 18375 3896 18420 3924
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20864 3896 20913 3924
rect 20864 3884 20870 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 22741 3927 22799 3933
rect 22741 3924 22753 3927
rect 21416 3896 22753 3924
rect 21416 3884 21422 3896
rect 22741 3893 22753 3896
rect 22787 3893 22799 3927
rect 22741 3887 22799 3893
rect 1104 3834 23276 3856
rect 1104 3782 8379 3834
rect 8431 3782 8443 3834
rect 8495 3782 8507 3834
rect 8559 3782 8571 3834
rect 8623 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 15904 3834
rect 15956 3782 15968 3834
rect 16020 3782 23276 3834
rect 1104 3760 23276 3782
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 12434 3720 12440 3732
rect 11195 3692 12440 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12529 3723 12587 3729
rect 12529 3689 12541 3723
rect 12575 3720 12587 3723
rect 15933 3723 15991 3729
rect 15933 3720 15945 3723
rect 12575 3692 15945 3720
rect 12575 3689 12587 3692
rect 12529 3683 12587 3689
rect 15933 3689 15945 3692
rect 15979 3689 15991 3723
rect 16114 3720 16120 3732
rect 16075 3692 16120 3720
rect 15933 3683 15991 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16485 3723 16543 3729
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 17218 3720 17224 3732
rect 16531 3692 17224 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 18414 3720 18420 3732
rect 17328 3692 18420 3720
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 13081 3655 13139 3661
rect 13081 3652 13093 3655
rect 9272 3624 13093 3652
rect 9272 3612 9278 3624
rect 13081 3621 13093 3624
rect 13127 3621 13139 3655
rect 13538 3652 13544 3664
rect 13499 3624 13544 3652
rect 13081 3615 13139 3621
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 13630 3612 13636 3664
rect 13688 3652 13694 3664
rect 13688 3624 13733 3652
rect 13688 3612 13694 3624
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 17328 3652 17356 3692
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 21634 3680 21640 3732
rect 21692 3720 21698 3732
rect 22741 3723 22799 3729
rect 22741 3720 22753 3723
rect 21692 3692 22753 3720
rect 21692 3680 21698 3692
rect 22741 3689 22753 3692
rect 22787 3689 22799 3723
rect 22741 3683 22799 3689
rect 17402 3661 17408 3664
rect 13872 3624 17356 3652
rect 13872 3612 13878 3624
rect 17396 3615 17408 3661
rect 17460 3652 17466 3664
rect 20901 3655 20959 3661
rect 20901 3652 20913 3655
rect 17460 3624 17496 3652
rect 18708 3624 20913 3652
rect 17402 3612 17408 3615
rect 17460 3612 17466 3624
rect 11514 3584 11520 3596
rect 11475 3556 11520 3584
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 14550 3584 14556 3596
rect 12667 3556 14044 3584
rect 14511 3556 14556 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 11609 3479 11667 3485
rect 11624 3380 11652 3479
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 12802 3516 12808 3528
rect 11940 3488 12808 3516
rect 11940 3476 11946 3488
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 13722 3516 13728 3528
rect 13683 3488 13728 3516
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 12161 3451 12219 3457
rect 12161 3417 12173 3451
rect 12207 3448 12219 3451
rect 13814 3448 13820 3460
rect 12207 3420 13820 3448
rect 12207 3417 12219 3420
rect 12161 3411 12219 3417
rect 13814 3408 13820 3420
rect 13872 3408 13878 3460
rect 14016 3448 14044 3556
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 15010 3584 15016 3596
rect 14691 3556 15016 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3584 15623 3587
rect 15930 3584 15936 3596
rect 15611 3556 15936 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 18708 3584 18736 3624
rect 20901 3621 20913 3624
rect 20947 3621 20959 3655
rect 20901 3615 20959 3621
rect 19242 3593 19248 3596
rect 19236 3584 19248 3593
rect 16540 3556 18736 3584
rect 19203 3556 19248 3584
rect 16540 3544 16546 3556
rect 19236 3547 19248 3556
rect 19242 3544 19248 3547
rect 19300 3544 19306 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 21361 3587 21419 3593
rect 21361 3584 21373 3587
rect 20772 3556 21373 3584
rect 20772 3544 20778 3556
rect 21361 3553 21373 3556
rect 21407 3553 21419 3587
rect 21361 3547 21419 3553
rect 21628 3587 21686 3593
rect 21628 3553 21640 3587
rect 21674 3584 21686 3587
rect 21910 3584 21916 3596
rect 21674 3556 21916 3584
rect 21674 3553 21686 3556
rect 21628 3547 21686 3553
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 14734 3516 14740 3528
rect 14695 3488 14740 3516
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 14884 3488 16589 3516
rect 14884 3476 14890 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 15933 3451 15991 3457
rect 14016 3420 15884 3448
rect 12894 3380 12900 3392
rect 11624 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13081 3383 13139 3389
rect 13081 3349 13093 3383
rect 13127 3380 13139 3383
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 13127 3352 13185 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 14185 3383 14243 3389
rect 14185 3349 14197 3383
rect 14231 3380 14243 3383
rect 14366 3380 14372 3392
rect 14231 3352 14372 3380
rect 14231 3349 14243 3352
rect 14185 3343 14243 3349
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 15562 3340 15568 3392
rect 15620 3380 15626 3392
rect 15749 3383 15807 3389
rect 15749 3380 15761 3383
rect 15620 3352 15761 3380
rect 15620 3340 15626 3352
rect 15749 3349 15761 3352
rect 15795 3349 15807 3383
rect 15856 3380 15884 3420
rect 15933 3417 15945 3451
rect 15979 3448 15991 3451
rect 16114 3448 16120 3460
rect 15979 3420 16120 3448
rect 15979 3417 15991 3420
rect 15933 3411 15991 3417
rect 16114 3408 16120 3420
rect 16172 3408 16178 3460
rect 16390 3408 16396 3460
rect 16448 3448 16454 3460
rect 16684 3448 16712 3479
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 17092 3488 17141 3516
rect 17092 3476 17098 3488
rect 17129 3485 17141 3488
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18966 3516 18972 3528
rect 18380 3488 18972 3516
rect 18380 3476 18386 3488
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 16448 3420 16712 3448
rect 16448 3408 16454 3420
rect 18414 3408 18420 3460
rect 18472 3448 18478 3460
rect 18472 3420 18736 3448
rect 18472 3408 18478 3420
rect 18509 3383 18567 3389
rect 18509 3380 18521 3383
rect 15856 3352 18521 3380
rect 15749 3343 15807 3349
rect 18509 3349 18521 3352
rect 18555 3380 18567 3383
rect 18598 3380 18604 3392
rect 18555 3352 18604 3380
rect 18555 3349 18567 3352
rect 18509 3343 18567 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 18708 3380 18736 3420
rect 19150 3380 19156 3392
rect 18708 3352 19156 3380
rect 19150 3340 19156 3352
rect 19208 3380 19214 3392
rect 20349 3383 20407 3389
rect 20349 3380 20361 3383
rect 19208 3352 20361 3380
rect 19208 3340 19214 3352
rect 20349 3349 20361 3352
rect 20395 3349 20407 3383
rect 20349 3343 20407 3349
rect 1104 3290 23276 3312
rect 1104 3238 4680 3290
rect 4732 3238 4744 3290
rect 4796 3238 4808 3290
rect 4860 3238 4872 3290
rect 4924 3238 12078 3290
rect 12130 3238 12142 3290
rect 12194 3238 12206 3290
rect 12258 3238 12270 3290
rect 12322 3238 19475 3290
rect 19527 3238 19539 3290
rect 19591 3238 19603 3290
rect 19655 3238 19667 3290
rect 19719 3238 23276 3290
rect 1104 3216 23276 3238
rect 13265 3179 13323 3185
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 15102 3176 15108 3188
rect 13311 3148 15108 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 15470 3176 15476 3188
rect 15335 3148 15476 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 17402 3176 17408 3188
rect 15580 3148 17408 3176
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 14090 3108 14096 3120
rect 11572 3080 14096 3108
rect 11572 3068 11578 3080
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14274 3108 14280 3120
rect 14235 3080 14280 3108
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 15010 3108 15016 3120
rect 14568 3080 15016 3108
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 12802 3000 12808 3052
rect 12860 3040 12866 3052
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 12860 3012 13921 3040
rect 12860 3000 12866 3012
rect 13909 3009 13921 3012
rect 13955 3040 13967 3043
rect 14568 3040 14596 3080
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 14734 3040 14740 3052
rect 13955 3012 14596 3040
rect 14695 3012 14740 3040
rect 13955 3009 13967 3012
rect 13909 3003 13967 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3040 14979 3043
rect 15378 3040 15384 3052
rect 14967 3012 15384 3040
rect 14967 3009 14979 3012
rect 14921 3003 14979 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2972 1823 2975
rect 2406 2972 2412 2984
rect 1811 2944 2412 2972
rect 1811 2941 1823 2944
rect 1765 2935 1823 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2507 2975 2565 2981
rect 2507 2941 2519 2975
rect 2553 2941 2565 2975
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 2507 2935 2565 2941
rect 2516 2904 2544 2935
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 13633 2975 13691 2981
rect 6052 2944 12204 2972
rect 6052 2932 6058 2944
rect 12176 2904 12204 2944
rect 13633 2941 13645 2975
rect 13679 2972 13691 2975
rect 15580 2972 15608 3148
rect 17402 3136 17408 3148
rect 17460 3176 17466 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17460 3148 17693 3176
rect 17460 3136 17466 3148
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 19150 3136 19156 3188
rect 19208 3136 19214 3188
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19300 3148 19625 3176
rect 19300 3136 19306 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 19613 3139 19671 3145
rect 19720 3148 21680 3176
rect 15838 3068 15844 3120
rect 15896 3108 15902 3120
rect 16206 3108 16212 3120
rect 15896 3080 16212 3108
rect 15896 3068 15902 3080
rect 16206 3068 16212 3080
rect 16264 3068 16270 3120
rect 19168 3108 19196 3136
rect 19720 3108 19748 3148
rect 19168 3080 19748 3108
rect 21652 3108 21680 3148
rect 21910 3136 21916 3188
rect 21968 3176 21974 3188
rect 22097 3179 22155 3185
rect 22097 3176 22109 3179
rect 21968 3148 22109 3176
rect 21968 3136 21974 3148
rect 22097 3145 22109 3148
rect 22143 3145 22155 3179
rect 22097 3139 22155 3145
rect 22557 3111 22615 3117
rect 22557 3108 22569 3111
rect 21652 3080 22569 3108
rect 22557 3077 22569 3080
rect 22603 3077 22615 3111
rect 22557 3071 22615 3077
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16022 3040 16028 3052
rect 15979 3012 16028 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 16298 3040 16304 3052
rect 16259 3012 16304 3040
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 20714 3040 20720 3052
rect 17460 3012 18368 3040
rect 20675 3012 20720 3040
rect 17460 3000 17466 3012
rect 13679 2944 15608 2972
rect 15657 2975 15715 2981
rect 13679 2941 13691 2944
rect 13633 2935 13691 2941
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 15746 2972 15752 2984
rect 15703 2944 15752 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 16574 2981 16580 2984
rect 16568 2972 16580 2981
rect 16040 2944 16580 2972
rect 14645 2907 14703 2913
rect 14645 2904 14657 2907
rect 2516 2876 9076 2904
rect 12176 2876 14657 2904
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 1728 2808 2697 2836
rect 1728 2796 1734 2808
rect 2685 2805 2697 2808
rect 2731 2805 2743 2839
rect 9048 2836 9076 2876
rect 14645 2873 14657 2876
rect 14691 2873 14703 2907
rect 16040 2904 16068 2944
rect 16568 2935 16580 2944
rect 16574 2932 16580 2935
rect 16632 2932 16638 2984
rect 17586 2972 17592 2984
rect 16776 2944 17592 2972
rect 16776 2904 16804 2944
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18340 2972 18368 3012
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 19242 2972 19248 2984
rect 18340 2944 19248 2972
rect 18233 2935 18291 2941
rect 14645 2867 14703 2873
rect 15672 2876 16068 2904
rect 16316 2876 16804 2904
rect 11974 2836 11980 2848
rect 9048 2808 11980 2836
rect 2685 2799 2743 2805
rect 11974 2796 11980 2808
rect 12032 2836 12038 2848
rect 13630 2836 13636 2848
rect 12032 2808 13636 2836
rect 12032 2796 12038 2808
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 15672 2836 15700 2876
rect 13771 2808 15700 2836
rect 15749 2839 15807 2845
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 15749 2805 15761 2839
rect 15795 2836 15807 2839
rect 16316 2836 16344 2876
rect 17034 2864 17040 2916
rect 17092 2904 17098 2916
rect 18246 2904 18274 2935
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 21450 2972 21456 2984
rect 20027 2944 21456 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 21450 2932 21456 2944
rect 21508 2972 21514 2984
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 21508 2944 22385 2972
rect 21508 2932 21514 2944
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 18322 2904 18328 2916
rect 17092 2876 18328 2904
rect 17092 2864 17098 2876
rect 18322 2864 18328 2876
rect 18380 2864 18386 2916
rect 18500 2907 18558 2913
rect 18500 2873 18512 2907
rect 18546 2873 18558 2907
rect 18500 2867 18558 2873
rect 20257 2907 20315 2913
rect 20257 2873 20269 2907
rect 20303 2873 20315 2907
rect 20257 2867 20315 2873
rect 15795 2808 16344 2836
rect 15795 2805 15807 2808
rect 15749 2799 15807 2805
rect 16390 2796 16396 2848
rect 16448 2836 16454 2848
rect 18524 2836 18552 2867
rect 19058 2836 19064 2848
rect 16448 2808 19064 2836
rect 16448 2796 16454 2808
rect 19058 2796 19064 2808
rect 19116 2796 19122 2848
rect 20272 2836 20300 2867
rect 20898 2864 20904 2916
rect 20956 2913 20962 2916
rect 20956 2907 21020 2913
rect 20956 2873 20974 2907
rect 21008 2873 21020 2907
rect 20956 2867 21020 2873
rect 20956 2864 20962 2867
rect 22554 2836 22560 2848
rect 20272 2808 22560 2836
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 1104 2746 23276 2768
rect 1104 2694 8379 2746
rect 8431 2694 8443 2746
rect 8495 2694 8507 2746
rect 8559 2694 8571 2746
rect 8623 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 15904 2746
rect 15956 2694 15968 2746
rect 16020 2694 23276 2746
rect 1104 2672 23276 2694
rect 13354 2632 13360 2644
rect 13315 2604 13360 2632
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 13817 2635 13875 2641
rect 13817 2601 13829 2635
rect 13863 2632 13875 2635
rect 14829 2635 14887 2641
rect 13863 2604 14688 2632
rect 13863 2601 13875 2604
rect 13817 2595 13875 2601
rect 11790 2524 11796 2576
rect 11848 2564 11854 2576
rect 11848 2536 13952 2564
rect 11848 2524 11854 2536
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2465 13783 2499
rect 13725 2459 13783 2465
rect 13740 2360 13768 2459
rect 13924 2437 13952 2536
rect 14660 2496 14688 2604
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 15654 2632 15660 2644
rect 14875 2604 15660 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2601 16267 2635
rect 16209 2595 16267 2601
rect 16669 2635 16727 2641
rect 16669 2601 16681 2635
rect 16715 2632 16727 2635
rect 17402 2632 17408 2644
rect 16715 2604 17408 2632
rect 16715 2601 16727 2604
rect 16669 2595 16727 2601
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 15286 2564 15292 2576
rect 14783 2536 15292 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 15654 2496 15660 2508
rect 14660 2468 15339 2496
rect 15615 2468 15660 2496
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2397 13967 2431
rect 15010 2428 15016 2440
rect 14971 2400 15016 2428
rect 13909 2391 13967 2397
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15311 2428 15339 2468
rect 15654 2456 15660 2468
rect 15712 2456 15718 2508
rect 16224 2496 16252 2595
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 17589 2635 17647 2641
rect 17589 2601 17601 2635
rect 17635 2632 17647 2635
rect 17635 2604 19012 2632
rect 17635 2601 17647 2604
rect 17589 2595 17647 2601
rect 16577 2567 16635 2573
rect 16577 2533 16589 2567
rect 16623 2564 16635 2567
rect 18414 2564 18420 2576
rect 16623 2536 18420 2564
rect 16623 2533 16635 2536
rect 16577 2527 16635 2533
rect 18414 2524 18420 2536
rect 18472 2524 18478 2576
rect 18598 2573 18604 2576
rect 18592 2564 18604 2573
rect 18559 2536 18604 2564
rect 18592 2527 18604 2536
rect 18598 2524 18604 2527
rect 18656 2524 18662 2576
rect 18984 2564 19012 2604
rect 19058 2592 19064 2644
rect 19116 2632 19122 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 19116 2604 19717 2632
rect 19116 2592 19122 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 20073 2635 20131 2641
rect 20073 2601 20085 2635
rect 20119 2632 20131 2635
rect 20254 2632 20260 2644
rect 20119 2604 20260 2632
rect 20119 2601 20131 2604
rect 20073 2595 20131 2601
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 20533 2635 20591 2641
rect 20533 2632 20545 2635
rect 20496 2604 20545 2632
rect 20496 2592 20502 2604
rect 20533 2601 20545 2604
rect 20579 2601 20591 2635
rect 20533 2595 20591 2601
rect 22557 2635 22615 2641
rect 22557 2601 22569 2635
rect 22603 2601 22615 2635
rect 22557 2595 22615 2601
rect 20898 2564 20904 2576
rect 18984 2536 20904 2564
rect 20898 2524 20904 2536
rect 20956 2564 20962 2576
rect 22572 2564 22600 2595
rect 20956 2536 22600 2564
rect 20956 2524 20962 2536
rect 16298 2496 16304 2508
rect 16224 2468 16304 2496
rect 16298 2456 16304 2468
rect 16356 2456 16362 2508
rect 16942 2496 16948 2508
rect 16855 2468 16948 2496
rect 16758 2428 16764 2440
rect 15311 2400 16764 2428
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 16868 2437 16896 2468
rect 16942 2456 16948 2468
rect 17000 2496 17006 2508
rect 18322 2496 18328 2508
rect 17000 2468 17816 2496
rect 18283 2468 18328 2496
rect 17000 2456 17006 2468
rect 17788 2440 17816 2468
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19392 2468 20453 2496
rect 19392 2456 19398 2468
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 20441 2459 20499 2465
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20772 2468 21189 2496
rect 20772 2456 20778 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 21433 2499 21491 2505
rect 21433 2496 21445 2499
rect 21177 2459 21235 2465
rect 21284 2468 21445 2496
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2397 16911 2431
rect 17678 2428 17684 2440
rect 17639 2400 17684 2428
rect 16853 2391 16911 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 20625 2431 20683 2437
rect 17828 2400 17873 2428
rect 17828 2388 17834 2400
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 20990 2428 20996 2440
rect 20671 2400 20996 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 21284 2428 21312 2468
rect 21433 2465 21445 2468
rect 21479 2465 21491 2499
rect 21433 2459 21491 2465
rect 21192 2400 21312 2428
rect 17586 2360 17592 2372
rect 13740 2332 17592 2360
rect 17586 2320 17592 2332
rect 17644 2320 17650 2372
rect 20806 2320 20812 2372
rect 20864 2360 20870 2372
rect 21192 2360 21220 2400
rect 20864 2332 21220 2360
rect 20864 2320 20870 2332
rect 14369 2295 14427 2301
rect 14369 2261 14381 2295
rect 14415 2292 14427 2295
rect 14458 2292 14464 2304
rect 14415 2264 14464 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 15841 2295 15899 2301
rect 15841 2261 15853 2295
rect 15887 2292 15899 2295
rect 16574 2292 16580 2304
rect 15887 2264 16580 2292
rect 15887 2261 15899 2264
rect 15841 2255 15899 2261
rect 16574 2252 16580 2264
rect 16632 2252 16638 2304
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2292 17279 2295
rect 19978 2292 19984 2304
rect 17267 2264 19984 2292
rect 17267 2261 17279 2264
rect 17221 2255 17279 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 1104 2202 23276 2224
rect 1104 2150 4680 2202
rect 4732 2150 4744 2202
rect 4796 2150 4808 2202
rect 4860 2150 4872 2202
rect 4924 2150 12078 2202
rect 12130 2150 12142 2202
rect 12194 2150 12206 2202
rect 12258 2150 12270 2202
rect 12322 2150 19475 2202
rect 19527 2150 19539 2202
rect 19591 2150 19603 2202
rect 19655 2150 19667 2202
rect 19719 2150 23276 2202
rect 1104 2128 23276 2150
rect 16298 2048 16304 2100
rect 16356 2088 16362 2100
rect 18690 2088 18696 2100
rect 16356 2060 18696 2088
rect 16356 2048 16362 2060
rect 18690 2048 18696 2060
rect 18748 2048 18754 2100
rect 17678 1912 17684 1964
rect 17736 1952 17742 1964
rect 20806 1952 20812 1964
rect 17736 1924 20812 1952
rect 17736 1912 17742 1924
rect 20806 1912 20812 1924
rect 20864 1912 20870 1964
rect 17310 1300 17316 1352
rect 17368 1340 17374 1352
rect 19334 1340 19340 1352
rect 17368 1312 19340 1340
rect 17368 1300 17374 1312
rect 19334 1300 19340 1312
rect 19392 1300 19398 1352
<< via1 >>
rect 9956 21904 10008 21956
rect 16948 21904 17000 21956
rect 11060 21836 11112 21888
rect 13728 21836 13780 21888
rect 18328 21836 18380 21888
rect 20444 21836 20496 21888
rect 4680 21734 4732 21786
rect 4744 21734 4796 21786
rect 4808 21734 4860 21786
rect 4872 21734 4924 21786
rect 12078 21734 12130 21786
rect 12142 21734 12194 21786
rect 12206 21734 12258 21786
rect 12270 21734 12322 21786
rect 19475 21734 19527 21786
rect 19539 21734 19591 21786
rect 19603 21734 19655 21786
rect 19667 21734 19719 21786
rect 1492 21632 1544 21684
rect 9956 21675 10008 21684
rect 9956 21641 9965 21675
rect 9965 21641 9999 21675
rect 9999 21641 10008 21675
rect 9956 21632 10008 21641
rect 16396 21632 16448 21684
rect 19248 21632 19300 21684
rect 16764 21564 16816 21616
rect 21824 21564 21876 21616
rect 2596 21539 2648 21548
rect 2596 21505 2605 21539
rect 2605 21505 2639 21539
rect 2639 21505 2648 21539
rect 2596 21496 2648 21505
rect 5540 21496 5592 21548
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 16580 21496 16632 21548
rect 21456 21496 21508 21548
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 4160 21428 4212 21480
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 2596 21360 2648 21412
rect 3792 21360 3844 21412
rect 9956 21428 10008 21480
rect 10416 21428 10468 21480
rect 12164 21428 12216 21480
rect 14832 21471 14884 21480
rect 14832 21437 14841 21471
rect 14841 21437 14875 21471
rect 14875 21437 14884 21471
rect 14832 21428 14884 21437
rect 15476 21428 15528 21480
rect 18236 21428 18288 21480
rect 18328 21471 18380 21480
rect 18328 21437 18337 21471
rect 18337 21437 18371 21471
rect 18371 21437 18380 21471
rect 18328 21428 18380 21437
rect 18788 21428 18840 21480
rect 6460 21360 6512 21412
rect 7748 21360 7800 21412
rect 8852 21403 8904 21412
rect 8852 21369 8861 21403
rect 8861 21369 8895 21403
rect 8895 21369 8904 21403
rect 8852 21360 8904 21369
rect 11704 21360 11756 21412
rect 14464 21360 14516 21412
rect 19892 21428 19944 21480
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 22284 21428 22336 21480
rect 1952 21335 2004 21344
rect 1952 21301 1961 21335
rect 1961 21301 1995 21335
rect 1995 21301 2004 21335
rect 1952 21292 2004 21301
rect 2504 21292 2556 21344
rect 2964 21335 3016 21344
rect 2964 21301 2973 21335
rect 2973 21301 3007 21335
rect 3007 21301 3016 21335
rect 2964 21292 3016 21301
rect 3332 21335 3384 21344
rect 3332 21301 3341 21335
rect 3341 21301 3375 21335
rect 3375 21301 3384 21335
rect 3332 21292 3384 21301
rect 3424 21335 3476 21344
rect 3424 21301 3433 21335
rect 3433 21301 3467 21335
rect 3467 21301 3476 21335
rect 4068 21335 4120 21344
rect 3424 21292 3476 21301
rect 4068 21301 4077 21335
rect 4077 21301 4111 21335
rect 4111 21301 4120 21335
rect 4068 21292 4120 21301
rect 4436 21335 4488 21344
rect 4436 21301 4445 21335
rect 4445 21301 4479 21335
rect 4479 21301 4488 21335
rect 4436 21292 4488 21301
rect 4528 21335 4580 21344
rect 4528 21301 4537 21335
rect 4537 21301 4571 21335
rect 4571 21301 4580 21335
rect 5264 21335 5316 21344
rect 4528 21292 4580 21301
rect 5264 21301 5273 21335
rect 5273 21301 5307 21335
rect 5307 21301 5316 21335
rect 5264 21292 5316 21301
rect 5816 21335 5868 21344
rect 5816 21301 5825 21335
rect 5825 21301 5859 21335
rect 5859 21301 5868 21335
rect 5816 21292 5868 21301
rect 5908 21292 5960 21344
rect 6920 21335 6972 21344
rect 6920 21301 6929 21335
rect 6929 21301 6963 21335
rect 6963 21301 6972 21335
rect 6920 21292 6972 21301
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 8668 21292 8720 21344
rect 8760 21335 8812 21344
rect 8760 21301 8769 21335
rect 8769 21301 8803 21335
rect 8803 21301 8812 21335
rect 8760 21292 8812 21301
rect 12256 21292 12308 21344
rect 12900 21292 12952 21344
rect 13728 21292 13780 21344
rect 19340 21360 19392 21412
rect 15568 21292 15620 21344
rect 16212 21292 16264 21344
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 16948 21335 17000 21344
rect 16948 21301 16957 21335
rect 16957 21301 16991 21335
rect 16991 21301 17000 21335
rect 16948 21292 17000 21301
rect 20352 21360 20404 21412
rect 20260 21335 20312 21344
rect 20260 21301 20269 21335
rect 20269 21301 20303 21335
rect 20303 21301 20312 21335
rect 20260 21292 20312 21301
rect 21916 21360 21968 21412
rect 21548 21335 21600 21344
rect 21548 21301 21557 21335
rect 21557 21301 21591 21335
rect 21591 21301 21600 21335
rect 21548 21292 21600 21301
rect 21640 21335 21692 21344
rect 21640 21301 21649 21335
rect 21649 21301 21683 21335
rect 21683 21301 21692 21335
rect 21640 21292 21692 21301
rect 23204 21292 23256 21344
rect 8379 21190 8431 21242
rect 8443 21190 8495 21242
rect 8507 21190 8559 21242
rect 8571 21190 8623 21242
rect 15776 21190 15828 21242
rect 15840 21190 15892 21242
rect 15904 21190 15956 21242
rect 15968 21190 16020 21242
rect 296 21088 348 21140
rect 4068 21088 4120 21140
rect 7380 21088 7432 21140
rect 8852 21088 8904 21140
rect 9036 21088 9088 21140
rect 16488 21088 16540 21140
rect 19156 21088 19208 21140
rect 2964 21020 3016 21072
rect 3424 20952 3476 21004
rect 1492 20884 1544 20936
rect 4344 20884 4396 20936
rect 5448 21020 5500 21072
rect 5172 20952 5224 21004
rect 7748 21020 7800 21072
rect 8668 21020 8720 21072
rect 13728 21020 13780 21072
rect 6460 20952 6512 21004
rect 6736 20952 6788 21004
rect 10048 20995 10100 21004
rect 10048 20961 10057 20995
rect 10057 20961 10091 20995
rect 10091 20961 10100 20995
rect 10048 20952 10100 20961
rect 12256 20952 12308 21004
rect 13176 20952 13228 21004
rect 3976 20816 4028 20868
rect 3332 20791 3384 20800
rect 3332 20757 3341 20791
rect 3341 20757 3375 20791
rect 3375 20757 3384 20791
rect 3332 20748 3384 20757
rect 4252 20748 4304 20800
rect 10416 20884 10468 20936
rect 14648 20952 14700 21004
rect 17316 20952 17368 21004
rect 18052 21020 18104 21072
rect 18236 21020 18288 21072
rect 20352 21088 20404 21140
rect 20260 21020 20312 21072
rect 21640 21020 21692 21072
rect 19800 20952 19852 21004
rect 20628 20952 20680 21004
rect 14924 20884 14976 20936
rect 18788 20884 18840 20936
rect 19156 20927 19208 20936
rect 19156 20893 19165 20927
rect 19165 20893 19199 20927
rect 19199 20893 19208 20927
rect 19156 20884 19208 20893
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 6828 20748 6880 20800
rect 12256 20816 12308 20868
rect 9772 20748 9824 20800
rect 12532 20748 12584 20800
rect 14004 20748 14056 20800
rect 14464 20791 14516 20800
rect 14464 20757 14473 20791
rect 14473 20757 14507 20791
rect 14507 20757 14516 20791
rect 14464 20748 14516 20757
rect 15200 20748 15252 20800
rect 19340 20748 19392 20800
rect 20168 20748 20220 20800
rect 21548 20748 21600 20800
rect 4680 20646 4732 20698
rect 4744 20646 4796 20698
rect 4808 20646 4860 20698
rect 4872 20646 4924 20698
rect 12078 20646 12130 20698
rect 12142 20646 12194 20698
rect 12206 20646 12258 20698
rect 12270 20646 12322 20698
rect 19475 20646 19527 20698
rect 19539 20646 19591 20698
rect 19603 20646 19655 20698
rect 19667 20646 19719 20698
rect 3424 20544 3476 20596
rect 3608 20544 3660 20596
rect 4436 20544 4488 20596
rect 6460 20587 6512 20596
rect 6460 20553 6469 20587
rect 6469 20553 6503 20587
rect 6503 20553 6512 20587
rect 6460 20544 6512 20553
rect 7748 20544 7800 20596
rect 8760 20544 8812 20596
rect 11704 20544 11756 20596
rect 14648 20587 14700 20596
rect 14648 20553 14657 20587
rect 14657 20553 14691 20587
rect 14691 20553 14700 20587
rect 14648 20544 14700 20553
rect 1400 20340 1452 20392
rect 3056 20340 3108 20392
rect 2320 20272 2372 20324
rect 4528 20340 4580 20392
rect 5908 20340 5960 20392
rect 6736 20340 6788 20392
rect 5632 20272 5684 20324
rect 6368 20272 6420 20324
rect 13176 20408 13228 20460
rect 19248 20544 19300 20596
rect 19800 20544 19852 20596
rect 16948 20476 17000 20528
rect 19156 20476 19208 20528
rect 7380 20340 7432 20392
rect 7840 20340 7892 20392
rect 9036 20340 9088 20392
rect 10232 20340 10284 20392
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 11980 20340 12032 20392
rect 12808 20340 12860 20392
rect 14464 20340 14516 20392
rect 10140 20272 10192 20324
rect 11520 20272 11572 20324
rect 12440 20272 12492 20324
rect 848 20204 900 20256
rect 5264 20204 5316 20256
rect 5448 20204 5500 20256
rect 14556 20272 14608 20324
rect 16764 20408 16816 20460
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 19432 20408 19484 20460
rect 19892 20408 19944 20460
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 20444 20408 20496 20460
rect 14924 20383 14976 20392
rect 14924 20349 14933 20383
rect 14933 20349 14967 20383
rect 14967 20349 14976 20383
rect 15200 20383 15252 20392
rect 14924 20340 14976 20349
rect 15200 20349 15234 20383
rect 15234 20349 15252 20383
rect 15200 20340 15252 20349
rect 16212 20340 16264 20392
rect 18052 20383 18104 20392
rect 15292 20272 15344 20324
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 19156 20272 19208 20324
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 17960 20204 18012 20256
rect 19984 20272 20036 20324
rect 20260 20272 20312 20324
rect 20904 20340 20956 20392
rect 21548 20340 21600 20392
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 24032 20272 24084 20324
rect 19708 20247 19760 20256
rect 19708 20213 19717 20247
rect 19717 20213 19751 20247
rect 19751 20213 19760 20247
rect 19708 20204 19760 20213
rect 21732 20204 21784 20256
rect 22928 20204 22980 20256
rect 8379 20102 8431 20154
rect 8443 20102 8495 20154
rect 8507 20102 8559 20154
rect 8571 20102 8623 20154
rect 15776 20102 15828 20154
rect 15840 20102 15892 20154
rect 15904 20102 15956 20154
rect 15968 20102 16020 20154
rect 2136 20000 2188 20052
rect 4160 20000 4212 20052
rect 6920 20000 6972 20052
rect 9864 20000 9916 20052
rect 10140 20000 10192 20052
rect 11612 20000 11664 20052
rect 11980 20000 12032 20052
rect 12072 20000 12124 20052
rect 13084 20000 13136 20052
rect 13728 20000 13780 20052
rect 14004 20043 14056 20052
rect 14004 20009 14013 20043
rect 14013 20009 14047 20043
rect 14047 20009 14056 20043
rect 14004 20000 14056 20009
rect 14556 20000 14608 20052
rect 19156 20043 19208 20052
rect 4436 19932 4488 19984
rect 5080 19932 5132 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 2780 19864 2832 19916
rect 3148 19864 3200 19916
rect 3608 19864 3660 19916
rect 4068 19796 4120 19848
rect 5632 19864 5684 19916
rect 5816 19932 5868 19984
rect 8576 19932 8628 19984
rect 9220 19864 9272 19916
rect 9864 19907 9916 19916
rect 9864 19873 9873 19907
rect 9873 19873 9907 19907
rect 9907 19873 9916 19907
rect 9864 19864 9916 19873
rect 6828 19839 6880 19848
rect 3240 19728 3292 19780
rect 3884 19728 3936 19780
rect 5908 19728 5960 19780
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 7840 19796 7892 19848
rect 8944 19796 8996 19848
rect 2320 19660 2372 19712
rect 5080 19660 5132 19712
rect 5448 19660 5500 19712
rect 7288 19660 7340 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 8208 19660 8260 19712
rect 8300 19660 8352 19712
rect 9680 19660 9732 19712
rect 10232 19796 10284 19848
rect 10692 19907 10744 19916
rect 10692 19873 10726 19907
rect 10726 19873 10744 19907
rect 10692 19864 10744 19873
rect 11244 19864 11296 19916
rect 11980 19864 12032 19916
rect 12532 19932 12584 19984
rect 16304 19932 16356 19984
rect 19156 20009 19165 20043
rect 19165 20009 19199 20043
rect 19199 20009 19208 20043
rect 19156 20000 19208 20009
rect 19432 19932 19484 19984
rect 19800 19975 19852 19984
rect 19800 19941 19809 19975
rect 19809 19941 19843 19975
rect 19843 19941 19852 19975
rect 19800 19932 19852 19941
rect 15016 19864 15068 19916
rect 19340 19864 19392 19916
rect 14188 19839 14240 19848
rect 14188 19805 14197 19839
rect 14197 19805 14231 19839
rect 14231 19805 14240 19839
rect 14188 19796 14240 19805
rect 14832 19796 14884 19848
rect 14924 19796 14976 19848
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 17500 19796 17552 19848
rect 18788 19796 18840 19848
rect 21364 19864 21416 19916
rect 21640 19907 21692 19916
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 22008 19864 22060 19916
rect 22652 19864 22704 19916
rect 19892 19796 19944 19848
rect 20444 19796 20496 19848
rect 21456 19796 21508 19848
rect 21732 19839 21784 19848
rect 11612 19660 11664 19712
rect 12440 19660 12492 19712
rect 12716 19660 12768 19712
rect 13084 19660 13136 19712
rect 16488 19728 16540 19780
rect 17408 19703 17460 19712
rect 17408 19669 17417 19703
rect 17417 19669 17451 19703
rect 17451 19669 17460 19703
rect 17408 19660 17460 19669
rect 20812 19728 20864 19780
rect 21180 19728 21232 19780
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 19892 19660 19944 19712
rect 21364 19660 21416 19712
rect 4680 19558 4732 19610
rect 4744 19558 4796 19610
rect 4808 19558 4860 19610
rect 4872 19558 4924 19610
rect 12078 19558 12130 19610
rect 12142 19558 12194 19610
rect 12206 19558 12258 19610
rect 12270 19558 12322 19610
rect 19475 19558 19527 19610
rect 19539 19558 19591 19610
rect 19603 19558 19655 19610
rect 19667 19558 19719 19610
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 2412 19252 2464 19304
rect 3056 19295 3108 19304
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 3332 19295 3384 19304
rect 3332 19261 3366 19295
rect 3366 19261 3384 19295
rect 3332 19252 3384 19261
rect 2228 19184 2280 19236
rect 4528 19456 4580 19508
rect 4344 19320 4396 19372
rect 4528 19320 4580 19372
rect 6644 19456 6696 19508
rect 7840 19456 7892 19508
rect 8852 19456 8904 19508
rect 4988 19388 5040 19440
rect 6552 19388 6604 19440
rect 5540 19320 5592 19372
rect 6460 19320 6512 19372
rect 10416 19456 10468 19508
rect 12532 19456 12584 19508
rect 10508 19388 10560 19440
rect 11152 19388 11204 19440
rect 4436 19252 4488 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 5264 19184 5316 19236
rect 8300 19252 8352 19304
rect 14188 19456 14240 19508
rect 15292 19456 15344 19508
rect 8484 19184 8536 19236
rect 10048 19252 10100 19304
rect 13636 19320 13688 19372
rect 8668 19184 8720 19236
rect 8760 19184 8812 19236
rect 4712 19159 4764 19168
rect 4712 19125 4721 19159
rect 4721 19125 4755 19159
rect 4755 19125 4764 19159
rect 4712 19116 4764 19125
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 5816 19116 5868 19168
rect 6828 19116 6880 19168
rect 8116 19116 8168 19168
rect 12992 19252 13044 19304
rect 13728 19295 13780 19304
rect 13728 19261 13737 19295
rect 13737 19261 13771 19295
rect 13771 19261 13780 19295
rect 13728 19252 13780 19261
rect 14924 19388 14976 19440
rect 14648 19320 14700 19372
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 15016 19320 15068 19372
rect 17132 19388 17184 19440
rect 19340 19456 19392 19508
rect 20260 19456 20312 19508
rect 20628 19456 20680 19508
rect 20076 19388 20128 19440
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 16120 19320 16172 19372
rect 19800 19320 19852 19372
rect 17040 19252 17092 19304
rect 17500 19252 17552 19304
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 19064 19252 19116 19304
rect 20904 19252 20956 19304
rect 12900 19227 12952 19236
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 12348 19116 12400 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12900 19193 12909 19227
rect 12909 19193 12943 19227
rect 12943 19193 12952 19227
rect 12900 19184 12952 19193
rect 12440 19116 12492 19125
rect 14464 19116 14516 19168
rect 15016 19116 15068 19168
rect 15292 19116 15344 19168
rect 18788 19184 18840 19236
rect 16304 19159 16356 19168
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 16304 19116 16356 19125
rect 16672 19159 16724 19168
rect 16672 19125 16681 19159
rect 16681 19125 16715 19159
rect 16715 19125 16724 19159
rect 16672 19116 16724 19125
rect 17684 19116 17736 19168
rect 17868 19116 17920 19168
rect 20168 19227 20220 19236
rect 20168 19193 20177 19227
rect 20177 19193 20211 19227
rect 20211 19193 20220 19227
rect 20168 19184 20220 19193
rect 19156 19116 19208 19168
rect 21732 19252 21784 19304
rect 21272 19116 21324 19168
rect 21640 19116 21692 19168
rect 8379 19014 8431 19066
rect 8443 19014 8495 19066
rect 8507 19014 8559 19066
rect 8571 19014 8623 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 15904 19014 15956 19066
rect 15968 19014 16020 19066
rect 2228 18844 2280 18896
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 2412 18776 2464 18828
rect 3700 18776 3752 18828
rect 4712 18912 4764 18964
rect 6644 18912 6696 18964
rect 7932 18912 7984 18964
rect 5724 18844 5776 18896
rect 5264 18776 5316 18828
rect 5448 18819 5500 18828
rect 5448 18785 5457 18819
rect 5457 18785 5491 18819
rect 5491 18785 5500 18819
rect 5448 18776 5500 18785
rect 7380 18844 7432 18896
rect 8852 18912 8904 18964
rect 9864 18912 9916 18964
rect 10692 18912 10744 18964
rect 8208 18887 8260 18896
rect 8208 18853 8242 18887
rect 8242 18853 8260 18887
rect 8208 18844 8260 18853
rect 8300 18844 8352 18896
rect 17868 18912 17920 18964
rect 18788 18955 18840 18964
rect 18788 18921 18797 18955
rect 18797 18921 18831 18955
rect 18831 18921 18840 18955
rect 18788 18912 18840 18921
rect 11980 18844 12032 18896
rect 4988 18708 5040 18760
rect 2228 18640 2280 18692
rect 1768 18572 1820 18624
rect 4344 18640 4396 18692
rect 9496 18776 9548 18828
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10784 18776 10836 18828
rect 11612 18776 11664 18828
rect 12532 18776 12584 18828
rect 7564 18708 7616 18760
rect 10232 18751 10284 18760
rect 5080 18615 5132 18624
rect 5080 18581 5089 18615
rect 5089 18581 5123 18615
rect 5123 18581 5132 18615
rect 5080 18572 5132 18581
rect 6460 18615 6512 18624
rect 6460 18581 6469 18615
rect 6469 18581 6503 18615
rect 6503 18581 6512 18615
rect 6460 18572 6512 18581
rect 6736 18572 6788 18624
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 8208 18572 8260 18624
rect 8668 18572 8720 18624
rect 9588 18572 9640 18624
rect 10140 18572 10192 18624
rect 13268 18776 13320 18828
rect 14188 18776 14240 18828
rect 15384 18819 15436 18828
rect 15384 18785 15393 18819
rect 15393 18785 15427 18819
rect 15427 18785 15436 18819
rect 15384 18776 15436 18785
rect 16488 18776 16540 18828
rect 17500 18776 17552 18828
rect 14832 18708 14884 18760
rect 19524 18776 19576 18828
rect 21640 18844 21692 18896
rect 19340 18708 19392 18760
rect 19892 18708 19944 18760
rect 18696 18640 18748 18692
rect 22744 18776 22796 18828
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 13544 18615 13596 18624
rect 13544 18581 13553 18615
rect 13553 18581 13587 18615
rect 13587 18581 13596 18615
rect 13544 18572 13596 18581
rect 14740 18572 14792 18624
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 18604 18572 18656 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 22652 18615 22704 18624
rect 22652 18581 22661 18615
rect 22661 18581 22695 18615
rect 22695 18581 22704 18615
rect 22652 18572 22704 18581
rect 4680 18470 4732 18522
rect 4744 18470 4796 18522
rect 4808 18470 4860 18522
rect 4872 18470 4924 18522
rect 12078 18470 12130 18522
rect 12142 18470 12194 18522
rect 12206 18470 12258 18522
rect 12270 18470 12322 18522
rect 19475 18470 19527 18522
rect 19539 18470 19591 18522
rect 19603 18470 19655 18522
rect 19667 18470 19719 18522
rect 4988 18368 5040 18420
rect 8944 18368 8996 18420
rect 9588 18368 9640 18420
rect 11612 18411 11664 18420
rect 11612 18377 11621 18411
rect 11621 18377 11655 18411
rect 11655 18377 11664 18411
rect 11612 18368 11664 18377
rect 12440 18368 12492 18420
rect 14464 18368 14516 18420
rect 19248 18368 19300 18420
rect 19340 18368 19392 18420
rect 4068 18300 4120 18352
rect 4344 18300 4396 18352
rect 2320 18275 2372 18284
rect 2320 18241 2329 18275
rect 2329 18241 2363 18275
rect 2363 18241 2372 18275
rect 2320 18232 2372 18241
rect 8300 18300 8352 18352
rect 9312 18300 9364 18352
rect 12992 18300 13044 18352
rect 14740 18300 14792 18352
rect 17960 18300 18012 18352
rect 12900 18232 12952 18284
rect 14832 18232 14884 18284
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 17500 18232 17552 18284
rect 18052 18275 18104 18284
rect 18052 18241 18061 18275
rect 18061 18241 18095 18275
rect 18095 18241 18104 18275
rect 18052 18232 18104 18241
rect 19156 18232 19208 18284
rect 19432 18232 19484 18284
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 2412 18164 2464 18216
rect 3608 18096 3660 18148
rect 4160 18164 4212 18216
rect 8300 18207 8352 18216
rect 8300 18173 8309 18207
rect 8309 18173 8343 18207
rect 8343 18173 8352 18207
rect 8300 18164 8352 18173
rect 9864 18164 9916 18216
rect 4804 18096 4856 18148
rect 10324 18164 10376 18216
rect 11704 18164 11756 18216
rect 13084 18164 13136 18216
rect 15936 18164 15988 18216
rect 17684 18164 17736 18216
rect 22008 18368 22060 18420
rect 22100 18300 22152 18352
rect 20812 18232 20864 18284
rect 22560 18232 22612 18284
rect 20076 18207 20128 18216
rect 3700 18071 3752 18080
rect 3700 18037 3709 18071
rect 3709 18037 3743 18071
rect 3743 18037 3752 18071
rect 3700 18028 3752 18037
rect 5816 18028 5868 18080
rect 6000 18071 6052 18080
rect 6000 18037 6009 18071
rect 6009 18037 6043 18071
rect 6043 18037 6052 18071
rect 6000 18028 6052 18037
rect 7012 18028 7064 18080
rect 9588 18028 9640 18080
rect 10968 18096 11020 18148
rect 14280 18096 14332 18148
rect 15752 18096 15804 18148
rect 16304 18096 16356 18148
rect 11612 18028 11664 18080
rect 14372 18028 14424 18080
rect 14464 18028 14516 18080
rect 15108 18071 15160 18080
rect 15108 18037 15117 18071
rect 15117 18037 15151 18071
rect 15151 18037 15160 18071
rect 15108 18028 15160 18037
rect 15384 18028 15436 18080
rect 16396 18028 16448 18080
rect 16764 18096 16816 18148
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20536 18164 20588 18216
rect 18788 18096 18840 18148
rect 17132 18071 17184 18080
rect 17132 18037 17141 18071
rect 17141 18037 17175 18071
rect 17175 18037 17184 18071
rect 17132 18028 17184 18037
rect 18052 18028 18104 18080
rect 20996 18071 21048 18080
rect 20996 18037 21005 18071
rect 21005 18037 21039 18071
rect 21039 18037 21048 18071
rect 20996 18028 21048 18037
rect 21732 18028 21784 18080
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 8379 17926 8431 17978
rect 8443 17926 8495 17978
rect 8507 17926 8559 17978
rect 8571 17926 8623 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 15904 17926 15956 17978
rect 15968 17926 16020 17978
rect 2320 17824 2372 17876
rect 3608 17867 3660 17876
rect 3608 17833 3617 17867
rect 3617 17833 3651 17867
rect 3651 17833 3660 17867
rect 3608 17824 3660 17833
rect 5448 17824 5500 17876
rect 6920 17824 6972 17876
rect 9496 17824 9548 17876
rect 9956 17824 10008 17876
rect 11428 17824 11480 17876
rect 11704 17867 11756 17876
rect 11704 17833 11713 17867
rect 11713 17833 11747 17867
rect 11747 17833 11756 17867
rect 11704 17824 11756 17833
rect 11888 17824 11940 17876
rect 13636 17824 13688 17876
rect 14280 17867 14332 17876
rect 14280 17833 14289 17867
rect 14289 17833 14323 17867
rect 14323 17833 14332 17867
rect 14280 17824 14332 17833
rect 14648 17824 14700 17876
rect 15660 17824 15712 17876
rect 16856 17824 16908 17876
rect 18052 17824 18104 17876
rect 18788 17867 18840 17876
rect 18788 17833 18797 17867
rect 18797 17833 18831 17867
rect 18831 17833 18840 17867
rect 18788 17824 18840 17833
rect 20996 17824 21048 17876
rect 1676 17731 1728 17740
rect 1676 17697 1685 17731
rect 1685 17697 1719 17731
rect 1719 17697 1728 17731
rect 1676 17688 1728 17697
rect 2136 17688 2188 17740
rect 10416 17756 10468 17808
rect 12348 17756 12400 17808
rect 13084 17756 13136 17808
rect 2320 17688 2372 17740
rect 4252 17731 4304 17740
rect 4252 17697 4261 17731
rect 4261 17697 4295 17731
rect 4295 17697 4304 17731
rect 4252 17688 4304 17697
rect 5080 17731 5132 17740
rect 5080 17697 5114 17731
rect 5114 17697 5132 17731
rect 5080 17688 5132 17697
rect 6276 17688 6328 17740
rect 9312 17688 9364 17740
rect 9772 17688 9824 17740
rect 11796 17688 11848 17740
rect 12624 17688 12676 17740
rect 14004 17688 14056 17740
rect 14096 17688 14148 17740
rect 16120 17756 16172 17808
rect 17592 17756 17644 17808
rect 19340 17756 19392 17808
rect 22652 17756 22704 17808
rect 14556 17688 14608 17740
rect 4436 17620 4488 17672
rect 6368 17620 6420 17672
rect 4160 17552 4212 17604
rect 4528 17552 4580 17604
rect 8760 17552 8812 17604
rect 9220 17620 9272 17672
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 10324 17620 10376 17629
rect 10232 17552 10284 17604
rect 3700 17484 3752 17536
rect 6092 17484 6144 17536
rect 6276 17484 6328 17536
rect 7472 17484 7524 17536
rect 7932 17484 7984 17536
rect 11428 17484 11480 17536
rect 11704 17484 11756 17536
rect 18972 17688 19024 17740
rect 20076 17688 20128 17740
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 17408 17663 17460 17672
rect 17408 17629 17417 17663
rect 17417 17629 17451 17663
rect 17451 17629 17460 17663
rect 17408 17620 17460 17629
rect 19892 17620 19944 17672
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 20996 17620 21048 17672
rect 21272 17620 21324 17672
rect 16304 17552 16356 17604
rect 15568 17484 15620 17536
rect 19800 17552 19852 17604
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 20812 17484 20864 17536
rect 4680 17382 4732 17434
rect 4744 17382 4796 17434
rect 4808 17382 4860 17434
rect 4872 17382 4924 17434
rect 12078 17382 12130 17434
rect 12142 17382 12194 17434
rect 12206 17382 12258 17434
rect 12270 17382 12322 17434
rect 19475 17382 19527 17434
rect 19539 17382 19591 17434
rect 19603 17382 19655 17434
rect 19667 17382 19719 17434
rect 6092 17280 6144 17332
rect 3700 17212 3752 17264
rect 4528 17212 4580 17264
rect 4620 17212 4672 17264
rect 6368 17212 6420 17264
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 3608 17144 3660 17196
rect 2780 17076 2832 17128
rect 3700 17076 3752 17128
rect 4252 17076 4304 17128
rect 5540 17144 5592 17196
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 6736 17144 6788 17196
rect 11980 17280 12032 17332
rect 8300 17144 8352 17196
rect 3148 17008 3200 17060
rect 3976 17008 4028 17060
rect 4068 17008 4120 17060
rect 7840 17076 7892 17128
rect 7932 17076 7984 17128
rect 11888 17212 11940 17264
rect 12256 17212 12308 17264
rect 14004 17255 14056 17264
rect 14004 17221 14013 17255
rect 14013 17221 14047 17255
rect 14047 17221 14056 17255
rect 14004 17212 14056 17221
rect 15108 17212 15160 17264
rect 16580 17212 16632 17264
rect 17132 17212 17184 17264
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 17960 17212 18012 17264
rect 18880 17212 18932 17264
rect 19892 17144 19944 17196
rect 20996 17280 21048 17332
rect 21640 17323 21692 17332
rect 21640 17289 21649 17323
rect 21649 17289 21683 17323
rect 21683 17289 21692 17323
rect 21640 17280 21692 17289
rect 22744 17144 22796 17196
rect 23388 17144 23440 17196
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 11428 17076 11480 17128
rect 12072 17076 12124 17128
rect 13268 17076 13320 17128
rect 14372 17076 14424 17128
rect 14832 17076 14884 17128
rect 15108 17119 15160 17128
rect 15108 17085 15117 17119
rect 15117 17085 15151 17119
rect 15151 17085 15160 17119
rect 15108 17076 15160 17085
rect 7472 17008 7524 17060
rect 2320 16940 2372 16992
rect 4252 16983 4304 16992
rect 4252 16949 4261 16983
rect 4261 16949 4295 16983
rect 4295 16949 4304 16983
rect 4252 16940 4304 16949
rect 4988 16940 5040 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 7656 16940 7708 16992
rect 9036 17008 9088 17060
rect 9128 17008 9180 17060
rect 8668 16940 8720 16992
rect 9864 16940 9916 16992
rect 11060 17008 11112 17060
rect 11428 16940 11480 16992
rect 12992 17008 13044 17060
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 20168 17076 20220 17128
rect 20812 17076 20864 17128
rect 20904 17076 20956 17128
rect 15568 17008 15620 17060
rect 16764 17008 16816 17060
rect 19248 17008 19300 17060
rect 21364 17008 21416 17060
rect 22100 17008 22152 17060
rect 14096 16940 14148 16992
rect 16212 16940 16264 16992
rect 17132 16983 17184 16992
rect 17132 16949 17141 16983
rect 17141 16949 17175 16983
rect 17175 16949 17184 16983
rect 17132 16940 17184 16949
rect 18236 16983 18288 16992
rect 18236 16949 18245 16983
rect 18245 16949 18279 16983
rect 18279 16949 18288 16983
rect 18236 16940 18288 16949
rect 18512 16940 18564 16992
rect 19800 16940 19852 16992
rect 19984 16940 20036 16992
rect 22008 16940 22060 16992
rect 8379 16838 8431 16890
rect 8443 16838 8495 16890
rect 8507 16838 8559 16890
rect 8571 16838 8623 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 15904 16838 15956 16890
rect 15968 16838 16020 16890
rect 2780 16736 2832 16788
rect 3148 16736 3200 16788
rect 3608 16736 3660 16788
rect 4252 16736 4304 16788
rect 5264 16736 5316 16788
rect 2964 16668 3016 16720
rect 2044 16600 2096 16652
rect 3424 16600 3476 16652
rect 4068 16600 4120 16652
rect 9128 16736 9180 16788
rect 9404 16736 9456 16788
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 11428 16736 11480 16788
rect 6000 16668 6052 16720
rect 7748 16668 7800 16720
rect 7932 16668 7984 16720
rect 8852 16668 8904 16720
rect 10048 16668 10100 16720
rect 10324 16668 10376 16720
rect 10600 16668 10652 16720
rect 12072 16736 12124 16788
rect 13544 16736 13596 16788
rect 14096 16736 14148 16788
rect 16304 16736 16356 16788
rect 16488 16736 16540 16788
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4988 16600 5040 16652
rect 8668 16600 8720 16652
rect 9128 16600 9180 16652
rect 9404 16600 9456 16652
rect 4620 16532 4672 16541
rect 6276 16575 6328 16584
rect 4252 16464 4304 16516
rect 5172 16464 5224 16516
rect 3424 16396 3476 16448
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 10968 16600 11020 16652
rect 11980 16643 12032 16652
rect 11980 16609 12014 16643
rect 12014 16609 12032 16643
rect 11980 16600 12032 16609
rect 12256 16600 12308 16652
rect 14464 16600 14516 16652
rect 7380 16396 7432 16448
rect 9404 16464 9456 16516
rect 13636 16532 13688 16584
rect 15016 16668 15068 16720
rect 17592 16736 17644 16788
rect 18972 16736 19024 16788
rect 19800 16736 19852 16788
rect 22192 16736 22244 16788
rect 14648 16643 14700 16652
rect 14648 16609 14657 16643
rect 14657 16609 14691 16643
rect 14691 16609 14700 16643
rect 15292 16643 15344 16652
rect 14648 16600 14700 16609
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 16580 16600 16632 16652
rect 17684 16668 17736 16720
rect 19892 16668 19944 16720
rect 19248 16600 19300 16652
rect 19432 16600 19484 16652
rect 13268 16464 13320 16516
rect 14740 16464 14792 16516
rect 17408 16532 17460 16584
rect 19340 16575 19392 16584
rect 19340 16541 19349 16575
rect 19349 16541 19383 16575
rect 19383 16541 19392 16575
rect 21640 16668 21692 16720
rect 19340 16532 19392 16541
rect 20444 16532 20496 16584
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 9680 16396 9732 16448
rect 9864 16396 9916 16448
rect 17500 16396 17552 16448
rect 18052 16396 18104 16448
rect 18420 16396 18472 16448
rect 18788 16396 18840 16448
rect 19892 16396 19944 16448
rect 21548 16396 21600 16448
rect 4680 16294 4732 16346
rect 4744 16294 4796 16346
rect 4808 16294 4860 16346
rect 4872 16294 4924 16346
rect 12078 16294 12130 16346
rect 12142 16294 12194 16346
rect 12206 16294 12258 16346
rect 12270 16294 12322 16346
rect 19475 16294 19527 16346
rect 19539 16294 19591 16346
rect 19603 16294 19655 16346
rect 19667 16294 19719 16346
rect 2780 16192 2832 16244
rect 3424 16235 3476 16244
rect 3424 16201 3433 16235
rect 3433 16201 3467 16235
rect 3467 16201 3476 16235
rect 3424 16192 3476 16201
rect 5632 16124 5684 16176
rect 4528 16099 4580 16108
rect 4528 16065 4540 16099
rect 4540 16065 4574 16099
rect 4574 16065 4580 16099
rect 4528 16056 4580 16065
rect 6092 16056 6144 16108
rect 2688 15920 2740 15972
rect 3700 15920 3752 15972
rect 5724 15988 5776 16040
rect 6368 16056 6420 16108
rect 10324 16124 10376 16176
rect 12624 16235 12676 16244
rect 12624 16201 12633 16235
rect 12633 16201 12667 16235
rect 12667 16201 12676 16235
rect 12624 16192 12676 16201
rect 17132 16192 17184 16244
rect 22560 16192 22612 16244
rect 7196 16056 7248 16108
rect 7656 16056 7708 16108
rect 6736 15988 6788 16040
rect 1860 15852 1912 15904
rect 3608 15852 3660 15904
rect 4344 15852 4396 15904
rect 4896 15852 4948 15904
rect 5172 15852 5224 15904
rect 6276 15852 6328 15904
rect 7196 15852 7248 15904
rect 7932 15852 7984 15904
rect 11060 16056 11112 16108
rect 13268 16124 13320 16176
rect 19708 16124 19760 16176
rect 8852 15988 8904 16040
rect 10692 15988 10744 16040
rect 13636 16056 13688 16108
rect 13820 16099 13872 16108
rect 13820 16065 13832 16099
rect 13832 16065 13866 16099
rect 13866 16065 13872 16099
rect 13820 16056 13872 16065
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 14280 16056 14332 16108
rect 14096 16031 14148 16040
rect 14096 15997 14105 16031
rect 14105 15997 14139 16031
rect 14139 15997 14148 16031
rect 14096 15988 14148 15997
rect 15292 15988 15344 16040
rect 20904 16056 20956 16108
rect 16764 15988 16816 16040
rect 8668 15895 8720 15904
rect 8668 15861 8677 15895
rect 8677 15861 8711 15895
rect 8711 15861 8720 15895
rect 8668 15852 8720 15861
rect 8852 15852 8904 15904
rect 10416 15852 10468 15904
rect 12072 15920 12124 15972
rect 11244 15852 11296 15904
rect 11428 15895 11480 15904
rect 11428 15861 11437 15895
rect 11437 15861 11471 15895
rect 11471 15861 11480 15895
rect 11428 15852 11480 15861
rect 11704 15852 11756 15904
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 13176 15852 13228 15904
rect 16488 15920 16540 15972
rect 17868 15988 17920 16040
rect 20812 15988 20864 16040
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 16764 15852 16816 15904
rect 17500 15852 17552 15904
rect 19340 15920 19392 15972
rect 19248 15852 19300 15904
rect 20996 15852 21048 15904
rect 21548 15920 21600 15972
rect 22560 15852 22612 15904
rect 8379 15750 8431 15802
rect 8443 15750 8495 15802
rect 8507 15750 8559 15802
rect 8571 15750 8623 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 15904 15750 15956 15802
rect 15968 15750 16020 15802
rect 3608 15648 3660 15700
rect 4528 15648 4580 15700
rect 8852 15648 8904 15700
rect 1860 15580 1912 15632
rect 3700 15580 3752 15632
rect 2964 15512 3016 15564
rect 4252 15512 4304 15564
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 4252 15376 4304 15428
rect 4712 15580 4764 15632
rect 9128 15648 9180 15700
rect 10692 15648 10744 15700
rect 2688 15308 2740 15360
rect 4896 15512 4948 15564
rect 6000 15512 6052 15564
rect 6368 15512 6420 15564
rect 6828 15512 6880 15564
rect 4712 15444 4764 15496
rect 5632 15444 5684 15496
rect 6092 15444 6144 15496
rect 7380 15555 7432 15564
rect 7380 15521 7414 15555
rect 7414 15521 7432 15555
rect 7380 15512 7432 15521
rect 7932 15512 7984 15564
rect 10876 15580 10928 15632
rect 12532 15648 12584 15700
rect 14096 15648 14148 15700
rect 14372 15648 14424 15700
rect 9864 15512 9916 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 10968 15555 11020 15564
rect 6736 15308 6788 15360
rect 9128 15444 9180 15496
rect 10416 15444 10468 15496
rect 10968 15521 10977 15555
rect 10977 15521 11011 15555
rect 11011 15521 11020 15555
rect 10968 15512 11020 15521
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 11612 15512 11664 15564
rect 12072 15512 12124 15564
rect 12256 15444 12308 15496
rect 13268 15512 13320 15564
rect 15016 15555 15068 15564
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 10600 15308 10652 15360
rect 12716 15308 12768 15360
rect 13084 15444 13136 15496
rect 13452 15308 13504 15360
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 19156 15648 19208 15700
rect 19340 15691 19392 15700
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 20352 15648 20404 15700
rect 15660 15512 15712 15564
rect 19708 15580 19760 15632
rect 15752 15487 15804 15496
rect 15752 15453 15764 15487
rect 15764 15453 15798 15487
rect 15798 15453 15804 15487
rect 15752 15444 15804 15453
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 17868 15512 17920 15564
rect 18052 15512 18104 15564
rect 18696 15512 18748 15564
rect 20996 15512 21048 15564
rect 16856 15376 16908 15428
rect 16764 15308 16816 15360
rect 17132 15351 17184 15360
rect 17132 15317 17141 15351
rect 17141 15317 17175 15351
rect 17175 15317 17184 15351
rect 17132 15308 17184 15317
rect 20812 15444 20864 15496
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 19800 15308 19852 15360
rect 20812 15308 20864 15360
rect 4680 15206 4732 15258
rect 4744 15206 4796 15258
rect 4808 15206 4860 15258
rect 4872 15206 4924 15258
rect 12078 15206 12130 15258
rect 12142 15206 12194 15258
rect 12206 15206 12258 15258
rect 12270 15206 12322 15258
rect 19475 15206 19527 15258
rect 19539 15206 19591 15258
rect 19603 15206 19655 15258
rect 19667 15206 19719 15258
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 8852 15104 8904 15156
rect 8944 15104 8996 15156
rect 4988 14968 5040 15020
rect 11980 15104 12032 15156
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 15016 15147 15068 15156
rect 12440 15104 12492 15113
rect 15016 15113 15025 15147
rect 15025 15113 15059 15147
rect 15059 15113 15068 15147
rect 15016 15104 15068 15113
rect 15292 15104 15344 15156
rect 15476 15104 15528 15156
rect 12624 15036 12676 15088
rect 4252 14900 4304 14952
rect 4436 14900 4488 14952
rect 5172 14900 5224 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 8484 14900 8536 14952
rect 10600 14900 10652 14952
rect 12256 14968 12308 15020
rect 14464 15036 14516 15088
rect 10968 14943 11020 14952
rect 10968 14909 10991 14943
rect 10991 14909 11020 14943
rect 10968 14900 11020 14909
rect 12348 14900 12400 14952
rect 13084 14900 13136 14952
rect 14740 14968 14792 15020
rect 17408 15011 17460 15020
rect 17408 14977 17417 15011
rect 17417 14977 17451 15011
rect 17451 14977 17460 15011
rect 17408 14968 17460 14977
rect 20996 15104 21048 15156
rect 21180 15147 21232 15156
rect 21180 15113 21189 15147
rect 21189 15113 21223 15147
rect 21223 15113 21232 15147
rect 21180 15104 21232 15113
rect 17684 15036 17736 15088
rect 18328 15036 18380 15088
rect 14556 14900 14608 14952
rect 16212 14900 16264 14952
rect 19984 14968 20036 15020
rect 20444 14968 20496 15020
rect 21916 14968 21968 15020
rect 18144 14900 18196 14952
rect 18788 14900 18840 14952
rect 19156 14900 19208 14952
rect 19432 14900 19484 14952
rect 19708 14900 19760 14952
rect 20996 14900 21048 14952
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 3056 14832 3108 14884
rect 5816 14832 5868 14884
rect 6368 14832 6420 14884
rect 7288 14832 7340 14884
rect 9680 14832 9732 14884
rect 1400 14807 1452 14816
rect 1400 14773 1409 14807
rect 1409 14773 1443 14807
rect 1443 14773 1452 14807
rect 1400 14764 1452 14773
rect 2964 14764 3016 14816
rect 3700 14764 3752 14816
rect 4620 14807 4672 14816
rect 4620 14773 4635 14807
rect 4635 14773 4669 14807
rect 4669 14773 4672 14807
rect 6000 14807 6052 14816
rect 4620 14764 4672 14773
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 6092 14764 6144 14816
rect 8024 14764 8076 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 10232 14764 10284 14816
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 11520 14764 11572 14816
rect 12164 14764 12216 14816
rect 16304 14875 16356 14884
rect 16304 14841 16313 14875
rect 16313 14841 16347 14875
rect 16347 14841 16356 14875
rect 16304 14832 16356 14841
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 14832 14807 14884 14816
rect 12808 14764 12860 14773
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 15476 14764 15528 14816
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 18696 14832 18748 14884
rect 18880 14875 18932 14884
rect 18880 14841 18889 14875
rect 18889 14841 18923 14875
rect 18923 14841 18932 14875
rect 18880 14832 18932 14841
rect 17684 14764 17736 14816
rect 21548 14832 21600 14884
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 21640 14764 21692 14816
rect 22008 14764 22060 14816
rect 8379 14662 8431 14714
rect 8443 14662 8495 14714
rect 8507 14662 8559 14714
rect 8571 14662 8623 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 15904 14662 15956 14714
rect 15968 14662 16020 14714
rect 1400 14560 1452 14612
rect 2872 14492 2924 14544
rect 8852 14560 8904 14612
rect 9128 14560 9180 14612
rect 1768 14424 1820 14476
rect 3424 14467 3476 14476
rect 3424 14433 3433 14467
rect 3433 14433 3467 14467
rect 3467 14433 3476 14467
rect 3424 14424 3476 14433
rect 3056 14331 3108 14340
rect 3056 14297 3065 14331
rect 3065 14297 3099 14331
rect 3099 14297 3108 14331
rect 3056 14288 3108 14297
rect 4344 14288 4396 14340
rect 8576 14492 8628 14544
rect 10324 14560 10376 14612
rect 10876 14560 10928 14612
rect 12440 14560 12492 14612
rect 12716 14560 12768 14612
rect 10232 14492 10284 14544
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 4068 14263 4120 14272
rect 4068 14229 4077 14263
rect 4077 14229 4111 14263
rect 4111 14229 4120 14263
rect 4068 14220 4120 14229
rect 4252 14220 4304 14272
rect 4988 14220 5040 14272
rect 8208 14424 8260 14476
rect 9128 14424 9180 14476
rect 9956 14424 10008 14476
rect 12532 14424 12584 14476
rect 13636 14424 13688 14476
rect 13912 14424 13964 14476
rect 19340 14560 19392 14612
rect 15200 14492 15252 14544
rect 17776 14492 17828 14544
rect 8852 14399 8904 14408
rect 6368 14288 6420 14340
rect 8852 14365 8861 14399
rect 8861 14365 8895 14399
rect 8895 14365 8904 14399
rect 8852 14356 8904 14365
rect 6828 14220 6880 14272
rect 8024 14263 8076 14272
rect 8024 14229 8033 14263
rect 8033 14229 8067 14263
rect 8067 14229 8076 14263
rect 8024 14220 8076 14229
rect 8576 14220 8628 14272
rect 8852 14220 8904 14272
rect 10968 14288 11020 14340
rect 14464 14399 14516 14408
rect 14464 14365 14473 14399
rect 14473 14365 14507 14399
rect 14507 14365 14516 14399
rect 15752 14467 15804 14476
rect 15752 14433 15761 14467
rect 15761 14433 15795 14467
rect 15795 14433 15804 14467
rect 16488 14467 16540 14476
rect 15752 14424 15804 14433
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 18052 14467 18104 14476
rect 18052 14433 18086 14467
rect 18086 14433 18104 14467
rect 18328 14492 18380 14544
rect 22008 14560 22060 14612
rect 18052 14424 18104 14433
rect 14464 14356 14516 14365
rect 12440 14288 12492 14340
rect 16580 14356 16632 14408
rect 16856 14356 16908 14408
rect 17684 14356 17736 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 19156 14356 19208 14408
rect 20812 14492 20864 14544
rect 10600 14220 10652 14272
rect 11520 14220 11572 14272
rect 17408 14288 17460 14340
rect 19248 14288 19300 14340
rect 20444 14356 20496 14408
rect 20996 14424 21048 14476
rect 21272 14424 21324 14476
rect 20720 14356 20772 14408
rect 20904 14356 20956 14408
rect 13452 14220 13504 14272
rect 13912 14263 13964 14272
rect 13912 14229 13921 14263
rect 13921 14229 13955 14263
rect 13955 14229 13964 14263
rect 13912 14220 13964 14229
rect 14740 14220 14792 14272
rect 15108 14220 15160 14272
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 18420 14220 18472 14272
rect 19340 14220 19392 14272
rect 20904 14220 20956 14272
rect 21916 14220 21968 14272
rect 4680 14118 4732 14170
rect 4744 14118 4796 14170
rect 4808 14118 4860 14170
rect 4872 14118 4924 14170
rect 12078 14118 12130 14170
rect 12142 14118 12194 14170
rect 12206 14118 12258 14170
rect 12270 14118 12322 14170
rect 19475 14118 19527 14170
rect 19539 14118 19591 14170
rect 19603 14118 19655 14170
rect 19667 14118 19719 14170
rect 1768 14016 1820 14068
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 3424 14016 3476 14068
rect 4252 14016 4304 14068
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 9864 14016 9916 14068
rect 10048 14016 10100 14068
rect 11428 14016 11480 14068
rect 12440 14016 12492 14068
rect 6644 13948 6696 14000
rect 6920 13948 6972 14000
rect 9680 13991 9732 14000
rect 9680 13957 9689 13991
rect 9689 13957 9723 13991
rect 9723 13957 9732 13991
rect 14464 14016 14516 14068
rect 16120 14016 16172 14068
rect 19156 14016 19208 14068
rect 21272 14016 21324 14068
rect 9680 13948 9732 13957
rect 15568 13948 15620 14000
rect 16028 13948 16080 14000
rect 4620 13880 4672 13932
rect 4896 13923 4948 13932
rect 4896 13889 4905 13923
rect 4905 13889 4939 13923
rect 4939 13889 4948 13923
rect 4896 13880 4948 13889
rect 6368 13880 6420 13932
rect 6092 13812 6144 13864
rect 10416 13880 10468 13932
rect 9956 13855 10008 13864
rect 4068 13744 4120 13796
rect 4252 13787 4304 13796
rect 4252 13753 4261 13787
rect 4261 13753 4295 13787
rect 4295 13753 4304 13787
rect 4252 13744 4304 13753
rect 5908 13744 5960 13796
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 10140 13812 10192 13864
rect 10324 13812 10376 13864
rect 10692 13812 10744 13864
rect 11428 13880 11480 13932
rect 11888 13880 11940 13932
rect 12532 13880 12584 13932
rect 17868 13880 17920 13932
rect 11520 13812 11572 13864
rect 11612 13812 11664 13864
rect 12716 13812 12768 13864
rect 15108 13812 15160 13864
rect 3148 13719 3200 13728
rect 3148 13685 3157 13719
rect 3157 13685 3191 13719
rect 3191 13685 3200 13719
rect 3148 13676 3200 13685
rect 4436 13676 4488 13728
rect 4620 13719 4672 13728
rect 4620 13685 4629 13719
rect 4629 13685 4663 13719
rect 4663 13685 4672 13719
rect 4620 13676 4672 13685
rect 6828 13676 6880 13728
rect 9772 13744 9824 13796
rect 10600 13744 10652 13796
rect 11888 13787 11940 13796
rect 7840 13719 7892 13728
rect 7840 13685 7849 13719
rect 7849 13685 7883 13719
rect 7883 13685 7892 13719
rect 7840 13676 7892 13685
rect 8208 13676 8260 13728
rect 10048 13676 10100 13728
rect 11060 13719 11112 13728
rect 11060 13685 11069 13719
rect 11069 13685 11103 13719
rect 11103 13685 11112 13719
rect 11060 13676 11112 13685
rect 11888 13753 11897 13787
rect 11897 13753 11931 13787
rect 11931 13753 11940 13787
rect 11888 13744 11940 13753
rect 19984 13880 20036 13932
rect 22836 13880 22888 13932
rect 18696 13812 18748 13864
rect 19156 13812 19208 13864
rect 19800 13812 19852 13864
rect 12164 13676 12216 13728
rect 12983 13676 13035 13728
rect 17868 13744 17920 13796
rect 18328 13787 18380 13796
rect 13820 13676 13872 13728
rect 16764 13676 16816 13728
rect 18328 13753 18340 13787
rect 18340 13753 18380 13787
rect 21456 13812 21508 13864
rect 18328 13744 18380 13753
rect 21640 13744 21692 13796
rect 18052 13676 18104 13728
rect 18972 13676 19024 13728
rect 19708 13676 19760 13728
rect 19984 13676 20036 13728
rect 20536 13676 20588 13728
rect 22192 13719 22244 13728
rect 22192 13685 22201 13719
rect 22201 13685 22235 13719
rect 22235 13685 22244 13719
rect 22192 13676 22244 13685
rect 8379 13574 8431 13626
rect 8443 13574 8495 13626
rect 8507 13574 8559 13626
rect 8571 13574 8623 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 15904 13574 15956 13626
rect 15968 13574 16020 13626
rect 1860 13515 1912 13524
rect 1860 13481 1869 13515
rect 1869 13481 1903 13515
rect 1903 13481 1912 13515
rect 1860 13472 1912 13481
rect 3148 13472 3200 13524
rect 4160 13472 4212 13524
rect 5908 13515 5960 13524
rect 5908 13481 5917 13515
rect 5917 13481 5951 13515
rect 5951 13481 5960 13515
rect 5908 13472 5960 13481
rect 10416 13472 10468 13524
rect 4620 13404 4672 13456
rect 5540 13404 5592 13456
rect 6092 13404 6144 13456
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 6644 13404 6696 13456
rect 6900 13404 6952 13456
rect 7564 13404 7616 13456
rect 8024 13404 8076 13456
rect 8116 13404 8168 13456
rect 8576 13404 8628 13456
rect 2688 13268 2740 13320
rect 3976 13268 4028 13320
rect 4528 13311 4580 13320
rect 4528 13277 4537 13311
rect 4537 13277 4571 13311
rect 4571 13277 4580 13311
rect 4528 13268 4580 13277
rect 3240 13200 3292 13252
rect 3516 13200 3568 13252
rect 7932 13336 7984 13388
rect 11060 13404 11112 13456
rect 11888 13472 11940 13524
rect 10048 13379 10100 13388
rect 8024 13268 8076 13320
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 11796 13336 11848 13388
rect 9496 13200 9548 13252
rect 9956 13200 10008 13252
rect 7932 13132 7984 13184
rect 8116 13175 8168 13184
rect 8116 13141 8125 13175
rect 8125 13141 8159 13175
rect 8159 13141 8168 13175
rect 8116 13132 8168 13141
rect 8944 13132 8996 13184
rect 10416 13268 10468 13320
rect 11428 13132 11480 13184
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 12716 13404 12768 13456
rect 13084 13404 13136 13456
rect 13820 13404 13872 13456
rect 14924 13404 14976 13456
rect 16580 13472 16632 13524
rect 17408 13472 17460 13524
rect 19984 13472 20036 13524
rect 20352 13472 20404 13524
rect 22192 13472 22244 13524
rect 15108 13336 15160 13388
rect 16856 13336 16908 13388
rect 17776 13336 17828 13388
rect 18972 13336 19024 13388
rect 17776 13200 17828 13252
rect 15016 13175 15068 13184
rect 15016 13141 15025 13175
rect 15025 13141 15059 13175
rect 15059 13141 15068 13175
rect 15016 13132 15068 13141
rect 15568 13132 15620 13184
rect 16764 13132 16816 13184
rect 18880 13132 18932 13184
rect 21916 13404 21968 13456
rect 19800 13336 19852 13388
rect 20352 13336 20404 13388
rect 19708 13268 19760 13320
rect 20904 13268 20956 13320
rect 22836 13132 22888 13184
rect 4680 13030 4732 13082
rect 4744 13030 4796 13082
rect 4808 13030 4860 13082
rect 4872 13030 4924 13082
rect 12078 13030 12130 13082
rect 12142 13030 12194 13082
rect 12206 13030 12258 13082
rect 12270 13030 12322 13082
rect 19475 13030 19527 13082
rect 19539 13030 19591 13082
rect 19603 13030 19655 13082
rect 19667 13030 19719 13082
rect 1676 12903 1728 12912
rect 1676 12869 1685 12903
rect 1685 12869 1719 12903
rect 1719 12869 1728 12903
rect 1676 12860 1728 12869
rect 1584 12724 1636 12776
rect 9496 12971 9548 12980
rect 5540 12860 5592 12912
rect 8852 12860 8904 12912
rect 2688 12724 2740 12776
rect 5724 12792 5776 12844
rect 6368 12792 6420 12844
rect 7840 12792 7892 12844
rect 4896 12724 4948 12776
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 8116 12724 8168 12776
rect 8576 12792 8628 12844
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 10416 12835 10468 12844
rect 2872 12656 2924 12708
rect 9220 12724 9272 12776
rect 9496 12724 9548 12776
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 11612 12792 11664 12844
rect 13268 12928 13320 12980
rect 16856 12928 16908 12980
rect 13636 12860 13688 12912
rect 14464 12860 14516 12912
rect 14924 12792 14976 12844
rect 15108 12792 15160 12844
rect 17408 12835 17460 12844
rect 17408 12801 17417 12835
rect 17417 12801 17451 12835
rect 17451 12801 17460 12835
rect 17408 12792 17460 12801
rect 18972 12928 19024 12980
rect 20628 12928 20680 12980
rect 19708 12860 19760 12912
rect 22284 12860 22336 12912
rect 21640 12835 21692 12844
rect 10692 12767 10744 12776
rect 10692 12733 10726 12767
rect 10726 12733 10744 12767
rect 10692 12724 10744 12733
rect 12440 12724 12492 12776
rect 12716 12724 12768 12776
rect 13452 12724 13504 12776
rect 18052 12767 18104 12776
rect 10324 12656 10376 12708
rect 11244 12656 11296 12708
rect 11428 12656 11480 12708
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 18328 12724 18380 12776
rect 18696 12767 18748 12776
rect 18696 12733 18705 12767
rect 18705 12733 18739 12767
rect 18739 12733 18748 12767
rect 18696 12724 18748 12733
rect 21640 12801 21649 12835
rect 21649 12801 21683 12835
rect 21683 12801 21692 12835
rect 21640 12792 21692 12801
rect 22100 12792 22152 12844
rect 21732 12724 21784 12776
rect 21916 12724 21968 12776
rect 22376 12724 22428 12776
rect 15568 12656 15620 12708
rect 4068 12588 4120 12640
rect 8024 12588 8076 12640
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 8944 12588 8996 12597
rect 11060 12588 11112 12640
rect 13268 12588 13320 12640
rect 13636 12588 13688 12640
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 16764 12588 16816 12640
rect 17776 12656 17828 12708
rect 18972 12699 19024 12708
rect 18972 12665 19006 12699
rect 19006 12665 19024 12699
rect 18972 12656 19024 12665
rect 17224 12588 17276 12640
rect 18420 12631 18472 12640
rect 18420 12597 18429 12631
rect 18429 12597 18463 12631
rect 18463 12597 18472 12631
rect 18420 12588 18472 12597
rect 18880 12588 18932 12640
rect 20812 12656 20864 12708
rect 19708 12588 19760 12640
rect 21548 12631 21600 12640
rect 21548 12597 21557 12631
rect 21557 12597 21591 12631
rect 21591 12597 21600 12631
rect 21548 12588 21600 12597
rect 8379 12486 8431 12538
rect 8443 12486 8495 12538
rect 8507 12486 8559 12538
rect 8571 12486 8623 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 15904 12486 15956 12538
rect 15968 12486 16020 12538
rect 3608 12427 3660 12436
rect 3608 12393 3617 12427
rect 3617 12393 3651 12427
rect 3651 12393 3660 12427
rect 3608 12384 3660 12393
rect 4896 12384 4948 12436
rect 5264 12384 5316 12436
rect 5448 12384 5500 12436
rect 8852 12384 8904 12436
rect 9956 12384 10008 12436
rect 10968 12384 11020 12436
rect 2780 12316 2832 12368
rect 7196 12316 7248 12368
rect 7564 12316 7616 12368
rect 7932 12316 7984 12368
rect 8208 12316 8260 12368
rect 12808 12384 12860 12436
rect 12624 12316 12676 12368
rect 13176 12359 13228 12368
rect 13176 12325 13185 12359
rect 13185 12325 13219 12359
rect 13219 12325 13228 12359
rect 13176 12316 13228 12325
rect 15200 12384 15252 12436
rect 15384 12316 15436 12368
rect 15568 12316 15620 12368
rect 18328 12384 18380 12436
rect 19248 12384 19300 12436
rect 19984 12384 20036 12436
rect 17408 12316 17460 12368
rect 1584 12291 1636 12300
rect 1584 12257 1593 12291
rect 1593 12257 1627 12291
rect 1627 12257 1636 12291
rect 1584 12248 1636 12257
rect 4344 12248 4396 12300
rect 3056 12180 3108 12232
rect 4620 12180 4672 12232
rect 5724 12180 5776 12232
rect 2688 12112 2740 12164
rect 3976 12112 4028 12164
rect 4896 12112 4948 12164
rect 3240 12044 3292 12096
rect 4436 12044 4488 12096
rect 5264 12044 5316 12096
rect 6552 12248 6604 12300
rect 6828 12248 6880 12300
rect 7288 12291 7340 12300
rect 7288 12257 7322 12291
rect 7322 12257 7340 12291
rect 7288 12248 7340 12257
rect 8024 12248 8076 12300
rect 8852 12291 8904 12300
rect 8852 12257 8861 12291
rect 8861 12257 8895 12291
rect 8895 12257 8904 12291
rect 8852 12248 8904 12257
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 10324 12180 10376 12232
rect 10968 12248 11020 12300
rect 13084 12248 13136 12300
rect 13360 12248 13412 12300
rect 14096 12248 14148 12300
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 15752 12248 15804 12300
rect 17868 12316 17920 12368
rect 18420 12316 18472 12368
rect 18696 12248 18748 12300
rect 20720 12316 20772 12368
rect 20352 12248 20404 12300
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 20996 12248 21048 12300
rect 8852 12112 8904 12164
rect 9680 12112 9732 12164
rect 11888 12112 11940 12164
rect 6276 12044 6328 12096
rect 8024 12044 8076 12096
rect 8576 12044 8628 12096
rect 11336 12044 11388 12096
rect 12440 12044 12492 12096
rect 13084 12044 13136 12096
rect 15384 12180 15436 12232
rect 19800 12180 19852 12232
rect 20076 12223 20128 12232
rect 20076 12189 20085 12223
rect 20085 12189 20119 12223
rect 20119 12189 20128 12223
rect 20076 12180 20128 12189
rect 14280 12112 14332 12164
rect 16488 12112 16540 12164
rect 18512 12112 18564 12164
rect 19708 12112 19760 12164
rect 14464 12044 14516 12096
rect 15476 12044 15528 12096
rect 18144 12044 18196 12096
rect 18788 12044 18840 12096
rect 20628 12044 20680 12096
rect 22192 12044 22244 12096
rect 4680 11942 4732 11994
rect 4744 11942 4796 11994
rect 4808 11942 4860 11994
rect 4872 11942 4924 11994
rect 12078 11942 12130 11994
rect 12142 11942 12194 11994
rect 12206 11942 12258 11994
rect 12270 11942 12322 11994
rect 19475 11942 19527 11994
rect 19539 11942 19591 11994
rect 19603 11942 19655 11994
rect 19667 11942 19719 11994
rect 2780 11840 2832 11892
rect 4804 11772 4856 11824
rect 3976 11704 4028 11756
rect 4528 11704 4580 11756
rect 4896 11704 4948 11756
rect 5264 11840 5316 11892
rect 8576 11840 8628 11892
rect 8944 11840 8996 11892
rect 10048 11840 10100 11892
rect 10692 11840 10744 11892
rect 14556 11840 14608 11892
rect 15660 11840 15712 11892
rect 19340 11840 19392 11892
rect 20168 11840 20220 11892
rect 20720 11840 20772 11892
rect 21640 11840 21692 11892
rect 9956 11772 10008 11824
rect 10416 11772 10468 11824
rect 12532 11772 12584 11824
rect 15844 11772 15896 11824
rect 6828 11704 6880 11756
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 1492 11679 1544 11688
rect 1492 11645 1501 11679
rect 1501 11645 1535 11679
rect 1535 11645 1544 11679
rect 1492 11636 1544 11645
rect 4068 11636 4120 11688
rect 7748 11636 7800 11688
rect 11152 11636 11204 11688
rect 14188 11704 14240 11756
rect 14464 11704 14516 11756
rect 13084 11636 13136 11688
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 16028 11772 16080 11824
rect 16396 11704 16448 11756
rect 18880 11772 18932 11824
rect 19064 11772 19116 11824
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 17776 11704 17828 11756
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 15200 11636 15252 11688
rect 3056 11568 3108 11620
rect 3424 11568 3476 11620
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 4436 11500 4488 11552
rect 4804 11543 4856 11552
rect 4804 11509 4813 11543
rect 4813 11509 4847 11543
rect 4847 11509 4856 11543
rect 4804 11500 4856 11509
rect 6552 11568 6604 11620
rect 6920 11568 6972 11620
rect 7104 11568 7156 11620
rect 8024 11568 8076 11620
rect 11888 11568 11940 11620
rect 7564 11500 7616 11552
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 10048 11500 10100 11552
rect 11520 11500 11572 11552
rect 12256 11500 12308 11552
rect 14648 11568 14700 11620
rect 15016 11568 15068 11620
rect 13912 11500 13964 11552
rect 14280 11500 14332 11552
rect 14556 11500 14608 11552
rect 14924 11500 14976 11552
rect 17868 11636 17920 11688
rect 19156 11636 19208 11688
rect 19616 11704 19668 11756
rect 19800 11747 19852 11756
rect 19800 11713 19809 11747
rect 19809 11713 19843 11747
rect 19843 11713 19852 11747
rect 19800 11704 19852 11713
rect 18512 11568 18564 11620
rect 16212 11500 16264 11552
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 16764 11500 16816 11552
rect 17132 11500 17184 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 18696 11500 18748 11552
rect 20260 11500 20312 11552
rect 21272 11636 21324 11688
rect 22652 11568 22704 11620
rect 8379 11398 8431 11450
rect 8443 11398 8495 11450
rect 8507 11398 8559 11450
rect 8571 11398 8623 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 15904 11398 15956 11450
rect 15968 11398 16020 11450
rect 3056 11296 3108 11348
rect 3700 11296 3752 11348
rect 5264 11296 5316 11348
rect 5448 11296 5500 11348
rect 6276 11296 6328 11348
rect 8852 11296 8904 11348
rect 9680 11296 9732 11348
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 13544 11296 13596 11348
rect 15568 11296 15620 11348
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 4804 11228 4856 11280
rect 4436 11203 4488 11212
rect 3516 11092 3568 11144
rect 3332 10956 3384 11008
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 4896 11160 4948 11212
rect 5724 11160 5776 11212
rect 6368 11160 6420 11212
rect 7564 11203 7616 11212
rect 7564 11169 7598 11203
rect 7598 11169 7616 11203
rect 7564 11160 7616 11169
rect 9128 11228 9180 11280
rect 12440 11228 12492 11280
rect 12992 11228 13044 11280
rect 4712 11135 4764 11144
rect 4344 11024 4396 11076
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 4528 11024 4580 11076
rect 6552 11024 6604 11076
rect 8760 11092 8812 11144
rect 11796 11160 11848 11212
rect 12256 11203 12308 11212
rect 12256 11169 12265 11203
rect 12265 11169 12299 11203
rect 12299 11169 12308 11203
rect 12256 11160 12308 11169
rect 12900 11160 12952 11212
rect 13360 11160 13412 11212
rect 16304 11228 16356 11280
rect 16580 11228 16632 11280
rect 17040 11228 17092 11280
rect 15568 11160 15620 11212
rect 16488 11160 16540 11212
rect 17408 11296 17460 11348
rect 19800 11339 19852 11348
rect 19800 11305 19809 11339
rect 19809 11305 19843 11339
rect 19843 11305 19852 11339
rect 19800 11296 19852 11305
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 22192 11228 22244 11280
rect 10416 11092 10468 11144
rect 12716 11092 12768 11144
rect 7012 10956 7064 11008
rect 8024 10956 8076 11008
rect 9956 11024 10008 11076
rect 14648 11024 14700 11076
rect 15016 11024 15068 11076
rect 15200 11024 15252 11076
rect 9864 10956 9916 11008
rect 12808 10956 12860 11008
rect 13728 10956 13780 11008
rect 13912 10956 13964 11008
rect 16672 11092 16724 11144
rect 17868 11092 17920 11144
rect 18236 11092 18288 11144
rect 18420 11135 18472 11144
rect 18420 11101 18432 11135
rect 18432 11101 18466 11135
rect 18466 11101 18472 11135
rect 18696 11135 18748 11144
rect 18420 11092 18472 11101
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 21272 11203 21324 11212
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 15936 10956 15988 11008
rect 17040 10999 17092 11008
rect 17040 10965 17049 10999
rect 17049 10965 17083 10999
rect 17083 10965 17092 10999
rect 17040 10956 17092 10965
rect 17500 10999 17552 11008
rect 17500 10965 17509 10999
rect 17509 10965 17543 10999
rect 17543 10965 17552 10999
rect 17500 10956 17552 10965
rect 18236 10956 18288 11008
rect 18512 10956 18564 11008
rect 18604 10956 18656 11008
rect 19156 10956 19208 11008
rect 4680 10854 4732 10906
rect 4744 10854 4796 10906
rect 4808 10854 4860 10906
rect 4872 10854 4924 10906
rect 12078 10854 12130 10906
rect 12142 10854 12194 10906
rect 12206 10854 12258 10906
rect 12270 10854 12322 10906
rect 19475 10854 19527 10906
rect 19539 10854 19591 10906
rect 19603 10854 19655 10906
rect 19667 10854 19719 10906
rect 3516 10752 3568 10804
rect 4436 10752 4488 10804
rect 6368 10795 6420 10804
rect 6368 10761 6377 10795
rect 6377 10761 6411 10795
rect 6411 10761 6420 10795
rect 6368 10752 6420 10761
rect 1492 10616 1544 10668
rect 4896 10616 4948 10668
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 4528 10548 4580 10600
rect 6184 10548 6236 10600
rect 5540 10480 5592 10532
rect 3424 10412 3476 10464
rect 6184 10412 6236 10464
rect 7472 10752 7524 10804
rect 9680 10684 9732 10736
rect 9956 10659 10008 10668
rect 9956 10625 9965 10659
rect 9965 10625 9999 10659
rect 9999 10625 10008 10659
rect 9956 10616 10008 10625
rect 11520 10616 11572 10668
rect 8944 10548 8996 10600
rect 7380 10480 7432 10532
rect 8024 10480 8076 10532
rect 9680 10548 9732 10600
rect 10784 10548 10836 10600
rect 12440 10548 12492 10600
rect 17040 10752 17092 10804
rect 17408 10752 17460 10804
rect 20260 10752 20312 10804
rect 20996 10752 21048 10804
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 17040 10616 17092 10668
rect 17224 10616 17276 10668
rect 8208 10412 8260 10464
rect 8944 10412 8996 10464
rect 9312 10412 9364 10464
rect 9588 10412 9640 10464
rect 9956 10412 10008 10464
rect 12532 10480 12584 10532
rect 14188 10548 14240 10600
rect 12716 10480 12768 10532
rect 10784 10412 10836 10464
rect 10968 10412 11020 10464
rect 11888 10412 11940 10464
rect 14924 10548 14976 10600
rect 16212 10591 16264 10600
rect 16212 10557 16246 10591
rect 16246 10557 16264 10591
rect 16212 10548 16264 10557
rect 16488 10548 16540 10600
rect 18236 10684 18288 10736
rect 19064 10684 19116 10736
rect 19248 10684 19300 10736
rect 18052 10616 18104 10668
rect 17500 10548 17552 10600
rect 18328 10548 18380 10600
rect 18788 10548 18840 10600
rect 20076 10548 20128 10600
rect 20628 10548 20680 10600
rect 22008 10548 22060 10600
rect 15016 10480 15068 10532
rect 19340 10480 19392 10532
rect 21180 10523 21232 10532
rect 21180 10489 21189 10523
rect 21189 10489 21223 10523
rect 21223 10489 21232 10523
rect 21180 10480 21232 10489
rect 14648 10412 14700 10464
rect 17132 10412 17184 10464
rect 17224 10412 17276 10464
rect 18052 10412 18104 10464
rect 18328 10412 18380 10464
rect 19616 10412 19668 10464
rect 19892 10412 19944 10464
rect 20260 10412 20312 10464
rect 21548 10412 21600 10464
rect 8379 10310 8431 10362
rect 8443 10310 8495 10362
rect 8507 10310 8559 10362
rect 8571 10310 8623 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 15904 10310 15956 10362
rect 15968 10310 16020 10362
rect 2596 10208 2648 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 6920 10208 6972 10260
rect 4436 10183 4488 10192
rect 1492 10072 1544 10124
rect 2780 10072 2832 10124
rect 4436 10149 4470 10183
rect 4470 10149 4488 10183
rect 4436 10140 4488 10149
rect 6276 10140 6328 10192
rect 7012 10140 7064 10192
rect 8944 10208 8996 10260
rect 9680 10140 9732 10192
rect 10140 10140 10192 10192
rect 10416 10208 10468 10260
rect 13452 10208 13504 10260
rect 15292 10208 15344 10260
rect 16212 10208 16264 10260
rect 3056 10072 3108 10124
rect 3332 10072 3384 10124
rect 6552 10072 6604 10124
rect 6920 10072 6972 10124
rect 8208 10115 8260 10124
rect 8208 10081 8231 10115
rect 8231 10081 8260 10115
rect 8208 10072 8260 10081
rect 10416 10072 10468 10124
rect 13728 10140 13780 10192
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 14648 10140 14700 10192
rect 16396 10140 16448 10192
rect 16580 10140 16632 10192
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 19800 10140 19852 10192
rect 20812 10140 20864 10192
rect 12716 10047 12768 10056
rect 11888 9936 11940 9988
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 14464 10072 14516 10124
rect 16948 10072 17000 10124
rect 17776 10072 17828 10124
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 18788 10072 18840 10124
rect 19616 10072 19668 10124
rect 20444 10072 20496 10124
rect 20996 10072 21048 10124
rect 21456 10072 21508 10124
rect 14188 9936 14240 9988
rect 15292 9936 15344 9988
rect 3332 9868 3384 9920
rect 8852 9868 8904 9920
rect 9956 9868 10008 9920
rect 12440 9868 12492 9920
rect 12992 9868 13044 9920
rect 14924 9911 14976 9920
rect 14924 9877 14933 9911
rect 14933 9877 14967 9911
rect 14967 9877 14976 9911
rect 14924 9868 14976 9877
rect 15108 9868 15160 9920
rect 16212 9868 16264 9920
rect 17500 10004 17552 10056
rect 18052 10004 18104 10056
rect 19248 10004 19300 10056
rect 22652 10004 22704 10056
rect 17224 9911 17276 9920
rect 17224 9877 17233 9911
rect 17233 9877 17267 9911
rect 17267 9877 17276 9911
rect 17224 9868 17276 9877
rect 18236 9868 18288 9920
rect 20720 9936 20772 9988
rect 21272 9936 21324 9988
rect 19340 9868 19392 9920
rect 19892 9868 19944 9920
rect 4680 9766 4732 9818
rect 4744 9766 4796 9818
rect 4808 9766 4860 9818
rect 4872 9766 4924 9818
rect 12078 9766 12130 9818
rect 12142 9766 12194 9818
rect 12206 9766 12258 9818
rect 12270 9766 12322 9818
rect 19475 9766 19527 9818
rect 19539 9766 19591 9818
rect 19603 9766 19655 9818
rect 19667 9766 19719 9818
rect 3976 9664 4028 9716
rect 2780 9639 2832 9648
rect 2780 9605 2789 9639
rect 2789 9605 2823 9639
rect 2823 9605 2832 9639
rect 2780 9596 2832 9605
rect 4528 9596 4580 9648
rect 6276 9664 6328 9716
rect 7196 9664 7248 9716
rect 9680 9664 9732 9716
rect 15016 9664 15068 9716
rect 16580 9664 16632 9716
rect 18144 9664 18196 9716
rect 18696 9664 18748 9716
rect 20628 9664 20680 9716
rect 20996 9664 21048 9716
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 5540 9528 5592 9580
rect 8760 9596 8812 9648
rect 11796 9639 11848 9648
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 12716 9596 12768 9648
rect 13728 9596 13780 9648
rect 15108 9596 15160 9648
rect 16396 9596 16448 9648
rect 16948 9639 17000 9648
rect 16948 9605 16957 9639
rect 16957 9605 16991 9639
rect 16991 9605 17000 9639
rect 16948 9596 17000 9605
rect 5908 9528 5960 9580
rect 3332 9503 3384 9512
rect 3332 9469 3366 9503
rect 3366 9469 3384 9503
rect 3332 9460 3384 9469
rect 4896 9460 4948 9512
rect 5264 9460 5316 9512
rect 7196 9528 7248 9580
rect 7656 9528 7708 9580
rect 8208 9528 8260 9580
rect 8392 9571 8444 9580
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 1492 9392 1544 9444
rect 3700 9392 3752 9444
rect 5264 9324 5316 9376
rect 5724 9392 5776 9444
rect 7932 9460 7984 9512
rect 8116 9460 8168 9512
rect 10232 9528 10284 9580
rect 16304 9528 16356 9580
rect 18236 9596 18288 9648
rect 19156 9596 19208 9648
rect 9864 9460 9916 9512
rect 10968 9460 11020 9512
rect 12624 9460 12676 9512
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 13360 9460 13412 9512
rect 13820 9460 13872 9512
rect 7656 9392 7708 9444
rect 8852 9392 8904 9444
rect 9496 9392 9548 9444
rect 9680 9392 9732 9444
rect 9772 9392 9824 9444
rect 6828 9324 6880 9376
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10508 9392 10560 9444
rect 11152 9392 11204 9444
rect 12348 9392 12400 9444
rect 15108 9392 15160 9444
rect 10692 9324 10744 9376
rect 13912 9324 13964 9376
rect 14372 9324 14424 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 15292 9503 15344 9512
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 16948 9460 17000 9512
rect 19340 9528 19392 9580
rect 19708 9528 19760 9580
rect 19800 9528 19852 9580
rect 20720 9528 20772 9580
rect 21272 9528 21324 9580
rect 16396 9392 16448 9444
rect 16580 9392 16632 9444
rect 18604 9503 18656 9512
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 17868 9367 17920 9376
rect 17868 9333 17877 9367
rect 17877 9333 17911 9367
rect 17911 9333 17920 9367
rect 17868 9324 17920 9333
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 18420 9392 18472 9444
rect 19432 9460 19484 9512
rect 19984 9460 20036 9512
rect 22652 9392 22704 9444
rect 8379 9222 8431 9274
rect 8443 9222 8495 9274
rect 8507 9222 8559 9274
rect 8571 9222 8623 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 15904 9222 15956 9274
rect 15968 9222 16020 9274
rect 2412 9120 2464 9172
rect 3332 9120 3384 9172
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 4344 9120 4396 9172
rect 4896 9120 4948 9172
rect 5356 9120 5408 9172
rect 6092 9120 6144 9172
rect 7748 9120 7800 9172
rect 1952 9052 2004 9104
rect 2780 8984 2832 9036
rect 5264 9052 5316 9104
rect 6184 8984 6236 9036
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 2964 8916 3016 8968
rect 3976 8916 4028 8968
rect 3608 8780 3660 8832
rect 3700 8780 3752 8832
rect 6828 8916 6880 8968
rect 9312 9120 9364 9172
rect 9772 9120 9824 9172
rect 10416 9120 10468 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 14188 9120 14240 9172
rect 17224 9120 17276 9172
rect 17868 9120 17920 9172
rect 22652 9163 22704 9172
rect 8208 8959 8260 8968
rect 6184 8848 6236 8900
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8576 8916 8628 8968
rect 9036 8916 9088 8968
rect 10048 8848 10100 8900
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 11152 9052 11204 9104
rect 12348 9052 12400 9104
rect 14372 9052 14424 9104
rect 14464 9052 14516 9104
rect 16304 9052 16356 9104
rect 22652 9129 22661 9163
rect 22661 9129 22695 9163
rect 22695 9129 22704 9163
rect 22652 9120 22704 9129
rect 22192 9052 22244 9104
rect 10692 8984 10744 9036
rect 13268 8984 13320 9036
rect 13452 8984 13504 9036
rect 15844 9027 15896 9036
rect 15844 8993 15853 9027
rect 15853 8993 15887 9027
rect 15887 8993 15896 9027
rect 15844 8984 15896 8993
rect 16396 8984 16448 9036
rect 16580 8984 16632 9036
rect 17316 8984 17368 9036
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 11888 8916 11940 8968
rect 11336 8848 11388 8900
rect 12900 8916 12952 8968
rect 16304 8916 16356 8968
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 7748 8780 7800 8832
rect 8024 8780 8076 8832
rect 8208 8780 8260 8832
rect 9036 8780 9088 8832
rect 11796 8780 11848 8832
rect 12716 8780 12768 8832
rect 12900 8780 12952 8832
rect 15108 8780 15160 8832
rect 15292 8780 15344 8832
rect 15568 8780 15620 8832
rect 16396 8780 16448 8832
rect 17132 8780 17184 8832
rect 17868 8823 17920 8832
rect 17868 8789 17877 8823
rect 17877 8789 17911 8823
rect 17911 8789 17920 8823
rect 17868 8780 17920 8789
rect 18144 8984 18196 9036
rect 18236 8916 18288 8968
rect 18512 8916 18564 8968
rect 19340 8984 19392 9036
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 20076 8916 20128 8968
rect 19708 8848 19760 8900
rect 19800 8848 19852 8900
rect 19984 8780 20036 8832
rect 20628 8780 20680 8832
rect 22376 8780 22428 8832
rect 23020 8780 23072 8832
rect 4680 8678 4732 8730
rect 4744 8678 4796 8730
rect 4808 8678 4860 8730
rect 4872 8678 4924 8730
rect 12078 8678 12130 8730
rect 12142 8678 12194 8730
rect 12206 8678 12258 8730
rect 12270 8678 12322 8730
rect 19475 8678 19527 8730
rect 19539 8678 19591 8730
rect 19603 8678 19655 8730
rect 19667 8678 19719 8730
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 5080 8576 5132 8628
rect 2320 8508 2372 8560
rect 3148 8440 3200 8492
rect 3700 8440 3752 8492
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 7012 8508 7064 8560
rect 8576 8576 8628 8628
rect 9036 8576 9088 8628
rect 15108 8576 15160 8628
rect 15384 8576 15436 8628
rect 15844 8576 15896 8628
rect 8484 8508 8536 8560
rect 9128 8508 9180 8560
rect 8024 8440 8076 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8392 8440 8444 8492
rect 9496 8440 9548 8492
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 5540 8372 5592 8424
rect 5724 8372 5776 8424
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 9680 8508 9732 8560
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 11336 8551 11388 8560
rect 11336 8517 11345 8551
rect 11345 8517 11379 8551
rect 11379 8517 11388 8551
rect 11336 8508 11388 8517
rect 13084 8508 13136 8560
rect 10784 8440 10836 8492
rect 11244 8440 11296 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 9680 8372 9732 8381
rect 6552 8304 6604 8356
rect 6092 8236 6144 8288
rect 8300 8304 8352 8356
rect 11796 8372 11848 8424
rect 12808 8415 12860 8424
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 13452 8372 13504 8424
rect 15568 8483 15620 8492
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 17960 8440 18012 8492
rect 18604 8576 18656 8628
rect 18420 8508 18472 8560
rect 22192 8619 22244 8628
rect 15016 8415 15068 8424
rect 15016 8381 15025 8415
rect 15025 8381 15059 8415
rect 15059 8381 15068 8415
rect 15016 8372 15068 8381
rect 15292 8372 15344 8424
rect 12624 8304 12676 8356
rect 12716 8304 12768 8356
rect 10048 8236 10100 8288
rect 10232 8236 10284 8288
rect 10968 8236 11020 8288
rect 11152 8236 11204 8288
rect 11244 8236 11296 8288
rect 12900 8236 12952 8288
rect 13084 8236 13136 8288
rect 13820 8304 13872 8356
rect 14556 8304 14608 8356
rect 14188 8236 14240 8288
rect 17408 8372 17460 8424
rect 17776 8372 17828 8424
rect 18788 8483 18840 8492
rect 18788 8449 18797 8483
rect 18797 8449 18831 8483
rect 18831 8449 18840 8483
rect 22192 8585 22201 8619
rect 22201 8585 22235 8619
rect 22235 8585 22244 8619
rect 22192 8576 22244 8585
rect 22376 8508 22428 8560
rect 18788 8440 18840 8449
rect 19064 8372 19116 8424
rect 20168 8372 20220 8424
rect 20720 8372 20772 8424
rect 22284 8372 22336 8424
rect 17500 8304 17552 8356
rect 18052 8304 18104 8356
rect 19248 8304 19300 8356
rect 20352 8304 20404 8356
rect 20628 8304 20680 8356
rect 17132 8236 17184 8288
rect 20076 8236 20128 8288
rect 8379 8134 8431 8186
rect 8443 8134 8495 8186
rect 8507 8134 8559 8186
rect 8571 8134 8623 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 15904 8134 15956 8186
rect 15968 8134 16020 8186
rect 5448 8032 5500 8084
rect 6000 8032 6052 8084
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 7012 8075 7064 8084
rect 7012 8041 7021 8075
rect 7021 8041 7055 8075
rect 7055 8041 7064 8075
rect 7012 8032 7064 8041
rect 7748 8032 7800 8084
rect 8760 8032 8812 8084
rect 9036 8075 9088 8084
rect 9036 8041 9045 8075
rect 9045 8041 9079 8075
rect 9079 8041 9088 8075
rect 9036 8032 9088 8041
rect 8024 7964 8076 8016
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 5080 7896 5132 7948
rect 5908 7896 5960 7948
rect 4160 7828 4212 7880
rect 7012 7896 7064 7948
rect 7564 7896 7616 7948
rect 7748 7896 7800 7948
rect 8668 7964 8720 8016
rect 11152 7964 11204 8016
rect 11244 7896 11296 7948
rect 6644 7760 6696 7812
rect 8024 7871 8076 7880
rect 7564 7803 7616 7812
rect 7564 7769 7573 7803
rect 7573 7769 7607 7803
rect 7607 7769 7616 7803
rect 7564 7760 7616 7769
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 9680 7871 9732 7880
rect 9680 7837 9689 7871
rect 9689 7837 9723 7871
rect 9723 7837 9732 7871
rect 9680 7828 9732 7837
rect 12624 8032 12676 8084
rect 13360 8032 13412 8084
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 17408 8032 17460 8084
rect 13268 8007 13320 8016
rect 13268 7973 13302 8007
rect 13302 7973 13320 8007
rect 13268 7964 13320 7973
rect 14188 7896 14240 7948
rect 15476 7964 15528 8016
rect 16488 7964 16540 8016
rect 18328 8032 18380 8084
rect 19248 8032 19300 8084
rect 17868 7964 17920 8016
rect 15660 7896 15712 7948
rect 16580 7871 16632 7880
rect 8484 7692 8536 7744
rect 9404 7760 9456 7812
rect 11060 7803 11112 7812
rect 11060 7769 11069 7803
rect 11069 7769 11103 7803
rect 11103 7769 11112 7803
rect 11060 7760 11112 7769
rect 10968 7692 11020 7744
rect 12900 7692 12952 7744
rect 16580 7837 16589 7871
rect 16589 7837 16623 7871
rect 16623 7837 16632 7871
rect 16580 7828 16632 7837
rect 17132 7828 17184 7880
rect 17224 7692 17276 7744
rect 19064 7964 19116 8016
rect 19156 7964 19208 8016
rect 21272 8007 21324 8016
rect 21272 7973 21281 8007
rect 21281 7973 21315 8007
rect 21315 7973 21324 8007
rect 21272 7964 21324 7973
rect 17960 7692 18012 7744
rect 20996 7939 21048 7948
rect 20996 7905 21005 7939
rect 21005 7905 21039 7939
rect 21039 7905 21048 7939
rect 20996 7896 21048 7905
rect 21180 7896 21232 7948
rect 19156 7828 19208 7880
rect 19432 7760 19484 7812
rect 22652 7828 22704 7880
rect 19800 7692 19852 7744
rect 19892 7692 19944 7744
rect 22192 7692 22244 7744
rect 4680 7590 4732 7642
rect 4744 7590 4796 7642
rect 4808 7590 4860 7642
rect 4872 7590 4924 7642
rect 12078 7590 12130 7642
rect 12142 7590 12194 7642
rect 12206 7590 12258 7642
rect 12270 7590 12322 7642
rect 19475 7590 19527 7642
rect 19539 7590 19591 7642
rect 19603 7590 19655 7642
rect 19667 7590 19719 7642
rect 5540 7488 5592 7540
rect 6184 7488 6236 7540
rect 6092 7420 6144 7472
rect 3884 7352 3936 7404
rect 4988 7352 5040 7404
rect 7012 7420 7064 7472
rect 7564 7488 7616 7540
rect 8024 7488 8076 7540
rect 3792 7284 3844 7336
rect 7564 7352 7616 7404
rect 8484 7420 8536 7472
rect 12716 7420 12768 7472
rect 9772 7352 9824 7404
rect 7012 7327 7064 7336
rect 7012 7293 7029 7327
rect 7029 7293 7063 7327
rect 7063 7293 7064 7327
rect 7012 7284 7064 7293
rect 7104 7216 7156 7268
rect 4528 7148 4580 7200
rect 6276 7148 6328 7200
rect 9680 7284 9732 7336
rect 10048 7284 10100 7336
rect 11152 7352 11204 7404
rect 12532 7352 12584 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 13268 7488 13320 7540
rect 15200 7488 15252 7540
rect 14464 7420 14516 7472
rect 16948 7488 17000 7540
rect 19156 7488 19208 7540
rect 18420 7420 18472 7472
rect 8024 7216 8076 7268
rect 10232 7216 10284 7268
rect 11060 7216 11112 7268
rect 11336 7284 11388 7336
rect 9128 7148 9180 7200
rect 11244 7148 11296 7200
rect 11612 7148 11664 7200
rect 12900 7216 12952 7268
rect 13360 7284 13412 7336
rect 14924 7352 14976 7404
rect 16120 7352 16172 7404
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 14740 7284 14792 7336
rect 15108 7327 15160 7336
rect 15108 7293 15117 7327
rect 15117 7293 15151 7327
rect 15151 7293 15160 7327
rect 15108 7284 15160 7293
rect 16948 7284 17000 7336
rect 18236 7284 18288 7336
rect 18696 7284 18748 7336
rect 19064 7284 19116 7336
rect 22744 7284 22796 7336
rect 14924 7216 14976 7268
rect 20720 7216 20772 7268
rect 22468 7259 22520 7268
rect 22468 7225 22477 7259
rect 22477 7225 22511 7259
rect 22511 7225 22520 7259
rect 22468 7216 22520 7225
rect 15108 7148 15160 7200
rect 18512 7148 18564 7200
rect 20076 7148 20128 7200
rect 20444 7148 20496 7200
rect 20996 7148 21048 7200
rect 8379 7046 8431 7098
rect 8443 7046 8495 7098
rect 8507 7046 8559 7098
rect 8571 7046 8623 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 15904 7046 15956 7098
rect 15968 7046 16020 7098
rect 4528 6987 4580 6996
rect 4528 6953 4537 6987
rect 4537 6953 4571 6987
rect 4571 6953 4580 6987
rect 4528 6944 4580 6953
rect 5816 6944 5868 6996
rect 6920 6987 6972 6996
rect 6920 6953 6929 6987
rect 6929 6953 6963 6987
rect 6963 6953 6972 6987
rect 6920 6944 6972 6953
rect 4436 6876 4488 6928
rect 5080 6876 5132 6928
rect 9864 6944 9916 6996
rect 9588 6876 9640 6928
rect 6368 6808 6420 6860
rect 7380 6808 7432 6860
rect 8024 6851 8076 6860
rect 8024 6817 8033 6851
rect 8033 6817 8067 6851
rect 8067 6817 8076 6851
rect 8024 6808 8076 6817
rect 8300 6808 8352 6860
rect 8760 6808 8812 6860
rect 9680 6808 9732 6860
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 4252 6740 4304 6792
rect 5632 6740 5684 6792
rect 5540 6715 5592 6724
rect 5540 6681 5549 6715
rect 5549 6681 5583 6715
rect 5583 6681 5592 6715
rect 5540 6672 5592 6681
rect 6828 6672 6880 6724
rect 7564 6740 7616 6792
rect 7748 6740 7800 6792
rect 8208 6672 8260 6724
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 8392 6672 8444 6724
rect 9404 6740 9456 6792
rect 10876 6944 10928 6996
rect 10968 6944 11020 6996
rect 22744 6944 22796 6996
rect 10232 6876 10284 6928
rect 10048 6808 10100 6860
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 11612 6808 11664 6860
rect 11980 6740 12032 6792
rect 12716 6808 12768 6860
rect 13360 6808 13412 6860
rect 14832 6808 14884 6860
rect 15108 6808 15160 6860
rect 17408 6808 17460 6860
rect 18512 6808 18564 6860
rect 19800 6851 19852 6860
rect 19800 6817 19809 6851
rect 19809 6817 19843 6851
rect 19843 6817 19852 6851
rect 19800 6808 19852 6817
rect 20812 6808 20864 6860
rect 20996 6808 21048 6860
rect 12900 6740 12952 6792
rect 9680 6604 9732 6656
rect 12624 6672 12676 6724
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 12532 6604 12584 6613
rect 13268 6740 13320 6792
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 17224 6740 17276 6792
rect 17500 6740 17552 6792
rect 18788 6740 18840 6792
rect 19708 6740 19760 6792
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 19064 6672 19116 6724
rect 13820 6604 13872 6656
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 16948 6604 17000 6656
rect 19340 6604 19392 6656
rect 20904 6604 20956 6656
rect 21088 6604 21140 6656
rect 4680 6502 4732 6554
rect 4744 6502 4796 6554
rect 4808 6502 4860 6554
rect 4872 6502 4924 6554
rect 12078 6502 12130 6554
rect 12142 6502 12194 6554
rect 12206 6502 12258 6554
rect 12270 6502 12322 6554
rect 19475 6502 19527 6554
rect 19539 6502 19591 6554
rect 19603 6502 19655 6554
rect 19667 6502 19719 6554
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 7656 6443 7708 6452
rect 7656 6409 7665 6443
rect 7665 6409 7699 6443
rect 7699 6409 7708 6443
rect 7656 6400 7708 6409
rect 7748 6400 7800 6452
rect 8208 6400 8260 6452
rect 8760 6400 8812 6452
rect 9312 6400 9364 6452
rect 11336 6400 11388 6452
rect 12532 6400 12584 6452
rect 23020 6400 23072 6452
rect 6092 6307 6144 6316
rect 6092 6273 6101 6307
rect 6101 6273 6135 6307
rect 6135 6273 6144 6307
rect 6092 6264 6144 6273
rect 7472 6264 7524 6316
rect 5448 6196 5500 6248
rect 10140 6332 10192 6384
rect 8208 6307 8260 6316
rect 8208 6273 8217 6307
rect 8217 6273 8251 6307
rect 8251 6273 8260 6307
rect 8208 6264 8260 6273
rect 9404 6264 9456 6316
rect 8300 6196 8352 6248
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 10600 6332 10652 6384
rect 17408 6375 17460 6384
rect 17408 6341 17417 6375
rect 17417 6341 17451 6375
rect 17451 6341 17460 6375
rect 17408 6332 17460 6341
rect 18420 6375 18472 6384
rect 18420 6341 18429 6375
rect 18429 6341 18463 6375
rect 18463 6341 18472 6375
rect 18420 6332 18472 6341
rect 18788 6332 18840 6384
rect 20720 6332 20772 6384
rect 10416 6264 10468 6316
rect 12256 6264 12308 6316
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 15660 6264 15712 6316
rect 17040 6264 17092 6316
rect 20076 6264 20128 6316
rect 9128 6171 9180 6180
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 10784 6196 10836 6248
rect 11796 6196 11848 6248
rect 13268 6196 13320 6248
rect 14372 6239 14424 6248
rect 10600 6128 10652 6180
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 11152 6060 11204 6112
rect 11980 6060 12032 6112
rect 13636 6128 13688 6180
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 14648 6171 14700 6180
rect 14648 6137 14682 6171
rect 14682 6137 14700 6171
rect 14648 6128 14700 6137
rect 13176 6060 13228 6112
rect 14280 6060 14332 6112
rect 15476 6060 15528 6112
rect 17132 6060 17184 6112
rect 17500 6060 17552 6112
rect 18144 6196 18196 6248
rect 18696 6196 18748 6248
rect 19340 6196 19392 6248
rect 19800 6128 19852 6180
rect 21088 6196 21140 6248
rect 21272 6196 21324 6248
rect 22376 6196 22428 6248
rect 19984 6060 20036 6112
rect 20812 6128 20864 6180
rect 22560 6128 22612 6180
rect 21088 6103 21140 6112
rect 21088 6069 21097 6103
rect 21097 6069 21131 6103
rect 21131 6069 21140 6103
rect 21088 6060 21140 6069
rect 22744 6103 22796 6112
rect 22744 6069 22753 6103
rect 22753 6069 22787 6103
rect 22787 6069 22796 6103
rect 22744 6060 22796 6069
rect 8379 5958 8431 6010
rect 8443 5958 8495 6010
rect 8507 5958 8559 6010
rect 8571 5958 8623 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 15904 5958 15956 6010
rect 15968 5958 16020 6010
rect 5724 5856 5776 5908
rect 6092 5856 6144 5908
rect 6736 5856 6788 5908
rect 7932 5856 7984 5908
rect 8116 5856 8168 5908
rect 9956 5856 10008 5908
rect 10048 5856 10100 5908
rect 11244 5856 11296 5908
rect 11336 5856 11388 5908
rect 12992 5856 13044 5908
rect 13636 5899 13688 5908
rect 13636 5865 13645 5899
rect 13645 5865 13679 5899
rect 13679 5865 13688 5899
rect 13636 5856 13688 5865
rect 14464 5856 14516 5908
rect 18052 5856 18104 5908
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 21640 5856 21692 5908
rect 9772 5788 9824 5840
rect 9864 5788 9916 5840
rect 7288 5720 7340 5772
rect 10232 5720 10284 5772
rect 10416 5720 10468 5772
rect 11980 5720 12032 5772
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 9312 5652 9364 5704
rect 8760 5584 8812 5636
rect 12992 5720 13044 5772
rect 14280 5763 14332 5772
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 14280 5720 14332 5729
rect 14556 5720 14608 5772
rect 16488 5763 16540 5772
rect 16488 5729 16497 5763
rect 16497 5729 16531 5763
rect 16531 5729 16540 5763
rect 16488 5720 16540 5729
rect 17040 5720 17092 5772
rect 19156 5763 19208 5772
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 16672 5652 16724 5704
rect 16948 5652 17000 5704
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 19156 5729 19165 5763
rect 19165 5729 19199 5763
rect 19199 5729 19208 5763
rect 19156 5720 19208 5729
rect 20076 5720 20128 5772
rect 20904 5763 20956 5772
rect 19616 5652 19668 5704
rect 13820 5516 13872 5568
rect 15568 5516 15620 5568
rect 16764 5516 16816 5568
rect 18420 5584 18472 5636
rect 19248 5584 19300 5636
rect 19800 5627 19852 5636
rect 19800 5593 19809 5627
rect 19809 5593 19843 5627
rect 19843 5593 19852 5627
rect 19800 5584 19852 5593
rect 18144 5516 18196 5568
rect 18788 5559 18840 5568
rect 18788 5525 18797 5559
rect 18797 5525 18831 5559
rect 18831 5525 18840 5559
rect 18788 5516 18840 5525
rect 18972 5516 19024 5568
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 21088 5720 21140 5772
rect 21916 5763 21968 5772
rect 21916 5729 21925 5763
rect 21925 5729 21959 5763
rect 21959 5729 21968 5763
rect 21916 5720 21968 5729
rect 20812 5652 20864 5704
rect 21548 5652 21600 5704
rect 20720 5516 20772 5568
rect 21548 5516 21600 5568
rect 4680 5414 4732 5466
rect 4744 5414 4796 5466
rect 4808 5414 4860 5466
rect 4872 5414 4924 5466
rect 12078 5414 12130 5466
rect 12142 5414 12194 5466
rect 12206 5414 12258 5466
rect 12270 5414 12322 5466
rect 19475 5414 19527 5466
rect 19539 5414 19591 5466
rect 19603 5414 19655 5466
rect 19667 5414 19719 5466
rect 7472 5355 7524 5364
rect 7472 5321 7481 5355
rect 7481 5321 7515 5355
rect 7515 5321 7524 5355
rect 7472 5312 7524 5321
rect 10784 5312 10836 5364
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 11244 5312 11296 5364
rect 14372 5312 14424 5364
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 16764 5312 16816 5364
rect 17316 5312 17368 5364
rect 19156 5312 19208 5364
rect 21548 5312 21600 5364
rect 22560 5355 22612 5364
rect 22560 5321 22569 5355
rect 22569 5321 22603 5355
rect 22603 5321 22612 5355
rect 22560 5312 22612 5321
rect 8852 5244 8904 5296
rect 13452 5244 13504 5296
rect 7840 5176 7892 5228
rect 10600 5219 10652 5228
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 10600 5176 10652 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 11336 5176 11388 5228
rect 11612 5219 11664 5228
rect 11612 5185 11621 5219
rect 11621 5185 11655 5219
rect 11655 5185 11664 5219
rect 11612 5176 11664 5185
rect 11888 5176 11940 5228
rect 11980 5176 12032 5228
rect 17960 5244 18012 5296
rect 18512 5244 18564 5296
rect 7196 5108 7248 5160
rect 11796 5108 11848 5160
rect 8668 5040 8720 5092
rect 11336 5040 11388 5092
rect 12992 5108 13044 5160
rect 16764 5176 16816 5228
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 19064 5244 19116 5296
rect 18696 5176 18748 5228
rect 14280 5108 14332 5160
rect 18788 5108 18840 5160
rect 19340 5108 19392 5160
rect 19984 5108 20036 5160
rect 9496 4972 9548 5024
rect 12256 4972 12308 5024
rect 14464 5040 14516 5092
rect 15476 5083 15528 5092
rect 15476 5049 15488 5083
rect 15488 5049 15528 5083
rect 15476 5040 15528 5049
rect 15568 5040 15620 5092
rect 21088 5108 21140 5160
rect 21272 5108 21324 5160
rect 15016 4972 15068 5024
rect 22100 5040 22152 5092
rect 17132 4972 17184 5024
rect 19064 4972 19116 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20812 5015 20864 5024
rect 20812 4981 20821 5015
rect 20821 4981 20855 5015
rect 20855 4981 20864 5015
rect 20812 4972 20864 4981
rect 8379 4870 8431 4922
rect 8443 4870 8495 4922
rect 8507 4870 8559 4922
rect 8571 4870 8623 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 15904 4870 15956 4922
rect 15968 4870 16020 4922
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 10324 4811 10376 4820
rect 10324 4777 10333 4811
rect 10333 4777 10367 4811
rect 10367 4777 10376 4811
rect 10324 4768 10376 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 12532 4768 12584 4820
rect 12808 4768 12860 4820
rect 14832 4768 14884 4820
rect 16212 4768 16264 4820
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 11704 4632 11756 4684
rect 12348 4675 12400 4684
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 11888 4564 11940 4616
rect 12348 4641 12357 4675
rect 12357 4641 12391 4675
rect 12391 4641 12400 4675
rect 12348 4632 12400 4641
rect 13820 4700 13872 4752
rect 14924 4700 14976 4752
rect 16948 4768 17000 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 22100 4768 22152 4820
rect 16672 4700 16724 4752
rect 20812 4700 20864 4752
rect 15660 4632 15712 4684
rect 15844 4632 15896 4684
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14924 4564 14976 4616
rect 15200 4564 15252 4616
rect 18972 4632 19024 4684
rect 19892 4632 19944 4684
rect 21364 4675 21416 4684
rect 21364 4641 21398 4675
rect 21398 4641 21416 4675
rect 21364 4632 21416 4641
rect 18512 4564 18564 4616
rect 19156 4564 19208 4616
rect 19800 4564 19852 4616
rect 15568 4496 15620 4548
rect 20720 4564 20772 4616
rect 21088 4607 21140 4616
rect 21088 4573 21097 4607
rect 21097 4573 21131 4607
rect 21131 4573 21140 4607
rect 21088 4564 21140 4573
rect 14096 4428 14148 4480
rect 14280 4428 14332 4480
rect 14556 4428 14608 4480
rect 15292 4428 15344 4480
rect 15752 4428 15804 4480
rect 16672 4428 16724 4480
rect 16948 4428 17000 4480
rect 19340 4428 19392 4480
rect 20904 4496 20956 4548
rect 22284 4428 22336 4480
rect 4680 4326 4732 4378
rect 4744 4326 4796 4378
rect 4808 4326 4860 4378
rect 4872 4326 4924 4378
rect 12078 4326 12130 4378
rect 12142 4326 12194 4378
rect 12206 4326 12258 4378
rect 12270 4326 12322 4378
rect 19475 4326 19527 4378
rect 19539 4326 19591 4378
rect 19603 4326 19655 4378
rect 19667 4326 19719 4378
rect 10232 4224 10284 4276
rect 14004 4224 14056 4276
rect 9588 4156 9640 4208
rect 10508 4156 10560 4208
rect 11796 4156 11848 4208
rect 12624 4156 12676 4208
rect 14280 4224 14332 4276
rect 16212 4224 16264 4276
rect 23204 4224 23256 4276
rect 11704 4088 11756 4140
rect 14004 4088 14056 4140
rect 17776 4156 17828 4208
rect 19524 4156 19576 4208
rect 14372 4088 14424 4140
rect 15660 4088 15712 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 17408 4088 17460 4140
rect 18512 4088 18564 4140
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 19064 4088 19116 4097
rect 11060 4020 11112 4072
rect 15200 4020 15252 4072
rect 15292 4020 15344 4072
rect 16948 4020 17000 4072
rect 18972 4020 19024 4072
rect 20720 4020 20772 4072
rect 21640 4063 21692 4072
rect 21640 4029 21674 4063
rect 21674 4029 21692 4063
rect 21640 4020 21692 4029
rect 12440 3952 12492 4004
rect 11428 3884 11480 3936
rect 11520 3884 11572 3936
rect 13820 3952 13872 4004
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 13084 3927 13136 3936
rect 13084 3893 13093 3927
rect 13093 3893 13127 3927
rect 13127 3893 13136 3927
rect 13084 3884 13136 3893
rect 13268 3884 13320 3936
rect 14648 3884 14700 3936
rect 14924 3995 14976 4004
rect 14924 3961 14958 3995
rect 14958 3961 14976 3995
rect 14924 3952 14976 3961
rect 15108 3952 15160 4004
rect 19156 3952 19208 4004
rect 15568 3884 15620 3936
rect 15660 3884 15712 3936
rect 16580 3884 16632 3936
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 18420 3927 18472 3936
rect 18420 3893 18429 3927
rect 18429 3893 18463 3927
rect 18463 3893 18472 3927
rect 18420 3884 18472 3893
rect 20812 3884 20864 3936
rect 21364 3884 21416 3936
rect 8379 3782 8431 3834
rect 8443 3782 8495 3834
rect 8507 3782 8559 3834
rect 8571 3782 8623 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 15904 3782 15956 3834
rect 15968 3782 16020 3834
rect 12440 3680 12492 3732
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 17224 3680 17276 3732
rect 9220 3612 9272 3664
rect 13544 3655 13596 3664
rect 13544 3621 13553 3655
rect 13553 3621 13587 3655
rect 13587 3621 13596 3655
rect 13544 3612 13596 3621
rect 13636 3655 13688 3664
rect 13636 3621 13645 3655
rect 13645 3621 13679 3655
rect 13679 3621 13688 3655
rect 13636 3612 13688 3621
rect 13820 3612 13872 3664
rect 18420 3680 18472 3732
rect 21640 3680 21692 3732
rect 17408 3655 17460 3664
rect 17408 3621 17442 3655
rect 17442 3621 17460 3655
rect 17408 3612 17460 3621
rect 11520 3587 11572 3596
rect 11520 3553 11529 3587
rect 11529 3553 11563 3587
rect 11563 3553 11572 3587
rect 11520 3544 11572 3553
rect 14556 3587 14608 3596
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 11888 3476 11940 3528
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 13820 3408 13872 3460
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15016 3544 15068 3596
rect 15936 3544 15988 3596
rect 16488 3544 16540 3596
rect 19248 3587 19300 3596
rect 19248 3553 19282 3587
rect 19282 3553 19300 3587
rect 19248 3544 19300 3553
rect 20720 3544 20772 3596
rect 21916 3544 21968 3596
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 14832 3476 14884 3528
rect 12900 3340 12952 3392
rect 14372 3340 14424 3392
rect 15568 3340 15620 3392
rect 16120 3408 16172 3460
rect 16396 3408 16448 3460
rect 17040 3476 17092 3528
rect 18328 3476 18380 3528
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 18420 3408 18472 3460
rect 18604 3340 18656 3392
rect 19156 3340 19208 3392
rect 4680 3238 4732 3290
rect 4744 3238 4796 3290
rect 4808 3238 4860 3290
rect 4872 3238 4924 3290
rect 12078 3238 12130 3290
rect 12142 3238 12194 3290
rect 12206 3238 12258 3290
rect 12270 3238 12322 3290
rect 19475 3238 19527 3290
rect 19539 3238 19591 3290
rect 19603 3238 19655 3290
rect 19667 3238 19719 3290
rect 15108 3136 15160 3188
rect 15476 3136 15528 3188
rect 11520 3068 11572 3120
rect 14096 3068 14148 3120
rect 14280 3111 14332 3120
rect 14280 3077 14289 3111
rect 14289 3077 14323 3111
rect 14323 3077 14332 3111
rect 14280 3068 14332 3077
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 12808 3000 12860 3052
rect 15016 3068 15068 3120
rect 14740 3043 14792 3052
rect 14740 3009 14749 3043
rect 14749 3009 14783 3043
rect 14783 3009 14792 3043
rect 14740 3000 14792 3009
rect 15384 3000 15436 3052
rect 2412 2932 2464 2984
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 6000 2932 6052 2984
rect 17408 3136 17460 3188
rect 19156 3136 19208 3188
rect 19248 3136 19300 3188
rect 15844 3068 15896 3120
rect 16212 3068 16264 3120
rect 21916 3136 21968 3188
rect 16028 3000 16080 3052
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 17408 3000 17460 3052
rect 20720 3043 20772 3052
rect 15752 2932 15804 2984
rect 16580 2975 16632 2984
rect 1676 2796 1728 2848
rect 16580 2941 16614 2975
rect 16614 2941 16632 2975
rect 16580 2932 16632 2941
rect 17592 2932 17644 2984
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 11980 2796 12032 2848
rect 13636 2796 13688 2848
rect 17040 2864 17092 2916
rect 19248 2932 19300 2984
rect 21456 2932 21508 2984
rect 18328 2864 18380 2916
rect 16396 2796 16448 2848
rect 19064 2796 19116 2848
rect 20904 2864 20956 2916
rect 22560 2796 22612 2848
rect 8379 2694 8431 2746
rect 8443 2694 8495 2746
rect 8507 2694 8559 2746
rect 8571 2694 8623 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 15904 2694 15956 2746
rect 15968 2694 16020 2746
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 13360 2592 13412 2601
rect 11796 2524 11848 2576
rect 15660 2592 15712 2644
rect 15292 2524 15344 2576
rect 15660 2499 15712 2508
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 15660 2465 15669 2499
rect 15669 2465 15703 2499
rect 15703 2465 15712 2499
rect 15660 2456 15712 2465
rect 17408 2592 17460 2644
rect 18420 2524 18472 2576
rect 18604 2567 18656 2576
rect 18604 2533 18638 2567
rect 18638 2533 18656 2567
rect 18604 2524 18656 2533
rect 19064 2592 19116 2644
rect 20260 2592 20312 2644
rect 20444 2592 20496 2644
rect 20904 2524 20956 2576
rect 16304 2456 16356 2508
rect 16764 2388 16816 2440
rect 16948 2456 17000 2508
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 19340 2456 19392 2508
rect 20720 2456 20772 2508
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 20996 2388 21048 2440
rect 17592 2320 17644 2372
rect 20812 2320 20864 2372
rect 14464 2252 14516 2304
rect 16580 2252 16632 2304
rect 19984 2252 20036 2304
rect 4680 2150 4732 2202
rect 4744 2150 4796 2202
rect 4808 2150 4860 2202
rect 4872 2150 4924 2202
rect 12078 2150 12130 2202
rect 12142 2150 12194 2202
rect 12206 2150 12258 2202
rect 12270 2150 12322 2202
rect 19475 2150 19527 2202
rect 19539 2150 19591 2202
rect 19603 2150 19655 2202
rect 19667 2150 19719 2202
rect 16304 2048 16356 2100
rect 18696 2048 18748 2100
rect 17684 1912 17736 1964
rect 20812 1912 20864 1964
rect 17316 1300 17368 1352
rect 19340 1300 19392 1352
<< metal2 >>
rect 294 23920 350 24400
rect 846 23920 902 24400
rect 1490 23920 1546 24400
rect 2134 23920 2190 24400
rect 2778 23920 2834 24400
rect 3422 23920 3478 24400
rect 4066 23920 4122 24400
rect 4710 23920 4766 24400
rect 5354 23920 5410 24400
rect 5998 23920 6054 24400
rect 6642 23920 6698 24400
rect 7286 23920 7342 24400
rect 7930 23920 7986 24400
rect 8574 23920 8630 24400
rect 9218 23920 9274 24400
rect 9862 23920 9918 24400
rect 10506 23920 10562 24400
rect 11150 23920 11206 24400
rect 11794 23920 11850 24400
rect 12438 23920 12494 24400
rect 13082 23920 13138 24400
rect 13726 23920 13782 24400
rect 14370 23920 14426 24400
rect 15014 23920 15070 24400
rect 15658 23920 15714 24400
rect 16302 23920 16358 24400
rect 16946 23920 17002 24400
rect 17590 23920 17646 24400
rect 18234 23920 18290 24400
rect 18878 23920 18934 24400
rect 19522 23920 19578 24400
rect 20166 23920 20222 24400
rect 20350 24032 20406 24041
rect 20350 23967 20406 23976
rect 308 21146 336 23920
rect 296 21140 348 21146
rect 296 21082 348 21088
rect 860 20262 888 23920
rect 1504 21690 1532 23920
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 21049 1440 21422
rect 1952 21344 2004 21350
rect 1952 21286 2004 21292
rect 1398 21040 1454 21049
rect 1398 20975 1454 20984
rect 1492 20936 1544 20942
rect 1412 20884 1492 20890
rect 1412 20878 1544 20884
rect 1412 20862 1532 20878
rect 1412 20398 1440 20862
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 848 20256 900 20262
rect 848 20198 900 20204
rect 1412 19922 1440 20334
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1780 18737 1808 18770
rect 1766 18728 1822 18737
rect 1766 18663 1822 18672
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1780 18222 1808 18566
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1674 17776 1730 17785
rect 1674 17711 1676 17720
rect 1728 17711 1730 17720
rect 1676 17682 1728 17688
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1872 15638 1900 15846
rect 1860 15632 1912 15638
rect 1860 15574 1912 15580
rect 1872 15026 1900 15574
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 14618 1440 14758
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1768 14476 1820 14482
rect 1872 14464 1900 14962
rect 1820 14436 1900 14464
rect 1768 14418 1820 14424
rect 1780 14074 1808 14418
rect 1858 14376 1914 14385
rect 1858 14311 1914 14320
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 1872 13530 1900 14311
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1676 12912 1728 12918
rect 1674 12880 1676 12889
rect 1728 12880 1730 12889
rect 1674 12815 1730 12824
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1596 12306 1624 12718
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 11218 1532 11630
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1504 10674 1532 11154
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 10130 1532 10610
rect 1492 10124 1544 10130
rect 1412 10084 1492 10112
rect 1412 9586 1440 10084
rect 1492 10066 1544 10072
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 9081 1532 9386
rect 1964 9110 1992 21286
rect 2148 20058 2176 23920
rect 2792 23066 2820 23920
rect 2792 23038 2912 23066
rect 2594 21584 2650 21593
rect 2594 21519 2596 21528
rect 2648 21519 2650 21528
rect 2596 21490 2648 21496
rect 2596 21412 2648 21418
rect 2596 21354 2648 21360
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2136 20052 2188 20058
rect 2136 19994 2188 20000
rect 2332 19718 2360 20266
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2240 18902 2268 19178
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 2424 18834 2452 19246
rect 2412 18828 2464 18834
rect 2332 18788 2412 18816
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2148 17202 2176 17682
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2044 16652 2096 16658
rect 2148 16640 2176 17138
rect 2096 16612 2176 16640
rect 2044 16594 2096 16600
rect 2240 10033 2268 18634
rect 2332 18290 2360 18788
rect 2412 18770 2464 18776
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2332 17882 2360 18226
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2332 16998 2360 17682
rect 2320 16992 2372 16998
rect 2320 16934 2372 16940
rect 2226 10024 2282 10033
rect 2226 9959 2282 9968
rect 2424 9178 2452 18158
rect 2516 12209 2544 21286
rect 2608 17649 2636 21354
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19514 2820 19858
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2594 17640 2650 17649
rect 2594 17575 2650 17584
rect 2778 17232 2834 17241
rect 2778 17167 2834 17176
rect 2792 17134 2820 17167
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2792 16697 2820 16730
rect 2778 16688 2834 16697
rect 2778 16623 2834 16632
rect 2780 16244 2832 16250
rect 2884 16232 2912 23038
rect 3436 22386 3464 23920
rect 4080 23066 4108 23920
rect 3896 23038 4108 23066
rect 4724 23066 4752 23920
rect 4724 23038 5028 23066
rect 3436 22358 3556 22386
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 2976 21078 3004 21286
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 3344 20806 3372 21286
rect 3436 21010 3464 21286
rect 3424 21004 3476 21010
rect 3424 20946 3476 20952
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 3068 19310 3096 20334
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2962 17640 3018 17649
rect 2962 17575 3018 17584
rect 2976 16726 3004 17575
rect 3160 17184 3188 19858
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3068 17156 3188 17184
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 3068 16674 3096 17156
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3160 16794 3188 17002
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3068 16646 3188 16674
rect 2832 16204 2912 16232
rect 2780 16186 2832 16192
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15366 2728 15914
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2502 12200 2558 12209
rect 2502 12135 2558 12144
rect 2608 10266 2636 13330
rect 2700 13326 2728 15302
rect 2976 14822 3004 15506
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2884 14074 2912 14486
rect 3068 14346 3096 14826
rect 3160 14498 3188 16646
rect 3252 15042 3280 19722
rect 3344 19310 3372 20742
rect 3436 20602 3464 20946
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3436 16454 3464 16594
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16250 3464 16390
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3344 15201 3372 15438
rect 3330 15192 3386 15201
rect 3330 15127 3386 15136
rect 3252 15014 3372 15042
rect 3160 14470 3280 14498
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13530 3188 13670
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 3252 13258 3280 14470
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2700 12170 2728 12718
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2792 11898 2820 12310
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2792 9654 2820 10066
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 1952 9104 2004 9110
rect 1490 9072 1546 9081
rect 1952 9046 2004 9052
rect 2792 9042 2820 9590
rect 1490 9007 1546 9016
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2332 8566 2360 8910
rect 2884 8634 2912 12650
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2962 11656 3018 11665
rect 3068 11626 3096 12174
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 2962 11591 3018 11600
rect 3056 11620 3108 11626
rect 2976 8974 3004 11591
rect 3056 11562 3108 11568
rect 3068 11354 3096 11562
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 3068 9586 3096 10066
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 3160 8498 3188 11494
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3252 8430 3280 12038
rect 3344 11121 3372 15014
rect 3422 14512 3478 14521
rect 3422 14447 3424 14456
rect 3476 14447 3478 14456
rect 3424 14418 3476 14424
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3436 13410 3464 14010
rect 3528 13818 3556 22358
rect 3792 21412 3844 21418
rect 3792 21354 3844 21360
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3620 19922 3648 20538
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 3620 17882 3648 18090
rect 3712 18086 3740 18770
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3620 17202 3648 17818
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3712 17270 3740 17478
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3700 17128 3752 17134
rect 3606 17096 3662 17105
rect 3662 17076 3700 17082
rect 3662 17070 3752 17076
rect 3662 17054 3740 17070
rect 3606 17031 3662 17040
rect 3620 16794 3648 17031
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3620 15706 3648 15846
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3712 15638 3740 15914
rect 3700 15632 3752 15638
rect 3700 15574 3752 15580
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3712 13938 3740 14758
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3528 13790 3740 13818
rect 3436 13382 3648 13410
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3528 12322 3556 13194
rect 3620 12442 3648 13382
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3528 12294 3648 12322
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3330 11112 3386 11121
rect 3330 11047 3386 11056
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10606 3372 10950
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10130 3372 10542
rect 3436 10470 3464 11562
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11150 3556 11494
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3528 10810 3556 11086
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3344 9518 3372 9862
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3344 9178 3372 9454
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3620 8838 3648 12294
rect 3712 11354 3740 13790
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3698 11112 3754 11121
rect 3698 11047 3754 11056
rect 3712 9450 3740 11047
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3712 8498 3740 8774
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 2502 7984 2558 7993
rect 2502 7919 2504 7928
rect 2556 7919 2558 7928
rect 2504 7890 2556 7896
rect 1950 3088 2006 3097
rect 1950 3023 1952 3032
rect 2004 3023 2006 3032
rect 1952 2994 2004 3000
rect 2412 2984 2464 2990
rect 2516 2972 2544 7890
rect 3804 7342 3832 21354
rect 3896 19786 3924 23038
rect 4654 21788 4950 21808
rect 4710 21786 4734 21788
rect 4790 21786 4814 21788
rect 4870 21786 4894 21788
rect 4732 21734 4734 21786
rect 4796 21734 4808 21786
rect 4870 21734 4872 21786
rect 4710 21732 4734 21734
rect 4790 21732 4814 21734
rect 4870 21732 4894 21734
rect 4654 21712 4950 21732
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4068 21344 4120 21350
rect 3974 21312 4030 21321
rect 4068 21286 4120 21292
rect 3974 21247 4030 21256
rect 3988 20874 4016 21247
rect 4080 21146 4108 21286
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 4172 20210 4200 21422
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 3988 20182 4200 20210
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3988 19666 4016 20182
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3896 19638 4016 19666
rect 3896 16946 3924 19638
rect 4080 18358 4108 19790
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 4172 18222 4200 19994
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4264 17746 4292 20742
rect 4356 19378 4384 20878
rect 4448 20602 4476 21286
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4448 19990 4476 20538
rect 4540 20398 4568 21286
rect 4654 20700 4950 20720
rect 4710 20698 4734 20700
rect 4790 20698 4814 20700
rect 4870 20698 4894 20700
rect 4732 20646 4734 20698
rect 4796 20646 4808 20698
rect 4870 20646 4872 20698
rect 4710 20644 4734 20646
rect 4790 20644 4814 20646
rect 4870 20644 4894 20646
rect 4654 20624 4950 20644
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 4540 19514 4568 20334
rect 4654 19612 4950 19632
rect 4710 19610 4734 19612
rect 4790 19610 4814 19612
rect 4870 19610 4894 19612
rect 4732 19558 4734 19610
rect 4796 19558 4808 19610
rect 4870 19558 4872 19610
rect 4710 19556 4734 19558
rect 4790 19556 4814 19558
rect 4870 19556 4894 19558
rect 4654 19536 4950 19556
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 5000 19446 5028 23038
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5092 19990 5120 21422
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 4988 19440 5040 19446
rect 4988 19382 5040 19388
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 4448 18873 4476 19246
rect 4434 18864 4490 18873
rect 4434 18799 4490 18808
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4356 18358 4384 18634
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 4172 17184 4200 17546
rect 3988 17156 4200 17184
rect 3988 17066 4016 17156
rect 4252 17128 4304 17134
rect 4250 17096 4252 17105
rect 4304 17096 4306 17105
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 4068 17060 4120 17066
rect 4250 17031 4306 17040
rect 4068 17002 4120 17008
rect 4080 16946 4108 17002
rect 4252 16992 4304 16998
rect 3896 16918 4016 16946
rect 4080 16918 4200 16946
rect 4252 16934 4304 16940
rect 3882 16824 3938 16833
rect 3882 16759 3938 16768
rect 3896 7410 3924 16759
rect 3988 13326 4016 16918
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4080 14278 4108 16594
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4080 13802 4108 14214
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4172 13530 4200 16918
rect 4264 16794 4292 16934
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4264 15570 4292 16458
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4264 14958 4292 15370
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4356 14793 4384 15846
rect 4448 15688 4476 17614
rect 4540 17610 4568 19314
rect 5092 19310 5120 19654
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 18970 4752 19110
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4654 18524 4950 18544
rect 4710 18522 4734 18524
rect 4790 18522 4814 18524
rect 4870 18522 4894 18524
rect 4732 18470 4734 18522
rect 4796 18470 4808 18522
rect 4870 18470 4872 18522
rect 4710 18468 4734 18470
rect 4790 18468 4814 18470
rect 4870 18468 4894 18470
rect 4654 18448 4950 18468
rect 5000 18426 5028 18702
rect 5080 18624 5132 18630
rect 5078 18592 5080 18601
rect 5132 18592 5134 18601
rect 5078 18527 5134 18536
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4816 18057 4844 18090
rect 4802 18048 4858 18057
rect 4802 17983 4858 17992
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 4528 17604 4580 17610
rect 4528 17546 4580 17552
rect 4654 17436 4950 17456
rect 4710 17434 4734 17436
rect 4790 17434 4814 17436
rect 4870 17434 4894 17436
rect 4732 17382 4734 17434
rect 4796 17382 4808 17434
rect 4870 17382 4872 17434
rect 4710 17380 4734 17382
rect 4790 17380 4814 17382
rect 4870 17380 4894 17382
rect 4654 17360 4950 17380
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4540 16114 4568 17206
rect 4632 16590 4660 17206
rect 4986 17096 5042 17105
rect 4986 17031 5042 17040
rect 5000 16998 5028 17031
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5092 16833 5120 17682
rect 5078 16824 5134 16833
rect 5078 16759 5134 16768
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4654 16348 4950 16368
rect 4710 16346 4734 16348
rect 4790 16346 4814 16348
rect 4870 16346 4894 16348
rect 4732 16294 4734 16346
rect 4796 16294 4808 16346
rect 4870 16294 4872 16346
rect 4710 16292 4734 16294
rect 4790 16292 4814 16294
rect 4870 16292 4894 16294
rect 4654 16272 4950 16292
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4896 15904 4948 15910
rect 4710 15872 4766 15881
rect 4896 15846 4948 15852
rect 4710 15807 4766 15816
rect 4528 15700 4580 15706
rect 4448 15660 4528 15688
rect 4528 15642 4580 15648
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4342 14784 4398 14793
rect 4342 14719 4398 14728
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 14074 4292 14214
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4250 13832 4306 13841
rect 4250 13767 4252 13776
rect 4304 13767 4306 13776
rect 4252 13738 4304 13744
rect 4250 13696 4306 13705
rect 4250 13631 4306 13640
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4158 13424 4214 13433
rect 4158 13359 4214 13368
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3976 12164 4028 12170
rect 4080 12152 4108 12582
rect 4028 12124 4108 12152
rect 3976 12106 4028 12112
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 9722 4016 11698
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3988 8974 4016 9658
rect 4080 9178 4108 11630
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4172 7886 4200 13359
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 4264 6798 4292 13631
rect 4356 12306 4384 14282
rect 4448 13734 4476 14894
rect 4540 13920 4568 15642
rect 4724 15638 4752 15807
rect 4908 15745 4936 15846
rect 4894 15736 4950 15745
rect 4894 15671 4950 15680
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4724 15502 4752 15574
rect 4908 15570 4936 15671
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4654 15260 4950 15280
rect 4710 15258 4734 15260
rect 4790 15258 4814 15260
rect 4870 15258 4894 15260
rect 4732 15206 4734 15258
rect 4796 15206 4808 15258
rect 4870 15206 4872 15258
rect 4710 15204 4734 15206
rect 4790 15204 4814 15206
rect 4870 15204 4894 15206
rect 4654 15184 4950 15204
rect 5000 15026 5028 16594
rect 5184 16522 5212 20946
rect 5276 20262 5304 21286
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5276 18834 5304 19178
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16794 5304 16934
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5078 16144 5134 16153
rect 5078 16079 5134 16088
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4620 14816 4672 14822
rect 4618 14784 4620 14793
rect 4672 14784 4674 14793
rect 4618 14719 4674 14728
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4654 14172 4950 14192
rect 4710 14170 4734 14172
rect 4790 14170 4814 14172
rect 4870 14170 4894 14172
rect 4732 14118 4734 14170
rect 4796 14118 4808 14170
rect 4870 14118 4872 14170
rect 4710 14116 4734 14118
rect 4790 14116 4814 14118
rect 4870 14116 4894 14118
rect 4654 14096 4950 14116
rect 4894 13968 4950 13977
rect 4620 13932 4672 13938
rect 4540 13892 4620 13920
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4540 13326 4568 13892
rect 4894 13903 4896 13912
rect 4620 13874 4672 13880
rect 4948 13903 4950 13912
rect 4896 13874 4948 13880
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 13462 4660 13670
rect 4620 13456 4672 13462
rect 4620 13398 4672 13404
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4654 13084 4950 13104
rect 4710 13082 4734 13084
rect 4790 13082 4814 13084
rect 4870 13082 4894 13084
rect 4732 13030 4734 13082
rect 4796 13030 4808 13082
rect 4870 13030 4872 13082
rect 4710 13028 4734 13030
rect 4790 13028 4814 13030
rect 4870 13028 4894 13030
rect 4654 13008 4950 13028
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4908 12442 4936 12718
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4620 12232 4672 12238
rect 4540 12192 4620 12220
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11558 4476 12038
rect 4540 11762 4568 12192
rect 4620 12174 4672 12180
rect 4908 12170 4936 12378
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4654 11996 4950 12016
rect 4710 11994 4734 11996
rect 4790 11994 4814 11996
rect 4870 11994 4894 11996
rect 4732 11942 4734 11994
rect 4796 11942 4808 11994
rect 4870 11942 4872 11994
rect 4710 11940 4734 11942
rect 4790 11940 4814 11942
rect 4870 11940 4894 11942
rect 4654 11920 4950 11940
rect 4804 11824 4856 11830
rect 4802 11792 4804 11801
rect 4856 11792 4858 11801
rect 4528 11756 4580 11762
rect 4802 11727 4858 11736
rect 4896 11756 4948 11762
rect 4528 11698 4580 11704
rect 4896 11698 4948 11704
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4540 11370 4568 11698
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4540 11342 4752 11370
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4356 9178 4384 11018
rect 4448 10810 4476 11154
rect 4724 11150 4752 11342
rect 4816 11286 4844 11494
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4908 11218 4936 11698
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4712 11144 4764 11150
rect 4908 11121 4936 11154
rect 4712 11086 4764 11092
rect 4894 11112 4950 11121
rect 4528 11076 4580 11082
rect 4894 11047 4950 11056
rect 4528 11018 4580 11024
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4448 10198 4476 10746
rect 4540 10606 4568 11018
rect 4654 10908 4950 10928
rect 4710 10906 4734 10908
rect 4790 10906 4814 10908
rect 4870 10906 4894 10908
rect 4732 10854 4734 10906
rect 4796 10854 4808 10906
rect 4870 10854 4872 10906
rect 4710 10852 4734 10854
rect 4790 10852 4814 10854
rect 4870 10852 4894 10854
rect 4654 10832 4950 10852
rect 4894 10704 4950 10713
rect 4894 10639 4896 10648
rect 4948 10639 4950 10648
rect 4896 10610 4948 10616
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4434 10024 4490 10033
rect 4434 9959 4490 9968
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4448 6934 4476 9959
rect 4540 9654 4568 10542
rect 4654 9820 4950 9840
rect 4710 9818 4734 9820
rect 4790 9818 4814 9820
rect 4870 9818 4894 9820
rect 4732 9766 4734 9818
rect 4796 9766 4808 9818
rect 4870 9766 4872 9818
rect 4710 9764 4734 9766
rect 4790 9764 4814 9766
rect 4870 9764 4894 9766
rect 4654 9744 4950 9764
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 9178 4936 9454
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4654 8732 4950 8752
rect 4710 8730 4734 8732
rect 4790 8730 4814 8732
rect 4870 8730 4894 8732
rect 4732 8678 4734 8730
rect 4796 8678 4808 8730
rect 4870 8678 4872 8730
rect 4710 8676 4734 8678
rect 4790 8676 4814 8678
rect 4870 8676 4894 8678
rect 4654 8656 4950 8676
rect 4654 7644 4950 7664
rect 4710 7642 4734 7644
rect 4790 7642 4814 7644
rect 4870 7642 4894 7644
rect 4732 7590 4734 7642
rect 4796 7590 4808 7642
rect 4870 7590 4872 7642
rect 4710 7588 4734 7590
rect 4790 7588 4814 7590
rect 4870 7588 4894 7590
rect 4654 7568 4950 7588
rect 5000 7410 5028 14214
rect 5092 8634 5120 16079
rect 5184 15994 5212 16458
rect 5184 15966 5304 15994
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 14958 5212 15846
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5170 14784 5226 14793
rect 5170 14719 5226 14728
rect 5184 13841 5212 14719
rect 5170 13832 5226 13841
rect 5170 13767 5226 13776
rect 5170 13696 5226 13705
rect 5170 13631 5226 13640
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5078 8528 5134 8537
rect 5184 8498 5212 13631
rect 5276 12753 5304 15966
rect 5368 13161 5396 23920
rect 6012 23066 6040 23920
rect 6012 23038 6224 23066
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5448 21072 5500 21078
rect 5448 21014 5500 21020
rect 5460 20262 5488 21014
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5460 18986 5488 19654
rect 5552 19378 5580 21490
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5632 20324 5684 20330
rect 5632 20266 5684 20272
rect 5644 19922 5672 20266
rect 5828 19990 5856 21286
rect 5920 20398 5948 21286
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5920 19786 5948 20334
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 5998 19680 6054 19689
rect 5998 19615 6054 19624
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5460 18958 5580 18986
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5460 17882 5488 18770
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5552 17762 5580 18958
rect 5736 18902 5764 19110
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5828 18086 5856 19110
rect 6012 18170 6040 19615
rect 5920 18142 6040 18170
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5460 17734 5580 17762
rect 5460 14793 5488 17734
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5446 14784 5502 14793
rect 5446 14719 5502 14728
rect 5552 13546 5580 17138
rect 5722 16552 5778 16561
rect 5722 16487 5778 16496
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5644 15881 5672 16118
rect 5736 16046 5764 16487
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5630 15872 5686 15881
rect 5630 15807 5686 15816
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5460 13518 5580 13546
rect 5354 13152 5410 13161
rect 5354 13087 5410 13096
rect 5460 12764 5488 13518
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 12918 5580 13398
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5262 12744 5318 12753
rect 5460 12736 5580 12764
rect 5262 12679 5318 12688
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5276 12186 5304 12378
rect 5276 12158 5396 12186
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5276 11898 5304 12038
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5276 9518 5304 11290
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 9110 5304 9318
rect 5368 9178 5396 12158
rect 5460 11354 5488 12378
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 10690 5580 12736
rect 5460 10662 5580 10690
rect 5460 9466 5488 10662
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10266 5580 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5552 9586 5580 10202
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5460 9438 5580 9466
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5354 8800 5410 8809
rect 5354 8735 5410 8744
rect 5368 8498 5396 8735
rect 5078 8463 5134 8472
rect 5172 8492 5224 8498
rect 5092 7954 5120 8463
rect 5172 8434 5224 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5552 8430 5580 9438
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 7002 4568 7142
rect 4528 6996 4580 7002
rect 4528 6938 4580 6944
rect 5092 6934 5120 7890
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4654 6556 4950 6576
rect 4710 6554 4734 6556
rect 4790 6554 4814 6556
rect 4870 6554 4894 6556
rect 4732 6502 4734 6554
rect 4796 6502 4808 6554
rect 4870 6502 4872 6554
rect 4710 6500 4734 6502
rect 4790 6500 4814 6502
rect 4870 6500 4894 6502
rect 4654 6480 4950 6500
rect 5460 6254 5488 8026
rect 5538 7712 5594 7721
rect 5538 7647 5594 7656
rect 5552 7546 5580 7647
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5644 6882 5672 15438
rect 5816 14884 5868 14890
rect 5816 14826 5868 14832
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5736 12238 5764 12786
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 9450 5764 11154
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5552 6854 5672 6882
rect 5552 6730 5580 6854
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5644 6458 5672 6734
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5736 5914 5764 8366
rect 5828 7002 5856 14826
rect 5920 13977 5948 18142
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 6012 16833 6040 18022
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 17338 6132 17478
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 5998 16824 6054 16833
rect 5998 16759 6054 16768
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6012 15570 6040 16662
rect 6104 16114 6132 17070
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 6012 14822 6040 15506
rect 6104 15502 6132 16050
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 5906 13968 5962 13977
rect 5906 13903 5962 13912
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 13530 5948 13738
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5906 13152 5962 13161
rect 5906 13087 5962 13096
rect 5920 9586 5948 13087
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5906 8256 5962 8265
rect 5906 8191 5962 8200
rect 5920 7954 5948 8191
rect 6012 8090 6040 14758
rect 6104 14482 6132 14758
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 13462 6132 13806
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6090 13288 6146 13297
rect 6090 13223 6146 13232
rect 6104 9178 6132 13223
rect 6196 10606 6224 23038
rect 6460 21412 6512 21418
rect 6460 21354 6512 21360
rect 6472 21010 6500 21354
rect 6460 21004 6512 21010
rect 6460 20946 6512 20952
rect 6472 20602 6500 20946
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6288 17542 6316 17682
rect 6380 17678 6408 20266
rect 6656 19514 6684 23920
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6748 20398 6776 20946
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6840 19854 6868 20742
rect 6932 20058 6960 21286
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6552 19440 6604 19446
rect 6552 19382 6604 19388
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6472 18630 6500 19314
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 6288 17048 6316 17478
rect 6380 17270 6408 17614
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 6288 17020 6500 17048
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6288 15994 6316 16526
rect 6366 16144 6422 16153
rect 6366 16079 6368 16088
rect 6420 16079 6422 16088
rect 6368 16050 6420 16056
rect 6288 15966 6408 15994
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6288 12345 6316 15846
rect 6380 15570 6408 15966
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6368 14884 6420 14890
rect 6368 14826 6420 14832
rect 6380 14346 6408 14826
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6380 12850 6408 13874
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6274 12336 6330 12345
rect 6274 12271 6330 12280
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6288 11354 6316 12038
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6196 9042 6224 10406
rect 6288 10198 6316 11290
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6380 10810 6408 11154
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6366 10704 6422 10713
rect 6366 10639 6422 10648
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6090 8528 6146 8537
rect 6090 8463 6146 8472
rect 6104 8430 6132 8463
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6104 7562 6132 8230
rect 6012 7534 6132 7562
rect 6196 7546 6224 8842
rect 6184 7540 6236 7546
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 4654 5468 4950 5488
rect 4710 5466 4734 5468
rect 4790 5466 4814 5468
rect 4870 5466 4894 5468
rect 4732 5414 4734 5466
rect 4796 5414 4808 5466
rect 4870 5414 4872 5466
rect 4710 5412 4734 5414
rect 4790 5412 4814 5414
rect 4870 5412 4894 5414
rect 4654 5392 4950 5412
rect 4654 4380 4950 4400
rect 4710 4378 4734 4380
rect 4790 4378 4814 4380
rect 4870 4378 4894 4380
rect 4732 4326 4734 4378
rect 4796 4326 4808 4378
rect 4870 4326 4872 4378
rect 4710 4324 4734 4326
rect 4790 4324 4814 4326
rect 4870 4324 4894 4326
rect 4654 4304 4950 4324
rect 4654 3292 4950 3312
rect 4710 3290 4734 3292
rect 4790 3290 4814 3292
rect 4870 3290 4894 3292
rect 4732 3238 4734 3290
rect 4796 3238 4808 3290
rect 4870 3238 4872 3290
rect 4710 3236 4734 3238
rect 4790 3236 4814 3238
rect 4870 3236 4894 3238
rect 4654 3216 4950 3236
rect 6012 2990 6040 7534
rect 6184 7482 6236 7488
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6104 6322 6132 7414
rect 6288 7206 6316 9658
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6380 6866 6408 10639
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6104 5914 6132 6258
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6472 5710 6500 17020
rect 6564 13308 6592 19382
rect 6840 19174 6868 19790
rect 7300 19718 7328 23920
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7392 21146 7420 21286
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7392 20398 7420 21082
rect 7760 21078 7788 21354
rect 7748 21072 7800 21078
rect 7748 21014 7800 21020
rect 7760 20602 7788 21014
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7852 19854 7880 20334
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 6828 19168 6880 19174
rect 6656 19128 6828 19156
rect 6656 18970 6684 19128
rect 6828 19110 6880 19116
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 7380 18896 7432 18902
rect 7300 18856 7380 18884
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 17202 6776 18566
rect 7010 18456 7066 18465
rect 7010 18391 7066 18400
rect 7024 18086 7052 18391
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6748 15366 6776 15982
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6656 13462 6684 13942
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6564 13280 6684 13308
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6564 11626 6592 12242
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6564 10130 6592 11018
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 8362 6592 8774
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6550 8256 6606 8265
rect 6550 8191 6606 8200
rect 6564 8090 6592 8191
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6656 7818 6684 13280
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6748 5914 6776 15302
rect 6840 14958 6868 15506
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14278 6868 14894
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 14113 6868 14214
rect 6826 14104 6882 14113
rect 6826 14039 6882 14048
rect 6840 13852 6868 14039
rect 6932 14006 6960 17818
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6840 13824 6960 13852
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 12782 6868 13670
rect 6932 13462 6960 13824
rect 6900 13456 6960 13462
rect 6952 13416 6960 13456
rect 6900 13398 6952 13404
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12306 6868 12718
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6840 11762 6868 12242
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6840 10577 6868 11086
rect 6826 10568 6882 10577
rect 6826 10503 6882 10512
rect 6932 10266 6960 11562
rect 7024 11014 7052 18022
rect 7194 16144 7250 16153
rect 7194 16079 7196 16088
rect 7248 16079 7250 16088
rect 7196 16050 7248 16056
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15745 7236 15846
rect 7194 15736 7250 15745
rect 7194 15671 7250 15680
rect 7300 14890 7328 18856
rect 7380 18838 7432 18844
rect 7576 18766 7604 19654
rect 7852 19514 7880 19790
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7944 18970 7972 23920
rect 8588 21672 8616 23920
rect 8220 21644 8616 21672
rect 8220 20040 8248 21644
rect 9034 21584 9090 21593
rect 9034 21519 9090 21528
rect 8852 21412 8904 21418
rect 8852 21354 8904 21360
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8353 21244 8649 21264
rect 8409 21242 8433 21244
rect 8489 21242 8513 21244
rect 8569 21242 8593 21244
rect 8431 21190 8433 21242
rect 8495 21190 8507 21242
rect 8569 21190 8571 21242
rect 8409 21188 8433 21190
rect 8489 21188 8513 21190
rect 8569 21188 8593 21190
rect 8353 21168 8649 21188
rect 8680 21078 8708 21286
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8772 20602 8800 21286
rect 8864 21146 8892 21354
rect 9048 21146 9076 21519
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8353 20156 8649 20176
rect 8409 20154 8433 20156
rect 8489 20154 8513 20156
rect 8569 20154 8593 20156
rect 8431 20102 8433 20154
rect 8495 20102 8507 20154
rect 8569 20102 8571 20154
rect 8409 20100 8433 20102
rect 8489 20100 8513 20102
rect 8569 20100 8593 20102
rect 8353 20080 8649 20100
rect 8220 20012 8524 20040
rect 8114 19816 8170 19825
rect 8114 19751 8170 19760
rect 8128 19174 8156 19751
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8220 19553 8248 19654
rect 8206 19544 8262 19553
rect 8206 19479 8262 19488
rect 8312 19310 8340 19654
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8116 19168 8168 19174
rect 8312 19156 8340 19246
rect 8496 19242 8524 20012
rect 8576 19984 8628 19990
rect 8576 19926 8628 19932
rect 8588 19825 8616 19926
rect 8574 19816 8630 19825
rect 8574 19751 8630 19760
rect 8772 19242 8800 20538
rect 8864 20482 8892 21082
rect 8864 20454 9076 20482
rect 9048 20398 9076 20454
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9232 19922 9260 23920
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8956 19689 8984 19790
rect 9680 19712 9732 19718
rect 8942 19680 8998 19689
rect 9680 19654 9732 19660
rect 8942 19615 8998 19624
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8116 19110 8168 19116
rect 8220 19128 8340 19156
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8220 18902 8248 19128
rect 8353 19068 8649 19088
rect 8409 19066 8433 19068
rect 8489 19066 8513 19068
rect 8569 19066 8593 19068
rect 8431 19014 8433 19066
rect 8495 19014 8507 19066
rect 8569 19014 8571 19066
rect 8409 19012 8433 19014
rect 8489 19012 8513 19014
rect 8569 19012 8593 19014
rect 8353 18992 8649 19012
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8220 18170 8248 18566
rect 8312 18358 8340 18838
rect 8680 18630 8708 19178
rect 8864 18970 8892 19450
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 9692 18834 9720 19654
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9402 18728 9458 18737
rect 9402 18663 9458 18672
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8300 18216 8352 18222
rect 8220 18164 8300 18170
rect 8220 18158 8352 18164
rect 8220 18142 8340 18158
rect 7930 17776 7986 17785
rect 8220 17762 8248 18142
rect 8353 17980 8649 18000
rect 8409 17978 8433 17980
rect 8489 17978 8513 17980
rect 8569 17978 8593 17980
rect 8431 17926 8433 17978
rect 8495 17926 8507 17978
rect 8569 17926 8571 17978
rect 8409 17924 8433 17926
rect 8489 17924 8513 17926
rect 8569 17924 8593 17926
rect 8353 17904 8649 17924
rect 8220 17734 8340 17762
rect 7930 17711 7986 17720
rect 7944 17542 7972 17711
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7484 17066 7512 17478
rect 8312 17202 8340 17734
rect 8760 17604 8812 17610
rect 8760 17546 8812 17552
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7392 15570 7420 16390
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 9081 6868 9318
rect 6826 9072 6882 9081
rect 6826 9007 6882 9016
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 6730 6868 8910
rect 6932 7002 6960 10066
rect 7024 8673 7052 10134
rect 7010 8664 7066 8673
rect 7010 8599 7066 8608
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7024 8090 7052 8502
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 7024 7478 7052 7890
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 7012 7336 7064 7342
rect 7010 7304 7012 7313
rect 7064 7304 7066 7313
rect 7116 7274 7144 11562
rect 7208 9722 7236 12310
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7010 7239 7066 7248
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 7208 5166 7236 9522
rect 7300 5778 7328 12242
rect 7392 10690 7420 15506
rect 7484 12050 7512 17002
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 16114 7696 16934
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7576 12374 7604 13398
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7484 12022 7604 12050
rect 7470 11928 7526 11937
rect 7470 11863 7526 11872
rect 7484 10810 7512 11863
rect 7576 11665 7604 12022
rect 7562 11656 7618 11665
rect 7562 11591 7618 11600
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7576 11218 7604 11494
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7392 10662 7512 10690
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7392 6866 7420 10474
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7484 6322 7512 10662
rect 7576 7954 7604 11154
rect 7668 9586 7696 16050
rect 7760 11778 7788 16662
rect 7852 13734 7880 17070
rect 7944 16726 7972 17070
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8353 16892 8649 16912
rect 8409 16890 8433 16892
rect 8489 16890 8513 16892
rect 8569 16890 8593 16892
rect 8431 16838 8433 16890
rect 8495 16838 8507 16890
rect 8569 16838 8571 16890
rect 8409 16836 8433 16838
rect 8489 16836 8513 16838
rect 8569 16836 8593 16838
rect 8353 16816 8649 16836
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 8298 16688 8354 16697
rect 8680 16658 8708 16934
rect 8298 16623 8354 16632
rect 8668 16652 8720 16658
rect 8022 16008 8078 16017
rect 8022 15943 8078 15952
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7944 15570 7972 15846
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 8036 14822 8064 15943
rect 8312 15892 8340 16623
rect 8668 16594 8720 16600
rect 8772 16538 8800 17546
rect 8852 16720 8904 16726
rect 8850 16688 8852 16697
rect 8904 16688 8906 16697
rect 8850 16623 8906 16632
rect 8680 16510 8800 16538
rect 8680 15994 8708 16510
rect 8850 16144 8906 16153
rect 8850 16079 8906 16088
rect 8864 16046 8892 16079
rect 8852 16040 8904 16046
rect 8680 15966 8800 15994
rect 8852 15982 8904 15988
rect 8220 15864 8340 15892
rect 8668 15904 8720 15910
rect 8220 15688 8248 15864
rect 8668 15846 8720 15852
rect 8353 15804 8649 15824
rect 8409 15802 8433 15804
rect 8489 15802 8513 15804
rect 8569 15802 8593 15804
rect 8431 15750 8433 15802
rect 8495 15750 8507 15802
rect 8569 15750 8571 15802
rect 8409 15748 8433 15750
rect 8489 15748 8513 15750
rect 8569 15748 8593 15750
rect 8353 15728 8649 15748
rect 8220 15660 8340 15688
rect 8312 14906 8340 15660
rect 8484 15360 8536 15366
rect 8482 15328 8484 15337
rect 8536 15328 8538 15337
rect 8482 15263 8538 15272
rect 8496 14958 8524 15263
rect 8128 14878 8340 14906
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 8036 13462 8064 14214
rect 8128 13462 8156 14878
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14482 8248 14758
rect 8353 14716 8649 14736
rect 8409 14714 8433 14716
rect 8489 14714 8513 14716
rect 8569 14714 8593 14716
rect 8431 14662 8433 14714
rect 8495 14662 8507 14714
rect 8569 14662 8571 14714
rect 8409 14660 8433 14662
rect 8489 14660 8513 14662
rect 8569 14660 8593 14662
rect 8353 14640 8649 14660
rect 8576 14544 8628 14550
rect 8574 14512 8576 14521
rect 8628 14512 8630 14521
rect 8208 14476 8260 14482
rect 8574 14447 8630 14456
rect 8208 14418 8260 14424
rect 8588 14278 8616 14447
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 13190 7972 13330
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 8036 12889 8064 13262
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8022 12880 8078 12889
rect 7840 12844 7892 12850
rect 8022 12815 8078 12824
rect 7840 12786 7892 12792
rect 7852 11937 7880 12786
rect 8128 12782 8156 13126
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7838 11928 7894 11937
rect 7838 11863 7894 11872
rect 7760 11750 7880 11778
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7562 7848 7618 7857
rect 7562 7783 7564 7792
rect 7616 7783 7618 7792
rect 7564 7754 7616 7760
rect 7562 7576 7618 7585
rect 7562 7511 7564 7520
rect 7616 7511 7618 7520
rect 7564 7482 7616 7488
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7576 6798 7604 7346
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7576 5817 7604 6598
rect 7668 6458 7696 9386
rect 7760 9178 7788 11630
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7760 8090 7788 8774
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7313 7788 7890
rect 7746 7304 7802 7313
rect 7746 7239 7802 7248
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6458 7788 6734
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7562 5808 7618 5817
rect 7288 5772 7340 5778
rect 7562 5743 7618 5752
rect 7288 5714 7340 5720
rect 7470 5400 7526 5409
rect 7470 5335 7472 5344
rect 7524 5335 7526 5344
rect 7472 5306 7524 5312
rect 7852 5234 7880 11750
rect 7944 9602 7972 12310
rect 8036 12306 8064 12582
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11626 8064 12038
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8036 10538 8064 10950
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7944 9574 8064 9602
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 5914 7972 9454
rect 8036 8838 8064 9574
rect 8128 9518 8156 12718
rect 8220 12374 8248 13670
rect 8353 13628 8649 13648
rect 8409 13626 8433 13628
rect 8489 13626 8513 13628
rect 8569 13626 8593 13628
rect 8431 13574 8433 13626
rect 8495 13574 8507 13626
rect 8569 13574 8571 13626
rect 8409 13572 8433 13574
rect 8489 13572 8513 13574
rect 8569 13572 8593 13574
rect 8353 13552 8649 13572
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8588 12850 8616 13398
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8353 12540 8649 12560
rect 8409 12538 8433 12540
rect 8489 12538 8513 12540
rect 8569 12538 8593 12540
rect 8431 12486 8433 12538
rect 8495 12486 8507 12538
rect 8569 12486 8571 12538
rect 8409 12484 8433 12486
rect 8489 12484 8513 12486
rect 8569 12484 8593 12486
rect 8353 12464 8649 12484
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8588 11898 8616 12038
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8353 11452 8649 11472
rect 8409 11450 8433 11452
rect 8489 11450 8513 11452
rect 8569 11450 8593 11452
rect 8431 11398 8433 11450
rect 8495 11398 8507 11450
rect 8569 11398 8571 11450
rect 8409 11396 8433 11398
rect 8489 11396 8513 11398
rect 8569 11396 8593 11398
rect 8353 11376 8649 11396
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10130 8248 10406
rect 8353 10364 8649 10384
rect 8409 10362 8433 10364
rect 8489 10362 8513 10364
rect 8569 10362 8593 10364
rect 8431 10310 8433 10362
rect 8495 10310 8507 10362
rect 8569 10310 8571 10362
rect 8409 10308 8433 10310
rect 8489 10308 8513 10310
rect 8569 10308 8593 10310
rect 8353 10288 8649 10308
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8390 9752 8446 9761
rect 8390 9687 8446 9696
rect 8404 9586 8432 9687
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8022 8664 8078 8673
rect 8022 8599 8078 8608
rect 8036 8498 8064 8599
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8024 8016 8076 8022
rect 8022 7984 8024 7993
rect 8076 7984 8078 7993
rect 8022 7919 8078 7928
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8036 7546 8064 7822
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8022 7440 8078 7449
rect 8022 7375 8078 7384
rect 8036 7274 8064 7375
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8022 6896 8078 6905
rect 8022 6831 8024 6840
rect 8076 6831 8078 6840
rect 8024 6802 8076 6808
rect 8128 5914 8156 9318
rect 8220 8974 8248 9522
rect 8353 9276 8649 9296
rect 8409 9274 8433 9276
rect 8489 9274 8513 9276
rect 8569 9274 8593 9276
rect 8431 9222 8433 9274
rect 8495 9222 8507 9274
rect 8569 9222 8571 9274
rect 8409 9220 8433 9222
rect 8489 9220 8513 9222
rect 8569 9220 8593 9222
rect 8353 9200 8649 9220
rect 8298 9072 8354 9081
rect 8298 9007 8354 9016
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8208 8832 8260 8838
rect 8206 8800 8208 8809
rect 8260 8800 8262 8809
rect 8206 8735 8262 8744
rect 8206 8664 8262 8673
rect 8206 8599 8262 8608
rect 8220 8498 8248 8599
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8312 8362 8340 9007
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8482 8800 8538 8809
rect 8482 8735 8538 8744
rect 8496 8566 8524 8735
rect 8588 8634 8616 8910
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8484 8560 8536 8566
rect 8390 8528 8446 8537
rect 8484 8502 8536 8508
rect 8390 8463 8392 8472
rect 8444 8463 8446 8472
rect 8392 8434 8444 8440
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8353 8188 8649 8208
rect 8409 8186 8433 8188
rect 8489 8186 8513 8188
rect 8569 8186 8593 8188
rect 8431 8134 8433 8186
rect 8495 8134 8507 8186
rect 8569 8134 8571 8186
rect 8409 8132 8433 8134
rect 8489 8132 8513 8134
rect 8569 8132 8593 8134
rect 8353 8112 8649 8132
rect 8680 8022 8708 15846
rect 8772 12753 8800 15966
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 15706 8892 15846
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8956 15162 8984 18362
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 9324 18193 9352 18294
rect 9310 18184 9366 18193
rect 9310 18119 9366 18128
rect 9312 17740 9364 17746
rect 9312 17682 9364 17688
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8864 14618 8892 15098
rect 8852 14612 8904 14618
rect 8904 14572 8984 14600
rect 8852 14554 8904 14560
rect 8852 14408 8904 14414
rect 8850 14376 8852 14385
rect 8904 14376 8906 14385
rect 8850 14311 8906 14320
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 12918 8892 14214
rect 8956 13190 8984 14572
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8758 12744 8814 12753
rect 8758 12679 8814 12688
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8864 12442 8892 12582
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8850 12336 8906 12345
rect 8850 12271 8852 12280
rect 8904 12271 8906 12280
rect 8852 12242 8904 12248
rect 8850 12200 8906 12209
rect 8850 12135 8852 12144
rect 8904 12135 8906 12144
rect 8852 12106 8904 12112
rect 8956 12050 8984 12582
rect 8864 12022 8984 12050
rect 8864 11801 8892 12022
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8850 11792 8906 11801
rect 8850 11727 8906 11736
rect 8850 11520 8906 11529
rect 8850 11455 8906 11464
rect 8864 11354 8892 11455
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8772 9654 8800 11086
rect 8956 10606 8984 11834
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8956 10266 8984 10406
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9048 10146 9076 17002
rect 9140 16794 9168 17002
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9140 15706 9168 16594
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 14618 9168 15438
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9140 13025 9168 14418
rect 9126 13016 9182 13025
rect 9126 12951 9182 12960
rect 9232 12782 9260 17614
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9218 12336 9274 12345
rect 9218 12271 9274 12280
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8956 10118 9076 10146
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8864 9450 8892 9862
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8864 8922 8892 9386
rect 8772 8894 8892 8922
rect 8772 8242 8800 8894
rect 8956 8344 8984 10118
rect 9140 10044 9168 11222
rect 9048 10016 9168 10044
rect 9048 8974 9076 10016
rect 9126 9480 9182 9489
rect 9126 9415 9182 9424
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8634 9076 8774
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8566 9168 9415
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 8956 8316 9045 8344
rect 9017 8276 9045 8316
rect 8956 8248 9045 8276
rect 8772 8214 8892 8242
rect 8758 8120 8814 8129
rect 8758 8055 8760 8064
rect 8812 8055 8814 8064
rect 8760 8026 8812 8032
rect 8668 8016 8720 8022
rect 8206 7984 8262 7993
rect 8668 7958 8720 7964
rect 8206 7919 8262 7928
rect 8220 7886 8248 7919
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8484 7744 8536 7750
rect 8482 7712 8484 7721
rect 8536 7712 8538 7721
rect 8482 7647 8538 7656
rect 8482 7576 8538 7585
rect 8482 7511 8538 7520
rect 8496 7478 8524 7511
rect 8484 7472 8536 7478
rect 8298 7440 8354 7449
rect 8220 7398 8298 7426
rect 8220 6730 8248 7398
rect 8484 7414 8536 7420
rect 8298 7375 8354 7384
rect 8353 7100 8649 7120
rect 8409 7098 8433 7100
rect 8489 7098 8513 7100
rect 8569 7098 8593 7100
rect 8431 7046 8433 7098
rect 8495 7046 8507 7098
rect 8569 7046 8571 7098
rect 8409 7044 8433 7046
rect 8489 7044 8513 7046
rect 8569 7044 8593 7046
rect 8353 7024 8649 7044
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8220 6322 8248 6394
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8220 5710 8248 6258
rect 8312 6254 8340 6802
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8404 6361 8432 6666
rect 8390 6352 8446 6361
rect 8390 6287 8446 6296
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8353 6012 8649 6032
rect 8409 6010 8433 6012
rect 8489 6010 8513 6012
rect 8569 6010 8593 6012
rect 8431 5958 8433 6010
rect 8495 5958 8507 6010
rect 8569 5958 8571 6010
rect 8409 5956 8433 5958
rect 8489 5956 8513 5958
rect 8569 5956 8593 5958
rect 8353 5936 8649 5956
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 8680 5098 8708 7958
rect 8864 6882 8892 8214
rect 8772 6866 8892 6882
rect 8760 6860 8892 6866
rect 8812 6854 8892 6860
rect 8760 6802 8812 6808
rect 8956 6780 8984 8248
rect 9034 8120 9090 8129
rect 9034 8055 9036 8064
rect 9088 8055 9090 8064
rect 9036 8026 9088 8032
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 8864 6752 8984 6780
rect 9034 6760 9090 6769
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8772 5642 8800 6394
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8864 5302 8892 6752
rect 9034 6695 9090 6704
rect 9048 6254 9076 6695
rect 9140 6304 9168 7142
rect 9232 7041 9260 12271
rect 9324 12209 9352 17682
rect 9416 16794 9444 18663
rect 9508 17882 9536 18770
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9600 18426 9628 18566
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9588 18080 9640 18086
rect 9678 18048 9734 18057
rect 9640 18028 9678 18034
rect 9588 18022 9678 18028
rect 9600 18006 9678 18022
rect 9678 17983 9734 17992
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9784 17746 9812 20742
rect 9876 20058 9904 23920
rect 9956 21956 10008 21962
rect 9956 21898 10008 21904
rect 9968 21690 9996 21898
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9876 18970 9904 19858
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9876 18222 9904 18906
rect 9864 18216 9916 18222
rect 9968 18193 9996 21422
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 10060 19310 10088 20946
rect 10428 20942 10456 21422
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10428 20398 10456 20878
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10152 20058 10180 20266
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10244 19854 10272 20334
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10244 18766 10272 19790
rect 10414 19544 10470 19553
rect 10414 19479 10416 19488
rect 10468 19479 10470 19488
rect 10416 19450 10468 19456
rect 10520 19446 10548 23920
rect 11164 23066 11192 23920
rect 11164 23038 11376 23066
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10508 19440 10560 19446
rect 10508 19382 10560 19388
rect 10704 19174 10732 19858
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10414 19000 10470 19009
rect 10704 18970 10732 19110
rect 10414 18935 10470 18944
rect 10692 18964 10744 18970
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 9864 18158 9916 18164
rect 9954 18184 10010 18193
rect 9954 18119 10010 18128
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9864 16992 9916 16998
rect 9968 16980 9996 17818
rect 9916 16952 9996 16980
rect 9864 16934 9916 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 10048 16720 10100 16726
rect 9862 16688 9918 16697
rect 9404 16652 9456 16658
rect 9862 16623 9918 16632
rect 9968 16680 10048 16708
rect 9404 16594 9456 16600
rect 9416 16522 9444 16594
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9310 12200 9366 12209
rect 9310 12135 9366 12144
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 9178 9352 10406
rect 9416 9908 9444 16458
rect 9876 16454 9904 16623
rect 9680 16448 9732 16454
rect 9678 16416 9680 16425
rect 9864 16448 9916 16454
rect 9732 16416 9734 16425
rect 9864 16390 9916 16396
rect 9678 16351 9734 16360
rect 9770 16280 9826 16289
rect 9770 16215 9826 16224
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9692 14006 9720 14826
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9784 13802 9812 16215
rect 9864 15564 9916 15570
rect 9968 15552 9996 16680
rect 10048 16662 10100 16668
rect 9916 15524 9996 15552
rect 10048 15564 10100 15570
rect 9864 15506 9916 15512
rect 10048 15506 10100 15512
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9508 12986 9536 13194
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 10044 9536 12718
rect 9600 10470 9628 13359
rect 9876 12782 9904 14010
rect 9968 13870 9996 14418
rect 10060 14074 10088 15506
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10046 13968 10102 13977
rect 10152 13954 10180 18566
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10336 17678 10364 18158
rect 10428 17814 10456 18935
rect 10692 18906 10744 18912
rect 10796 18834 10824 19110
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10414 17640 10470 17649
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10244 16164 10272 17546
rect 10336 17134 10364 17614
rect 10414 17575 10470 17584
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10336 16726 10364 17070
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10324 16176 10376 16182
rect 10244 16136 10324 16164
rect 10244 15065 10272 16136
rect 10324 16118 10376 16124
rect 10428 15910 10456 17575
rect 10782 17096 10838 17105
rect 10782 17031 10838 17040
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 10612 16425 10640 16662
rect 10598 16416 10654 16425
rect 10598 16351 10654 16360
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10230 15056 10286 15065
rect 10230 14991 10286 15000
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10244 14550 10272 14758
rect 10336 14618 10364 14758
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10322 14376 10378 14385
rect 10322 14311 10378 14320
rect 10152 13926 10272 13954
rect 10046 13903 10102 13912
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9968 13258 9996 13806
rect 10060 13734 10088 13903
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9954 12472 10010 12481
rect 9784 12416 9954 12424
rect 9784 12396 9956 12416
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11354 9720 12106
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9680 10736 9732 10742
rect 9678 10704 9680 10713
rect 9732 10704 9734 10713
rect 9678 10639 9734 10648
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9692 10198 9720 10542
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9692 10062 9720 10134
rect 9680 10056 9732 10062
rect 9508 10016 9628 10044
rect 9416 9880 9536 9908
rect 9508 9602 9536 9880
rect 9416 9574 9536 9602
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9310 9072 9366 9081
rect 9310 9007 9366 9016
rect 9218 7032 9274 7041
rect 9218 6967 9274 6976
rect 9324 6458 9352 9007
rect 9416 7818 9444 9574
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 8498 9536 9386
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9600 7562 9628 10016
rect 9680 9998 9732 10004
rect 9784 9761 9812 12396
rect 10008 12407 10010 12416
rect 9956 12378 10008 12384
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 12209 9904 12242
rect 9862 12200 9918 12209
rect 9862 12135 9918 12144
rect 9954 11928 10010 11937
rect 10060 11898 10088 13330
rect 9954 11863 10010 11872
rect 10048 11892 10100 11898
rect 9968 11830 9996 11863
rect 10048 11834 10100 11840
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 11558 10088 11698
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9876 11014 9904 11494
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9968 10674 9996 11018
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10060 10554 10088 11494
rect 10152 11354 10180 13806
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9876 10526 10088 10554
rect 9770 9752 9826 9761
rect 9680 9716 9732 9722
rect 9770 9687 9826 9696
rect 9680 9658 9732 9664
rect 9692 9450 9720 9658
rect 9876 9625 9904 10526
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 9926 9996 10406
rect 10244 10282 10272 13926
rect 10336 13870 10364 14311
rect 10428 13938 10456 15438
rect 10612 15366 10640 16351
rect 10690 16144 10746 16153
rect 10690 16079 10746 16088
rect 10704 16046 10732 16079
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10704 15706 10732 15982
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10612 14958 10640 15302
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10506 14784 10562 14793
rect 10506 14719 10562 14728
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10428 13530 10456 13874
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12850 10456 13262
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10336 12238 10364 12650
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10428 11830 10456 12786
rect 10416 11824 10468 11830
rect 10322 11792 10378 11801
rect 10416 11766 10468 11772
rect 10322 11727 10378 11736
rect 10060 10254 10272 10282
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9862 9616 9918 9625
rect 9862 9551 9918 9560
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9784 9178 9812 9386
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9876 8956 9904 9454
rect 9784 8928 9904 8956
rect 9784 8650 9812 8928
rect 9784 8622 9904 8650
rect 9680 8560 9732 8566
rect 9732 8520 9812 8548
rect 9680 8502 9732 8508
rect 9680 8424 9732 8430
rect 9678 8392 9680 8401
rect 9732 8392 9734 8401
rect 9678 8327 9734 8336
rect 9692 7886 9720 8327
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9508 7534 9628 7562
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9416 6322 9444 6734
rect 9404 6316 9456 6322
rect 9140 6276 9260 6304
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9126 6216 9182 6225
rect 9126 6151 9128 6160
rect 9180 6151 9182 6160
rect 9128 6122 9180 6128
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8353 4924 8649 4944
rect 8409 4922 8433 4924
rect 8489 4922 8513 4924
rect 8569 4922 8593 4924
rect 8431 4870 8433 4922
rect 8495 4870 8507 4922
rect 8569 4870 8571 4922
rect 8409 4868 8433 4870
rect 8489 4868 8513 4870
rect 8569 4868 8593 4870
rect 8353 4848 8649 4868
rect 8353 3836 8649 3856
rect 8409 3834 8433 3836
rect 8489 3834 8513 3836
rect 8569 3834 8593 3836
rect 8431 3782 8433 3834
rect 8495 3782 8507 3834
rect 8569 3782 8571 3834
rect 8409 3780 8433 3782
rect 8489 3780 8513 3782
rect 8569 3780 8593 3782
rect 8353 3760 8649 3780
rect 9232 3670 9260 6276
rect 9404 6258 9456 6264
rect 9310 5944 9366 5953
rect 9310 5879 9366 5888
rect 9324 5710 9352 5879
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9416 5273 9444 6258
rect 9402 5264 9458 5273
rect 9402 5199 9458 5208
rect 9508 5030 9536 7534
rect 9586 7440 9642 7449
rect 9586 7375 9642 7384
rect 9600 7018 9628 7375
rect 9692 7342 9720 7822
rect 9784 7410 9812 8520
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9680 7336 9732 7342
rect 9876 7290 9904 8622
rect 9680 7278 9732 7284
rect 9784 7262 9904 7290
rect 9600 6990 9720 7018
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9600 4214 9628 6870
rect 9692 6866 9720 6990
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9680 6656 9732 6662
rect 9678 6624 9680 6633
rect 9732 6624 9734 6633
rect 9678 6559 9734 6568
rect 9784 5846 9812 7262
rect 9862 7032 9918 7041
rect 9862 6967 9864 6976
rect 9916 6967 9918 6976
rect 9864 6938 9916 6944
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 5846 9904 6802
rect 9968 5914 9996 9862
rect 10060 8906 10088 10254
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10152 9382 10180 10134
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10140 9376 10192 9382
rect 10244 9353 10272 9522
rect 10140 9318 10192 9324
rect 10230 9344 10286 9353
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10046 8800 10102 8809
rect 10046 8735 10102 8744
rect 10060 8294 10088 8735
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10060 6866 10088 7278
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10152 6390 10180 9318
rect 10230 9279 10286 9288
rect 10230 9072 10286 9081
rect 10230 9007 10286 9016
rect 10244 8974 10272 9007
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 8129 10272 8230
rect 10230 8120 10286 8129
rect 10230 8055 10286 8064
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 6934 10272 7210
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5914 10088 6054
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 10230 5808 10286 5817
rect 10230 5743 10232 5752
rect 10284 5743 10286 5752
rect 10232 5714 10284 5720
rect 9862 4856 9918 4865
rect 10336 4826 10364 11727
rect 10428 11150 10456 11766
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10428 10266 10456 11086
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10428 9178 10456 10066
rect 10520 9450 10548 14719
rect 10612 14278 10640 14894
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 13802 10640 14214
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10704 12782 10732 13806
rect 10796 13308 10824 17031
rect 10980 16658 11008 18090
rect 11072 17241 11100 21830
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11058 17232 11114 17241
rect 11058 17167 11114 17176
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11072 16794 11100 17002
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10876 15632 10928 15638
rect 10876 15574 10928 15580
rect 10888 14618 10916 15574
rect 10980 15570 11008 16594
rect 11058 16552 11114 16561
rect 11058 16487 11114 16496
rect 11072 16114 11100 16487
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10980 14346 11008 14894
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 11072 13818 11100 15506
rect 10980 13790 11100 13818
rect 10796 13280 10916 13308
rect 10782 12880 10838 12889
rect 10782 12815 10838 12824
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10598 12336 10654 12345
rect 10598 12271 10654 12280
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 6322 10456 6802
rect 10612 6390 10640 12271
rect 10704 11898 10732 12718
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10796 10606 10824 12815
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9042 10732 9318
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10690 8664 10746 8673
rect 10796 8650 10824 10406
rect 10746 8622 10824 8650
rect 10690 8599 10746 8608
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10428 5778 10456 6258
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10612 5234 10640 6122
rect 10704 5234 10732 8599
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10796 6254 10824 8434
rect 10888 7002 10916 13280
rect 10980 12442 11008 13790
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13462 11100 13670
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11060 12640 11112 12646
rect 11058 12608 11060 12617
rect 11112 12608 11114 12617
rect 11058 12543 11114 12552
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10980 10554 11008 12242
rect 11164 11694 11192 19382
rect 11256 16017 11284 19858
rect 11242 16008 11298 16017
rect 11242 15943 11298 15952
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 12714 11284 15846
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11242 12336 11298 12345
rect 11242 12271 11298 12280
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10980 10526 11100 10554
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 9518 11008 10406
rect 10968 9512 11020 9518
rect 11072 9489 11100 10526
rect 10968 9454 11020 9460
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11164 9353 11192 9386
rect 11150 9344 11206 9353
rect 11150 9279 11206 9288
rect 11256 9194 11284 12271
rect 11348 12209 11376 23038
rect 11704 21412 11756 21418
rect 11704 21354 11756 21360
rect 11716 20602 11744 21354
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11520 20324 11572 20330
rect 11520 20266 11572 20272
rect 11426 18864 11482 18873
rect 11426 18799 11482 18808
rect 11440 17882 11468 18799
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11440 17134 11468 17478
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11440 16794 11468 16934
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 14074 11468 15846
rect 11532 15144 11560 20266
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11624 19718 11652 19994
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11624 18426 11652 18770
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11716 18222 11744 19110
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11624 16697 11652 18022
rect 11716 17882 11744 18158
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11808 17746 11836 23920
rect 12052 21788 12348 21808
rect 12108 21786 12132 21788
rect 12188 21786 12212 21788
rect 12268 21786 12292 21788
rect 12130 21734 12132 21786
rect 12194 21734 12206 21786
rect 12268 21734 12270 21786
rect 12108 21732 12132 21734
rect 12188 21732 12212 21734
rect 12268 21732 12292 21734
rect 12052 21712 12348 21732
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 12176 20788 12204 21422
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12268 21010 12296 21286
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12268 20874 12296 20946
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 11992 20760 12204 20788
rect 11992 20398 12020 20760
rect 12052 20700 12348 20720
rect 12108 20698 12132 20700
rect 12188 20698 12212 20700
rect 12268 20698 12292 20700
rect 12130 20646 12132 20698
rect 12194 20646 12206 20698
rect 12268 20646 12270 20698
rect 12108 20644 12132 20646
rect 12188 20644 12212 20646
rect 12268 20644 12292 20646
rect 12052 20624 12348 20644
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11992 20058 12020 20334
rect 12452 20330 12480 23920
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12084 19938 12112 19994
rect 12544 19990 12572 20742
rect 12808 20392 12860 20398
rect 12714 20360 12770 20369
rect 12808 20334 12860 20340
rect 12714 20295 12770 20304
rect 11992 19922 12112 19938
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 11980 19916 12112 19922
rect 12032 19910 12112 19916
rect 11980 19858 12032 19864
rect 12438 19816 12494 19825
rect 12438 19751 12494 19760
rect 12452 19718 12480 19751
rect 12728 19718 12756 20295
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12052 19612 12348 19632
rect 12108 19610 12132 19612
rect 12188 19610 12212 19612
rect 12268 19610 12292 19612
rect 12130 19558 12132 19610
rect 12194 19558 12206 19610
rect 12268 19558 12270 19610
rect 12108 19556 12132 19558
rect 12188 19556 12212 19558
rect 12268 19556 12292 19558
rect 12052 19536 12348 19556
rect 12530 19544 12586 19553
rect 12530 19479 12532 19488
rect 12584 19479 12586 19488
rect 12532 19450 12584 19456
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11610 16688 11666 16697
rect 11610 16623 11666 16632
rect 11716 16538 11744 17478
rect 11900 17270 11928 17818
rect 11992 17338 12020 18838
rect 12360 18612 12388 19110
rect 12452 18737 12480 19110
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12438 18728 12494 18737
rect 12438 18663 12494 18672
rect 12360 18584 12480 18612
rect 12052 18524 12348 18544
rect 12108 18522 12132 18524
rect 12188 18522 12212 18524
rect 12268 18522 12292 18524
rect 12130 18470 12132 18522
rect 12194 18470 12206 18522
rect 12268 18470 12270 18522
rect 12108 18468 12132 18470
rect 12188 18468 12212 18470
rect 12268 18468 12292 18470
rect 12052 18448 12348 18468
rect 12452 18426 12480 18584
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12452 18306 12480 18362
rect 12544 18329 12572 18770
rect 12360 18278 12480 18306
rect 12530 18320 12586 18329
rect 12360 17814 12388 18278
rect 12530 18255 12586 18264
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12052 17436 12348 17456
rect 12108 17434 12132 17436
rect 12188 17434 12212 17436
rect 12268 17434 12292 17436
rect 12130 17382 12132 17434
rect 12194 17382 12206 17434
rect 12268 17382 12270 17434
rect 12108 17380 12132 17382
rect 12188 17380 12212 17382
rect 12268 17380 12292 17382
rect 12052 17360 12348 17380
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12084 16794 12112 17070
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12268 16658 12296 17206
rect 12636 17202 12664 17682
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 11716 16510 11836 16538
rect 11610 16008 11666 16017
rect 11610 15943 11666 15952
rect 11624 15570 11652 15943
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11532 15116 11652 15144
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14278 11560 14758
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11428 13932 11480 13938
rect 11428 13874 11480 13880
rect 11440 13190 11468 13874
rect 11624 13870 11652 15116
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11334 12200 11390 12209
rect 11334 12135 11390 12144
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11121 11376 12038
rect 11334 11112 11390 11121
rect 11334 11047 11390 11056
rect 11334 10024 11390 10033
rect 11334 9959 11390 9968
rect 11348 9217 11376 9959
rect 10980 9166 11284 9194
rect 11334 9208 11390 9217
rect 10980 8294 11008 9166
rect 11334 9143 11390 9152
rect 11152 9104 11204 9110
rect 11072 9064 11152 9092
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10966 8120 11022 8129
rect 10966 8055 11022 8064
rect 10980 7750 11008 8055
rect 11072 7818 11100 9064
rect 11152 9046 11204 9052
rect 11242 9072 11298 9081
rect 11242 9007 11298 9016
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8294 11192 8910
rect 11256 8498 11284 9007
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11348 8566 11376 8842
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11164 8022 11192 8230
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11256 7954 11284 8230
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11072 7274 11100 7754
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10966 7032 11022 7041
rect 10876 6996 10928 7002
rect 10966 6967 10968 6976
rect 10876 6938 10928 6944
rect 11020 6967 11022 6976
rect 10968 6938 11020 6944
rect 10784 6248 10836 6254
rect 11164 6202 11192 7346
rect 11256 7206 11284 7890
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11348 6458 11376 7278
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 10784 6190 10836 6196
rect 10796 5370 10824 6190
rect 11072 6174 11192 6202
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 9862 4791 9864 4800
rect 9916 4791 9918 4800
rect 10324 4820 10376 4826
rect 9864 4762 9916 4768
rect 10324 4762 10376 4768
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10244 4282 10272 4626
rect 10508 4616 10560 4622
rect 10704 4604 10732 5170
rect 10560 4576 10732 4604
rect 10508 4558 10560 4564
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10520 4214 10548 4558
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 11072 4078 11100 6174
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5370 11192 6054
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11256 5370 11284 5850
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11348 5234 11376 5850
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 11348 4826 11376 5034
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11440 3942 11468 12650
rect 11532 11558 11560 13806
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 8809 11560 10610
rect 11518 8800 11574 8809
rect 11518 8735 11574 8744
rect 11624 7585 11652 12786
rect 11716 11937 11744 15846
rect 11808 14906 11836 16510
rect 11992 15162 12020 16594
rect 12052 16348 12348 16368
rect 12108 16346 12132 16348
rect 12188 16346 12212 16348
rect 12268 16346 12292 16348
rect 12130 16294 12132 16346
rect 12194 16294 12206 16346
rect 12268 16294 12270 16346
rect 12108 16292 12132 16294
rect 12188 16292 12212 16294
rect 12268 16292 12292 16294
rect 12052 16272 12348 16292
rect 12624 16244 12676 16250
rect 12268 16204 12624 16232
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 12084 15570 12112 15914
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12268 15502 12296 16204
rect 12624 16186 12676 16192
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12052 15260 12348 15280
rect 12108 15258 12132 15260
rect 12188 15258 12212 15260
rect 12268 15258 12292 15260
rect 12130 15206 12132 15258
rect 12194 15206 12206 15258
rect 12268 15206 12270 15258
rect 12108 15204 12132 15206
rect 12188 15204 12212 15206
rect 12268 15204 12292 15206
rect 12052 15184 12348 15204
rect 12452 15162 12480 15982
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12544 15609 12572 15642
rect 12530 15600 12586 15609
rect 12530 15535 12586 15544
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12268 14906 12296 14962
rect 11808 14878 12296 14906
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 11992 14226 12020 14878
rect 12164 14816 12216 14822
rect 12162 14784 12164 14793
rect 12216 14784 12218 14793
rect 12162 14719 12218 14728
rect 12360 14385 12388 14894
rect 12452 14618 12480 15098
rect 12624 15088 12676 15094
rect 12624 15030 12676 15036
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12346 14376 12402 14385
rect 12346 14311 12402 14320
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 11900 14198 12020 14226
rect 11900 13938 11928 14198
rect 12052 14172 12348 14192
rect 12108 14170 12132 14172
rect 12188 14170 12212 14172
rect 12268 14170 12292 14172
rect 12130 14118 12132 14170
rect 12194 14118 12206 14170
rect 12268 14118 12270 14170
rect 12108 14116 12132 14118
rect 12188 14116 12212 14118
rect 12268 14116 12292 14118
rect 12052 14096 12348 14116
rect 12452 14074 12480 14282
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12544 13938 12572 14418
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12636 13818 12664 15030
rect 12728 14618 12756 15302
rect 12820 14906 12848 20334
rect 12912 19242 12940 21286
rect 13096 20058 13124 23920
rect 13740 21894 13768 23920
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 21078 13768 21286
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13188 20466 13216 20946
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13096 19394 13124 19654
rect 13004 19366 13124 19394
rect 13004 19310 13032 19366
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12990 18456 13046 18465
rect 12990 18391 13046 18400
rect 13004 18358 13032 18391
rect 12992 18352 13044 18358
rect 12898 18320 12954 18329
rect 12992 18294 13044 18300
rect 12898 18255 12900 18264
rect 12952 18255 12954 18264
rect 12900 18226 12952 18232
rect 13084 18216 13136 18222
rect 13188 18204 13216 20402
rect 13740 20058 13768 21014
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 14016 20058 14044 20742
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14200 19854 14228 21490
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14200 19514 14228 19790
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 13634 19408 13690 19417
rect 13634 19343 13636 19352
rect 13688 19343 13690 19352
rect 13636 19314 13688 19320
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 18630 13308 18770
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13136 18176 13216 18204
rect 13084 18158 13136 18164
rect 13096 17814 13124 18158
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 13280 17134 13308 18566
rect 13268 17128 13320 17134
rect 12990 17096 13046 17105
rect 13268 17070 13320 17076
rect 12990 17031 12992 17040
rect 13044 17031 13046 17040
rect 12992 17002 13044 17008
rect 13556 16794 13584 18566
rect 13648 17882 13676 19314
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13648 16590 13676 17818
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13280 16182 13308 16458
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 16017 13676 16050
rect 13634 16008 13690 16017
rect 13634 15943 13690 15952
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13096 15502 13124 15846
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13096 14958 13124 15438
rect 13084 14952 13136 14958
rect 12820 14878 13032 14906
rect 13084 14894 13136 14900
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 12544 13790 12664 13818
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 11900 13530 11928 13738
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 12176 13394 12204 13670
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11808 12986 11836 13330
rect 11886 13288 11942 13297
rect 11886 13223 11942 13232
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11794 12744 11850 12753
rect 11794 12679 11850 12688
rect 11702 11928 11758 11937
rect 11702 11863 11758 11872
rect 11808 11812 11836 12679
rect 11900 12170 11928 13223
rect 12052 13084 12348 13104
rect 12108 13082 12132 13084
rect 12188 13082 12212 13084
rect 12268 13082 12292 13084
rect 12130 13030 12132 13082
rect 12194 13030 12206 13082
rect 12268 13030 12270 13082
rect 12108 13028 12132 13030
rect 12188 13028 12212 13030
rect 12268 13028 12292 13030
rect 12052 13008 12348 13028
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 12452 12102 12480 12718
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12052 11996 12348 12016
rect 12108 11994 12132 11996
rect 12188 11994 12212 11996
rect 12268 11994 12292 11996
rect 12130 11942 12132 11994
rect 12194 11942 12206 11994
rect 12268 11942 12270 11994
rect 12108 11940 12132 11942
rect 12188 11940 12212 11942
rect 12268 11940 12292 11942
rect 12052 11920 12348 11940
rect 12544 11914 12572 13790
rect 12728 13462 12756 13806
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12624 12368 12676 12374
rect 12624 12310 12676 12316
rect 11716 11784 11836 11812
rect 12452 11886 12572 11914
rect 11610 7576 11666 7585
rect 11610 7511 11666 7520
rect 11612 7200 11664 7206
rect 11518 7168 11574 7177
rect 11612 7142 11664 7148
rect 11518 7103 11574 7112
rect 11532 3942 11560 7103
rect 11624 6866 11652 7142
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11624 5234 11652 6802
rect 11716 6633 11744 11784
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11900 11354 11928 11562
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12268 11218 12296 11494
rect 12452 11286 12480 11886
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 11808 9654 11836 11154
rect 12052 10908 12348 10928
rect 12108 10906 12132 10908
rect 12188 10906 12212 10908
rect 12268 10906 12292 10908
rect 12130 10854 12132 10906
rect 12194 10854 12206 10906
rect 12268 10854 12270 10906
rect 12108 10852 12132 10854
rect 12188 10852 12212 10854
rect 12268 10852 12292 10854
rect 12052 10832 12348 10852
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 11888 10464 11940 10470
rect 12452 10441 12480 10542
rect 12544 10538 12572 11766
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 11888 10406 11940 10412
rect 12438 10432 12494 10441
rect 11900 9994 11928 10406
rect 12438 10367 12494 10376
rect 12530 10296 12586 10305
rect 12530 10231 12586 10240
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 11900 8974 11928 9930
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12052 9820 12348 9840
rect 12108 9818 12132 9820
rect 12188 9818 12212 9820
rect 12268 9818 12292 9820
rect 12130 9766 12132 9818
rect 12194 9766 12206 9818
rect 12268 9766 12270 9818
rect 12108 9764 12132 9766
rect 12188 9764 12212 9766
rect 12268 9764 12292 9766
rect 12052 9744 12348 9764
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 12360 9110 12388 9386
rect 12348 9104 12400 9110
rect 12348 9046 12400 9052
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8430 11836 8774
rect 11900 8498 11928 8910
rect 12052 8732 12348 8752
rect 12108 8730 12132 8732
rect 12188 8730 12212 8732
rect 12268 8730 12292 8732
rect 12130 8678 12132 8730
rect 12194 8678 12206 8730
rect 12268 8678 12270 8730
rect 12108 8676 12132 8678
rect 12188 8676 12212 8678
rect 12268 8676 12292 8678
rect 12052 8656 12348 8676
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11796 6656 11848 6662
rect 11702 6624 11758 6633
rect 11796 6598 11848 6604
rect 11702 6559 11758 6568
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11716 4690 11744 6559
rect 11808 6254 11836 6598
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5166 11836 6190
rect 11900 5234 11928 8434
rect 12052 7644 12348 7664
rect 12108 7642 12132 7644
rect 12188 7642 12212 7644
rect 12268 7642 12292 7644
rect 12130 7590 12132 7642
rect 12194 7590 12206 7642
rect 12268 7590 12270 7642
rect 12108 7588 12132 7590
rect 12188 7588 12212 7590
rect 12268 7588 12292 7590
rect 12052 7568 12348 7588
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 6304 12020 6734
rect 12052 6556 12348 6576
rect 12108 6554 12132 6556
rect 12188 6554 12212 6556
rect 12268 6554 12292 6556
rect 12130 6502 12132 6554
rect 12194 6502 12206 6554
rect 12268 6502 12270 6554
rect 12108 6500 12132 6502
rect 12188 6500 12212 6502
rect 12268 6500 12292 6502
rect 12052 6480 12348 6500
rect 12256 6316 12308 6322
rect 11992 6276 12204 6304
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5778 12020 6054
rect 12176 5817 12204 6276
rect 12256 6258 12308 6264
rect 12162 5808 12218 5817
rect 11980 5772 12032 5778
rect 12162 5743 12218 5752
rect 11980 5714 12032 5720
rect 11992 5234 12020 5714
rect 12268 5710 12296 6258
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12052 5468 12348 5488
rect 12108 5466 12132 5468
rect 12188 5466 12212 5468
rect 12268 5466 12292 5468
rect 12130 5414 12132 5466
rect 12194 5414 12206 5466
rect 12268 5414 12270 5466
rect 12108 5412 12132 5414
rect 12188 5412 12212 5414
rect 12268 5412 12292 5414
rect 12052 5392 12348 5412
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 11704 4684 11756 4690
rect 12268 4672 12296 4966
rect 12348 4684 12400 4690
rect 12268 4644 12348 4672
rect 11704 4626 11756 4632
rect 12348 4626 12400 4632
rect 11716 4146 11744 4626
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11532 3126 11560 3538
rect 11808 3534 11836 4150
rect 11900 3534 11928 4558
rect 12052 4380 12348 4400
rect 12108 4378 12132 4380
rect 12188 4378 12212 4380
rect 12268 4378 12292 4380
rect 12130 4326 12132 4378
rect 12194 4326 12206 4378
rect 12268 4326 12270 4378
rect 12108 4324 12132 4326
rect 12188 4324 12212 4326
rect 12268 4324 12292 4326
rect 12052 4304 12348 4324
rect 12452 4010 12480 9862
rect 12544 7410 12572 10231
rect 12636 9625 12664 12310
rect 12728 11150 12756 12718
rect 12820 12442 12848 14758
rect 13004 13818 13032 14878
rect 12912 13790 13032 13818
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12912 11370 12940 13790
rect 12983 13728 13035 13734
rect 12983 13670 13035 13676
rect 13004 12073 13032 13670
rect 13096 13462 13124 14894
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13096 12306 13124 13398
rect 13188 12481 13216 15846
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13280 12986 13308 15506
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 14521 13492 15302
rect 13542 15192 13598 15201
rect 13542 15127 13598 15136
rect 13450 14512 13506 14521
rect 13450 14447 13506 14456
rect 13452 14272 13504 14278
rect 13372 14232 13452 14260
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13174 12472 13230 12481
rect 13174 12407 13230 12416
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13188 12209 13216 12310
rect 13174 12200 13230 12209
rect 13096 12158 13174 12186
rect 13096 12102 13124 12158
rect 13174 12135 13230 12144
rect 13084 12096 13136 12102
rect 12990 12064 13046 12073
rect 13084 12038 13136 12044
rect 12990 11999 13046 12008
rect 13174 11928 13230 11937
rect 13174 11863 13230 11872
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12820 11342 12940 11370
rect 12716 11144 12768 11150
rect 12820 11121 12848 11342
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12716 11086 12768 11092
rect 12806 11112 12862 11121
rect 12728 10538 12756 11086
rect 12806 11047 12862 11056
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12728 10062 12756 10474
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12728 9654 12756 9998
rect 12716 9648 12768 9654
rect 12622 9616 12678 9625
rect 12716 9590 12768 9596
rect 12622 9551 12678 9560
rect 12728 9518 12756 9590
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12636 9194 12664 9454
rect 12636 9166 12756 9194
rect 12728 8838 12756 9166
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 8362 12756 8774
rect 12820 8514 12848 10950
rect 12912 9738 12940 11154
rect 13004 9926 13032 11222
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12912 9710 13032 9738
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12912 8838 12940 8910
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12820 8486 12940 8514
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12636 8090 12664 8298
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12714 7576 12770 7585
rect 12714 7511 12770 7520
rect 12728 7478 12756 7511
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 6458 12572 6598
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12636 6066 12664 6666
rect 12728 6322 12756 6802
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12636 6038 12756 6066
rect 12728 5409 12756 6038
rect 12714 5400 12770 5409
rect 12714 5335 12770 5344
rect 12622 5264 12678 5273
rect 12622 5199 12678 5208
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12440 3732 12492 3738
rect 12544 3720 12572 4762
rect 12636 4214 12664 5199
rect 12820 4826 12848 8366
rect 12912 8294 12940 8486
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7410 12940 7686
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12898 7304 12954 7313
rect 12898 7239 12900 7248
rect 12952 7239 12954 7248
rect 12900 7210 12952 7216
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12912 6361 12940 6734
rect 12898 6352 12954 6361
rect 12898 6287 12954 6296
rect 13004 5914 13032 9710
rect 13096 8566 13124 11630
rect 13188 11529 13216 11863
rect 13174 11520 13230 11529
rect 13174 11455 13230 11464
rect 13174 11112 13230 11121
rect 13174 11047 13230 11056
rect 13188 9353 13216 11047
rect 13174 9344 13230 9353
rect 13174 9279 13230 9288
rect 13280 9160 13308 12582
rect 13372 12306 13400 14232
rect 13452 14214 13504 14220
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13372 11218 13400 12242
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13464 11098 13492 12718
rect 13556 11354 13584 15127
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13648 12918 13676 14418
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 13648 12646 13676 12854
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13634 12472 13690 12481
rect 13634 12407 13690 12416
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13372 11070 13492 11098
rect 13542 11112 13598 11121
rect 13372 10305 13400 11070
rect 13542 11047 13598 11056
rect 13358 10296 13414 10305
rect 13358 10231 13414 10240
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13372 9178 13400 9454
rect 13188 9132 13308 9160
rect 13360 9172 13412 9178
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13096 6089 13124 8230
rect 13188 6118 13216 9132
rect 13360 9114 13412 9120
rect 13464 9042 13492 10202
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13280 8022 13308 8978
rect 13358 8528 13414 8537
rect 13358 8463 13360 8472
rect 13412 8463 13414 8472
rect 13360 8434 13412 8440
rect 13372 8090 13400 8434
rect 13464 8430 13492 8978
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13280 7546 13308 7958
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13372 7342 13400 8026
rect 13450 7576 13506 7585
rect 13450 7511 13506 7520
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13372 7041 13400 7278
rect 13358 7032 13414 7041
rect 13358 6967 13414 6976
rect 13372 6866 13400 6967
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13268 6792 13320 6798
rect 13464 6746 13492 7511
rect 13268 6734 13320 6740
rect 13280 6254 13308 6734
rect 13372 6718 13492 6746
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13176 6112 13228 6118
rect 13082 6080 13138 6089
rect 13372 6100 13400 6718
rect 13176 6054 13228 6060
rect 13280 6072 13400 6100
rect 13082 6015 13138 6024
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12898 5536 12954 5545
rect 12898 5471 12954 5480
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12492 3692 12572 3720
rect 12440 3674 12492 3680
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 2464 2944 2544 2972
rect 5080 2984 5132 2990
rect 2412 2926 2464 2932
rect 5080 2926 5132 2932
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1688 480 1716 2790
rect 4654 2204 4950 2224
rect 4710 2202 4734 2204
rect 4790 2202 4814 2204
rect 4870 2202 4894 2204
rect 4732 2150 4734 2202
rect 4796 2150 4808 2202
rect 4870 2150 4872 2202
rect 4710 2148 4734 2150
rect 4790 2148 4814 2150
rect 4870 2148 4894 2150
rect 4654 2128 4950 2148
rect 5092 480 5120 2926
rect 8353 2748 8649 2768
rect 8409 2746 8433 2748
rect 8489 2746 8513 2748
rect 8569 2746 8593 2748
rect 8431 2694 8433 2746
rect 8495 2694 8507 2746
rect 8569 2694 8571 2746
rect 8409 2692 8433 2694
rect 8489 2692 8513 2694
rect 8569 2692 8593 2694
rect 8353 2672 8649 2692
rect 11808 2582 11836 3470
rect 12052 3292 12348 3312
rect 12108 3290 12132 3292
rect 12188 3290 12212 3292
rect 12268 3290 12292 3292
rect 12130 3238 12132 3290
rect 12194 3238 12206 3290
rect 12268 3238 12270 3290
rect 12108 3236 12132 3238
rect 12188 3236 12212 3238
rect 12268 3236 12292 3238
rect 12052 3216 12348 3236
rect 12820 3058 12848 3470
rect 12912 3398 12940 5471
rect 13004 5166 13032 5714
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13280 3942 13308 6072
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 13464 4622 13492 5238
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13004 3641 13032 3878
rect 12990 3632 13046 3641
rect 12990 3567 13046 3576
rect 12900 3392 12952 3398
rect 13096 3369 13124 3878
rect 13556 3670 13584 11047
rect 13648 7528 13676 12407
rect 13740 11014 13768 19246
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14016 17270 14044 17682
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 14108 17116 14136 17682
rect 14016 17088 14136 17116
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13832 15337 13860 16050
rect 13818 15328 13874 15337
rect 13818 15263 13874 15272
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13924 14278 13952 14418
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13462 13860 13670
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13832 12322 13860 13398
rect 13924 12481 13952 14214
rect 14016 13433 14044 17088
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16794 14136 16934
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14108 15706 14136 15982
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14200 13818 14228 18770
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14292 17882 14320 18090
rect 14384 18086 14412 23920
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14476 20806 14504 21354
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14476 20398 14504 20742
rect 14660 20602 14688 20946
rect 14844 20777 14872 21422
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14830 20768 14886 20777
rect 14830 20703 14886 20712
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 14464 20392 14516 20398
rect 14464 20334 14516 20340
rect 14556 20324 14608 20330
rect 14556 20266 14608 20272
rect 14568 20058 14596 20266
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14660 19378 14688 20538
rect 14936 20398 14964 20878
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14936 19854 14964 20334
rect 15028 19922 15056 23920
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20398 15240 20742
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 14844 19378 14872 19790
rect 15014 19544 15070 19553
rect 15014 19479 15070 19488
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18426 14504 19110
rect 14844 18766 14872 19314
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14752 18358 14780 18566
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14844 18290 14872 18702
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14830 18184 14886 18193
rect 14830 18119 14886 18128
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14280 16108 14332 16114
rect 14384 16096 14412 17070
rect 14476 16658 14504 18022
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14568 16538 14596 17682
rect 14660 16658 14688 17818
rect 14844 17134 14872 18119
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14332 16068 14412 16096
rect 14280 16050 14332 16056
rect 14384 15706 14412 16068
rect 14476 16510 14596 16538
rect 14738 16552 14794 16561
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14476 15094 14504 16510
rect 14738 16487 14740 16496
rect 14792 16487 14794 16496
rect 14740 16458 14792 16464
rect 14936 15858 14964 19382
rect 15028 19378 15056 19479
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15016 19168 15068 19174
rect 15212 19156 15240 20334
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15304 19514 15332 20266
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15068 19128 15240 19156
rect 15292 19168 15344 19174
rect 15016 19110 15068 19116
rect 15292 19110 15344 19116
rect 15304 19009 15332 19110
rect 15290 19000 15346 19009
rect 15290 18935 15346 18944
rect 15396 18834 15424 19790
rect 15384 18828 15436 18834
rect 15304 18788 15384 18816
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15120 17270 15148 18022
rect 15304 17678 15332 18788
rect 15384 18770 15436 18776
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 15108 17128 15160 17134
rect 15304 17116 15332 17614
rect 15160 17088 15332 17116
rect 15108 17070 15160 17076
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15106 16688 15162 16697
rect 14660 15830 14964 15858
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14464 15088 14516 15094
rect 14384 15048 14464 15076
rect 14200 13790 14320 13818
rect 14002 13424 14058 13433
rect 14002 13359 14058 13368
rect 14186 13424 14242 13433
rect 14186 13359 14242 13368
rect 14002 12608 14058 12617
rect 14002 12543 14058 12552
rect 13910 12472 13966 12481
rect 13910 12407 13966 12416
rect 13832 12294 13952 12322
rect 13818 12200 13874 12209
rect 13818 12135 13874 12144
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13740 9654 13768 10134
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13740 8616 13768 9590
rect 13832 9518 13860 12135
rect 13924 11558 13952 12294
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13924 10305 13952 10950
rect 13910 10296 13966 10305
rect 13910 10231 13966 10240
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13740 8588 13860 8616
rect 13832 8362 13860 8588
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13648 7500 13768 7528
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 5914 13676 6122
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13634 5536 13690 5545
rect 13634 5471 13690 5480
rect 13648 3670 13676 5471
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 13740 3534 13768 7500
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 5681 13860 6598
rect 13818 5672 13874 5681
rect 13818 5607 13874 5616
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 4758 13860 5510
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13818 4176 13874 4185
rect 13818 4111 13874 4120
rect 13832 4010 13860 4111
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13832 3466 13860 3606
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 12900 3334 12952 3340
rect 13082 3360 13138 3369
rect 13082 3295 13138 3304
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 13636 2848 13688 2854
rect 13924 2836 13952 9318
rect 14016 4282 14044 12543
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14108 4486 14136 12242
rect 14200 11762 14228 13359
rect 14292 12345 14320 13790
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14292 12073 14320 12106
rect 14278 12064 14334 12073
rect 14278 11999 14334 12008
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 9994 14228 10542
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14200 9178 14228 9930
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 7954 14228 8230
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14292 6202 14320 11494
rect 14384 9382 14412 15048
rect 14464 15030 14516 15036
rect 14568 14958 14596 15302
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14476 14074 14504 14350
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14464 12912 14516 12918
rect 14462 12880 14464 12889
rect 14516 12880 14518 12889
rect 14462 12815 14518 12824
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11762 14504 12038
rect 14568 11898 14596 12582
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14476 10130 14504 11698
rect 14554 11656 14610 11665
rect 14660 11626 14688 15830
rect 15028 15570 15056 16662
rect 15304 16658 15332 17088
rect 15106 16623 15162 16632
rect 15292 16652 15344 16658
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15028 15162 15056 15506
rect 15120 15314 15148 16623
rect 15292 16594 15344 16600
rect 15304 16046 15332 16594
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15212 15473 15240 15846
rect 15198 15464 15254 15473
rect 15198 15399 15254 15408
rect 15120 15286 15240 15314
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14752 14278 14780 14962
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 12753 14780 14214
rect 14738 12744 14794 12753
rect 14738 12679 14794 12688
rect 14738 12336 14794 12345
rect 14738 12271 14794 12280
rect 14554 11591 14610 11600
rect 14648 11620 14700 11626
rect 14568 11558 14596 11591
rect 14648 11562 14700 11568
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14752 11370 14780 12271
rect 14568 11342 14780 11370
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14372 9104 14424 9110
rect 14464 9104 14516 9110
rect 14372 9046 14424 9052
rect 14462 9072 14464 9081
rect 14516 9072 14518 9081
rect 14384 8090 14412 9046
rect 14462 9007 14518 9016
rect 14568 8514 14596 11342
rect 14646 11112 14702 11121
rect 14646 11047 14648 11056
rect 14700 11047 14702 11056
rect 14648 11018 14700 11024
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14660 10198 14688 10406
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14568 8486 14688 8514
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14476 7313 14504 7414
rect 14462 7304 14518 7313
rect 14462 7239 14518 7248
rect 14370 7032 14426 7041
rect 14370 6967 14426 6976
rect 14384 6254 14412 6967
rect 14200 6174 14320 6202
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 14016 3641 14044 4082
rect 14002 3632 14058 3641
rect 14002 3567 14058 3576
rect 14200 3210 14228 6174
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5778 14320 6054
rect 14384 5896 14412 6190
rect 14464 5908 14516 5914
rect 14384 5868 14464 5896
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14292 5166 14320 5714
rect 14384 5370 14412 5868
rect 14464 5850 14516 5856
rect 14568 5778 14596 8298
rect 14660 7857 14688 8486
rect 14844 8129 14872 14758
rect 15212 14634 15240 15286
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15120 14606 15240 14634
rect 15120 14278 15148 14606
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15106 13968 15162 13977
rect 15106 13903 15162 13912
rect 15120 13870 15148 13903
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14936 12850 14964 13398
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 15028 11801 15056 13126
rect 15120 12850 15148 13330
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15212 12442 15240 14486
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15014 11792 15070 11801
rect 15014 11727 15070 11736
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14936 10606 14964 11494
rect 15028 11082 15056 11562
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15016 10532 15068 10538
rect 15016 10474 15068 10480
rect 15028 10441 15056 10474
rect 15014 10432 15070 10441
rect 15014 10367 15070 10376
rect 15120 10146 15148 11698
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15212 11257 15240 11630
rect 15198 11248 15254 11257
rect 15198 11183 15254 11192
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15028 10118 15148 10146
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9081 14964 9862
rect 15028 9722 15056 10118
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 15120 9654 15148 9862
rect 15108 9648 15160 9654
rect 15108 9590 15160 9596
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14922 9072 14978 9081
rect 14922 9007 14978 9016
rect 14830 8120 14886 8129
rect 14830 8055 14886 8064
rect 14646 7848 14702 7857
rect 14646 7783 14702 7792
rect 14844 7426 14872 8055
rect 14660 7398 14872 7426
rect 14936 7410 14964 9007
rect 15028 8430 15056 9318
rect 15120 8838 15148 9386
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 14924 7404 14976 7410
rect 14660 6186 14688 7398
rect 14924 7346 14976 7352
rect 15120 7342 15148 8570
rect 15212 7546 15240 11018
rect 15304 10266 15332 15098
rect 15396 12374 15424 18022
rect 15488 15162 15516 21422
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15580 17649 15608 21286
rect 15672 18873 15700 23920
rect 16960 21962 16988 23920
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 15750 21244 16046 21264
rect 15806 21242 15830 21244
rect 15886 21242 15910 21244
rect 15966 21242 15990 21244
rect 15828 21190 15830 21242
rect 15892 21190 15904 21242
rect 15966 21190 15968 21242
rect 15806 21188 15830 21190
rect 15886 21188 15910 21190
rect 15966 21188 15990 21190
rect 15750 21168 16046 21188
rect 15750 20156 16046 20176
rect 15806 20154 15830 20156
rect 15886 20154 15910 20156
rect 15966 20154 15990 20156
rect 15828 20102 15830 20154
rect 15892 20102 15904 20154
rect 15966 20102 15968 20154
rect 15806 20100 15830 20102
rect 15886 20100 15910 20102
rect 15966 20100 15990 20102
rect 15750 20080 16046 20100
rect 15750 19408 15806 19417
rect 16132 19378 16160 21490
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16224 20398 16252 21286
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 16224 19961 16252 20334
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16316 19990 16344 20198
rect 16304 19984 16356 19990
rect 16210 19952 16266 19961
rect 16304 19926 16356 19932
rect 16210 19887 16266 19896
rect 15750 19343 15752 19352
rect 15804 19343 15806 19352
rect 16120 19372 16172 19378
rect 15752 19314 15804 19320
rect 16120 19314 16172 19320
rect 15750 19068 16046 19088
rect 15806 19066 15830 19068
rect 15886 19066 15910 19068
rect 15966 19066 15990 19068
rect 15828 19014 15830 19066
rect 15892 19014 15904 19066
rect 15966 19014 15968 19066
rect 15806 19012 15830 19014
rect 15886 19012 15910 19014
rect 15966 19012 15990 19014
rect 15750 18992 16046 19012
rect 15658 18864 15714 18873
rect 15658 18799 15714 18808
rect 16132 18465 16160 19314
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16118 18456 16174 18465
rect 16118 18391 16174 18400
rect 15934 18320 15990 18329
rect 15934 18255 15990 18264
rect 16118 18320 16174 18329
rect 16118 18255 16174 18264
rect 16212 18284 16264 18290
rect 15948 18222 15976 18255
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15752 18148 15804 18154
rect 15672 18108 15752 18136
rect 15672 17882 15700 18108
rect 15752 18090 15804 18096
rect 15750 17980 16046 18000
rect 15806 17978 15830 17980
rect 15886 17978 15910 17980
rect 15966 17978 15990 17980
rect 15828 17926 15830 17978
rect 15892 17926 15904 17978
rect 15966 17926 15968 17978
rect 15806 17924 15830 17926
rect 15886 17924 15910 17926
rect 15966 17924 15990 17926
rect 15750 17904 16046 17924
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 16132 17814 16160 18255
rect 16212 18226 16264 18232
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 15566 17640 15622 17649
rect 15566 17575 15622 17584
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17066 15608 17478
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15488 12306 15516 14758
rect 15580 14006 15608 17002
rect 16224 16998 16252 18226
rect 16316 18154 16344 19110
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16408 18086 16436 21626
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16580 21548 16632 21554
rect 16580 21490 16632 21496
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16500 19786 16528 21082
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16500 18834 16528 19722
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 15750 16892 16046 16912
rect 15806 16890 15830 16892
rect 15886 16890 15910 16892
rect 15966 16890 15990 16892
rect 15828 16838 15830 16890
rect 15892 16838 15904 16890
rect 15966 16838 15968 16890
rect 15806 16836 15830 16838
rect 15886 16836 15910 16838
rect 15966 16836 15990 16838
rect 15750 16816 16046 16836
rect 16316 16794 16344 17546
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 15658 16008 15714 16017
rect 15658 15943 15714 15952
rect 15672 15570 15700 15943
rect 15750 15804 16046 15824
rect 15806 15802 15830 15804
rect 15886 15802 15910 15804
rect 15966 15802 15990 15804
rect 15828 15750 15830 15802
rect 15892 15750 15904 15802
rect 15966 15750 15968 15802
rect 15806 15748 15830 15750
rect 15886 15748 15910 15750
rect 15966 15748 15990 15750
rect 15750 15728 16046 15748
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15752 15496 15804 15502
rect 16028 15496 16080 15502
rect 15752 15438 15804 15444
rect 16026 15464 16028 15473
rect 16080 15464 16082 15473
rect 15764 15065 15792 15438
rect 16026 15399 16082 15408
rect 15750 15056 15806 15065
rect 15750 14991 15806 15000
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16302 14920 16358 14929
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15672 13841 15700 14758
rect 15750 14716 16046 14736
rect 15806 14714 15830 14716
rect 15886 14714 15910 14716
rect 15966 14714 15990 14716
rect 15828 14662 15830 14714
rect 15892 14662 15904 14714
rect 15966 14662 15968 14714
rect 15806 14660 15830 14662
rect 15886 14660 15910 14662
rect 15966 14660 15990 14662
rect 15750 14640 16046 14660
rect 15750 14512 15806 14521
rect 15750 14447 15752 14456
rect 15804 14447 15806 14456
rect 15752 14418 15804 14424
rect 16120 14272 16172 14278
rect 16118 14240 16120 14249
rect 16172 14240 16174 14249
rect 16118 14175 16174 14184
rect 16132 14074 16160 14175
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 14000 16080 14006
rect 16080 13948 16160 13954
rect 16028 13942 16160 13948
rect 16040 13926 16160 13942
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15750 13628 16046 13648
rect 15806 13626 15830 13628
rect 15886 13626 15910 13628
rect 15966 13626 15990 13628
rect 15828 13574 15830 13626
rect 15892 13574 15904 13626
rect 15966 13574 15968 13626
rect 15806 13572 15830 13574
rect 15886 13572 15910 13574
rect 15966 13572 15990 13574
rect 15750 13552 16046 13572
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15580 12714 15608 13126
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15580 12617 15608 12650
rect 15566 12608 15622 12617
rect 15566 12543 15622 12552
rect 15750 12540 16046 12560
rect 15806 12538 15830 12540
rect 15886 12538 15910 12540
rect 15966 12538 15990 12540
rect 15828 12486 15830 12538
rect 15892 12486 15904 12538
rect 15966 12486 15968 12538
rect 15806 12484 15830 12486
rect 15886 12484 15910 12486
rect 15966 12484 15990 12486
rect 15750 12464 16046 12484
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9518 15332 9930
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15304 8430 15332 8774
rect 15396 8634 15424 12174
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15488 8022 15516 12038
rect 15580 11354 15608 12310
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15658 11928 15714 11937
rect 15658 11863 15660 11872
rect 15712 11863 15714 11872
rect 15660 11834 15712 11840
rect 15764 11665 15792 12242
rect 15844 11824 15896 11830
rect 16028 11824 16080 11830
rect 15896 11784 16028 11812
rect 15844 11766 15896 11772
rect 16028 11766 16080 11772
rect 15750 11656 15806 11665
rect 15672 11614 15750 11642
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 10169 15608 11154
rect 15566 10160 15622 10169
rect 15566 10095 15622 10104
rect 15566 9344 15622 9353
rect 15566 9279 15622 9288
rect 15580 8838 15608 9279
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15566 8528 15622 8537
rect 15566 8463 15568 8472
rect 15620 8463 15622 8472
rect 15568 8434 15620 8440
rect 15476 8016 15528 8022
rect 15476 7958 15528 7964
rect 15672 7954 15700 11614
rect 15750 11591 15806 11600
rect 15750 11452 16046 11472
rect 15806 11450 15830 11452
rect 15886 11450 15910 11452
rect 15966 11450 15990 11452
rect 15828 11398 15830 11450
rect 15892 11398 15904 11450
rect 15966 11398 15968 11450
rect 15806 11396 15830 11398
rect 15886 11396 15910 11398
rect 15966 11396 15990 11398
rect 15750 11376 16046 11396
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10849 15976 10950
rect 15934 10840 15990 10849
rect 15934 10775 15990 10784
rect 15948 10674 15976 10775
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15750 10364 16046 10384
rect 15806 10362 15830 10364
rect 15886 10362 15910 10364
rect 15966 10362 15990 10364
rect 15828 10310 15830 10362
rect 15892 10310 15904 10362
rect 15966 10310 15968 10362
rect 15806 10308 15830 10310
rect 15886 10308 15910 10310
rect 15966 10308 15990 10310
rect 15750 10288 16046 10308
rect 15750 9276 16046 9296
rect 15806 9274 15830 9276
rect 15886 9274 15910 9276
rect 15966 9274 15990 9276
rect 15828 9222 15830 9274
rect 15892 9222 15904 9274
rect 15966 9222 15968 9274
rect 15806 9220 15830 9222
rect 15886 9220 15910 9222
rect 15966 9220 15990 9222
rect 15750 9200 16046 9220
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15856 8634 15884 8978
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15750 8188 16046 8208
rect 15806 8186 15830 8188
rect 15886 8186 15910 8188
rect 15966 8186 15990 8188
rect 15828 8134 15830 8186
rect 15892 8134 15904 8186
rect 15966 8134 15968 8186
rect 15806 8132 15830 8134
rect 15886 8132 15910 8134
rect 15966 8132 15990 8134
rect 15750 8112 16046 8132
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 16132 7698 16160 13926
rect 16224 11665 16252 14894
rect 16302 14855 16304 14864
rect 16356 14855 16358 14864
rect 16304 14826 16356 14832
rect 16408 14770 16436 18022
rect 16592 17270 16620 21490
rect 16776 20466 16804 21558
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16500 15978 16528 16730
rect 16592 16658 16620 17206
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16684 15201 16712 19110
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16776 18329 16804 18566
rect 16762 18320 16818 18329
rect 16762 18255 16818 18264
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16776 17218 16804 18090
rect 16868 17882 16896 21286
rect 16960 20777 16988 21286
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 16946 20768 17002 20777
rect 16946 20703 17002 20712
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 16776 17190 16896 17218
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16776 16046 16804 17002
rect 16868 16561 16896 17190
rect 16854 16552 16910 16561
rect 16854 16487 16910 16496
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16776 15366 16804 15846
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16670 15192 16726 15201
rect 16670 15127 16726 15136
rect 16316 14742 16436 14770
rect 16210 11656 16266 11665
rect 16210 11591 16266 11600
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 10606 16252 11494
rect 16316 11286 16344 14742
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16500 12170 16528 14418
rect 16868 14414 16896 15370
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16592 13530 16620 14350
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16776 13190 16804 13670
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16868 12986 16896 13330
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16764 12640 16816 12646
rect 16762 12608 16764 12617
rect 16816 12608 16818 12617
rect 16762 12543 16818 12552
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16408 11665 16436 11698
rect 16394 11656 16450 11665
rect 16394 11591 16450 11600
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16302 11112 16358 11121
rect 16302 11047 16358 11056
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16224 10266 16252 10542
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16316 10146 16344 11047
rect 16408 10198 16436 11494
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16500 10606 16528 11154
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16486 10432 16542 10441
rect 16486 10367 16542 10376
rect 16224 10118 16344 10146
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16224 9926 16252 10118
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16408 9654 16436 10134
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16210 9208 16266 9217
rect 16210 9143 16266 9152
rect 15396 7670 16160 7698
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4282 14320 4422
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14384 4146 14412 5306
rect 14476 5098 14504 5646
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14476 4622 14504 5034
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14646 4584 14702 4593
rect 14646 4519 14702 4528
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14462 4312 14518 4321
rect 14462 4247 14518 4256
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14108 3182 14228 3210
rect 14278 3224 14334 3233
rect 14108 3126 14136 3182
rect 14278 3159 14334 3168
rect 14292 3126 14320 3159
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14384 2961 14412 3334
rect 14370 2952 14426 2961
rect 14370 2887 14426 2896
rect 13688 2808 13952 2836
rect 13636 2790 13688 2796
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 8574 2408 8630 2417
rect 8574 2343 8630 2352
rect 8588 480 8616 2343
rect 11992 2088 12020 2790
rect 13358 2680 13414 2689
rect 13358 2615 13360 2624
rect 13412 2615 13414 2624
rect 13360 2586 13412 2592
rect 14476 2310 14504 4247
rect 14568 3720 14596 4422
rect 14660 3942 14688 4519
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14752 3754 14780 7278
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14844 5370 14872 6802
rect 14936 6662 14964 7210
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15198 7168 15254 7177
rect 15120 6866 15148 7142
rect 15198 7103 15254 7112
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14844 4826 14872 5306
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14936 4758 14964 6598
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14924 4616 14976 4622
rect 15028 4604 15056 4966
rect 15212 4729 15240 7103
rect 15290 6216 15346 6225
rect 15290 6151 15346 6160
rect 15198 4720 15254 4729
rect 15198 4655 15254 4664
rect 14976 4576 15056 4604
rect 15200 4616 15252 4622
rect 14924 4558 14976 4564
rect 15200 4558 15252 4564
rect 14936 4010 14964 4558
rect 15014 4448 15070 4457
rect 15014 4383 15070 4392
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14752 3726 14872 3754
rect 14568 3692 14688 3720
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14568 3505 14596 3538
rect 14660 3516 14688 3692
rect 14844 3534 14872 3726
rect 15028 3602 15056 4383
rect 15212 4078 15240 4558
rect 15304 4486 15332 6151
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14740 3528 14792 3534
rect 14554 3496 14610 3505
rect 14660 3488 14740 3516
rect 14740 3470 14792 3476
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14554 3431 14610 3440
rect 15120 3194 15148 3946
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15016 3120 15068 3126
rect 14738 3088 14794 3097
rect 15016 3062 15068 3068
rect 14738 3023 14740 3032
rect 14792 3023 14794 3032
rect 14740 2994 14792 3000
rect 15028 2446 15056 3062
rect 15304 2582 15332 4014
rect 15396 3058 15424 7670
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 15750 7100 16046 7120
rect 15806 7098 15830 7100
rect 15886 7098 15910 7100
rect 15966 7098 15990 7100
rect 15828 7046 15830 7098
rect 15892 7046 15904 7098
rect 15966 7046 15968 7098
rect 15806 7044 15830 7046
rect 15886 7044 15910 7046
rect 15966 7044 15990 7046
rect 15750 7024 16046 7044
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15672 6322 15700 6734
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15566 6080 15622 6089
rect 15488 5098 15516 6054
rect 15566 6015 15622 6024
rect 15580 5574 15608 6015
rect 15568 5568 15620 5574
rect 15672 5545 15700 6258
rect 15750 6012 16046 6032
rect 15806 6010 15830 6012
rect 15886 6010 15910 6012
rect 15966 6010 15990 6012
rect 15828 5958 15830 6010
rect 15892 5958 15904 6010
rect 15966 5958 15968 6010
rect 15806 5956 15830 5958
rect 15886 5956 15910 5958
rect 15966 5956 15990 5958
rect 15750 5936 16046 5956
rect 15568 5510 15620 5516
rect 15658 5536 15714 5545
rect 15658 5471 15714 5480
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15568 5092 15620 5098
rect 15568 5034 15620 5040
rect 15474 4720 15530 4729
rect 15474 4655 15530 4664
rect 15488 3194 15516 4655
rect 15580 4554 15608 5034
rect 15672 4690 15700 5471
rect 15750 4924 16046 4944
rect 15806 4922 15830 4924
rect 15886 4922 15910 4924
rect 15966 4922 15990 4924
rect 15828 4870 15830 4922
rect 15892 4870 15904 4922
rect 15966 4870 15968 4922
rect 15806 4868 15830 4870
rect 15886 4868 15910 4870
rect 15966 4868 15990 4870
rect 15750 4848 16046 4868
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15672 4146 15700 4626
rect 15752 4480 15804 4486
rect 15750 4448 15752 4457
rect 15804 4448 15806 4457
rect 15750 4383 15806 4392
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15566 4040 15622 4049
rect 15856 4026 15884 4626
rect 15566 3975 15622 3984
rect 15672 3998 15884 4026
rect 15580 3942 15608 3975
rect 15672 3942 15700 3998
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 14464 2304 14516 2310
rect 15028 2281 15056 2382
rect 14464 2246 14516 2252
rect 15014 2272 15070 2281
rect 12052 2204 12348 2224
rect 15014 2207 15070 2216
rect 12108 2202 12132 2204
rect 12188 2202 12212 2204
rect 12268 2202 12292 2204
rect 12130 2150 12132 2202
rect 12194 2150 12206 2202
rect 12268 2150 12270 2202
rect 12108 2148 12132 2150
rect 12188 2148 12212 2150
rect 12268 2148 12292 2150
rect 12052 2128 12348 2148
rect 11992 2060 12112 2088
rect 12084 480 12112 2060
rect 15580 480 15608 3334
rect 15672 2650 15700 3878
rect 15750 3836 16046 3856
rect 15806 3834 15830 3836
rect 15886 3834 15910 3836
rect 15966 3834 15990 3836
rect 15828 3782 15830 3834
rect 15892 3782 15904 3834
rect 15966 3782 15968 3834
rect 15806 3780 15830 3782
rect 15886 3780 15910 3782
rect 15966 3780 15990 3782
rect 15750 3760 16046 3780
rect 16132 3738 16160 7346
rect 16224 4826 16252 9143
rect 16316 9110 16344 9522
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16408 9042 16436 9386
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8401 16344 8910
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16302 8392 16358 8401
rect 16302 8327 16358 8336
rect 16408 7154 16436 8774
rect 16500 8022 16528 10367
rect 16592 10282 16620 11222
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16684 10441 16712 11086
rect 16670 10432 16726 10441
rect 16670 10367 16726 10376
rect 16592 10254 16712 10282
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16592 9722 16620 10134
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16592 9217 16620 9386
rect 16578 9208 16634 9217
rect 16578 9143 16634 9152
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16592 7886 16620 8978
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16316 7126 16436 7154
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16316 4457 16344 7126
rect 16394 6352 16450 6361
rect 16394 6287 16450 6296
rect 16302 4448 16358 4457
rect 16302 4383 16358 4392
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 15750 3632 15806 3641
rect 15934 3632 15990 3641
rect 15806 3590 15884 3618
rect 15750 3567 15806 3576
rect 15856 3126 15884 3590
rect 16224 3618 16252 4218
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 15934 3567 15936 3576
rect 15988 3567 15990 3576
rect 16040 3590 16252 3618
rect 15936 3538 15988 3544
rect 15844 3120 15896 3126
rect 15750 3088 15806 3097
rect 15844 3062 15896 3068
rect 16040 3058 16068 3590
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 15750 3023 15806 3032
rect 16028 3052 16080 3058
rect 15764 2990 15792 3023
rect 16028 2994 16080 3000
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 15750 2748 16046 2768
rect 15806 2746 15830 2748
rect 15886 2746 15910 2748
rect 15966 2746 15990 2748
rect 15828 2694 15830 2746
rect 15892 2694 15904 2746
rect 15966 2694 15968 2746
rect 15806 2692 15830 2694
rect 15886 2692 15910 2694
rect 15966 2692 15990 2694
rect 15750 2672 16046 2692
rect 16132 2666 16160 3402
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 16224 2825 16252 3062
rect 16316 3058 16344 4082
rect 16408 3466 16436 6287
rect 16684 5794 16712 10254
rect 16776 6905 16804 11494
rect 16762 6896 16818 6905
rect 16762 6831 16818 6840
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16592 5766 16712 5794
rect 16500 3602 16528 5714
rect 16592 4185 16620 5766
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16684 4758 16712 5646
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 5370 16804 5510
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16578 4176 16634 4185
rect 16578 4111 16634 4120
rect 16580 3936 16632 3942
rect 16684 3913 16712 4422
rect 16580 3878 16632 3884
rect 16670 3904 16726 3913
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16592 2990 16620 3878
rect 16670 3839 16726 3848
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16396 2848 16448 2854
rect 16210 2816 16266 2825
rect 16776 2836 16804 5170
rect 16396 2790 16448 2796
rect 16592 2808 16804 2836
rect 16210 2751 16266 2760
rect 16408 2666 16436 2790
rect 15660 2644 15712 2650
rect 16132 2638 16436 2666
rect 15660 2586 15712 2592
rect 15658 2544 15714 2553
rect 15658 2479 15660 2488
rect 15712 2479 15714 2488
rect 16304 2508 16356 2514
rect 15660 2450 15712 2456
rect 16304 2450 16356 2456
rect 16316 2106 16344 2450
rect 16592 2310 16620 2808
rect 16764 2440 16816 2446
rect 16868 2428 16896 12922
rect 16960 10130 16988 20470
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17144 19446 17172 20402
rect 17132 19440 17184 19446
rect 17132 19382 17184 19388
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17052 11286 17080 19246
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17144 17270 17172 18022
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17222 17232 17278 17241
rect 17222 17167 17278 17176
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17144 16250 17172 16934
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17144 11642 17172 15302
rect 17236 12646 17264 17167
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17144 11614 17264 11642
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17040 11280 17092 11286
rect 17040 11222 17092 11228
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10810 17080 10950
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16948 9648 17000 9654
rect 16946 9616 16948 9625
rect 17000 9616 17002 9625
rect 16946 9551 17002 9560
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16960 9353 16988 9454
rect 16946 9344 17002 9353
rect 16946 9279 17002 9288
rect 17052 9194 17080 10610
rect 17144 10470 17172 11494
rect 17236 10674 17264 11614
rect 17328 10826 17356 20946
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17420 18193 17448 19654
rect 17512 19310 17540 19790
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17512 18834 17540 19246
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17406 18184 17462 18193
rect 17406 18119 17462 18128
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17420 16590 17448 17614
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17512 16454 17540 18226
rect 17604 17814 17632 23920
rect 18248 23066 18276 23920
rect 18156 23038 18276 23066
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 18064 20398 18092 21014
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17696 18329 17724 19110
rect 17880 18970 17908 19110
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17972 18358 18000 20198
rect 18064 19310 18092 20334
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17960 18352 18012 18358
rect 17682 18320 17738 18329
rect 17960 18294 18012 18300
rect 18064 18290 18092 19246
rect 17682 18255 17738 18264
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17406 15056 17462 15065
rect 17406 14991 17408 15000
rect 17460 14991 17462 15000
rect 17408 14962 17460 14968
rect 17406 14512 17462 14521
rect 17406 14447 17462 14456
rect 17420 14346 17448 14447
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17420 12850 17448 13466
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17420 11354 17448 12310
rect 17512 11762 17540 15846
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 17500 11008 17552 11014
rect 17498 10976 17500 10985
rect 17552 10976 17554 10985
rect 17498 10911 17554 10920
rect 17328 10810 17448 10826
rect 17328 10804 17460 10810
rect 17328 10798 17408 10804
rect 17408 10746 17460 10752
rect 17604 10690 17632 16730
rect 17696 16726 17724 18158
rect 18064 18086 18092 18226
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17882 18092 18022
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 17696 15094 17724 16662
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17880 15570 17908 15982
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17696 14414 17724 14758
rect 17774 14648 17830 14657
rect 17774 14583 17830 14592
rect 17788 14550 17816 14583
rect 17776 14544 17828 14550
rect 17776 14486 17828 14492
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17776 14408 17828 14414
rect 17880 14396 17908 15506
rect 17828 14368 17908 14396
rect 17776 14350 17828 14356
rect 17880 13938 17908 14368
rect 17868 13932 17920 13938
rect 17788 13892 17868 13920
rect 17788 13394 17816 13892
rect 17868 13874 17920 13880
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17776 13252 17828 13258
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17420 10662 17632 10690
rect 17696 13212 17776 13240
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 10282 17264 10406
rect 16960 9166 17080 9194
rect 17144 10254 17264 10282
rect 16960 7546 16988 9166
rect 17144 9081 17172 10254
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17236 9178 17264 9862
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17130 9072 17186 9081
rect 17328 9042 17356 9318
rect 17130 9007 17186 9016
rect 17316 9036 17368 9042
rect 17144 8838 17172 9007
rect 17316 8978 17368 8984
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17328 8650 17356 8978
rect 17236 8622 17356 8650
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 7886 17172 8230
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17236 7750 17264 8622
rect 17420 8514 17448 10662
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17512 10062 17540 10542
rect 17590 10432 17646 10441
rect 17590 10367 17646 10376
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17604 9466 17632 10367
rect 17512 9438 17632 9466
rect 17512 9058 17540 9438
rect 17512 9030 17632 9058
rect 17328 8486 17448 8514
rect 17328 7993 17356 8486
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17420 8090 17448 8366
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17512 8265 17540 8298
rect 17498 8256 17554 8265
rect 17498 8191 17554 8200
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17314 7984 17370 7993
rect 17314 7919 17370 7928
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16960 7342 16988 7482
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16960 6361 16988 6598
rect 16946 6352 17002 6361
rect 16946 6287 17002 6296
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16946 6080 17002 6089
rect 16946 6015 17002 6024
rect 16960 5710 16988 6015
rect 17052 5778 17080 6258
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 17144 5710 17172 6054
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17144 5545 17172 5646
rect 17130 5536 17186 5545
rect 17052 5494 17130 5522
rect 16946 5264 17002 5273
rect 16946 5199 17002 5208
rect 16960 4826 16988 5199
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16960 4078 16988 4422
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16946 3768 17002 3777
rect 16946 3703 17002 3712
rect 16960 3505 16988 3703
rect 17052 3534 17080 5494
rect 17130 5471 17186 5480
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4321 17172 4966
rect 17130 4312 17186 4321
rect 17130 4247 17186 4256
rect 17236 3738 17264 6734
rect 17420 6390 17448 6802
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 17512 6118 17540 6734
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17040 3528 17092 3534
rect 16946 3496 17002 3505
rect 17040 3470 17092 3476
rect 16946 3431 17002 3440
rect 17052 2922 17080 3470
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 16816 2400 16896 2428
rect 16764 2382 16816 2388
rect 16580 2304 16632 2310
rect 16960 2281 16988 2450
rect 16580 2246 16632 2252
rect 16946 2272 17002 2281
rect 16946 2207 17002 2216
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 17328 1358 17356 5306
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17420 4146 17448 5170
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17420 3194 17448 3606
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17420 2650 17448 2994
rect 17604 2990 17632 9030
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17696 2530 17724 13212
rect 17880 13240 17908 13738
rect 17828 13212 17908 13240
rect 17776 13194 17828 13200
rect 17866 13016 17922 13025
rect 17866 12951 17922 12960
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17788 11762 17816 12650
rect 17880 12374 17908 12951
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11150 17908 11630
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10305 17908 11086
rect 17866 10296 17922 10305
rect 17866 10231 17922 10240
rect 17866 10160 17922 10169
rect 17776 10124 17828 10130
rect 17866 10095 17922 10104
rect 17776 10066 17828 10072
rect 17788 8430 17816 10066
rect 17880 9489 17908 10095
rect 17866 9480 17922 9489
rect 17866 9415 17922 9424
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17880 9178 17908 9318
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17880 8022 17908 8774
rect 17972 8498 18000 17206
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 15570 18092 16390
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 18156 14958 18184 23038
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18340 21486 18368 21830
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18248 21078 18276 21422
rect 18236 21072 18288 21078
rect 18236 21014 18288 21020
rect 18800 20942 18828 21422
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18788 19848 18840 19854
rect 18786 19816 18788 19825
rect 18840 19816 18842 19825
rect 18786 19751 18842 19760
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18800 18970 18828 19178
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18052 14476 18104 14482
rect 18104 14436 18184 14464
rect 18052 14418 18104 14424
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 18064 12782 18092 13670
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18050 12336 18106 12345
rect 18050 12271 18106 12280
rect 18064 11642 18092 12271
rect 18156 12102 18184 14436
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18064 11614 18184 11642
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 10674 18092 11494
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18052 10464 18104 10470
rect 18050 10432 18052 10441
rect 18104 10432 18106 10441
rect 18050 10367 18106 10376
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18064 8362 18092 9998
rect 18156 9722 18184 11614
rect 18248 11257 18276 16934
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18328 15088 18380 15094
rect 18328 15030 18380 15036
rect 18340 14793 18368 15030
rect 18326 14784 18382 14793
rect 18326 14719 18382 14728
rect 18326 14648 18382 14657
rect 18326 14583 18382 14592
rect 18340 14550 18368 14583
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18432 14278 18460 16390
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18340 12782 18368 13738
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18234 11248 18290 11257
rect 18234 11183 18290 11192
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18248 11014 18276 11086
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18234 10840 18290 10849
rect 18234 10775 18290 10784
rect 18248 10742 18276 10775
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18248 10130 18276 10678
rect 18340 10606 18368 12378
rect 18432 12374 18460 12582
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18524 12322 18552 16934
rect 18616 12481 18644 18566
rect 18708 16153 18736 18634
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 18800 17882 18828 18090
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18892 17270 18920 23920
rect 19246 23352 19302 23361
rect 19246 23287 19302 23296
rect 19154 22672 19210 22681
rect 19154 22607 19210 22616
rect 19168 21146 19196 22607
rect 19260 21690 19288 23287
rect 19536 21978 19564 23920
rect 20180 22522 20208 23920
rect 20088 22494 20208 22522
rect 19890 21992 19946 22001
rect 19536 21950 19840 21978
rect 19449 21788 19745 21808
rect 19505 21786 19529 21788
rect 19585 21786 19609 21788
rect 19665 21786 19689 21788
rect 19527 21734 19529 21786
rect 19591 21734 19603 21786
rect 19665 21734 19667 21786
rect 19505 21732 19529 21734
rect 19585 21732 19609 21734
rect 19665 21732 19689 21734
rect 19449 21712 19745 21732
rect 19248 21684 19300 21690
rect 19248 21626 19300 21632
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19246 21312 19302 21321
rect 19246 21247 19302 21256
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 19168 20534 19196 20878
rect 19260 20602 19288 21247
rect 19352 20806 19380 21354
rect 19812 21128 19840 21950
rect 19890 21927 19946 21936
rect 19904 21486 19932 21927
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19812 21100 19932 21128
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19449 20700 19745 20720
rect 19505 20698 19529 20700
rect 19585 20698 19609 20700
rect 19665 20698 19689 20700
rect 19527 20646 19529 20698
rect 19591 20646 19603 20698
rect 19665 20646 19667 20698
rect 19505 20644 19529 20646
rect 19585 20644 19609 20646
rect 19665 20644 19689 20646
rect 19449 20624 19745 20644
rect 19812 20602 19840 20946
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19156 20528 19208 20534
rect 19076 20476 19156 20482
rect 19076 20470 19208 20476
rect 19076 20454 19196 20470
rect 19432 20460 19484 20466
rect 19076 19310 19104 20454
rect 19432 20402 19484 20408
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19168 20058 19196 20266
rect 19246 20088 19302 20097
rect 19156 20052 19208 20058
rect 19246 20023 19302 20032
rect 19156 19994 19208 20000
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19168 18290 19196 19110
rect 19260 18426 19288 20023
rect 19444 19990 19472 20402
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19514 19380 19858
rect 19720 19825 19748 20198
rect 19812 19990 19840 20538
rect 19904 20466 19932 21100
rect 19982 20632 20038 20641
rect 19982 20567 20038 20576
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19996 20330 20024 20567
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19800 19984 19852 19990
rect 19800 19926 19852 19932
rect 19892 19848 19944 19854
rect 19706 19816 19762 19825
rect 19944 19796 20024 19802
rect 19892 19790 20024 19796
rect 19904 19774 20024 19790
rect 19706 19751 19762 19760
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19449 19612 19745 19632
rect 19505 19610 19529 19612
rect 19585 19610 19609 19612
rect 19665 19610 19689 19612
rect 19527 19558 19529 19610
rect 19591 19558 19603 19610
rect 19665 19558 19667 19610
rect 19505 19556 19529 19558
rect 19585 19556 19609 19558
rect 19665 19556 19689 19558
rect 19449 19536 19745 19556
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19352 19394 19380 19450
rect 19904 19417 19932 19654
rect 19890 19408 19946 19417
rect 19352 19366 19564 19394
rect 19536 18834 19564 19366
rect 19800 19372 19852 19378
rect 19890 19343 19946 19352
rect 19800 19314 19852 19320
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18426 19380 18702
rect 19449 18524 19745 18544
rect 19505 18522 19529 18524
rect 19585 18522 19609 18524
rect 19665 18522 19689 18524
rect 19527 18470 19529 18522
rect 19591 18470 19603 18522
rect 19665 18470 19667 18522
rect 19505 18468 19529 18470
rect 19585 18468 19609 18470
rect 19665 18468 19689 18470
rect 19449 18448 19745 18468
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19352 17814 19380 18362
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 18972 17740 19024 17746
rect 18972 17682 19024 17688
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18984 17134 19012 17682
rect 19064 17536 19116 17542
rect 19444 17524 19472 18226
rect 19812 17610 19840 19314
rect 19996 18850 20024 19774
rect 20088 19446 20116 22494
rect 20364 21418 20392 23967
rect 20810 23920 20866 24400
rect 21454 23920 21510 24400
rect 22098 23920 22154 24400
rect 22742 23920 22798 24400
rect 23386 23920 23442 24400
rect 24030 23920 24086 24400
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 20352 21412 20404 21418
rect 20352 21354 20404 21360
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20272 21078 20300 21286
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20260 21072 20312 21078
rect 20260 21014 20312 21020
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20180 20466 20208 20742
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20272 20330 20300 21014
rect 20260 20324 20312 20330
rect 20260 20266 20312 20272
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20166 19272 20222 19281
rect 20166 19207 20168 19216
rect 20220 19207 20222 19216
rect 20168 19178 20220 19184
rect 19904 18822 20024 18850
rect 19904 18766 19932 18822
rect 19892 18760 19944 18766
rect 20272 18714 20300 19450
rect 19892 18702 19944 18708
rect 19904 17678 19932 18702
rect 20180 18686 20300 18714
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20088 18057 20116 18158
rect 20074 18048 20130 18057
rect 20074 17983 20130 17992
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19064 17478 19116 17484
rect 19352 17496 19472 17524
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18984 16794 19012 17070
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18788 16448 18840 16454
rect 18786 16416 18788 16425
rect 18840 16416 18842 16425
rect 18786 16351 18842 16360
rect 18694 16144 18750 16153
rect 18694 16079 18750 16088
rect 18970 16144 19026 16153
rect 18970 16079 19026 16088
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18708 14890 18736 15506
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18708 13025 18736 13806
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 18708 12782 18736 12951
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18602 12472 18658 12481
rect 18800 12458 18828 14894
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18892 13569 18920 14826
rect 18984 13734 19012 16079
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18878 13560 18934 13569
rect 18878 13495 18934 13504
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12646 18920 13126
rect 18984 12986 19012 13330
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18984 12714 19012 12922
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18800 12430 19012 12458
rect 18602 12407 18658 12416
rect 18524 12294 18644 12322
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18524 11762 18552 12106
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18328 10464 18380 10470
rect 18432 10441 18460 11086
rect 18524 11014 18552 11562
rect 18616 11014 18644 12294
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18708 11762 18736 12242
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11150 18736 11494
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18328 10406 18380 10412
rect 18418 10432 18474 10441
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18248 9654 18276 9862
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 9042 18184 9318
rect 18234 9208 18290 9217
rect 18234 9143 18290 9152
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18248 8974 18276 9143
rect 18236 8968 18288 8974
rect 18142 8936 18198 8945
rect 18236 8910 18288 8916
rect 18142 8871 18198 8880
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 5302 18000 7686
rect 18156 6474 18184 8871
rect 18248 7342 18276 8910
rect 18340 8090 18368 10406
rect 18418 10367 18474 10376
rect 18418 10296 18474 10305
rect 18418 10231 18474 10240
rect 18432 9450 18460 10231
rect 18524 9489 18552 10950
rect 18708 9722 18736 11086
rect 18800 10606 18828 12038
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18604 9512 18656 9518
rect 18510 9480 18566 9489
rect 18420 9444 18472 9450
rect 18604 9454 18656 9460
rect 18510 9415 18566 9424
rect 18420 9386 18472 9392
rect 18432 9217 18460 9386
rect 18418 9208 18474 9217
rect 18418 9143 18474 9152
rect 18524 8974 18552 9415
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18432 8401 18460 8502
rect 18418 8392 18474 8401
rect 18418 8327 18474 8336
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18156 6446 18276 6474
rect 18142 6352 18198 6361
rect 18142 6287 18198 6296
rect 18156 6254 18184 6287
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17604 2502 17724 2530
rect 17604 2378 17632 2502
rect 17788 2446 17816 4150
rect 18064 3942 18092 5850
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 4826 18184 5510
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18248 4049 18276 6446
rect 18432 6390 18460 7414
rect 18524 7206 18552 8910
rect 18616 8634 18644 9454
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18800 8498 18828 10066
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18432 5642 18460 6326
rect 18524 5914 18552 6802
rect 18708 6254 18736 7278
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18800 6390 18828 6734
rect 18892 6497 18920 11766
rect 18984 9625 19012 12430
rect 19076 11830 19104 17478
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19260 16658 19288 17002
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19352 16590 19380 17496
rect 19449 17436 19745 17456
rect 19505 17434 19529 17436
rect 19585 17434 19609 17436
rect 19665 17434 19689 17436
rect 19527 17382 19529 17434
rect 19591 17382 19603 17434
rect 19665 17382 19667 17434
rect 19505 17380 19529 17382
rect 19585 17380 19609 17382
rect 19665 17380 19689 17382
rect 19449 17360 19745 17380
rect 19904 17202 19932 17614
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19812 16794 19840 16934
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19444 16436 19472 16594
rect 19352 16408 19472 16436
rect 19352 15978 19380 16408
rect 19449 16348 19745 16368
rect 19505 16346 19529 16348
rect 19585 16346 19609 16348
rect 19665 16346 19689 16348
rect 19527 16294 19529 16346
rect 19591 16294 19603 16346
rect 19665 16294 19667 16346
rect 19505 16292 19529 16294
rect 19585 16292 19609 16294
rect 19665 16292 19689 16294
rect 19449 16272 19745 16292
rect 19708 16176 19760 16182
rect 19812 16130 19840 16730
rect 19904 16726 19932 17138
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19760 16124 19840 16130
rect 19708 16118 19840 16124
rect 19720 16102 19840 16118
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19168 14958 19196 15642
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19260 14498 19288 15846
rect 19352 15706 19380 15914
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19708 15632 19760 15638
rect 19708 15574 19760 15580
rect 19720 15473 19748 15574
rect 19706 15464 19762 15473
rect 19706 15399 19762 15408
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19449 15260 19745 15280
rect 19505 15258 19529 15260
rect 19585 15258 19609 15260
rect 19665 15258 19689 15260
rect 19527 15206 19529 15258
rect 19591 15206 19603 15258
rect 19665 15206 19667 15258
rect 19505 15204 19529 15206
rect 19585 15204 19609 15206
rect 19665 15204 19689 15206
rect 19449 15184 19745 15204
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19708 14952 19760 14958
rect 19812 14940 19840 15302
rect 19760 14929 19840 14940
rect 19760 14920 19854 14929
rect 19760 14912 19798 14920
rect 19708 14894 19760 14900
rect 19338 14784 19394 14793
rect 19338 14719 19394 14728
rect 19352 14618 19380 14719
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19260 14470 19380 14498
rect 19156 14408 19208 14414
rect 19352 14385 19380 14470
rect 19156 14350 19208 14356
rect 19338 14376 19394 14385
rect 19168 14074 19196 14350
rect 19248 14340 19300 14346
rect 19338 14311 19394 14320
rect 19248 14282 19300 14288
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 19168 11694 19196 13806
rect 19260 12442 19288 14282
rect 19340 14272 19392 14278
rect 19444 14260 19472 14894
rect 19798 14855 19854 14864
rect 19444 14232 19840 14260
rect 19340 14214 19392 14220
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19352 11898 19380 14214
rect 19449 14172 19745 14192
rect 19505 14170 19529 14172
rect 19585 14170 19609 14172
rect 19665 14170 19689 14172
rect 19527 14118 19529 14170
rect 19591 14118 19603 14170
rect 19665 14118 19667 14170
rect 19505 14116 19529 14118
rect 19585 14116 19609 14118
rect 19665 14116 19689 14118
rect 19449 14096 19745 14116
rect 19812 13870 19840 14232
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19720 13326 19748 13670
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19449 13084 19745 13104
rect 19505 13082 19529 13084
rect 19585 13082 19609 13084
rect 19665 13082 19689 13084
rect 19527 13030 19529 13082
rect 19591 13030 19603 13082
rect 19665 13030 19667 13082
rect 19505 13028 19529 13030
rect 19585 13028 19609 13030
rect 19665 13028 19689 13030
rect 19449 13008 19745 13028
rect 19708 12912 19760 12918
rect 19628 12872 19708 12900
rect 19628 12617 19656 12872
rect 19708 12854 19760 12860
rect 19708 12640 19760 12646
rect 19614 12608 19670 12617
rect 19708 12582 19760 12588
rect 19614 12543 19670 12552
rect 19720 12170 19748 12582
rect 19812 12322 19840 13330
rect 19904 12481 19932 16390
rect 19996 15026 20024 16934
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19982 14920 20038 14929
rect 19982 14855 20038 14864
rect 19996 13938 20024 14855
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19996 13734 20024 13874
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19890 12472 19946 12481
rect 19996 12442 20024 13466
rect 20088 12753 20116 17682
rect 20180 17241 20208 18686
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20166 17232 20222 17241
rect 20166 17167 20222 17176
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20074 12744 20130 12753
rect 20074 12679 20130 12688
rect 20074 12608 20130 12617
rect 20074 12543 20130 12552
rect 19890 12407 19946 12416
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20088 12322 20116 12543
rect 19812 12294 19932 12322
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19449 11996 19745 12016
rect 19505 11994 19529 11996
rect 19585 11994 19609 11996
rect 19665 11994 19689 11996
rect 19527 11942 19529 11994
rect 19591 11942 19603 11994
rect 19665 11942 19667 11994
rect 19505 11940 19529 11942
rect 19585 11940 19609 11942
rect 19665 11940 19689 11942
rect 19449 11920 19745 11940
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19812 11762 19840 12174
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19156 11688 19208 11694
rect 19628 11665 19656 11698
rect 19156 11630 19208 11636
rect 19614 11656 19670 11665
rect 19670 11614 19748 11642
rect 19614 11591 19670 11600
rect 19338 11520 19394 11529
rect 19338 11455 19394 11464
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18970 9616 19026 9625
rect 18970 9551 19026 9560
rect 18970 9344 19026 9353
rect 18970 9279 19026 9288
rect 18878 6488 18934 6497
rect 18878 6423 18934 6432
rect 18788 6384 18840 6390
rect 18984 6338 19012 9279
rect 19076 8430 19104 10678
rect 19168 9738 19196 10950
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19260 10062 19288 10678
rect 19352 10538 19380 11455
rect 19720 11098 19748 11614
rect 19812 11354 19840 11698
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19720 11070 19840 11098
rect 19449 10908 19745 10928
rect 19505 10906 19529 10908
rect 19585 10906 19609 10908
rect 19665 10906 19689 10908
rect 19527 10854 19529 10906
rect 19591 10854 19603 10906
rect 19665 10854 19667 10906
rect 19505 10852 19529 10854
rect 19585 10852 19609 10854
rect 19665 10852 19689 10854
rect 19449 10832 19745 10852
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19628 10130 19656 10406
rect 19812 10282 19840 11070
rect 19904 10713 19932 12294
rect 19996 12294 20116 12322
rect 19890 10704 19946 10713
rect 19890 10639 19946 10648
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19720 10254 19840 10282
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19248 10056 19300 10062
rect 19720 10033 19748 10254
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19248 9998 19300 10004
rect 19706 10024 19762 10033
rect 19706 9959 19762 9968
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19168 9710 19288 9738
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19168 9217 19196 9590
rect 19154 9208 19210 9217
rect 19154 9143 19210 9152
rect 19260 8514 19288 9710
rect 19352 9586 19380 9862
rect 19449 9820 19745 9840
rect 19505 9818 19529 9820
rect 19585 9818 19609 9820
rect 19665 9818 19689 9820
rect 19527 9766 19529 9818
rect 19591 9766 19603 9818
rect 19665 9766 19667 9818
rect 19505 9764 19529 9766
rect 19585 9764 19609 9766
rect 19665 9764 19689 9766
rect 19449 9744 19745 9764
rect 19812 9586 19840 10134
rect 19904 10010 19932 10406
rect 19996 10112 20024 12294
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20088 10606 20116 12174
rect 20180 12073 20208 17070
rect 20272 12617 20300 18566
rect 20364 15706 20392 21082
rect 20456 20618 20484 21830
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20548 20777 20576 21422
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20534 20768 20590 20777
rect 20534 20703 20590 20712
rect 20456 20590 20576 20618
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 19854 20484 20402
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20548 18329 20576 20590
rect 20640 19514 20668 20946
rect 20824 19786 20852 23920
rect 21468 22522 21496 23920
rect 21376 22494 21496 22522
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20916 20398 20944 20878
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20626 19408 20682 19417
rect 20626 19343 20682 19352
rect 20534 18320 20590 18329
rect 20534 18255 20590 18264
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20364 13530 20392 15642
rect 20456 15026 20484 16526
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 20548 14634 20576 18158
rect 20456 14606 20576 14634
rect 20456 14521 20484 14606
rect 20442 14512 20498 14521
rect 20442 14447 20498 14456
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20364 13297 20392 13330
rect 20350 13288 20406 13297
rect 20350 13223 20406 13232
rect 20456 12889 20484 14350
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20442 12880 20498 12889
rect 20442 12815 20498 12824
rect 20548 12730 20576 13670
rect 20640 12986 20668 19343
rect 20916 19310 20944 20334
rect 21376 19922 21404 22494
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 21468 19854 21496 21490
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21560 20806 21588 21286
rect 21652 21078 21680 21286
rect 21640 21072 21692 21078
rect 21640 21014 21692 21020
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21560 20398 21588 20742
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21732 20256 21784 20262
rect 21732 20198 21784 20204
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 21183 19360 21211 19722
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21100 19332 21211 19360
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20824 17542 20852 18226
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 21008 17882 21036 18022
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20824 17134 20852 17478
rect 20916 17134 20944 17614
rect 21008 17338 21036 17614
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 21008 16946 21036 17274
rect 20916 16918 21036 16946
rect 20916 16590 20944 16918
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20916 16114 20944 16526
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20812 16040 20864 16046
rect 20864 15988 20944 15994
rect 20812 15982 20944 15988
rect 20824 15966 20944 15982
rect 20916 15502 20944 15966
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15570 21036 15846
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20824 15366 20852 15438
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20718 14648 20774 14657
rect 20718 14583 20774 14592
rect 20732 14414 20760 14583
rect 20824 14550 20852 15302
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20916 14414 20944 15438
rect 21008 15162 21036 15506
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 21008 14482 21036 14894
rect 21100 14600 21128 19332
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18766 21312 19110
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21284 17678 21312 18702
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21376 17066 21404 19654
rect 21652 19174 21680 19858
rect 21744 19854 21772 20198
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21744 19310 21772 19790
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18902 21680 19110
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 21730 18320 21786 18329
rect 21730 18255 21786 18264
rect 21744 18086 21772 18255
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 21364 17060 21416 17066
rect 21364 17002 21416 17008
rect 21652 16726 21680 17274
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21560 15978 21588 16390
rect 21548 15972 21600 15978
rect 21548 15914 21600 15920
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21192 15065 21220 15098
rect 21178 15056 21234 15065
rect 21178 14991 21234 15000
rect 21560 14890 21588 15914
rect 21836 15314 21864 21558
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 21744 15286 21864 15314
rect 21548 14884 21600 14890
rect 21548 14826 21600 14832
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21100 14572 21220 14600
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20916 14278 20944 14350
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 13326 20944 14214
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20364 12702 20576 12730
rect 20812 12708 20864 12714
rect 20258 12608 20314 12617
rect 20258 12543 20314 12552
rect 20364 12424 20392 12702
rect 20812 12650 20864 12656
rect 20272 12396 20392 12424
rect 20166 12064 20222 12073
rect 20166 11999 20222 12008
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 19996 10084 20116 10112
rect 19904 9982 20024 10010
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 9625 19932 9862
rect 19890 9616 19946 9625
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19800 9580 19852 9586
rect 19890 9551 19946 9560
rect 19800 9522 19852 9528
rect 19432 9512 19484 9518
rect 19430 9480 19432 9489
rect 19484 9480 19486 9489
rect 19430 9415 19486 9424
rect 19338 9072 19394 9081
rect 19338 9007 19340 9016
rect 19392 9007 19394 9016
rect 19340 8978 19392 8984
rect 19720 8906 19748 9522
rect 19812 8906 19840 9522
rect 19996 9518 20024 9982
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 20088 9081 20116 10084
rect 20074 9072 20130 9081
rect 20074 9007 20130 9016
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19449 8732 19745 8752
rect 19505 8730 19529 8732
rect 19585 8730 19609 8732
rect 19665 8730 19689 8732
rect 19527 8678 19529 8730
rect 19591 8678 19603 8730
rect 19665 8678 19667 8730
rect 19505 8676 19529 8678
rect 19585 8676 19609 8678
rect 19665 8676 19689 8678
rect 19449 8656 19745 8676
rect 19260 8486 19380 8514
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19076 8022 19104 8366
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19154 8120 19210 8129
rect 19260 8090 19288 8298
rect 19154 8055 19210 8064
rect 19248 8084 19300 8090
rect 19168 8022 19196 8055
rect 19248 8026 19300 8032
rect 19064 8016 19116 8022
rect 19064 7958 19116 7964
rect 19156 8016 19208 8022
rect 19352 7970 19380 8486
rect 19156 7958 19208 7964
rect 19076 7342 19104 7958
rect 19260 7942 19380 7970
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19168 7546 19196 7822
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19168 7410 19196 7482
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19260 6769 19288 7942
rect 19890 7848 19946 7857
rect 19352 7818 19472 7834
rect 19352 7812 19484 7818
rect 19352 7806 19432 7812
rect 19246 6760 19302 6769
rect 19064 6724 19116 6730
rect 19246 6695 19302 6704
rect 19064 6666 19116 6672
rect 18788 6326 18840 6332
rect 18892 6310 19012 6338
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 18524 5302 18552 5850
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4146 18552 4558
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18234 4040 18290 4049
rect 18234 3975 18290 3984
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18432 3738 18460 3878
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18340 2922 18368 3470
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18340 2514 18368 2858
rect 18432 2582 18460 3402
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 2582 18644 3334
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17696 1970 17724 2382
rect 18708 2106 18736 5170
rect 18800 5166 18828 5510
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18892 2553 18920 6310
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18984 4690 19012 5510
rect 19076 5409 19104 6666
rect 19352 6662 19380 7806
rect 19890 7783 19946 7792
rect 19432 7754 19484 7760
rect 19904 7750 19932 7783
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19449 7644 19745 7664
rect 19505 7642 19529 7644
rect 19585 7642 19609 7644
rect 19665 7642 19689 7644
rect 19527 7590 19529 7642
rect 19591 7590 19603 7642
rect 19665 7590 19667 7642
rect 19505 7588 19529 7590
rect 19585 7588 19609 7590
rect 19665 7588 19689 7590
rect 19449 7568 19745 7588
rect 19812 6984 19840 7686
rect 19720 6956 19840 6984
rect 19720 6798 19748 6956
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6254 19380 6598
rect 19449 6556 19745 6576
rect 19505 6554 19529 6556
rect 19585 6554 19609 6556
rect 19665 6554 19689 6556
rect 19527 6502 19529 6554
rect 19591 6502 19603 6554
rect 19665 6502 19667 6554
rect 19505 6500 19529 6502
rect 19585 6500 19609 6502
rect 19665 6500 19689 6502
rect 19449 6480 19745 6500
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19812 6186 19840 6802
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 19614 5944 19670 5953
rect 19614 5879 19670 5888
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 19062 5400 19118 5409
rect 19168 5370 19196 5714
rect 19628 5710 19656 5879
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19812 5642 19840 6122
rect 19904 5658 19932 6734
rect 19996 6361 20024 8774
rect 20088 8294 20116 8910
rect 20180 8430 20208 11834
rect 20272 11558 20300 12396
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 20272 10470 20300 10746
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20076 8288 20128 8294
rect 20272 8276 20300 10406
rect 20364 8362 20392 12242
rect 20534 12200 20590 12209
rect 20534 12135 20590 12144
rect 20442 12064 20498 12073
rect 20442 11999 20498 12008
rect 20456 10130 20484 11999
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20442 9616 20498 9625
rect 20442 9551 20498 9560
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20076 8230 20128 8236
rect 20180 8248 20300 8276
rect 20088 7206 20116 8230
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19982 6352 20038 6361
rect 19982 6287 20038 6296
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19984 6112 20036 6118
rect 19982 6080 19984 6089
rect 20036 6080 20038 6089
rect 19982 6015 20038 6024
rect 20088 5778 20116 6258
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19800 5636 19852 5642
rect 19904 5630 20024 5658
rect 19800 5578 19852 5584
rect 19062 5335 19118 5344
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 19064 5296 19116 5302
rect 19116 5244 19196 5250
rect 19064 5238 19196 5244
rect 19076 5222 19196 5238
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 19076 4146 19104 4966
rect 19168 4622 19196 5222
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18984 3534 19012 4014
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 19168 3398 19196 3946
rect 19260 3754 19288 5578
rect 19890 5536 19946 5545
rect 19449 5468 19745 5488
rect 19890 5471 19946 5480
rect 19505 5466 19529 5468
rect 19585 5466 19609 5468
rect 19665 5466 19689 5468
rect 19527 5414 19529 5466
rect 19591 5414 19603 5466
rect 19665 5414 19667 5466
rect 19505 5412 19529 5414
rect 19585 5412 19609 5414
rect 19665 5412 19689 5414
rect 19449 5392 19745 5412
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19352 4486 19380 5102
rect 19904 4690 19932 5471
rect 19996 5166 20024 5630
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19449 4380 19745 4400
rect 19505 4378 19529 4380
rect 19585 4378 19609 4380
rect 19665 4378 19689 4380
rect 19527 4326 19529 4378
rect 19591 4326 19603 4378
rect 19665 4326 19667 4378
rect 19505 4324 19529 4326
rect 19585 4324 19609 4326
rect 19665 4324 19689 4326
rect 19449 4304 19745 4324
rect 19524 4208 19576 4214
rect 19812 4196 19840 4558
rect 19576 4168 19840 4196
rect 19524 4150 19576 4156
rect 19260 3726 19380 3754
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19260 3194 19288 3538
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 19076 2650 19104 2790
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 18878 2544 18934 2553
rect 18878 2479 18934 2488
rect 18696 2100 18748 2106
rect 18696 2042 18748 2048
rect 17684 1964 17736 1970
rect 17684 1906 17736 1912
rect 19168 1578 19196 3130
rect 19260 2990 19288 3130
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19352 2514 19380 3726
rect 19449 3292 19745 3312
rect 19505 3290 19529 3292
rect 19585 3290 19609 3292
rect 19665 3290 19689 3292
rect 19527 3238 19529 3290
rect 19591 3238 19603 3290
rect 19665 3238 19667 3290
rect 19505 3236 19529 3238
rect 19585 3236 19609 3238
rect 19665 3236 19689 3238
rect 19449 3216 19745 3236
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19996 2310 20024 4966
rect 20180 3641 20208 8248
rect 20456 7290 20484 9551
rect 20364 7262 20484 7290
rect 20258 5672 20314 5681
rect 20258 5607 20314 5616
rect 20166 3632 20222 3641
rect 20166 3567 20222 3576
rect 20272 2650 20300 5607
rect 20364 2961 20392 7262
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20350 2952 20406 2961
rect 20350 2887 20406 2896
rect 20456 2650 20484 7142
rect 20548 4865 20576 12135
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 10606 20668 12038
rect 20732 11898 20760 12310
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20824 10198 20852 12650
rect 20916 12306 20944 13262
rect 21192 12356 21220 14572
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21284 14074 21312 14418
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21468 13870 21496 14758
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21652 13802 21680 14758
rect 21640 13796 21692 13802
rect 21640 13738 21692 13744
rect 21652 12850 21680 13738
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21454 12744 21510 12753
rect 21454 12679 21510 12688
rect 21192 12328 21404 12356
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20902 10840 20958 10849
rect 21008 10810 21036 12242
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21284 11218 21312 11630
rect 21272 11212 21324 11218
rect 21272 11154 21324 11160
rect 20902 10775 20958 10784
rect 20996 10804 21048 10810
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20720 9988 20772 9994
rect 20720 9930 20772 9936
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20640 8838 20668 9658
rect 20732 9586 20760 9930
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20732 8430 20760 9522
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20534 4856 20590 4865
rect 20534 4791 20590 4800
rect 20640 4321 20668 8298
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20732 6390 20760 7210
rect 20810 6896 20866 6905
rect 20810 6831 20812 6840
rect 20864 6831 20866 6840
rect 20812 6802 20864 6808
rect 20916 6746 20944 10775
rect 20996 10746 21048 10752
rect 21178 10568 21234 10577
rect 21178 10503 21180 10512
rect 21232 10503 21234 10512
rect 21180 10474 21232 10480
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 21008 9722 21036 10066
rect 21284 9994 21312 11154
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21284 9042 21312 9522
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20994 8256 21050 8265
rect 20994 8191 21050 8200
rect 21270 8256 21326 8265
rect 21270 8191 21326 8200
rect 21008 7954 21036 8191
rect 21284 8022 21312 8191
rect 21376 8129 21404 12328
rect 21468 10130 21496 12679
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21560 11665 21588 12582
rect 21652 11898 21680 12786
rect 21744 12782 21772 15286
rect 21928 15144 21956 21354
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22020 18737 22048 19858
rect 22006 18728 22062 18737
rect 22006 18663 22062 18672
rect 22112 18612 22140 23920
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22020 18584 22140 18612
rect 22020 18426 22048 18584
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 22112 17066 22140 18294
rect 22192 18080 22244 18086
rect 22296 18057 22324 21422
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22192 18022 22244 18028
rect 22282 18048 22338 18057
rect 22100 17060 22152 17066
rect 22100 17002 22152 17008
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21836 15116 21956 15144
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21546 11656 21602 11665
rect 21546 11591 21602 11600
rect 21836 11370 21864 15116
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21928 14278 21956 14962
rect 22020 14822 22048 16934
rect 22204 16794 22232 18022
rect 22282 17983 22338 17992
rect 22480 17377 22508 20334
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 22664 18630 22692 19858
rect 22756 18834 22784 23920
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22466 17368 22522 17377
rect 22466 17303 22522 17312
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22466 16688 22522 16697
rect 22466 16623 22522 16632
rect 22480 14958 22508 16623
rect 22572 16250 22600 18226
rect 22664 17814 22692 18566
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22572 15910 22600 16186
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 22020 14618 22048 14758
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21928 13462 21956 14214
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 13530 22232 13670
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 21916 13456 21968 13462
rect 21916 13398 21968 13404
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22100 12844 22152 12850
rect 22152 12804 22232 12832
rect 22100 12786 22152 12792
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 21744 11342 21864 11370
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21362 8120 21418 8129
rect 21362 8055 21418 8064
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21008 7585 21036 7890
rect 20994 7576 21050 7585
rect 20994 7511 21050 7520
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 21008 6866 21036 7142
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20824 6718 20944 6746
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20824 6186 20852 6718
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 20916 5778 20944 6598
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20812 5704 20864 5710
rect 20864 5652 20944 5658
rect 20812 5646 20944 5652
rect 20824 5630 20944 5646
rect 20720 5568 20772 5574
rect 20718 5536 20720 5545
rect 20772 5536 20774 5545
rect 20718 5471 20774 5480
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20824 4758 20852 4966
rect 20812 4752 20864 4758
rect 20812 4694 20864 4700
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20626 4312 20682 4321
rect 20626 4247 20682 4256
rect 20732 4078 20760 4558
rect 20916 4554 20944 5630
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20732 3602 20760 4014
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20732 3058 20760 3538
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20732 2514 20760 2994
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 20824 2378 20852 3878
rect 20904 2916 20956 2922
rect 20904 2858 20956 2864
rect 20916 2582 20944 2858
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 21008 2446 21036 6802
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 6254 21128 6598
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21100 5778 21128 6054
rect 21192 5817 21220 7890
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 21270 6896 21326 6905
rect 21270 6831 21326 6840
rect 21284 6254 21312 6831
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21178 5808 21234 5817
rect 21088 5772 21140 5778
rect 21178 5743 21234 5752
rect 21088 5714 21140 5720
rect 21284 5166 21312 6190
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21100 4622 21128 5102
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 21376 3942 21404 4626
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21468 2990 21496 7511
rect 21560 5710 21588 10406
rect 21744 9738 21772 11342
rect 21928 11132 21956 12718
rect 22204 12102 22232 12804
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22204 11286 22232 12038
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 21652 9710 21772 9738
rect 21836 11104 21956 11132
rect 21652 6066 21680 9710
rect 21652 6038 21772 6066
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21560 5370 21588 5510
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21652 4078 21680 5850
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 21652 3738 21680 4014
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21744 3097 21772 6038
rect 21836 3913 21864 11104
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 8809 22048 10542
rect 22296 10266 22324 12854
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22192 9104 22244 9110
rect 22192 9046 22244 9052
rect 22006 8800 22062 8809
rect 22006 8735 22062 8744
rect 22204 8634 22232 9046
rect 22388 8838 22416 12718
rect 22652 11620 22704 11626
rect 22652 11562 22704 11568
rect 22664 11354 22692 11562
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22664 10062 22692 11290
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22652 9444 22704 9450
rect 22652 9386 22704 9392
rect 22664 9178 22692 9386
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21822 3904 21878 3913
rect 21822 3839 21878 3848
rect 21928 3602 21956 5714
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 22112 4826 22140 5034
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22204 4162 22232 7686
rect 22296 4486 22324 8366
rect 22388 6254 22416 8502
rect 22664 7886 22692 9114
rect 22756 8537 22784 17138
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22848 13190 22876 13874
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22742 8528 22798 8537
rect 22742 8463 22798 8472
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22376 6248 22428 6254
rect 22480 6225 22508 7210
rect 22756 7002 22784 7278
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22756 6905 22784 6938
rect 22742 6896 22798 6905
rect 22742 6831 22798 6840
rect 22376 6190 22428 6196
rect 22466 6216 22522 6225
rect 22466 6151 22522 6160
rect 22560 6180 22612 6186
rect 22560 6122 22612 6128
rect 22572 5370 22600 6122
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 22756 5953 22784 6054
rect 22742 5944 22798 5953
rect 22742 5879 22798 5888
rect 22848 5545 22876 13126
rect 22940 6361 22968 20198
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 23032 6458 23060 8774
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 22926 6352 22982 6361
rect 22926 6287 22982 6296
rect 22834 5536 22890 5545
rect 22834 5471 22890 5480
rect 22560 5364 22612 5370
rect 22560 5306 22612 5312
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22204 4134 22416 4162
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21928 3194 21956 3538
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 21730 3088 21786 3097
rect 21730 3023 21786 3032
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 20812 2372 20864 2378
rect 20812 2314 20864 2320
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19449 2204 19745 2224
rect 19505 2202 19529 2204
rect 19585 2202 19609 2204
rect 19665 2202 19689 2204
rect 19527 2150 19529 2202
rect 19591 2150 19603 2202
rect 19665 2150 19667 2202
rect 19505 2148 19529 2150
rect 19585 2148 19609 2150
rect 19665 2148 19689 2150
rect 19449 2128 19745 2148
rect 20824 1970 20852 2314
rect 20812 1964 20864 1970
rect 20812 1906 20864 1912
rect 22388 1601 22416 4134
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 19076 1550 19196 1578
rect 22374 1592 22430 1601
rect 17316 1352 17368 1358
rect 17316 1294 17368 1300
rect 19076 480 19104 1550
rect 22374 1527 22430 1536
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 19352 921 19380 1294
rect 19338 912 19394 921
rect 19338 847 19394 856
rect 22572 480 22600 2790
rect 1674 0 1730 480
rect 5078 0 5134 480
rect 8574 0 8630 480
rect 12070 0 12126 480
rect 15566 0 15622 480
rect 19062 0 19118 480
rect 22558 0 22614 480
rect 23032 377 23060 6394
rect 23216 4282 23244 21286
rect 23400 17202 23428 23920
rect 24044 20330 24072 23920
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23204 4276 23256 4282
rect 23204 4218 23256 4224
rect 23018 368 23074 377
rect 23018 303 23074 312
<< via2 >>
rect 20350 23976 20406 24032
rect 1398 20984 1454 21040
rect 1766 18672 1822 18728
rect 1674 17740 1730 17776
rect 1674 17720 1676 17740
rect 1676 17720 1728 17740
rect 1728 17720 1730 17740
rect 1858 14320 1914 14376
rect 1674 12860 1676 12880
rect 1676 12860 1728 12880
rect 1728 12860 1730 12880
rect 1674 12824 1730 12860
rect 2594 21548 2650 21584
rect 2594 21528 2596 21548
rect 2596 21528 2648 21548
rect 2648 21528 2650 21548
rect 2226 9968 2282 10024
rect 2594 17584 2650 17640
rect 2778 17176 2834 17232
rect 2778 16632 2834 16688
rect 2962 17584 3018 17640
rect 2502 12144 2558 12200
rect 3330 15136 3386 15192
rect 1490 9016 1546 9072
rect 2962 11600 3018 11656
rect 3422 14476 3478 14512
rect 3422 14456 3424 14476
rect 3424 14456 3476 14476
rect 3476 14456 3478 14476
rect 3606 17040 3662 17096
rect 3330 11056 3386 11112
rect 3698 11056 3754 11112
rect 2502 7948 2558 7984
rect 2502 7928 2504 7948
rect 2504 7928 2556 7948
rect 2556 7928 2558 7948
rect 1950 3052 2006 3088
rect 1950 3032 1952 3052
rect 1952 3032 2004 3052
rect 2004 3032 2006 3052
rect 4654 21786 4710 21788
rect 4734 21786 4790 21788
rect 4814 21786 4870 21788
rect 4894 21786 4950 21788
rect 4654 21734 4680 21786
rect 4680 21734 4710 21786
rect 4734 21734 4744 21786
rect 4744 21734 4790 21786
rect 4814 21734 4860 21786
rect 4860 21734 4870 21786
rect 4894 21734 4924 21786
rect 4924 21734 4950 21786
rect 4654 21732 4710 21734
rect 4734 21732 4790 21734
rect 4814 21732 4870 21734
rect 4894 21732 4950 21734
rect 3974 21256 4030 21312
rect 4654 20698 4710 20700
rect 4734 20698 4790 20700
rect 4814 20698 4870 20700
rect 4894 20698 4950 20700
rect 4654 20646 4680 20698
rect 4680 20646 4710 20698
rect 4734 20646 4744 20698
rect 4744 20646 4790 20698
rect 4814 20646 4860 20698
rect 4860 20646 4870 20698
rect 4894 20646 4924 20698
rect 4924 20646 4950 20698
rect 4654 20644 4710 20646
rect 4734 20644 4790 20646
rect 4814 20644 4870 20646
rect 4894 20644 4950 20646
rect 4654 19610 4710 19612
rect 4734 19610 4790 19612
rect 4814 19610 4870 19612
rect 4894 19610 4950 19612
rect 4654 19558 4680 19610
rect 4680 19558 4710 19610
rect 4734 19558 4744 19610
rect 4744 19558 4790 19610
rect 4814 19558 4860 19610
rect 4860 19558 4870 19610
rect 4894 19558 4924 19610
rect 4924 19558 4950 19610
rect 4654 19556 4710 19558
rect 4734 19556 4790 19558
rect 4814 19556 4870 19558
rect 4894 19556 4950 19558
rect 4434 18808 4490 18864
rect 4250 17076 4252 17096
rect 4252 17076 4304 17096
rect 4304 17076 4306 17096
rect 4250 17040 4306 17076
rect 3882 16768 3938 16824
rect 4654 18522 4710 18524
rect 4734 18522 4790 18524
rect 4814 18522 4870 18524
rect 4894 18522 4950 18524
rect 4654 18470 4680 18522
rect 4680 18470 4710 18522
rect 4734 18470 4744 18522
rect 4744 18470 4790 18522
rect 4814 18470 4860 18522
rect 4860 18470 4870 18522
rect 4894 18470 4924 18522
rect 4924 18470 4950 18522
rect 4654 18468 4710 18470
rect 4734 18468 4790 18470
rect 4814 18468 4870 18470
rect 4894 18468 4950 18470
rect 5078 18572 5080 18592
rect 5080 18572 5132 18592
rect 5132 18572 5134 18592
rect 5078 18536 5134 18572
rect 4802 17992 4858 18048
rect 4654 17434 4710 17436
rect 4734 17434 4790 17436
rect 4814 17434 4870 17436
rect 4894 17434 4950 17436
rect 4654 17382 4680 17434
rect 4680 17382 4710 17434
rect 4734 17382 4744 17434
rect 4744 17382 4790 17434
rect 4814 17382 4860 17434
rect 4860 17382 4870 17434
rect 4894 17382 4924 17434
rect 4924 17382 4950 17434
rect 4654 17380 4710 17382
rect 4734 17380 4790 17382
rect 4814 17380 4870 17382
rect 4894 17380 4950 17382
rect 4986 17040 5042 17096
rect 5078 16768 5134 16824
rect 4654 16346 4710 16348
rect 4734 16346 4790 16348
rect 4814 16346 4870 16348
rect 4894 16346 4950 16348
rect 4654 16294 4680 16346
rect 4680 16294 4710 16346
rect 4734 16294 4744 16346
rect 4744 16294 4790 16346
rect 4814 16294 4860 16346
rect 4860 16294 4870 16346
rect 4894 16294 4924 16346
rect 4924 16294 4950 16346
rect 4654 16292 4710 16294
rect 4734 16292 4790 16294
rect 4814 16292 4870 16294
rect 4894 16292 4950 16294
rect 4710 15816 4766 15872
rect 4342 14728 4398 14784
rect 4250 13796 4306 13832
rect 4250 13776 4252 13796
rect 4252 13776 4304 13796
rect 4304 13776 4306 13796
rect 4250 13640 4306 13696
rect 4158 13368 4214 13424
rect 4894 15680 4950 15736
rect 4654 15258 4710 15260
rect 4734 15258 4790 15260
rect 4814 15258 4870 15260
rect 4894 15258 4950 15260
rect 4654 15206 4680 15258
rect 4680 15206 4710 15258
rect 4734 15206 4744 15258
rect 4744 15206 4790 15258
rect 4814 15206 4860 15258
rect 4860 15206 4870 15258
rect 4894 15206 4924 15258
rect 4924 15206 4950 15258
rect 4654 15204 4710 15206
rect 4734 15204 4790 15206
rect 4814 15204 4870 15206
rect 4894 15204 4950 15206
rect 5078 16088 5134 16144
rect 4618 14764 4620 14784
rect 4620 14764 4672 14784
rect 4672 14764 4674 14784
rect 4618 14728 4674 14764
rect 4654 14170 4710 14172
rect 4734 14170 4790 14172
rect 4814 14170 4870 14172
rect 4894 14170 4950 14172
rect 4654 14118 4680 14170
rect 4680 14118 4710 14170
rect 4734 14118 4744 14170
rect 4744 14118 4790 14170
rect 4814 14118 4860 14170
rect 4860 14118 4870 14170
rect 4894 14118 4924 14170
rect 4924 14118 4950 14170
rect 4654 14116 4710 14118
rect 4734 14116 4790 14118
rect 4814 14116 4870 14118
rect 4894 14116 4950 14118
rect 4894 13932 4950 13968
rect 4894 13912 4896 13932
rect 4896 13912 4948 13932
rect 4948 13912 4950 13932
rect 4654 13082 4710 13084
rect 4734 13082 4790 13084
rect 4814 13082 4870 13084
rect 4894 13082 4950 13084
rect 4654 13030 4680 13082
rect 4680 13030 4710 13082
rect 4734 13030 4744 13082
rect 4744 13030 4790 13082
rect 4814 13030 4860 13082
rect 4860 13030 4870 13082
rect 4894 13030 4924 13082
rect 4924 13030 4950 13082
rect 4654 13028 4710 13030
rect 4734 13028 4790 13030
rect 4814 13028 4870 13030
rect 4894 13028 4950 13030
rect 4654 11994 4710 11996
rect 4734 11994 4790 11996
rect 4814 11994 4870 11996
rect 4894 11994 4950 11996
rect 4654 11942 4680 11994
rect 4680 11942 4710 11994
rect 4734 11942 4744 11994
rect 4744 11942 4790 11994
rect 4814 11942 4860 11994
rect 4860 11942 4870 11994
rect 4894 11942 4924 11994
rect 4924 11942 4950 11994
rect 4654 11940 4710 11942
rect 4734 11940 4790 11942
rect 4814 11940 4870 11942
rect 4894 11940 4950 11942
rect 4802 11772 4804 11792
rect 4804 11772 4856 11792
rect 4856 11772 4858 11792
rect 4802 11736 4858 11772
rect 4894 11056 4950 11112
rect 4654 10906 4710 10908
rect 4734 10906 4790 10908
rect 4814 10906 4870 10908
rect 4894 10906 4950 10908
rect 4654 10854 4680 10906
rect 4680 10854 4710 10906
rect 4734 10854 4744 10906
rect 4744 10854 4790 10906
rect 4814 10854 4860 10906
rect 4860 10854 4870 10906
rect 4894 10854 4924 10906
rect 4924 10854 4950 10906
rect 4654 10852 4710 10854
rect 4734 10852 4790 10854
rect 4814 10852 4870 10854
rect 4894 10852 4950 10854
rect 4894 10668 4950 10704
rect 4894 10648 4896 10668
rect 4896 10648 4948 10668
rect 4948 10648 4950 10668
rect 4434 9968 4490 10024
rect 4654 9818 4710 9820
rect 4734 9818 4790 9820
rect 4814 9818 4870 9820
rect 4894 9818 4950 9820
rect 4654 9766 4680 9818
rect 4680 9766 4710 9818
rect 4734 9766 4744 9818
rect 4744 9766 4790 9818
rect 4814 9766 4860 9818
rect 4860 9766 4870 9818
rect 4894 9766 4924 9818
rect 4924 9766 4950 9818
rect 4654 9764 4710 9766
rect 4734 9764 4790 9766
rect 4814 9764 4870 9766
rect 4894 9764 4950 9766
rect 4654 8730 4710 8732
rect 4734 8730 4790 8732
rect 4814 8730 4870 8732
rect 4894 8730 4950 8732
rect 4654 8678 4680 8730
rect 4680 8678 4710 8730
rect 4734 8678 4744 8730
rect 4744 8678 4790 8730
rect 4814 8678 4860 8730
rect 4860 8678 4870 8730
rect 4894 8678 4924 8730
rect 4924 8678 4950 8730
rect 4654 8676 4710 8678
rect 4734 8676 4790 8678
rect 4814 8676 4870 8678
rect 4894 8676 4950 8678
rect 4654 7642 4710 7644
rect 4734 7642 4790 7644
rect 4814 7642 4870 7644
rect 4894 7642 4950 7644
rect 4654 7590 4680 7642
rect 4680 7590 4710 7642
rect 4734 7590 4744 7642
rect 4744 7590 4790 7642
rect 4814 7590 4860 7642
rect 4860 7590 4870 7642
rect 4894 7590 4924 7642
rect 4924 7590 4950 7642
rect 4654 7588 4710 7590
rect 4734 7588 4790 7590
rect 4814 7588 4870 7590
rect 4894 7588 4950 7590
rect 5170 14728 5226 14784
rect 5170 13776 5226 13832
rect 5170 13640 5226 13696
rect 5078 8472 5134 8528
rect 5998 19624 6054 19680
rect 5446 14728 5502 14784
rect 5722 16496 5778 16552
rect 5630 15816 5686 15872
rect 5354 13096 5410 13152
rect 5262 12688 5318 12744
rect 5354 8744 5410 8800
rect 4654 6554 4710 6556
rect 4734 6554 4790 6556
rect 4814 6554 4870 6556
rect 4894 6554 4950 6556
rect 4654 6502 4680 6554
rect 4680 6502 4710 6554
rect 4734 6502 4744 6554
rect 4744 6502 4790 6554
rect 4814 6502 4860 6554
rect 4860 6502 4870 6554
rect 4894 6502 4924 6554
rect 4924 6502 4950 6554
rect 4654 6500 4710 6502
rect 4734 6500 4790 6502
rect 4814 6500 4870 6502
rect 4894 6500 4950 6502
rect 5538 7656 5594 7712
rect 5998 16768 6054 16824
rect 5906 13912 5962 13968
rect 5906 13096 5962 13152
rect 5906 8200 5962 8256
rect 6090 13232 6146 13288
rect 6366 16108 6422 16144
rect 6366 16088 6368 16108
rect 6368 16088 6420 16108
rect 6420 16088 6422 16108
rect 6274 12280 6330 12336
rect 6366 10648 6422 10704
rect 6090 8472 6146 8528
rect 4654 5466 4710 5468
rect 4734 5466 4790 5468
rect 4814 5466 4870 5468
rect 4894 5466 4950 5468
rect 4654 5414 4680 5466
rect 4680 5414 4710 5466
rect 4734 5414 4744 5466
rect 4744 5414 4790 5466
rect 4814 5414 4860 5466
rect 4860 5414 4870 5466
rect 4894 5414 4924 5466
rect 4924 5414 4950 5466
rect 4654 5412 4710 5414
rect 4734 5412 4790 5414
rect 4814 5412 4870 5414
rect 4894 5412 4950 5414
rect 4654 4378 4710 4380
rect 4734 4378 4790 4380
rect 4814 4378 4870 4380
rect 4894 4378 4950 4380
rect 4654 4326 4680 4378
rect 4680 4326 4710 4378
rect 4734 4326 4744 4378
rect 4744 4326 4790 4378
rect 4814 4326 4860 4378
rect 4860 4326 4870 4378
rect 4894 4326 4924 4378
rect 4924 4326 4950 4378
rect 4654 4324 4710 4326
rect 4734 4324 4790 4326
rect 4814 4324 4870 4326
rect 4894 4324 4950 4326
rect 4654 3290 4710 3292
rect 4734 3290 4790 3292
rect 4814 3290 4870 3292
rect 4894 3290 4950 3292
rect 4654 3238 4680 3290
rect 4680 3238 4710 3290
rect 4734 3238 4744 3290
rect 4744 3238 4790 3290
rect 4814 3238 4860 3290
rect 4860 3238 4870 3290
rect 4894 3238 4924 3290
rect 4924 3238 4950 3290
rect 4654 3236 4710 3238
rect 4734 3236 4790 3238
rect 4814 3236 4870 3238
rect 4894 3236 4950 3238
rect 7010 18400 7066 18456
rect 6550 8200 6606 8256
rect 6826 14048 6882 14104
rect 6826 10512 6882 10568
rect 7194 16108 7250 16144
rect 7194 16088 7196 16108
rect 7196 16088 7248 16108
rect 7248 16088 7250 16108
rect 7194 15680 7250 15736
rect 9034 21528 9090 21584
rect 8353 21242 8409 21244
rect 8433 21242 8489 21244
rect 8513 21242 8569 21244
rect 8593 21242 8649 21244
rect 8353 21190 8379 21242
rect 8379 21190 8409 21242
rect 8433 21190 8443 21242
rect 8443 21190 8489 21242
rect 8513 21190 8559 21242
rect 8559 21190 8569 21242
rect 8593 21190 8623 21242
rect 8623 21190 8649 21242
rect 8353 21188 8409 21190
rect 8433 21188 8489 21190
rect 8513 21188 8569 21190
rect 8593 21188 8649 21190
rect 8353 20154 8409 20156
rect 8433 20154 8489 20156
rect 8513 20154 8569 20156
rect 8593 20154 8649 20156
rect 8353 20102 8379 20154
rect 8379 20102 8409 20154
rect 8433 20102 8443 20154
rect 8443 20102 8489 20154
rect 8513 20102 8559 20154
rect 8559 20102 8569 20154
rect 8593 20102 8623 20154
rect 8623 20102 8649 20154
rect 8353 20100 8409 20102
rect 8433 20100 8489 20102
rect 8513 20100 8569 20102
rect 8593 20100 8649 20102
rect 8114 19760 8170 19816
rect 8206 19488 8262 19544
rect 8574 19760 8630 19816
rect 8942 19624 8998 19680
rect 8353 19066 8409 19068
rect 8433 19066 8489 19068
rect 8513 19066 8569 19068
rect 8593 19066 8649 19068
rect 8353 19014 8379 19066
rect 8379 19014 8409 19066
rect 8433 19014 8443 19066
rect 8443 19014 8489 19066
rect 8513 19014 8559 19066
rect 8559 19014 8569 19066
rect 8593 19014 8623 19066
rect 8623 19014 8649 19066
rect 8353 19012 8409 19014
rect 8433 19012 8489 19014
rect 8513 19012 8569 19014
rect 8593 19012 8649 19014
rect 9402 18672 9458 18728
rect 7930 17720 7986 17776
rect 8353 17978 8409 17980
rect 8433 17978 8489 17980
rect 8513 17978 8569 17980
rect 8593 17978 8649 17980
rect 8353 17926 8379 17978
rect 8379 17926 8409 17978
rect 8433 17926 8443 17978
rect 8443 17926 8489 17978
rect 8513 17926 8559 17978
rect 8559 17926 8569 17978
rect 8593 17926 8623 17978
rect 8623 17926 8649 17978
rect 8353 17924 8409 17926
rect 8433 17924 8489 17926
rect 8513 17924 8569 17926
rect 8593 17924 8649 17926
rect 6826 9016 6882 9072
rect 7010 8608 7066 8664
rect 7010 7284 7012 7304
rect 7012 7284 7064 7304
rect 7064 7284 7066 7304
rect 7010 7248 7066 7284
rect 7470 11872 7526 11928
rect 7562 11600 7618 11656
rect 8353 16890 8409 16892
rect 8433 16890 8489 16892
rect 8513 16890 8569 16892
rect 8593 16890 8649 16892
rect 8353 16838 8379 16890
rect 8379 16838 8409 16890
rect 8433 16838 8443 16890
rect 8443 16838 8489 16890
rect 8513 16838 8559 16890
rect 8559 16838 8569 16890
rect 8593 16838 8623 16890
rect 8623 16838 8649 16890
rect 8353 16836 8409 16838
rect 8433 16836 8489 16838
rect 8513 16836 8569 16838
rect 8593 16836 8649 16838
rect 8298 16632 8354 16688
rect 8022 15952 8078 16008
rect 8850 16668 8852 16688
rect 8852 16668 8904 16688
rect 8904 16668 8906 16688
rect 8850 16632 8906 16668
rect 8850 16088 8906 16144
rect 8353 15802 8409 15804
rect 8433 15802 8489 15804
rect 8513 15802 8569 15804
rect 8593 15802 8649 15804
rect 8353 15750 8379 15802
rect 8379 15750 8409 15802
rect 8433 15750 8443 15802
rect 8443 15750 8489 15802
rect 8513 15750 8559 15802
rect 8559 15750 8569 15802
rect 8593 15750 8623 15802
rect 8623 15750 8649 15802
rect 8353 15748 8409 15750
rect 8433 15748 8489 15750
rect 8513 15748 8569 15750
rect 8593 15748 8649 15750
rect 8482 15308 8484 15328
rect 8484 15308 8536 15328
rect 8536 15308 8538 15328
rect 8482 15272 8538 15308
rect 8353 14714 8409 14716
rect 8433 14714 8489 14716
rect 8513 14714 8569 14716
rect 8593 14714 8649 14716
rect 8353 14662 8379 14714
rect 8379 14662 8409 14714
rect 8433 14662 8443 14714
rect 8443 14662 8489 14714
rect 8513 14662 8559 14714
rect 8559 14662 8569 14714
rect 8593 14662 8623 14714
rect 8623 14662 8649 14714
rect 8353 14660 8409 14662
rect 8433 14660 8489 14662
rect 8513 14660 8569 14662
rect 8593 14660 8649 14662
rect 8574 14492 8576 14512
rect 8576 14492 8628 14512
rect 8628 14492 8630 14512
rect 8574 14456 8630 14492
rect 8022 12824 8078 12880
rect 7838 11872 7894 11928
rect 7562 7812 7618 7848
rect 7562 7792 7564 7812
rect 7564 7792 7616 7812
rect 7616 7792 7618 7812
rect 7562 7540 7618 7576
rect 7562 7520 7564 7540
rect 7564 7520 7616 7540
rect 7616 7520 7618 7540
rect 7746 7248 7802 7304
rect 7562 5752 7618 5808
rect 7470 5364 7526 5400
rect 7470 5344 7472 5364
rect 7472 5344 7524 5364
rect 7524 5344 7526 5364
rect 8353 13626 8409 13628
rect 8433 13626 8489 13628
rect 8513 13626 8569 13628
rect 8593 13626 8649 13628
rect 8353 13574 8379 13626
rect 8379 13574 8409 13626
rect 8433 13574 8443 13626
rect 8443 13574 8489 13626
rect 8513 13574 8559 13626
rect 8559 13574 8569 13626
rect 8593 13574 8623 13626
rect 8623 13574 8649 13626
rect 8353 13572 8409 13574
rect 8433 13572 8489 13574
rect 8513 13572 8569 13574
rect 8593 13572 8649 13574
rect 8353 12538 8409 12540
rect 8433 12538 8489 12540
rect 8513 12538 8569 12540
rect 8593 12538 8649 12540
rect 8353 12486 8379 12538
rect 8379 12486 8409 12538
rect 8433 12486 8443 12538
rect 8443 12486 8489 12538
rect 8513 12486 8559 12538
rect 8559 12486 8569 12538
rect 8593 12486 8623 12538
rect 8623 12486 8649 12538
rect 8353 12484 8409 12486
rect 8433 12484 8489 12486
rect 8513 12484 8569 12486
rect 8593 12484 8649 12486
rect 8353 11450 8409 11452
rect 8433 11450 8489 11452
rect 8513 11450 8569 11452
rect 8593 11450 8649 11452
rect 8353 11398 8379 11450
rect 8379 11398 8409 11450
rect 8433 11398 8443 11450
rect 8443 11398 8489 11450
rect 8513 11398 8559 11450
rect 8559 11398 8569 11450
rect 8593 11398 8623 11450
rect 8623 11398 8649 11450
rect 8353 11396 8409 11398
rect 8433 11396 8489 11398
rect 8513 11396 8569 11398
rect 8593 11396 8649 11398
rect 8353 10362 8409 10364
rect 8433 10362 8489 10364
rect 8513 10362 8569 10364
rect 8593 10362 8649 10364
rect 8353 10310 8379 10362
rect 8379 10310 8409 10362
rect 8433 10310 8443 10362
rect 8443 10310 8489 10362
rect 8513 10310 8559 10362
rect 8559 10310 8569 10362
rect 8593 10310 8623 10362
rect 8623 10310 8649 10362
rect 8353 10308 8409 10310
rect 8433 10308 8489 10310
rect 8513 10308 8569 10310
rect 8593 10308 8649 10310
rect 8390 9696 8446 9752
rect 8022 8608 8078 8664
rect 8022 7964 8024 7984
rect 8024 7964 8076 7984
rect 8076 7964 8078 7984
rect 8022 7928 8078 7964
rect 8022 7384 8078 7440
rect 8022 6860 8078 6896
rect 8022 6840 8024 6860
rect 8024 6840 8076 6860
rect 8076 6840 8078 6860
rect 8353 9274 8409 9276
rect 8433 9274 8489 9276
rect 8513 9274 8569 9276
rect 8593 9274 8649 9276
rect 8353 9222 8379 9274
rect 8379 9222 8409 9274
rect 8433 9222 8443 9274
rect 8443 9222 8489 9274
rect 8513 9222 8559 9274
rect 8559 9222 8569 9274
rect 8593 9222 8623 9274
rect 8623 9222 8649 9274
rect 8353 9220 8409 9222
rect 8433 9220 8489 9222
rect 8513 9220 8569 9222
rect 8593 9220 8649 9222
rect 8298 9016 8354 9072
rect 8206 8780 8208 8800
rect 8208 8780 8260 8800
rect 8260 8780 8262 8800
rect 8206 8744 8262 8780
rect 8206 8608 8262 8664
rect 8482 8744 8538 8800
rect 8390 8492 8446 8528
rect 8390 8472 8392 8492
rect 8392 8472 8444 8492
rect 8444 8472 8446 8492
rect 8353 8186 8409 8188
rect 8433 8186 8489 8188
rect 8513 8186 8569 8188
rect 8593 8186 8649 8188
rect 8353 8134 8379 8186
rect 8379 8134 8409 8186
rect 8433 8134 8443 8186
rect 8443 8134 8489 8186
rect 8513 8134 8559 8186
rect 8559 8134 8569 8186
rect 8593 8134 8623 8186
rect 8623 8134 8649 8186
rect 8353 8132 8409 8134
rect 8433 8132 8489 8134
rect 8513 8132 8569 8134
rect 8593 8132 8649 8134
rect 9310 18128 9366 18184
rect 8850 14356 8852 14376
rect 8852 14356 8904 14376
rect 8904 14356 8906 14376
rect 8850 14320 8906 14356
rect 8758 12688 8814 12744
rect 8850 12300 8906 12336
rect 8850 12280 8852 12300
rect 8852 12280 8904 12300
rect 8904 12280 8906 12300
rect 8850 12164 8906 12200
rect 8850 12144 8852 12164
rect 8852 12144 8904 12164
rect 8904 12144 8906 12164
rect 8850 11736 8906 11792
rect 8850 11464 8906 11520
rect 9126 12960 9182 13016
rect 9218 12280 9274 12336
rect 9126 9424 9182 9480
rect 8758 8084 8814 8120
rect 8758 8064 8760 8084
rect 8760 8064 8812 8084
rect 8812 8064 8814 8084
rect 8206 7928 8262 7984
rect 8482 7692 8484 7712
rect 8484 7692 8536 7712
rect 8536 7692 8538 7712
rect 8482 7656 8538 7692
rect 8482 7520 8538 7576
rect 8298 7384 8354 7440
rect 8353 7098 8409 7100
rect 8433 7098 8489 7100
rect 8513 7098 8569 7100
rect 8593 7098 8649 7100
rect 8353 7046 8379 7098
rect 8379 7046 8409 7098
rect 8433 7046 8443 7098
rect 8443 7046 8489 7098
rect 8513 7046 8559 7098
rect 8559 7046 8569 7098
rect 8593 7046 8623 7098
rect 8623 7046 8649 7098
rect 8353 7044 8409 7046
rect 8433 7044 8489 7046
rect 8513 7044 8569 7046
rect 8593 7044 8649 7046
rect 8390 6296 8446 6352
rect 8353 6010 8409 6012
rect 8433 6010 8489 6012
rect 8513 6010 8569 6012
rect 8593 6010 8649 6012
rect 8353 5958 8379 6010
rect 8379 5958 8409 6010
rect 8433 5958 8443 6010
rect 8443 5958 8489 6010
rect 8513 5958 8559 6010
rect 8559 5958 8569 6010
rect 8593 5958 8623 6010
rect 8623 5958 8649 6010
rect 8353 5956 8409 5958
rect 8433 5956 8489 5958
rect 8513 5956 8569 5958
rect 8593 5956 8649 5958
rect 9034 8084 9090 8120
rect 9034 8064 9036 8084
rect 9036 8064 9088 8084
rect 9088 8064 9090 8084
rect 9034 6704 9090 6760
rect 9678 17992 9734 18048
rect 10414 19508 10470 19544
rect 10414 19488 10416 19508
rect 10416 19488 10468 19508
rect 10468 19488 10470 19508
rect 10414 18944 10470 19000
rect 9954 18128 10010 18184
rect 9862 16632 9918 16688
rect 9310 12144 9366 12200
rect 9678 16396 9680 16416
rect 9680 16396 9732 16416
rect 9732 16396 9734 16416
rect 9678 16360 9734 16396
rect 9770 16224 9826 16280
rect 9586 13368 9642 13424
rect 10046 13912 10102 13968
rect 10414 17584 10470 17640
rect 10782 17040 10838 17096
rect 10598 16360 10654 16416
rect 10230 15000 10286 15056
rect 10322 14320 10378 14376
rect 9954 12436 10010 12472
rect 9954 12416 9956 12436
rect 9956 12416 10008 12436
rect 10008 12416 10010 12436
rect 9678 10684 9680 10704
rect 9680 10684 9732 10704
rect 9732 10684 9734 10704
rect 9678 10648 9734 10684
rect 9310 9016 9366 9072
rect 9218 6976 9274 7032
rect 9862 12144 9918 12200
rect 9954 11872 10010 11928
rect 9770 9696 9826 9752
rect 10690 16088 10746 16144
rect 10506 14728 10562 14784
rect 10322 11736 10378 11792
rect 9862 9560 9918 9616
rect 9678 8372 9680 8392
rect 9680 8372 9732 8392
rect 9732 8372 9734 8392
rect 9678 8336 9734 8372
rect 9126 6180 9182 6216
rect 9126 6160 9128 6180
rect 9128 6160 9180 6180
rect 9180 6160 9182 6180
rect 8353 4922 8409 4924
rect 8433 4922 8489 4924
rect 8513 4922 8569 4924
rect 8593 4922 8649 4924
rect 8353 4870 8379 4922
rect 8379 4870 8409 4922
rect 8433 4870 8443 4922
rect 8443 4870 8489 4922
rect 8513 4870 8559 4922
rect 8559 4870 8569 4922
rect 8593 4870 8623 4922
rect 8623 4870 8649 4922
rect 8353 4868 8409 4870
rect 8433 4868 8489 4870
rect 8513 4868 8569 4870
rect 8593 4868 8649 4870
rect 8353 3834 8409 3836
rect 8433 3834 8489 3836
rect 8513 3834 8569 3836
rect 8593 3834 8649 3836
rect 8353 3782 8379 3834
rect 8379 3782 8409 3834
rect 8433 3782 8443 3834
rect 8443 3782 8489 3834
rect 8513 3782 8559 3834
rect 8559 3782 8569 3834
rect 8593 3782 8623 3834
rect 8623 3782 8649 3834
rect 8353 3780 8409 3782
rect 8433 3780 8489 3782
rect 8513 3780 8569 3782
rect 8593 3780 8649 3782
rect 9310 5888 9366 5944
rect 9402 5208 9458 5264
rect 9586 7384 9642 7440
rect 9678 6604 9680 6624
rect 9680 6604 9732 6624
rect 9732 6604 9734 6624
rect 9678 6568 9734 6604
rect 9862 6996 9918 7032
rect 9862 6976 9864 6996
rect 9864 6976 9916 6996
rect 9916 6976 9918 6996
rect 10046 8744 10102 8800
rect 10230 9288 10286 9344
rect 10230 9016 10286 9072
rect 10230 8064 10286 8120
rect 10230 5772 10286 5808
rect 10230 5752 10232 5772
rect 10232 5752 10284 5772
rect 10284 5752 10286 5772
rect 9862 4820 9918 4856
rect 11058 17176 11114 17232
rect 11058 16496 11114 16552
rect 10782 12824 10838 12880
rect 10598 12280 10654 12336
rect 10690 8608 10746 8664
rect 11058 12588 11060 12608
rect 11060 12588 11112 12608
rect 11112 12588 11114 12608
rect 11058 12552 11114 12588
rect 11242 15952 11298 16008
rect 11242 12280 11298 12336
rect 11058 9424 11114 9480
rect 11150 9288 11206 9344
rect 11426 18808 11482 18864
rect 12052 21786 12108 21788
rect 12132 21786 12188 21788
rect 12212 21786 12268 21788
rect 12292 21786 12348 21788
rect 12052 21734 12078 21786
rect 12078 21734 12108 21786
rect 12132 21734 12142 21786
rect 12142 21734 12188 21786
rect 12212 21734 12258 21786
rect 12258 21734 12268 21786
rect 12292 21734 12322 21786
rect 12322 21734 12348 21786
rect 12052 21732 12108 21734
rect 12132 21732 12188 21734
rect 12212 21732 12268 21734
rect 12292 21732 12348 21734
rect 12052 20698 12108 20700
rect 12132 20698 12188 20700
rect 12212 20698 12268 20700
rect 12292 20698 12348 20700
rect 12052 20646 12078 20698
rect 12078 20646 12108 20698
rect 12132 20646 12142 20698
rect 12142 20646 12188 20698
rect 12212 20646 12258 20698
rect 12258 20646 12268 20698
rect 12292 20646 12322 20698
rect 12322 20646 12348 20698
rect 12052 20644 12108 20646
rect 12132 20644 12188 20646
rect 12212 20644 12268 20646
rect 12292 20644 12348 20646
rect 12714 20304 12770 20360
rect 12438 19760 12494 19816
rect 12052 19610 12108 19612
rect 12132 19610 12188 19612
rect 12212 19610 12268 19612
rect 12292 19610 12348 19612
rect 12052 19558 12078 19610
rect 12078 19558 12108 19610
rect 12132 19558 12142 19610
rect 12142 19558 12188 19610
rect 12212 19558 12258 19610
rect 12258 19558 12268 19610
rect 12292 19558 12322 19610
rect 12322 19558 12348 19610
rect 12052 19556 12108 19558
rect 12132 19556 12188 19558
rect 12212 19556 12268 19558
rect 12292 19556 12348 19558
rect 12530 19508 12586 19544
rect 12530 19488 12532 19508
rect 12532 19488 12584 19508
rect 12584 19488 12586 19508
rect 11610 16632 11666 16688
rect 12438 18672 12494 18728
rect 12052 18522 12108 18524
rect 12132 18522 12188 18524
rect 12212 18522 12268 18524
rect 12292 18522 12348 18524
rect 12052 18470 12078 18522
rect 12078 18470 12108 18522
rect 12132 18470 12142 18522
rect 12142 18470 12188 18522
rect 12212 18470 12258 18522
rect 12258 18470 12268 18522
rect 12292 18470 12322 18522
rect 12322 18470 12348 18522
rect 12052 18468 12108 18470
rect 12132 18468 12188 18470
rect 12212 18468 12268 18470
rect 12292 18468 12348 18470
rect 12530 18264 12586 18320
rect 12052 17434 12108 17436
rect 12132 17434 12188 17436
rect 12212 17434 12268 17436
rect 12292 17434 12348 17436
rect 12052 17382 12078 17434
rect 12078 17382 12108 17434
rect 12132 17382 12142 17434
rect 12142 17382 12188 17434
rect 12212 17382 12258 17434
rect 12258 17382 12268 17434
rect 12292 17382 12322 17434
rect 12322 17382 12348 17434
rect 12052 17380 12108 17382
rect 12132 17380 12188 17382
rect 12212 17380 12268 17382
rect 12292 17380 12348 17382
rect 11610 15952 11666 16008
rect 11334 12144 11390 12200
rect 11334 11056 11390 11112
rect 11334 9968 11390 10024
rect 11334 9152 11390 9208
rect 10966 8064 11022 8120
rect 11242 9016 11298 9072
rect 10966 6996 11022 7032
rect 10966 6976 10968 6996
rect 10968 6976 11020 6996
rect 11020 6976 11022 6996
rect 9862 4800 9864 4820
rect 9864 4800 9916 4820
rect 9916 4800 9918 4820
rect 11518 8744 11574 8800
rect 12052 16346 12108 16348
rect 12132 16346 12188 16348
rect 12212 16346 12268 16348
rect 12292 16346 12348 16348
rect 12052 16294 12078 16346
rect 12078 16294 12108 16346
rect 12132 16294 12142 16346
rect 12142 16294 12188 16346
rect 12212 16294 12258 16346
rect 12258 16294 12268 16346
rect 12292 16294 12322 16346
rect 12322 16294 12348 16346
rect 12052 16292 12108 16294
rect 12132 16292 12188 16294
rect 12212 16292 12268 16294
rect 12292 16292 12348 16294
rect 12052 15258 12108 15260
rect 12132 15258 12188 15260
rect 12212 15258 12268 15260
rect 12292 15258 12348 15260
rect 12052 15206 12078 15258
rect 12078 15206 12108 15258
rect 12132 15206 12142 15258
rect 12142 15206 12188 15258
rect 12212 15206 12258 15258
rect 12258 15206 12268 15258
rect 12292 15206 12322 15258
rect 12322 15206 12348 15258
rect 12052 15204 12108 15206
rect 12132 15204 12188 15206
rect 12212 15204 12268 15206
rect 12292 15204 12348 15206
rect 12530 15544 12586 15600
rect 12162 14764 12164 14784
rect 12164 14764 12216 14784
rect 12216 14764 12218 14784
rect 12162 14728 12218 14764
rect 12346 14320 12402 14376
rect 12052 14170 12108 14172
rect 12132 14170 12188 14172
rect 12212 14170 12268 14172
rect 12292 14170 12348 14172
rect 12052 14118 12078 14170
rect 12078 14118 12108 14170
rect 12132 14118 12142 14170
rect 12142 14118 12188 14170
rect 12212 14118 12258 14170
rect 12258 14118 12268 14170
rect 12292 14118 12322 14170
rect 12322 14118 12348 14170
rect 12052 14116 12108 14118
rect 12132 14116 12188 14118
rect 12212 14116 12268 14118
rect 12292 14116 12348 14118
rect 12990 18400 13046 18456
rect 12898 18284 12954 18320
rect 12898 18264 12900 18284
rect 12900 18264 12952 18284
rect 12952 18264 12954 18284
rect 13634 19372 13690 19408
rect 13634 19352 13636 19372
rect 13636 19352 13688 19372
rect 13688 19352 13690 19372
rect 12990 17060 13046 17096
rect 12990 17040 12992 17060
rect 12992 17040 13044 17060
rect 13044 17040 13046 17060
rect 13634 15952 13690 16008
rect 11886 13232 11942 13288
rect 11794 12688 11850 12744
rect 11702 11872 11758 11928
rect 12052 13082 12108 13084
rect 12132 13082 12188 13084
rect 12212 13082 12268 13084
rect 12292 13082 12348 13084
rect 12052 13030 12078 13082
rect 12078 13030 12108 13082
rect 12132 13030 12142 13082
rect 12142 13030 12188 13082
rect 12212 13030 12258 13082
rect 12258 13030 12268 13082
rect 12292 13030 12322 13082
rect 12322 13030 12348 13082
rect 12052 13028 12108 13030
rect 12132 13028 12188 13030
rect 12212 13028 12268 13030
rect 12292 13028 12348 13030
rect 12052 11994 12108 11996
rect 12132 11994 12188 11996
rect 12212 11994 12268 11996
rect 12292 11994 12348 11996
rect 12052 11942 12078 11994
rect 12078 11942 12108 11994
rect 12132 11942 12142 11994
rect 12142 11942 12188 11994
rect 12212 11942 12258 11994
rect 12258 11942 12268 11994
rect 12292 11942 12322 11994
rect 12322 11942 12348 11994
rect 12052 11940 12108 11942
rect 12132 11940 12188 11942
rect 12212 11940 12268 11942
rect 12292 11940 12348 11942
rect 11610 7520 11666 7576
rect 11518 7112 11574 7168
rect 12052 10906 12108 10908
rect 12132 10906 12188 10908
rect 12212 10906 12268 10908
rect 12292 10906 12348 10908
rect 12052 10854 12078 10906
rect 12078 10854 12108 10906
rect 12132 10854 12142 10906
rect 12142 10854 12188 10906
rect 12212 10854 12258 10906
rect 12258 10854 12268 10906
rect 12292 10854 12322 10906
rect 12322 10854 12348 10906
rect 12052 10852 12108 10854
rect 12132 10852 12188 10854
rect 12212 10852 12268 10854
rect 12292 10852 12348 10854
rect 12438 10376 12494 10432
rect 12530 10240 12586 10296
rect 12052 9818 12108 9820
rect 12132 9818 12188 9820
rect 12212 9818 12268 9820
rect 12292 9818 12348 9820
rect 12052 9766 12078 9818
rect 12078 9766 12108 9818
rect 12132 9766 12142 9818
rect 12142 9766 12188 9818
rect 12212 9766 12258 9818
rect 12258 9766 12268 9818
rect 12292 9766 12322 9818
rect 12322 9766 12348 9818
rect 12052 9764 12108 9766
rect 12132 9764 12188 9766
rect 12212 9764 12268 9766
rect 12292 9764 12348 9766
rect 12052 8730 12108 8732
rect 12132 8730 12188 8732
rect 12212 8730 12268 8732
rect 12292 8730 12348 8732
rect 12052 8678 12078 8730
rect 12078 8678 12108 8730
rect 12132 8678 12142 8730
rect 12142 8678 12188 8730
rect 12212 8678 12258 8730
rect 12258 8678 12268 8730
rect 12292 8678 12322 8730
rect 12322 8678 12348 8730
rect 12052 8676 12108 8678
rect 12132 8676 12188 8678
rect 12212 8676 12268 8678
rect 12292 8676 12348 8678
rect 11702 6568 11758 6624
rect 12052 7642 12108 7644
rect 12132 7642 12188 7644
rect 12212 7642 12268 7644
rect 12292 7642 12348 7644
rect 12052 7590 12078 7642
rect 12078 7590 12108 7642
rect 12132 7590 12142 7642
rect 12142 7590 12188 7642
rect 12212 7590 12258 7642
rect 12258 7590 12268 7642
rect 12292 7590 12322 7642
rect 12322 7590 12348 7642
rect 12052 7588 12108 7590
rect 12132 7588 12188 7590
rect 12212 7588 12268 7590
rect 12292 7588 12348 7590
rect 12052 6554 12108 6556
rect 12132 6554 12188 6556
rect 12212 6554 12268 6556
rect 12292 6554 12348 6556
rect 12052 6502 12078 6554
rect 12078 6502 12108 6554
rect 12132 6502 12142 6554
rect 12142 6502 12188 6554
rect 12212 6502 12258 6554
rect 12258 6502 12268 6554
rect 12292 6502 12322 6554
rect 12322 6502 12348 6554
rect 12052 6500 12108 6502
rect 12132 6500 12188 6502
rect 12212 6500 12268 6502
rect 12292 6500 12348 6502
rect 12162 5752 12218 5808
rect 12052 5466 12108 5468
rect 12132 5466 12188 5468
rect 12212 5466 12268 5468
rect 12292 5466 12348 5468
rect 12052 5414 12078 5466
rect 12078 5414 12108 5466
rect 12132 5414 12142 5466
rect 12142 5414 12188 5466
rect 12212 5414 12258 5466
rect 12258 5414 12268 5466
rect 12292 5414 12322 5466
rect 12322 5414 12348 5466
rect 12052 5412 12108 5414
rect 12132 5412 12188 5414
rect 12212 5412 12268 5414
rect 12292 5412 12348 5414
rect 12052 4378 12108 4380
rect 12132 4378 12188 4380
rect 12212 4378 12268 4380
rect 12292 4378 12348 4380
rect 12052 4326 12078 4378
rect 12078 4326 12108 4378
rect 12132 4326 12142 4378
rect 12142 4326 12188 4378
rect 12212 4326 12258 4378
rect 12258 4326 12268 4378
rect 12292 4326 12322 4378
rect 12322 4326 12348 4378
rect 12052 4324 12108 4326
rect 12132 4324 12188 4326
rect 12212 4324 12268 4326
rect 12292 4324 12348 4326
rect 13542 15136 13598 15192
rect 13450 14456 13506 14512
rect 13174 12416 13230 12472
rect 13174 12144 13230 12200
rect 12990 12008 13046 12064
rect 13174 11872 13230 11928
rect 12806 11056 12862 11112
rect 12622 9560 12678 9616
rect 12714 7520 12770 7576
rect 12714 5344 12770 5400
rect 12622 5208 12678 5264
rect 12898 7268 12954 7304
rect 12898 7248 12900 7268
rect 12900 7248 12952 7268
rect 12952 7248 12954 7268
rect 12898 6296 12954 6352
rect 13174 11464 13230 11520
rect 13174 11056 13230 11112
rect 13174 9288 13230 9344
rect 13634 12416 13690 12472
rect 13542 11056 13598 11112
rect 13358 10240 13414 10296
rect 13358 8492 13414 8528
rect 13358 8472 13360 8492
rect 13360 8472 13412 8492
rect 13412 8472 13414 8492
rect 13450 7520 13506 7576
rect 13358 6976 13414 7032
rect 13082 6024 13138 6080
rect 12898 5480 12954 5536
rect 4654 2202 4710 2204
rect 4734 2202 4790 2204
rect 4814 2202 4870 2204
rect 4894 2202 4950 2204
rect 4654 2150 4680 2202
rect 4680 2150 4710 2202
rect 4734 2150 4744 2202
rect 4744 2150 4790 2202
rect 4814 2150 4860 2202
rect 4860 2150 4870 2202
rect 4894 2150 4924 2202
rect 4924 2150 4950 2202
rect 4654 2148 4710 2150
rect 4734 2148 4790 2150
rect 4814 2148 4870 2150
rect 4894 2148 4950 2150
rect 8353 2746 8409 2748
rect 8433 2746 8489 2748
rect 8513 2746 8569 2748
rect 8593 2746 8649 2748
rect 8353 2694 8379 2746
rect 8379 2694 8409 2746
rect 8433 2694 8443 2746
rect 8443 2694 8489 2746
rect 8513 2694 8559 2746
rect 8559 2694 8569 2746
rect 8593 2694 8623 2746
rect 8623 2694 8649 2746
rect 8353 2692 8409 2694
rect 8433 2692 8489 2694
rect 8513 2692 8569 2694
rect 8593 2692 8649 2694
rect 12052 3290 12108 3292
rect 12132 3290 12188 3292
rect 12212 3290 12268 3292
rect 12292 3290 12348 3292
rect 12052 3238 12078 3290
rect 12078 3238 12108 3290
rect 12132 3238 12142 3290
rect 12142 3238 12188 3290
rect 12212 3238 12258 3290
rect 12258 3238 12268 3290
rect 12292 3238 12322 3290
rect 12322 3238 12348 3290
rect 12052 3236 12108 3238
rect 12132 3236 12188 3238
rect 12212 3236 12268 3238
rect 12292 3236 12348 3238
rect 12990 3576 13046 3632
rect 13818 15272 13874 15328
rect 14830 20712 14886 20768
rect 15014 19488 15070 19544
rect 14830 18128 14886 18184
rect 14738 16516 14794 16552
rect 14738 16496 14740 16516
rect 14740 16496 14792 16516
rect 14792 16496 14794 16516
rect 15290 18944 15346 19000
rect 14002 13368 14058 13424
rect 14186 13368 14242 13424
rect 14002 12552 14058 12608
rect 13910 12416 13966 12472
rect 13818 12144 13874 12200
rect 13910 10240 13966 10296
rect 13634 5480 13690 5536
rect 13818 5616 13874 5672
rect 13818 4120 13874 4176
rect 13082 3304 13138 3360
rect 14278 12280 14334 12336
rect 14278 12008 14334 12064
rect 14462 12860 14464 12880
rect 14464 12860 14516 12880
rect 14516 12860 14518 12880
rect 14462 12824 14518 12860
rect 14554 11600 14610 11656
rect 15106 16632 15162 16688
rect 15198 15408 15254 15464
rect 14738 12688 14794 12744
rect 14738 12280 14794 12336
rect 14462 9052 14464 9072
rect 14464 9052 14516 9072
rect 14516 9052 14518 9072
rect 14462 9016 14518 9052
rect 14646 11076 14702 11112
rect 14646 11056 14648 11076
rect 14648 11056 14700 11076
rect 14700 11056 14702 11076
rect 14462 7248 14518 7304
rect 14370 6976 14426 7032
rect 14002 3576 14058 3632
rect 15106 13912 15162 13968
rect 15014 11736 15070 11792
rect 15014 10376 15070 10432
rect 15198 11192 15254 11248
rect 14922 9016 14978 9072
rect 14830 8064 14886 8120
rect 14646 7792 14702 7848
rect 15750 21242 15806 21244
rect 15830 21242 15886 21244
rect 15910 21242 15966 21244
rect 15990 21242 16046 21244
rect 15750 21190 15776 21242
rect 15776 21190 15806 21242
rect 15830 21190 15840 21242
rect 15840 21190 15886 21242
rect 15910 21190 15956 21242
rect 15956 21190 15966 21242
rect 15990 21190 16020 21242
rect 16020 21190 16046 21242
rect 15750 21188 15806 21190
rect 15830 21188 15886 21190
rect 15910 21188 15966 21190
rect 15990 21188 16046 21190
rect 15750 20154 15806 20156
rect 15830 20154 15886 20156
rect 15910 20154 15966 20156
rect 15990 20154 16046 20156
rect 15750 20102 15776 20154
rect 15776 20102 15806 20154
rect 15830 20102 15840 20154
rect 15840 20102 15886 20154
rect 15910 20102 15956 20154
rect 15956 20102 15966 20154
rect 15990 20102 16020 20154
rect 16020 20102 16046 20154
rect 15750 20100 15806 20102
rect 15830 20100 15886 20102
rect 15910 20100 15966 20102
rect 15990 20100 16046 20102
rect 15750 19372 15806 19408
rect 16210 19896 16266 19952
rect 15750 19352 15752 19372
rect 15752 19352 15804 19372
rect 15804 19352 15806 19372
rect 15750 19066 15806 19068
rect 15830 19066 15886 19068
rect 15910 19066 15966 19068
rect 15990 19066 16046 19068
rect 15750 19014 15776 19066
rect 15776 19014 15806 19066
rect 15830 19014 15840 19066
rect 15840 19014 15886 19066
rect 15910 19014 15956 19066
rect 15956 19014 15966 19066
rect 15990 19014 16020 19066
rect 16020 19014 16046 19066
rect 15750 19012 15806 19014
rect 15830 19012 15886 19014
rect 15910 19012 15966 19014
rect 15990 19012 16046 19014
rect 15658 18808 15714 18864
rect 16118 18400 16174 18456
rect 15934 18264 15990 18320
rect 16118 18264 16174 18320
rect 15750 17978 15806 17980
rect 15830 17978 15886 17980
rect 15910 17978 15966 17980
rect 15990 17978 16046 17980
rect 15750 17926 15776 17978
rect 15776 17926 15806 17978
rect 15830 17926 15840 17978
rect 15840 17926 15886 17978
rect 15910 17926 15956 17978
rect 15956 17926 15966 17978
rect 15990 17926 16020 17978
rect 16020 17926 16046 17978
rect 15750 17924 15806 17926
rect 15830 17924 15886 17926
rect 15910 17924 15966 17926
rect 15990 17924 16046 17926
rect 15566 17584 15622 17640
rect 15750 16890 15806 16892
rect 15830 16890 15886 16892
rect 15910 16890 15966 16892
rect 15990 16890 16046 16892
rect 15750 16838 15776 16890
rect 15776 16838 15806 16890
rect 15830 16838 15840 16890
rect 15840 16838 15886 16890
rect 15910 16838 15956 16890
rect 15956 16838 15966 16890
rect 15990 16838 16020 16890
rect 16020 16838 16046 16890
rect 15750 16836 15806 16838
rect 15830 16836 15886 16838
rect 15910 16836 15966 16838
rect 15990 16836 16046 16838
rect 15658 15952 15714 16008
rect 15750 15802 15806 15804
rect 15830 15802 15886 15804
rect 15910 15802 15966 15804
rect 15990 15802 16046 15804
rect 15750 15750 15776 15802
rect 15776 15750 15806 15802
rect 15830 15750 15840 15802
rect 15840 15750 15886 15802
rect 15910 15750 15956 15802
rect 15956 15750 15966 15802
rect 15990 15750 16020 15802
rect 16020 15750 16046 15802
rect 15750 15748 15806 15750
rect 15830 15748 15886 15750
rect 15910 15748 15966 15750
rect 15990 15748 16046 15750
rect 16026 15444 16028 15464
rect 16028 15444 16080 15464
rect 16080 15444 16082 15464
rect 16026 15408 16082 15444
rect 15750 15000 15806 15056
rect 15750 14714 15806 14716
rect 15830 14714 15886 14716
rect 15910 14714 15966 14716
rect 15990 14714 16046 14716
rect 15750 14662 15776 14714
rect 15776 14662 15806 14714
rect 15830 14662 15840 14714
rect 15840 14662 15886 14714
rect 15910 14662 15956 14714
rect 15956 14662 15966 14714
rect 15990 14662 16020 14714
rect 16020 14662 16046 14714
rect 15750 14660 15806 14662
rect 15830 14660 15886 14662
rect 15910 14660 15966 14662
rect 15990 14660 16046 14662
rect 15750 14476 15806 14512
rect 15750 14456 15752 14476
rect 15752 14456 15804 14476
rect 15804 14456 15806 14476
rect 16118 14220 16120 14240
rect 16120 14220 16172 14240
rect 16172 14220 16174 14240
rect 16118 14184 16174 14220
rect 15658 13776 15714 13832
rect 15750 13626 15806 13628
rect 15830 13626 15886 13628
rect 15910 13626 15966 13628
rect 15990 13626 16046 13628
rect 15750 13574 15776 13626
rect 15776 13574 15806 13626
rect 15830 13574 15840 13626
rect 15840 13574 15886 13626
rect 15910 13574 15956 13626
rect 15956 13574 15966 13626
rect 15990 13574 16020 13626
rect 16020 13574 16046 13626
rect 15750 13572 15806 13574
rect 15830 13572 15886 13574
rect 15910 13572 15966 13574
rect 15990 13572 16046 13574
rect 15566 12552 15622 12608
rect 15750 12538 15806 12540
rect 15830 12538 15886 12540
rect 15910 12538 15966 12540
rect 15990 12538 16046 12540
rect 15750 12486 15776 12538
rect 15776 12486 15806 12538
rect 15830 12486 15840 12538
rect 15840 12486 15886 12538
rect 15910 12486 15956 12538
rect 15956 12486 15966 12538
rect 15990 12486 16020 12538
rect 16020 12486 16046 12538
rect 15750 12484 15806 12486
rect 15830 12484 15886 12486
rect 15910 12484 15966 12486
rect 15990 12484 16046 12486
rect 15658 11892 15714 11928
rect 15658 11872 15660 11892
rect 15660 11872 15712 11892
rect 15712 11872 15714 11892
rect 15566 10104 15622 10160
rect 15566 9288 15622 9344
rect 15566 8492 15622 8528
rect 15566 8472 15568 8492
rect 15568 8472 15620 8492
rect 15620 8472 15622 8492
rect 15750 11600 15806 11656
rect 15750 11450 15806 11452
rect 15830 11450 15886 11452
rect 15910 11450 15966 11452
rect 15990 11450 16046 11452
rect 15750 11398 15776 11450
rect 15776 11398 15806 11450
rect 15830 11398 15840 11450
rect 15840 11398 15886 11450
rect 15910 11398 15956 11450
rect 15956 11398 15966 11450
rect 15990 11398 16020 11450
rect 16020 11398 16046 11450
rect 15750 11396 15806 11398
rect 15830 11396 15886 11398
rect 15910 11396 15966 11398
rect 15990 11396 16046 11398
rect 15934 10784 15990 10840
rect 15750 10362 15806 10364
rect 15830 10362 15886 10364
rect 15910 10362 15966 10364
rect 15990 10362 16046 10364
rect 15750 10310 15776 10362
rect 15776 10310 15806 10362
rect 15830 10310 15840 10362
rect 15840 10310 15886 10362
rect 15910 10310 15956 10362
rect 15956 10310 15966 10362
rect 15990 10310 16020 10362
rect 16020 10310 16046 10362
rect 15750 10308 15806 10310
rect 15830 10308 15886 10310
rect 15910 10308 15966 10310
rect 15990 10308 16046 10310
rect 15750 9274 15806 9276
rect 15830 9274 15886 9276
rect 15910 9274 15966 9276
rect 15990 9274 16046 9276
rect 15750 9222 15776 9274
rect 15776 9222 15806 9274
rect 15830 9222 15840 9274
rect 15840 9222 15886 9274
rect 15910 9222 15956 9274
rect 15956 9222 15966 9274
rect 15990 9222 16020 9274
rect 16020 9222 16046 9274
rect 15750 9220 15806 9222
rect 15830 9220 15886 9222
rect 15910 9220 15966 9222
rect 15990 9220 16046 9222
rect 15750 8186 15806 8188
rect 15830 8186 15886 8188
rect 15910 8186 15966 8188
rect 15990 8186 16046 8188
rect 15750 8134 15776 8186
rect 15776 8134 15806 8186
rect 15830 8134 15840 8186
rect 15840 8134 15886 8186
rect 15910 8134 15956 8186
rect 15956 8134 15966 8186
rect 15990 8134 16020 8186
rect 16020 8134 16046 8186
rect 15750 8132 15806 8134
rect 15830 8132 15886 8134
rect 15910 8132 15966 8134
rect 15990 8132 16046 8134
rect 16302 14884 16358 14920
rect 16302 14864 16304 14884
rect 16304 14864 16356 14884
rect 16356 14864 16358 14884
rect 16762 18264 16818 18320
rect 16946 20712 17002 20768
rect 16854 16496 16910 16552
rect 16670 15136 16726 15192
rect 16210 11600 16266 11656
rect 16762 12588 16764 12608
rect 16764 12588 16816 12608
rect 16816 12588 16818 12608
rect 16762 12552 16818 12588
rect 16394 11600 16450 11656
rect 16302 11056 16358 11112
rect 16486 10376 16542 10432
rect 16210 9152 16266 9208
rect 14646 4528 14702 4584
rect 14462 4256 14518 4312
rect 14278 3168 14334 3224
rect 14370 2896 14426 2952
rect 8574 2352 8630 2408
rect 13358 2644 13414 2680
rect 13358 2624 13360 2644
rect 13360 2624 13412 2644
rect 13412 2624 13414 2644
rect 15198 7112 15254 7168
rect 15290 6160 15346 6216
rect 15198 4664 15254 4720
rect 15014 4392 15070 4448
rect 14554 3440 14610 3496
rect 14738 3052 14794 3088
rect 14738 3032 14740 3052
rect 14740 3032 14792 3052
rect 14792 3032 14794 3052
rect 15750 7098 15806 7100
rect 15830 7098 15886 7100
rect 15910 7098 15966 7100
rect 15990 7098 16046 7100
rect 15750 7046 15776 7098
rect 15776 7046 15806 7098
rect 15830 7046 15840 7098
rect 15840 7046 15886 7098
rect 15910 7046 15956 7098
rect 15956 7046 15966 7098
rect 15990 7046 16020 7098
rect 16020 7046 16046 7098
rect 15750 7044 15806 7046
rect 15830 7044 15886 7046
rect 15910 7044 15966 7046
rect 15990 7044 16046 7046
rect 15566 6024 15622 6080
rect 15750 6010 15806 6012
rect 15830 6010 15886 6012
rect 15910 6010 15966 6012
rect 15990 6010 16046 6012
rect 15750 5958 15776 6010
rect 15776 5958 15806 6010
rect 15830 5958 15840 6010
rect 15840 5958 15886 6010
rect 15910 5958 15956 6010
rect 15956 5958 15966 6010
rect 15990 5958 16020 6010
rect 16020 5958 16046 6010
rect 15750 5956 15806 5958
rect 15830 5956 15886 5958
rect 15910 5956 15966 5958
rect 15990 5956 16046 5958
rect 15658 5480 15714 5536
rect 15474 4664 15530 4720
rect 15750 4922 15806 4924
rect 15830 4922 15886 4924
rect 15910 4922 15966 4924
rect 15990 4922 16046 4924
rect 15750 4870 15776 4922
rect 15776 4870 15806 4922
rect 15830 4870 15840 4922
rect 15840 4870 15886 4922
rect 15910 4870 15956 4922
rect 15956 4870 15966 4922
rect 15990 4870 16020 4922
rect 16020 4870 16046 4922
rect 15750 4868 15806 4870
rect 15830 4868 15886 4870
rect 15910 4868 15966 4870
rect 15990 4868 16046 4870
rect 15750 4428 15752 4448
rect 15752 4428 15804 4448
rect 15804 4428 15806 4448
rect 15750 4392 15806 4428
rect 15566 3984 15622 4040
rect 15014 2216 15070 2272
rect 12052 2202 12108 2204
rect 12132 2202 12188 2204
rect 12212 2202 12268 2204
rect 12292 2202 12348 2204
rect 12052 2150 12078 2202
rect 12078 2150 12108 2202
rect 12132 2150 12142 2202
rect 12142 2150 12188 2202
rect 12212 2150 12258 2202
rect 12258 2150 12268 2202
rect 12292 2150 12322 2202
rect 12322 2150 12348 2202
rect 12052 2148 12108 2150
rect 12132 2148 12188 2150
rect 12212 2148 12268 2150
rect 12292 2148 12348 2150
rect 15750 3834 15806 3836
rect 15830 3834 15886 3836
rect 15910 3834 15966 3836
rect 15990 3834 16046 3836
rect 15750 3782 15776 3834
rect 15776 3782 15806 3834
rect 15830 3782 15840 3834
rect 15840 3782 15886 3834
rect 15910 3782 15956 3834
rect 15956 3782 15966 3834
rect 15990 3782 16020 3834
rect 16020 3782 16046 3834
rect 15750 3780 15806 3782
rect 15830 3780 15886 3782
rect 15910 3780 15966 3782
rect 15990 3780 16046 3782
rect 16302 8336 16358 8392
rect 16670 10376 16726 10432
rect 16578 9152 16634 9208
rect 16394 6296 16450 6352
rect 16302 4392 16358 4448
rect 15750 3576 15806 3632
rect 15934 3596 15990 3632
rect 15934 3576 15936 3596
rect 15936 3576 15988 3596
rect 15988 3576 15990 3596
rect 15750 3032 15806 3088
rect 15750 2746 15806 2748
rect 15830 2746 15886 2748
rect 15910 2746 15966 2748
rect 15990 2746 16046 2748
rect 15750 2694 15776 2746
rect 15776 2694 15806 2746
rect 15830 2694 15840 2746
rect 15840 2694 15886 2746
rect 15910 2694 15956 2746
rect 15956 2694 15966 2746
rect 15990 2694 16020 2746
rect 16020 2694 16046 2746
rect 15750 2692 15806 2694
rect 15830 2692 15886 2694
rect 15910 2692 15966 2694
rect 15990 2692 16046 2694
rect 16762 6840 16818 6896
rect 16578 4120 16634 4176
rect 16670 3848 16726 3904
rect 16210 2760 16266 2816
rect 15658 2508 15714 2544
rect 15658 2488 15660 2508
rect 15660 2488 15712 2508
rect 15712 2488 15714 2508
rect 17222 17176 17278 17232
rect 16946 9596 16948 9616
rect 16948 9596 17000 9616
rect 17000 9596 17002 9616
rect 16946 9560 17002 9596
rect 16946 9288 17002 9344
rect 17406 18128 17462 18184
rect 17682 18264 17738 18320
rect 17406 15020 17462 15056
rect 17406 15000 17408 15020
rect 17408 15000 17460 15020
rect 17460 15000 17462 15020
rect 17406 14456 17462 14512
rect 17498 10956 17500 10976
rect 17500 10956 17552 10976
rect 17552 10956 17554 10976
rect 17498 10920 17554 10956
rect 17774 14592 17830 14648
rect 17130 9016 17186 9072
rect 17590 10376 17646 10432
rect 17498 8200 17554 8256
rect 17314 7928 17370 7984
rect 16946 6296 17002 6352
rect 16946 6024 17002 6080
rect 16946 5208 17002 5264
rect 16946 3712 17002 3768
rect 17130 5480 17186 5536
rect 17130 4256 17186 4312
rect 16946 3440 17002 3496
rect 16946 2216 17002 2272
rect 17866 12960 17922 13016
rect 17866 10240 17922 10296
rect 17866 10104 17922 10160
rect 17866 9424 17922 9480
rect 18786 19796 18788 19816
rect 18788 19796 18840 19816
rect 18840 19796 18842 19816
rect 18786 19760 18842 19796
rect 18050 12280 18106 12336
rect 18050 10412 18052 10432
rect 18052 10412 18104 10432
rect 18104 10412 18106 10432
rect 18050 10376 18106 10412
rect 18326 14728 18382 14784
rect 18326 14592 18382 14648
rect 18234 11192 18290 11248
rect 18234 10784 18290 10840
rect 19246 23296 19302 23352
rect 19154 22616 19210 22672
rect 19449 21786 19505 21788
rect 19529 21786 19585 21788
rect 19609 21786 19665 21788
rect 19689 21786 19745 21788
rect 19449 21734 19475 21786
rect 19475 21734 19505 21786
rect 19529 21734 19539 21786
rect 19539 21734 19585 21786
rect 19609 21734 19655 21786
rect 19655 21734 19665 21786
rect 19689 21734 19719 21786
rect 19719 21734 19745 21786
rect 19449 21732 19505 21734
rect 19529 21732 19585 21734
rect 19609 21732 19665 21734
rect 19689 21732 19745 21734
rect 19246 21256 19302 21312
rect 19890 21936 19946 21992
rect 19449 20698 19505 20700
rect 19529 20698 19585 20700
rect 19609 20698 19665 20700
rect 19689 20698 19745 20700
rect 19449 20646 19475 20698
rect 19475 20646 19505 20698
rect 19529 20646 19539 20698
rect 19539 20646 19585 20698
rect 19609 20646 19655 20698
rect 19655 20646 19665 20698
rect 19689 20646 19719 20698
rect 19719 20646 19745 20698
rect 19449 20644 19505 20646
rect 19529 20644 19585 20646
rect 19609 20644 19665 20646
rect 19689 20644 19745 20646
rect 19246 20032 19302 20088
rect 19982 20576 20038 20632
rect 19706 19760 19762 19816
rect 19449 19610 19505 19612
rect 19529 19610 19585 19612
rect 19609 19610 19665 19612
rect 19689 19610 19745 19612
rect 19449 19558 19475 19610
rect 19475 19558 19505 19610
rect 19529 19558 19539 19610
rect 19539 19558 19585 19610
rect 19609 19558 19655 19610
rect 19655 19558 19665 19610
rect 19689 19558 19719 19610
rect 19719 19558 19745 19610
rect 19449 19556 19505 19558
rect 19529 19556 19585 19558
rect 19609 19556 19665 19558
rect 19689 19556 19745 19558
rect 19890 19352 19946 19408
rect 19449 18522 19505 18524
rect 19529 18522 19585 18524
rect 19609 18522 19665 18524
rect 19689 18522 19745 18524
rect 19449 18470 19475 18522
rect 19475 18470 19505 18522
rect 19529 18470 19539 18522
rect 19539 18470 19585 18522
rect 19609 18470 19655 18522
rect 19655 18470 19665 18522
rect 19689 18470 19719 18522
rect 19719 18470 19745 18522
rect 19449 18468 19505 18470
rect 19529 18468 19585 18470
rect 19609 18468 19665 18470
rect 19689 18468 19745 18470
rect 20166 19236 20222 19272
rect 20166 19216 20168 19236
rect 20168 19216 20220 19236
rect 20220 19216 20222 19236
rect 20074 17992 20130 18048
rect 18786 16396 18788 16416
rect 18788 16396 18840 16416
rect 18840 16396 18842 16416
rect 18786 16360 18842 16396
rect 18694 16088 18750 16144
rect 18970 16088 19026 16144
rect 18694 12960 18750 13016
rect 18602 12416 18658 12472
rect 18878 13504 18934 13560
rect 18234 9152 18290 9208
rect 18142 8880 18198 8936
rect 18418 10376 18474 10432
rect 18418 10240 18474 10296
rect 18510 9424 18566 9480
rect 18418 9152 18474 9208
rect 18418 8336 18474 8392
rect 18142 6296 18198 6352
rect 19449 17434 19505 17436
rect 19529 17434 19585 17436
rect 19609 17434 19665 17436
rect 19689 17434 19745 17436
rect 19449 17382 19475 17434
rect 19475 17382 19505 17434
rect 19529 17382 19539 17434
rect 19539 17382 19585 17434
rect 19609 17382 19655 17434
rect 19655 17382 19665 17434
rect 19689 17382 19719 17434
rect 19719 17382 19745 17434
rect 19449 17380 19505 17382
rect 19529 17380 19585 17382
rect 19609 17380 19665 17382
rect 19689 17380 19745 17382
rect 19449 16346 19505 16348
rect 19529 16346 19585 16348
rect 19609 16346 19665 16348
rect 19689 16346 19745 16348
rect 19449 16294 19475 16346
rect 19475 16294 19505 16346
rect 19529 16294 19539 16346
rect 19539 16294 19585 16346
rect 19609 16294 19655 16346
rect 19655 16294 19665 16346
rect 19689 16294 19719 16346
rect 19719 16294 19745 16346
rect 19449 16292 19505 16294
rect 19529 16292 19585 16294
rect 19609 16292 19665 16294
rect 19689 16292 19745 16294
rect 19706 15408 19762 15464
rect 19449 15258 19505 15260
rect 19529 15258 19585 15260
rect 19609 15258 19665 15260
rect 19689 15258 19745 15260
rect 19449 15206 19475 15258
rect 19475 15206 19505 15258
rect 19529 15206 19539 15258
rect 19539 15206 19585 15258
rect 19609 15206 19655 15258
rect 19655 15206 19665 15258
rect 19689 15206 19719 15258
rect 19719 15206 19745 15258
rect 19449 15204 19505 15206
rect 19529 15204 19585 15206
rect 19609 15204 19665 15206
rect 19689 15204 19745 15206
rect 19338 14728 19394 14784
rect 19338 14320 19394 14376
rect 19798 14864 19854 14920
rect 19449 14170 19505 14172
rect 19529 14170 19585 14172
rect 19609 14170 19665 14172
rect 19689 14170 19745 14172
rect 19449 14118 19475 14170
rect 19475 14118 19505 14170
rect 19529 14118 19539 14170
rect 19539 14118 19585 14170
rect 19609 14118 19655 14170
rect 19655 14118 19665 14170
rect 19689 14118 19719 14170
rect 19719 14118 19745 14170
rect 19449 14116 19505 14118
rect 19529 14116 19585 14118
rect 19609 14116 19665 14118
rect 19689 14116 19745 14118
rect 19449 13082 19505 13084
rect 19529 13082 19585 13084
rect 19609 13082 19665 13084
rect 19689 13082 19745 13084
rect 19449 13030 19475 13082
rect 19475 13030 19505 13082
rect 19529 13030 19539 13082
rect 19539 13030 19585 13082
rect 19609 13030 19655 13082
rect 19655 13030 19665 13082
rect 19689 13030 19719 13082
rect 19719 13030 19745 13082
rect 19449 13028 19505 13030
rect 19529 13028 19585 13030
rect 19609 13028 19665 13030
rect 19689 13028 19745 13030
rect 19614 12552 19670 12608
rect 19982 14864 20038 14920
rect 19890 12416 19946 12472
rect 20166 17176 20222 17232
rect 20074 12688 20130 12744
rect 20074 12552 20130 12608
rect 19449 11994 19505 11996
rect 19529 11994 19585 11996
rect 19609 11994 19665 11996
rect 19689 11994 19745 11996
rect 19449 11942 19475 11994
rect 19475 11942 19505 11994
rect 19529 11942 19539 11994
rect 19539 11942 19585 11994
rect 19609 11942 19655 11994
rect 19655 11942 19665 11994
rect 19689 11942 19719 11994
rect 19719 11942 19745 11994
rect 19449 11940 19505 11942
rect 19529 11940 19585 11942
rect 19609 11940 19665 11942
rect 19689 11940 19745 11942
rect 19614 11600 19670 11656
rect 19338 11464 19394 11520
rect 18970 9560 19026 9616
rect 18970 9288 19026 9344
rect 18878 6432 18934 6488
rect 19449 10906 19505 10908
rect 19529 10906 19585 10908
rect 19609 10906 19665 10908
rect 19689 10906 19745 10908
rect 19449 10854 19475 10906
rect 19475 10854 19505 10906
rect 19529 10854 19539 10906
rect 19539 10854 19585 10906
rect 19609 10854 19655 10906
rect 19655 10854 19665 10906
rect 19689 10854 19719 10906
rect 19719 10854 19745 10906
rect 19449 10852 19505 10854
rect 19529 10852 19585 10854
rect 19609 10852 19665 10854
rect 19689 10852 19745 10854
rect 19890 10648 19946 10704
rect 19706 9968 19762 10024
rect 19154 9152 19210 9208
rect 19449 9818 19505 9820
rect 19529 9818 19585 9820
rect 19609 9818 19665 9820
rect 19689 9818 19745 9820
rect 19449 9766 19475 9818
rect 19475 9766 19505 9818
rect 19529 9766 19539 9818
rect 19539 9766 19585 9818
rect 19609 9766 19655 9818
rect 19655 9766 19665 9818
rect 19689 9766 19719 9818
rect 19719 9766 19745 9818
rect 19449 9764 19505 9766
rect 19529 9764 19585 9766
rect 19609 9764 19665 9766
rect 19689 9764 19745 9766
rect 20534 20712 20590 20768
rect 20626 19352 20682 19408
rect 20534 18264 20590 18320
rect 20442 14456 20498 14512
rect 20350 13232 20406 13288
rect 20442 12824 20498 12880
rect 20718 14592 20774 14648
rect 21730 18264 21786 18320
rect 21178 15000 21234 15056
rect 20258 12552 20314 12608
rect 20166 12008 20222 12064
rect 19890 9560 19946 9616
rect 19430 9460 19432 9480
rect 19432 9460 19484 9480
rect 19484 9460 19486 9480
rect 19430 9424 19486 9460
rect 19338 9036 19394 9072
rect 19338 9016 19340 9036
rect 19340 9016 19392 9036
rect 19392 9016 19394 9036
rect 20074 9016 20130 9072
rect 19449 8730 19505 8732
rect 19529 8730 19585 8732
rect 19609 8730 19665 8732
rect 19689 8730 19745 8732
rect 19449 8678 19475 8730
rect 19475 8678 19505 8730
rect 19529 8678 19539 8730
rect 19539 8678 19585 8730
rect 19609 8678 19655 8730
rect 19655 8678 19665 8730
rect 19689 8678 19719 8730
rect 19719 8678 19745 8730
rect 19449 8676 19505 8678
rect 19529 8676 19585 8678
rect 19609 8676 19665 8678
rect 19689 8676 19745 8678
rect 19154 8064 19210 8120
rect 19246 6704 19302 6760
rect 18234 3984 18290 4040
rect 19890 7792 19946 7848
rect 19449 7642 19505 7644
rect 19529 7642 19585 7644
rect 19609 7642 19665 7644
rect 19689 7642 19745 7644
rect 19449 7590 19475 7642
rect 19475 7590 19505 7642
rect 19529 7590 19539 7642
rect 19539 7590 19585 7642
rect 19609 7590 19655 7642
rect 19655 7590 19665 7642
rect 19689 7590 19719 7642
rect 19719 7590 19745 7642
rect 19449 7588 19505 7590
rect 19529 7588 19585 7590
rect 19609 7588 19665 7590
rect 19689 7588 19745 7590
rect 19449 6554 19505 6556
rect 19529 6554 19585 6556
rect 19609 6554 19665 6556
rect 19689 6554 19745 6556
rect 19449 6502 19475 6554
rect 19475 6502 19505 6554
rect 19529 6502 19539 6554
rect 19539 6502 19585 6554
rect 19609 6502 19655 6554
rect 19655 6502 19665 6554
rect 19689 6502 19719 6554
rect 19719 6502 19745 6554
rect 19449 6500 19505 6502
rect 19529 6500 19585 6502
rect 19609 6500 19665 6502
rect 19689 6500 19745 6502
rect 19614 5888 19670 5944
rect 19062 5344 19118 5400
rect 20534 12144 20590 12200
rect 20442 12008 20498 12064
rect 20442 9560 20498 9616
rect 19982 6296 20038 6352
rect 19982 6060 19984 6080
rect 19984 6060 20036 6080
rect 20036 6060 20038 6080
rect 19982 6024 20038 6060
rect 19890 5480 19946 5536
rect 19449 5466 19505 5468
rect 19529 5466 19585 5468
rect 19609 5466 19665 5468
rect 19689 5466 19745 5468
rect 19449 5414 19475 5466
rect 19475 5414 19505 5466
rect 19529 5414 19539 5466
rect 19539 5414 19585 5466
rect 19609 5414 19655 5466
rect 19655 5414 19665 5466
rect 19689 5414 19719 5466
rect 19719 5414 19745 5466
rect 19449 5412 19505 5414
rect 19529 5412 19585 5414
rect 19609 5412 19665 5414
rect 19689 5412 19745 5414
rect 19449 4378 19505 4380
rect 19529 4378 19585 4380
rect 19609 4378 19665 4380
rect 19689 4378 19745 4380
rect 19449 4326 19475 4378
rect 19475 4326 19505 4378
rect 19529 4326 19539 4378
rect 19539 4326 19585 4378
rect 19609 4326 19655 4378
rect 19655 4326 19665 4378
rect 19689 4326 19719 4378
rect 19719 4326 19745 4378
rect 19449 4324 19505 4326
rect 19529 4324 19585 4326
rect 19609 4324 19665 4326
rect 19689 4324 19745 4326
rect 18878 2488 18934 2544
rect 19449 3290 19505 3292
rect 19529 3290 19585 3292
rect 19609 3290 19665 3292
rect 19689 3290 19745 3292
rect 19449 3238 19475 3290
rect 19475 3238 19505 3290
rect 19529 3238 19539 3290
rect 19539 3238 19585 3290
rect 19609 3238 19655 3290
rect 19655 3238 19665 3290
rect 19689 3238 19719 3290
rect 19719 3238 19745 3290
rect 19449 3236 19505 3238
rect 19529 3236 19585 3238
rect 19609 3236 19665 3238
rect 19689 3236 19745 3238
rect 20258 5616 20314 5672
rect 20166 3576 20222 3632
rect 20350 2896 20406 2952
rect 21454 12688 21510 12744
rect 20902 10784 20958 10840
rect 20534 4800 20590 4856
rect 20810 6860 20866 6896
rect 20810 6840 20812 6860
rect 20812 6840 20864 6860
rect 20864 6840 20866 6860
rect 21178 10532 21234 10568
rect 21178 10512 21180 10532
rect 21180 10512 21232 10532
rect 21232 10512 21234 10532
rect 20994 8200 21050 8256
rect 21270 8200 21326 8256
rect 22006 18672 22062 18728
rect 21546 11600 21602 11656
rect 22282 17992 22338 18048
rect 22466 17312 22522 17368
rect 22466 16632 22522 16688
rect 21362 8064 21418 8120
rect 20994 7520 21050 7576
rect 20718 5516 20720 5536
rect 20720 5516 20772 5536
rect 20772 5516 20774 5536
rect 20718 5480 20774 5516
rect 20626 4256 20682 4312
rect 21454 7520 21510 7576
rect 21270 6840 21326 6896
rect 21178 5752 21234 5808
rect 22006 8744 22062 8800
rect 21822 3848 21878 3904
rect 22742 8472 22798 8528
rect 22742 6840 22798 6896
rect 22466 6160 22522 6216
rect 22742 5888 22798 5944
rect 22926 6296 22982 6352
rect 22834 5480 22890 5536
rect 21730 3032 21786 3088
rect 19449 2202 19505 2204
rect 19529 2202 19585 2204
rect 19609 2202 19665 2204
rect 19689 2202 19745 2204
rect 19449 2150 19475 2202
rect 19475 2150 19505 2202
rect 19529 2150 19539 2202
rect 19539 2150 19585 2202
rect 19609 2150 19655 2202
rect 19655 2150 19665 2202
rect 19689 2150 19719 2202
rect 19719 2150 19745 2202
rect 19449 2148 19505 2150
rect 19529 2148 19585 2150
rect 19609 2148 19665 2150
rect 19689 2148 19745 2150
rect 22374 1536 22430 1592
rect 19338 856 19394 912
rect 23018 312 23074 368
<< metal3 >>
rect 20345 24034 20411 24037
rect 23920 24034 24400 24064
rect 20345 24032 24400 24034
rect 20345 23976 20350 24032
rect 20406 23976 24400 24032
rect 20345 23974 24400 23976
rect 20345 23971 20411 23974
rect 23920 23944 24400 23974
rect 19241 23354 19307 23357
rect 23920 23354 24400 23384
rect 19241 23352 24400 23354
rect 19241 23296 19246 23352
rect 19302 23296 24400 23352
rect 19241 23294 24400 23296
rect 19241 23291 19307 23294
rect 23920 23264 24400 23294
rect 19149 22674 19215 22677
rect 23920 22674 24400 22704
rect 19149 22672 24400 22674
rect 19149 22616 19154 22672
rect 19210 22616 24400 22672
rect 19149 22614 24400 22616
rect 19149 22611 19215 22614
rect 23920 22584 24400 22614
rect 19885 21994 19951 21997
rect 23920 21994 24400 22024
rect 19885 21992 24400 21994
rect 19885 21936 19890 21992
rect 19946 21936 24400 21992
rect 19885 21934 24400 21936
rect 19885 21931 19951 21934
rect 23920 21904 24400 21934
rect 4642 21792 4962 21793
rect 4642 21728 4650 21792
rect 4714 21728 4730 21792
rect 4794 21728 4810 21792
rect 4874 21728 4890 21792
rect 4954 21728 4962 21792
rect 4642 21727 4962 21728
rect 12040 21792 12360 21793
rect 12040 21728 12048 21792
rect 12112 21728 12128 21792
rect 12192 21728 12208 21792
rect 12272 21728 12288 21792
rect 12352 21728 12360 21792
rect 12040 21727 12360 21728
rect 19437 21792 19757 21793
rect 19437 21728 19445 21792
rect 19509 21728 19525 21792
rect 19589 21728 19605 21792
rect 19669 21728 19685 21792
rect 19749 21728 19757 21792
rect 19437 21727 19757 21728
rect 2589 21586 2655 21589
rect 9029 21586 9095 21589
rect 2589 21584 9095 21586
rect 2589 21528 2594 21584
rect 2650 21528 9034 21584
rect 9090 21528 9095 21584
rect 2589 21526 9095 21528
rect 2589 21523 2655 21526
rect 9029 21523 9095 21526
rect 0 21314 480 21344
rect 3969 21314 4035 21317
rect 0 21312 4035 21314
rect 0 21256 3974 21312
rect 4030 21256 4035 21312
rect 0 21254 4035 21256
rect 0 21224 480 21254
rect 3969 21251 4035 21254
rect 19241 21314 19307 21317
rect 23920 21314 24400 21344
rect 19241 21312 24400 21314
rect 19241 21256 19246 21312
rect 19302 21256 24400 21312
rect 19241 21254 24400 21256
rect 19241 21251 19307 21254
rect 8341 21248 8661 21249
rect 8341 21184 8349 21248
rect 8413 21184 8429 21248
rect 8493 21184 8509 21248
rect 8573 21184 8589 21248
rect 8653 21184 8661 21248
rect 8341 21183 8661 21184
rect 15738 21248 16058 21249
rect 15738 21184 15746 21248
rect 15810 21184 15826 21248
rect 15890 21184 15906 21248
rect 15970 21184 15986 21248
rect 16050 21184 16058 21248
rect 23920 21224 24400 21254
rect 15738 21183 16058 21184
rect 1393 21042 1459 21045
rect 7598 21042 7604 21044
rect 1393 21040 7604 21042
rect 1393 20984 1398 21040
rect 1454 20984 7604 21040
rect 1393 20982 7604 20984
rect 1393 20979 1459 20982
rect 7598 20980 7604 20982
rect 7668 20980 7674 21044
rect 14825 20770 14891 20773
rect 16941 20772 17007 20773
rect 20529 20772 20595 20773
rect 14958 20770 14964 20772
rect 14825 20768 14964 20770
rect 14825 20712 14830 20768
rect 14886 20712 14964 20768
rect 14825 20710 14964 20712
rect 14825 20707 14891 20710
rect 14958 20708 14964 20710
rect 15028 20708 15034 20772
rect 16941 20768 16988 20772
rect 17052 20770 17058 20772
rect 20478 20770 20484 20772
rect 16941 20712 16946 20768
rect 16941 20708 16988 20712
rect 17052 20710 17098 20770
rect 20438 20710 20484 20770
rect 20548 20768 20595 20772
rect 20590 20712 20595 20768
rect 17052 20708 17058 20710
rect 20478 20708 20484 20710
rect 20548 20708 20595 20712
rect 16941 20707 17007 20708
rect 20529 20707 20595 20708
rect 4642 20704 4962 20705
rect 4642 20640 4650 20704
rect 4714 20640 4730 20704
rect 4794 20640 4810 20704
rect 4874 20640 4890 20704
rect 4954 20640 4962 20704
rect 4642 20639 4962 20640
rect 12040 20704 12360 20705
rect 12040 20640 12048 20704
rect 12112 20640 12128 20704
rect 12192 20640 12208 20704
rect 12272 20640 12288 20704
rect 12352 20640 12360 20704
rect 12040 20639 12360 20640
rect 19437 20704 19757 20705
rect 19437 20640 19445 20704
rect 19509 20640 19525 20704
rect 19589 20640 19605 20704
rect 19669 20640 19685 20704
rect 19749 20640 19757 20704
rect 19437 20639 19757 20640
rect 19977 20634 20043 20637
rect 23920 20634 24400 20664
rect 19977 20632 24400 20634
rect 19977 20576 19982 20632
rect 20038 20576 24400 20632
rect 19977 20574 24400 20576
rect 19977 20571 20043 20574
rect 23920 20544 24400 20574
rect 7598 20300 7604 20364
rect 7668 20362 7674 20364
rect 12709 20362 12775 20365
rect 7668 20360 12775 20362
rect 7668 20304 12714 20360
rect 12770 20304 12775 20360
rect 7668 20302 12775 20304
rect 7668 20300 7674 20302
rect 12709 20299 12775 20302
rect 8341 20160 8661 20161
rect 8341 20096 8349 20160
rect 8413 20096 8429 20160
rect 8493 20096 8509 20160
rect 8573 20096 8589 20160
rect 8653 20096 8661 20160
rect 8341 20095 8661 20096
rect 15738 20160 16058 20161
rect 15738 20096 15746 20160
rect 15810 20096 15826 20160
rect 15890 20096 15906 20160
rect 15970 20096 15986 20160
rect 16050 20096 16058 20160
rect 15738 20095 16058 20096
rect 19241 20090 19307 20093
rect 23920 20090 24400 20120
rect 19241 20088 24400 20090
rect 19241 20032 19246 20088
rect 19302 20032 24400 20088
rect 19241 20030 24400 20032
rect 19241 20027 19307 20030
rect 23920 20000 24400 20030
rect 5942 19892 5948 19956
rect 6012 19954 6018 19956
rect 16205 19954 16271 19957
rect 6012 19952 16271 19954
rect 6012 19896 16210 19952
rect 16266 19896 16271 19952
rect 6012 19894 16271 19896
rect 6012 19892 6018 19894
rect 16205 19891 16271 19894
rect 8109 19818 8175 19821
rect 8569 19818 8635 19821
rect 8109 19816 8635 19818
rect 8109 19760 8114 19816
rect 8170 19760 8574 19816
rect 8630 19760 8635 19816
rect 8109 19758 8635 19760
rect 8109 19755 8175 19758
rect 8569 19755 8635 19758
rect 12433 19818 12499 19821
rect 18781 19818 18847 19821
rect 12433 19816 18847 19818
rect 12433 19760 12438 19816
rect 12494 19760 18786 19816
rect 18842 19760 18847 19816
rect 12433 19758 18847 19760
rect 12433 19755 12499 19758
rect 18781 19755 18847 19758
rect 19701 19818 19767 19821
rect 20110 19818 20116 19820
rect 19701 19816 20116 19818
rect 19701 19760 19706 19816
rect 19762 19760 20116 19816
rect 19701 19758 20116 19760
rect 19701 19755 19767 19758
rect 20110 19756 20116 19758
rect 20180 19756 20186 19820
rect 5993 19682 6059 19685
rect 8937 19682 9003 19685
rect 5993 19680 9003 19682
rect 5993 19624 5998 19680
rect 6054 19624 8942 19680
rect 8998 19624 9003 19680
rect 5993 19622 9003 19624
rect 5993 19619 6059 19622
rect 8937 19619 9003 19622
rect 4642 19616 4962 19617
rect 4642 19552 4650 19616
rect 4714 19552 4730 19616
rect 4794 19552 4810 19616
rect 4874 19552 4890 19616
rect 4954 19552 4962 19616
rect 4642 19551 4962 19552
rect 12040 19616 12360 19617
rect 12040 19552 12048 19616
rect 12112 19552 12128 19616
rect 12192 19552 12208 19616
rect 12272 19552 12288 19616
rect 12352 19552 12360 19616
rect 12040 19551 12360 19552
rect 19437 19616 19757 19617
rect 19437 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19605 19616
rect 19669 19552 19685 19616
rect 19749 19552 19757 19616
rect 19437 19551 19757 19552
rect 8201 19546 8267 19549
rect 10409 19546 10475 19549
rect 8201 19544 10475 19546
rect 8201 19488 8206 19544
rect 8262 19488 10414 19544
rect 10470 19488 10475 19544
rect 8201 19486 10475 19488
rect 8201 19483 8267 19486
rect 10409 19483 10475 19486
rect 12525 19546 12591 19549
rect 15009 19546 15075 19549
rect 12525 19544 15075 19546
rect 12525 19488 12530 19544
rect 12586 19488 15014 19544
rect 15070 19488 15075 19544
rect 12525 19486 15075 19488
rect 12525 19483 12591 19486
rect 15009 19483 15075 19486
rect 13629 19410 13695 19413
rect 15745 19410 15811 19413
rect 13629 19408 15811 19410
rect 13629 19352 13634 19408
rect 13690 19352 15750 19408
rect 15806 19352 15811 19408
rect 13629 19350 15811 19352
rect 13629 19347 13695 19350
rect 15745 19347 15811 19350
rect 19885 19412 19951 19413
rect 19885 19408 19932 19412
rect 19996 19410 20002 19412
rect 20621 19410 20687 19413
rect 23920 19410 24400 19440
rect 19885 19352 19890 19408
rect 19885 19348 19932 19352
rect 19996 19350 20042 19410
rect 20621 19408 24400 19410
rect 20621 19352 20626 19408
rect 20682 19352 24400 19408
rect 20621 19350 24400 19352
rect 19996 19348 20002 19350
rect 19885 19347 19951 19348
rect 20621 19347 20687 19350
rect 23920 19320 24400 19350
rect 8886 19212 8892 19276
rect 8956 19274 8962 19276
rect 20161 19274 20227 19277
rect 8956 19272 20227 19274
rect 8956 19216 20166 19272
rect 20222 19216 20227 19272
rect 8956 19214 20227 19216
rect 8956 19212 8962 19214
rect 20161 19211 20227 19214
rect 8341 19072 8661 19073
rect 8341 19008 8349 19072
rect 8413 19008 8429 19072
rect 8493 19008 8509 19072
rect 8573 19008 8589 19072
rect 8653 19008 8661 19072
rect 8341 19007 8661 19008
rect 15738 19072 16058 19073
rect 15738 19008 15746 19072
rect 15810 19008 15826 19072
rect 15890 19008 15906 19072
rect 15970 19008 15986 19072
rect 16050 19008 16058 19072
rect 15738 19007 16058 19008
rect 10409 19002 10475 19005
rect 15285 19002 15351 19005
rect 10409 19000 15351 19002
rect 10409 18944 10414 19000
rect 10470 18944 15290 19000
rect 15346 18944 15351 19000
rect 10409 18942 15351 18944
rect 10409 18939 10475 18942
rect 15285 18939 15351 18942
rect 4429 18868 4495 18869
rect 4429 18864 4476 18868
rect 4540 18866 4546 18868
rect 11421 18866 11487 18869
rect 15653 18866 15719 18869
rect 4429 18808 4434 18864
rect 4429 18804 4476 18808
rect 4540 18806 4586 18866
rect 11421 18864 15719 18866
rect 11421 18808 11426 18864
rect 11482 18808 15658 18864
rect 15714 18808 15719 18864
rect 11421 18806 15719 18808
rect 4540 18804 4546 18806
rect 4429 18803 4495 18804
rect 11421 18803 11487 18806
rect 15653 18803 15719 18806
rect 1761 18730 1827 18733
rect 9397 18730 9463 18733
rect 12433 18730 12499 18733
rect 1761 18728 5136 18730
rect 1761 18672 1766 18728
rect 1822 18672 5136 18728
rect 1761 18670 5136 18672
rect 1761 18667 1827 18670
rect 5076 18597 5136 18670
rect 9397 18728 12499 18730
rect 9397 18672 9402 18728
rect 9458 18672 12438 18728
rect 12494 18672 12499 18728
rect 9397 18670 12499 18672
rect 9397 18667 9463 18670
rect 12433 18667 12499 18670
rect 22001 18730 22067 18733
rect 23920 18730 24400 18760
rect 22001 18728 24400 18730
rect 22001 18672 22006 18728
rect 22062 18672 24400 18728
rect 22001 18670 24400 18672
rect 22001 18667 22067 18670
rect 23920 18640 24400 18670
rect 5073 18594 5139 18597
rect 5206 18594 5212 18596
rect 5073 18592 5212 18594
rect 5073 18536 5078 18592
rect 5134 18536 5212 18592
rect 5073 18534 5212 18536
rect 5073 18531 5139 18534
rect 5206 18532 5212 18534
rect 5276 18532 5282 18596
rect 4642 18528 4962 18529
rect 4642 18464 4650 18528
rect 4714 18464 4730 18528
rect 4794 18464 4810 18528
rect 4874 18464 4890 18528
rect 4954 18464 4962 18528
rect 4642 18463 4962 18464
rect 12040 18528 12360 18529
rect 12040 18464 12048 18528
rect 12112 18464 12128 18528
rect 12192 18464 12208 18528
rect 12272 18464 12288 18528
rect 12352 18464 12360 18528
rect 12040 18463 12360 18464
rect 19437 18528 19757 18529
rect 19437 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19605 18528
rect 19669 18464 19685 18528
rect 19749 18464 19757 18528
rect 19437 18463 19757 18464
rect 7005 18458 7071 18461
rect 12985 18458 13051 18461
rect 16113 18458 16179 18461
rect 7005 18456 10058 18458
rect 7005 18400 7010 18456
rect 7066 18400 10058 18456
rect 7005 18398 10058 18400
rect 7005 18395 7071 18398
rect 9998 18322 10058 18398
rect 12985 18456 16179 18458
rect 12985 18400 12990 18456
rect 13046 18400 16118 18456
rect 16174 18400 16179 18456
rect 12985 18398 16179 18400
rect 12985 18395 13051 18398
rect 16113 18395 16179 18398
rect 12525 18322 12591 18325
rect 9998 18320 12591 18322
rect 9998 18264 12530 18320
rect 12586 18264 12591 18320
rect 9998 18262 12591 18264
rect 12525 18259 12591 18262
rect 12893 18322 12959 18325
rect 15929 18322 15995 18325
rect 12893 18320 15995 18322
rect 12893 18264 12898 18320
rect 12954 18264 15934 18320
rect 15990 18264 15995 18320
rect 12893 18262 15995 18264
rect 12893 18259 12959 18262
rect 15929 18259 15995 18262
rect 16113 18322 16179 18325
rect 16757 18322 16823 18325
rect 16113 18320 16823 18322
rect 16113 18264 16118 18320
rect 16174 18264 16762 18320
rect 16818 18264 16823 18320
rect 16113 18262 16823 18264
rect 16113 18259 16179 18262
rect 16757 18259 16823 18262
rect 17677 18324 17743 18325
rect 17677 18320 17724 18324
rect 17788 18322 17794 18324
rect 20529 18322 20595 18325
rect 20662 18322 20668 18324
rect 17677 18264 17682 18320
rect 17677 18260 17724 18264
rect 17788 18262 17834 18322
rect 20529 18320 20668 18322
rect 20529 18264 20534 18320
rect 20590 18264 20668 18320
rect 20529 18262 20668 18264
rect 17788 18260 17794 18262
rect 17677 18259 17743 18260
rect 20529 18259 20595 18262
rect 20662 18260 20668 18262
rect 20732 18322 20738 18324
rect 21725 18322 21791 18325
rect 20732 18320 21791 18322
rect 20732 18264 21730 18320
rect 21786 18264 21791 18320
rect 20732 18262 21791 18264
rect 20732 18260 20738 18262
rect 21725 18259 21791 18262
rect 9305 18186 9371 18189
rect 4800 18184 9371 18186
rect 4800 18128 9310 18184
rect 9366 18128 9371 18184
rect 4800 18126 9371 18128
rect 4800 18053 4860 18126
rect 9305 18123 9371 18126
rect 9622 18124 9628 18188
rect 9692 18186 9698 18188
rect 9949 18186 10015 18189
rect 9692 18184 10015 18186
rect 9692 18128 9954 18184
rect 10010 18128 10015 18184
rect 9692 18126 10015 18128
rect 9692 18124 9698 18126
rect 9949 18123 10015 18126
rect 14825 18186 14891 18189
rect 17401 18186 17467 18189
rect 14825 18184 17467 18186
rect 14825 18128 14830 18184
rect 14886 18128 17406 18184
rect 17462 18128 17467 18184
rect 14825 18126 17467 18128
rect 14825 18123 14891 18126
rect 17401 18123 17467 18126
rect 4286 17988 4292 18052
rect 4356 18050 4362 18052
rect 4797 18050 4863 18053
rect 4356 18048 4863 18050
rect 4356 17992 4802 18048
rect 4858 17992 4863 18048
rect 4356 17990 4863 17992
rect 4356 17988 4362 17990
rect 4797 17987 4863 17990
rect 9673 18050 9739 18053
rect 9806 18050 9812 18052
rect 9673 18048 9812 18050
rect 9673 17992 9678 18048
rect 9734 17992 9812 18048
rect 9673 17990 9812 17992
rect 9673 17987 9739 17990
rect 9806 17988 9812 17990
rect 9876 17988 9882 18052
rect 20069 18050 20135 18053
rect 20294 18050 20300 18052
rect 20069 18048 20300 18050
rect 20069 17992 20074 18048
rect 20130 17992 20300 18048
rect 20069 17990 20300 17992
rect 20069 17987 20135 17990
rect 20294 17988 20300 17990
rect 20364 17988 20370 18052
rect 22277 18050 22343 18053
rect 23920 18050 24400 18080
rect 22277 18048 24400 18050
rect 22277 17992 22282 18048
rect 22338 17992 24400 18048
rect 22277 17990 24400 17992
rect 22277 17987 22343 17990
rect 8341 17984 8661 17985
rect 8341 17920 8349 17984
rect 8413 17920 8429 17984
rect 8493 17920 8509 17984
rect 8573 17920 8589 17984
rect 8653 17920 8661 17984
rect 8341 17919 8661 17920
rect 15738 17984 16058 17985
rect 15738 17920 15746 17984
rect 15810 17920 15826 17984
rect 15890 17920 15906 17984
rect 15970 17920 15986 17984
rect 16050 17920 16058 17984
rect 23920 17960 24400 17990
rect 15738 17919 16058 17920
rect 1669 17778 1735 17781
rect 7925 17778 7991 17781
rect 1669 17776 7991 17778
rect 1669 17720 1674 17776
rect 1730 17720 7930 17776
rect 7986 17720 7991 17776
rect 1669 17718 7991 17720
rect 1669 17715 1735 17718
rect 7925 17715 7991 17718
rect 2589 17642 2655 17645
rect 2957 17642 3023 17645
rect 2589 17640 3023 17642
rect 2589 17584 2594 17640
rect 2650 17584 2962 17640
rect 3018 17584 3023 17640
rect 2589 17582 3023 17584
rect 2589 17579 2655 17582
rect 2957 17579 3023 17582
rect 10409 17642 10475 17645
rect 15561 17642 15627 17645
rect 10409 17640 15627 17642
rect 10409 17584 10414 17640
rect 10470 17584 15566 17640
rect 15622 17584 15627 17640
rect 10409 17582 15627 17584
rect 10409 17579 10475 17582
rect 15561 17579 15627 17582
rect 4642 17440 4962 17441
rect 4642 17376 4650 17440
rect 4714 17376 4730 17440
rect 4794 17376 4810 17440
rect 4874 17376 4890 17440
rect 4954 17376 4962 17440
rect 4642 17375 4962 17376
rect 12040 17440 12360 17441
rect 12040 17376 12048 17440
rect 12112 17376 12128 17440
rect 12192 17376 12208 17440
rect 12272 17376 12288 17440
rect 12352 17376 12360 17440
rect 12040 17375 12360 17376
rect 19437 17440 19757 17441
rect 19437 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19605 17440
rect 19669 17376 19685 17440
rect 19749 17376 19757 17440
rect 19437 17375 19757 17376
rect 22461 17370 22527 17373
rect 23920 17370 24400 17400
rect 22461 17368 24400 17370
rect 22461 17312 22466 17368
rect 22522 17312 24400 17368
rect 22461 17310 24400 17312
rect 22461 17307 22527 17310
rect 23920 17280 24400 17310
rect 2773 17234 2839 17237
rect 11053 17234 11119 17237
rect 2773 17232 11119 17234
rect 2773 17176 2778 17232
rect 2834 17176 11058 17232
rect 11114 17176 11119 17232
rect 2773 17174 11119 17176
rect 2773 17171 2839 17174
rect 11053 17171 11119 17174
rect 17217 17234 17283 17237
rect 20161 17234 20227 17237
rect 17217 17232 20227 17234
rect 17217 17176 17222 17232
rect 17278 17176 20166 17232
rect 20222 17176 20227 17232
rect 17217 17174 20227 17176
rect 17217 17171 17283 17174
rect 20161 17171 20227 17174
rect 3601 17098 3667 17101
rect 4245 17098 4311 17101
rect 3601 17096 4311 17098
rect 3601 17040 3606 17096
rect 3662 17040 4250 17096
rect 4306 17040 4311 17096
rect 3601 17038 4311 17040
rect 3601 17035 3667 17038
rect 4245 17035 4311 17038
rect 4470 17036 4476 17100
rect 4540 17098 4546 17100
rect 4981 17098 5047 17101
rect 4540 17096 5047 17098
rect 4540 17040 4986 17096
rect 5042 17040 5047 17096
rect 4540 17038 5047 17040
rect 4540 17036 4546 17038
rect 4981 17035 5047 17038
rect 10777 17098 10843 17101
rect 12985 17098 13051 17101
rect 10777 17096 13051 17098
rect 10777 17040 10782 17096
rect 10838 17040 12990 17096
rect 13046 17040 13051 17096
rect 10777 17038 13051 17040
rect 10777 17035 10843 17038
rect 12985 17035 13051 17038
rect 8341 16896 8661 16897
rect 8341 16832 8349 16896
rect 8413 16832 8429 16896
rect 8493 16832 8509 16896
rect 8573 16832 8589 16896
rect 8653 16832 8661 16896
rect 8341 16831 8661 16832
rect 15738 16896 16058 16897
rect 15738 16832 15746 16896
rect 15810 16832 15826 16896
rect 15890 16832 15906 16896
rect 15970 16832 15986 16896
rect 16050 16832 16058 16896
rect 15738 16831 16058 16832
rect 3877 16826 3943 16829
rect 5073 16826 5139 16829
rect 5993 16826 6059 16829
rect 3877 16824 6059 16826
rect 3877 16768 3882 16824
rect 3938 16768 5078 16824
rect 5134 16768 5998 16824
rect 6054 16768 6059 16824
rect 3877 16766 6059 16768
rect 3877 16763 3943 16766
rect 5073 16763 5139 16766
rect 5993 16763 6059 16766
rect 2773 16690 2839 16693
rect 8293 16690 8359 16693
rect 2773 16688 8359 16690
rect 2773 16632 2778 16688
rect 2834 16632 8298 16688
rect 8354 16632 8359 16688
rect 2773 16630 8359 16632
rect 2773 16627 2839 16630
rect 8293 16627 8359 16630
rect 8845 16690 8911 16693
rect 9857 16690 9923 16693
rect 8845 16688 9923 16690
rect 8845 16632 8850 16688
rect 8906 16632 9862 16688
rect 9918 16632 9923 16688
rect 8845 16630 9923 16632
rect 8845 16627 8911 16630
rect 9857 16627 9923 16630
rect 11605 16690 11671 16693
rect 15101 16690 15167 16693
rect 11605 16688 15167 16690
rect 11605 16632 11610 16688
rect 11666 16632 15106 16688
rect 15162 16632 15167 16688
rect 11605 16630 15167 16632
rect 11605 16627 11671 16630
rect 15101 16627 15167 16630
rect 22461 16690 22527 16693
rect 23920 16690 24400 16720
rect 22461 16688 24400 16690
rect 22461 16632 22466 16688
rect 22522 16632 24400 16688
rect 22461 16630 24400 16632
rect 22461 16627 22527 16630
rect 23920 16600 24400 16630
rect 5717 16554 5783 16557
rect 9254 16554 9260 16556
rect 5717 16552 9260 16554
rect 5717 16496 5722 16552
rect 5778 16496 9260 16552
rect 5717 16494 9260 16496
rect 5717 16491 5783 16494
rect 9254 16492 9260 16494
rect 9324 16554 9330 16556
rect 9622 16554 9628 16556
rect 9324 16494 9628 16554
rect 9324 16492 9330 16494
rect 9622 16492 9628 16494
rect 9692 16492 9698 16556
rect 11053 16554 11119 16557
rect 14733 16554 14799 16557
rect 16849 16554 16915 16557
rect 11053 16552 12496 16554
rect 11053 16496 11058 16552
rect 11114 16496 12496 16552
rect 11053 16494 12496 16496
rect 11053 16491 11119 16494
rect 9673 16418 9739 16421
rect 10593 16418 10659 16421
rect 9673 16416 10659 16418
rect 9673 16360 9678 16416
rect 9734 16360 10598 16416
rect 10654 16360 10659 16416
rect 9673 16358 10659 16360
rect 12436 16418 12496 16494
rect 14733 16552 16915 16554
rect 14733 16496 14738 16552
rect 14794 16496 16854 16552
rect 16910 16496 16915 16552
rect 14733 16494 16915 16496
rect 14733 16491 14799 16494
rect 16849 16491 16915 16494
rect 18781 16418 18847 16421
rect 12436 16416 18847 16418
rect 12436 16360 18786 16416
rect 18842 16360 18847 16416
rect 12436 16358 18847 16360
rect 9673 16355 9739 16358
rect 10593 16355 10659 16358
rect 18781 16355 18847 16358
rect 4642 16352 4962 16353
rect 4642 16288 4650 16352
rect 4714 16288 4730 16352
rect 4794 16288 4810 16352
rect 4874 16288 4890 16352
rect 4954 16288 4962 16352
rect 4642 16287 4962 16288
rect 12040 16352 12360 16353
rect 12040 16288 12048 16352
rect 12112 16288 12128 16352
rect 12192 16288 12208 16352
rect 12272 16288 12288 16352
rect 12352 16288 12360 16352
rect 12040 16287 12360 16288
rect 19437 16352 19757 16353
rect 19437 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19605 16352
rect 19669 16288 19685 16352
rect 19749 16288 19757 16352
rect 19437 16287 19757 16288
rect 9765 16284 9831 16285
rect 9765 16280 9812 16284
rect 9876 16282 9882 16284
rect 9765 16224 9770 16280
rect 9765 16220 9812 16224
rect 9876 16222 9922 16282
rect 9876 16220 9882 16222
rect 9765 16219 9831 16220
rect 5073 16146 5139 16149
rect 6361 16146 6427 16149
rect 5073 16144 6427 16146
rect 5073 16088 5078 16144
rect 5134 16088 6366 16144
rect 6422 16088 6427 16144
rect 5073 16086 6427 16088
rect 5073 16083 5139 16086
rect 6361 16083 6427 16086
rect 7189 16146 7255 16149
rect 8845 16146 8911 16149
rect 10685 16146 10751 16149
rect 7189 16144 10751 16146
rect 7189 16088 7194 16144
rect 7250 16088 8850 16144
rect 8906 16088 10690 16144
rect 10746 16088 10751 16144
rect 7189 16086 10751 16088
rect 7189 16083 7255 16086
rect 8845 16083 8911 16086
rect 10685 16083 10751 16086
rect 11094 16084 11100 16148
rect 11164 16146 11170 16148
rect 18689 16146 18755 16149
rect 11164 16144 18755 16146
rect 11164 16088 18694 16144
rect 18750 16088 18755 16144
rect 11164 16086 18755 16088
rect 11164 16084 11170 16086
rect 18689 16083 18755 16086
rect 18965 16146 19031 16149
rect 23920 16146 24400 16176
rect 18965 16144 24400 16146
rect 18965 16088 18970 16144
rect 19026 16088 24400 16144
rect 18965 16086 24400 16088
rect 18965 16083 19031 16086
rect 23920 16056 24400 16086
rect 8017 16010 8083 16013
rect 11237 16010 11303 16013
rect 8017 16008 11303 16010
rect 8017 15952 8022 16008
rect 8078 15952 11242 16008
rect 11298 15952 11303 16008
rect 8017 15950 11303 15952
rect 8017 15947 8083 15950
rect 11237 15947 11303 15950
rect 11605 16010 11671 16013
rect 13629 16010 13695 16013
rect 15653 16010 15719 16013
rect 11605 16008 15719 16010
rect 11605 15952 11610 16008
rect 11666 15952 13634 16008
rect 13690 15952 15658 16008
rect 15714 15952 15719 16008
rect 11605 15950 15719 15952
rect 11605 15947 11671 15950
rect 13629 15947 13695 15950
rect 15653 15947 15719 15950
rect 4705 15874 4771 15877
rect 5625 15874 5691 15877
rect 4705 15872 5691 15874
rect 4705 15816 4710 15872
rect 4766 15816 5630 15872
rect 5686 15816 5691 15872
rect 4705 15814 5691 15816
rect 4705 15811 4771 15814
rect 5625 15811 5691 15814
rect 8341 15808 8661 15809
rect 8341 15744 8349 15808
rect 8413 15744 8429 15808
rect 8493 15744 8509 15808
rect 8573 15744 8589 15808
rect 8653 15744 8661 15808
rect 8341 15743 8661 15744
rect 15738 15808 16058 15809
rect 15738 15744 15746 15808
rect 15810 15744 15826 15808
rect 15890 15744 15906 15808
rect 15970 15744 15986 15808
rect 16050 15744 16058 15808
rect 15738 15743 16058 15744
rect 4889 15738 4955 15741
rect 7189 15738 7255 15741
rect 4889 15736 7255 15738
rect 4889 15680 4894 15736
rect 4950 15680 7194 15736
rect 7250 15680 7255 15736
rect 4889 15678 7255 15680
rect 4889 15675 4955 15678
rect 7189 15675 7255 15678
rect 7966 15540 7972 15604
rect 8036 15602 8042 15604
rect 12525 15602 12591 15605
rect 8036 15600 12591 15602
rect 8036 15544 12530 15600
rect 12586 15544 12591 15600
rect 8036 15542 12591 15544
rect 8036 15540 8042 15542
rect 12525 15539 12591 15542
rect 15193 15466 15259 15469
rect 15510 15466 15516 15468
rect 15193 15464 15516 15466
rect 15193 15408 15198 15464
rect 15254 15408 15516 15464
rect 15193 15406 15516 15408
rect 15193 15403 15259 15406
rect 15510 15404 15516 15406
rect 15580 15466 15586 15468
rect 16021 15466 16087 15469
rect 15580 15464 16087 15466
rect 15580 15408 16026 15464
rect 16082 15408 16087 15464
rect 15580 15406 16087 15408
rect 15580 15404 15586 15406
rect 16021 15403 16087 15406
rect 19701 15466 19767 15469
rect 23920 15466 24400 15496
rect 19701 15464 24400 15466
rect 19701 15408 19706 15464
rect 19762 15408 24400 15464
rect 19701 15406 24400 15408
rect 19701 15403 19767 15406
rect 23920 15376 24400 15406
rect 8477 15330 8543 15333
rect 13813 15332 13879 15333
rect 9070 15330 9076 15332
rect 8477 15328 9076 15330
rect 8477 15272 8482 15328
rect 8538 15272 9076 15328
rect 8477 15270 9076 15272
rect 8477 15267 8543 15270
rect 9070 15268 9076 15270
rect 9140 15268 9146 15332
rect 13813 15328 13860 15332
rect 13924 15330 13930 15332
rect 13813 15272 13818 15328
rect 13813 15268 13860 15272
rect 13924 15270 13970 15330
rect 13924 15268 13930 15270
rect 13813 15267 13879 15268
rect 4642 15264 4962 15265
rect 0 15194 480 15224
rect 4642 15200 4650 15264
rect 4714 15200 4730 15264
rect 4794 15200 4810 15264
rect 4874 15200 4890 15264
rect 4954 15200 4962 15264
rect 4642 15199 4962 15200
rect 12040 15264 12360 15265
rect 12040 15200 12048 15264
rect 12112 15200 12128 15264
rect 12192 15200 12208 15264
rect 12272 15200 12288 15264
rect 12352 15200 12360 15264
rect 12040 15199 12360 15200
rect 19437 15264 19757 15265
rect 19437 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19605 15264
rect 19669 15200 19685 15264
rect 19749 15200 19757 15264
rect 19437 15199 19757 15200
rect 3325 15194 3391 15197
rect 0 15192 3391 15194
rect 0 15136 3330 15192
rect 3386 15136 3391 15192
rect 0 15134 3391 15136
rect 0 15104 480 15134
rect 3325 15131 3391 15134
rect 13537 15194 13603 15197
rect 16665 15194 16731 15197
rect 13537 15192 16731 15194
rect 13537 15136 13542 15192
rect 13598 15136 16670 15192
rect 16726 15136 16731 15192
rect 13537 15134 16731 15136
rect 13537 15131 13603 15134
rect 16665 15131 16731 15134
rect 10225 15060 10291 15061
rect 10174 15058 10180 15060
rect 10134 14998 10180 15058
rect 10244 15056 10291 15060
rect 10286 15000 10291 15056
rect 10174 14996 10180 14998
rect 10244 14996 10291 15000
rect 14774 14996 14780 15060
rect 14844 15058 14850 15060
rect 15745 15058 15811 15061
rect 14844 15056 15811 15058
rect 14844 15000 15750 15056
rect 15806 15000 15811 15056
rect 14844 14998 15811 15000
rect 14844 14996 14850 14998
rect 10225 14995 10291 14996
rect 15745 14995 15811 14998
rect 17401 15058 17467 15061
rect 21173 15058 21239 15061
rect 17401 15056 21239 15058
rect 17401 15000 17406 15056
rect 17462 15000 21178 15056
rect 21234 15000 21239 15056
rect 17401 14998 21239 15000
rect 17401 14995 17467 14998
rect 21173 14995 21239 14998
rect 8150 14860 8156 14924
rect 8220 14922 8226 14924
rect 16297 14922 16363 14925
rect 8220 14920 16363 14922
rect 8220 14864 16302 14920
rect 16358 14864 16363 14920
rect 8220 14862 16363 14864
rect 8220 14860 8226 14862
rect 16297 14859 16363 14862
rect 19793 14922 19859 14925
rect 19977 14922 20043 14925
rect 19793 14920 20043 14922
rect 19793 14864 19798 14920
rect 19854 14864 19982 14920
rect 20038 14864 20043 14920
rect 19793 14862 20043 14864
rect 19793 14859 19859 14862
rect 19977 14859 20043 14862
rect 4337 14786 4403 14789
rect 4470 14786 4476 14788
rect 4337 14784 4476 14786
rect 4337 14728 4342 14784
rect 4398 14728 4476 14784
rect 4337 14726 4476 14728
rect 4337 14723 4403 14726
rect 4470 14724 4476 14726
rect 4540 14786 4546 14788
rect 4613 14786 4679 14789
rect 4540 14784 4679 14786
rect 4540 14728 4618 14784
rect 4674 14728 4679 14784
rect 4540 14726 4679 14728
rect 4540 14724 4546 14726
rect 4613 14723 4679 14726
rect 5165 14786 5231 14789
rect 5441 14786 5507 14789
rect 5165 14784 5507 14786
rect 5165 14728 5170 14784
rect 5226 14728 5446 14784
rect 5502 14728 5507 14784
rect 5165 14726 5507 14728
rect 5165 14723 5231 14726
rect 5441 14723 5507 14726
rect 10501 14786 10567 14789
rect 12157 14786 12223 14789
rect 10501 14784 12223 14786
rect 10501 14728 10506 14784
rect 10562 14728 12162 14784
rect 12218 14728 12223 14784
rect 10501 14726 12223 14728
rect 10501 14723 10567 14726
rect 12157 14723 12223 14726
rect 18321 14786 18387 14789
rect 19333 14786 19399 14789
rect 23920 14786 24400 14816
rect 18321 14784 18522 14786
rect 18321 14728 18326 14784
rect 18382 14728 18522 14784
rect 18321 14726 18522 14728
rect 18321 14723 18387 14726
rect 8341 14720 8661 14721
rect 8341 14656 8349 14720
rect 8413 14656 8429 14720
rect 8493 14656 8509 14720
rect 8573 14656 8589 14720
rect 8653 14656 8661 14720
rect 8341 14655 8661 14656
rect 15738 14720 16058 14721
rect 15738 14656 15746 14720
rect 15810 14656 15826 14720
rect 15890 14656 15906 14720
rect 15970 14656 15986 14720
rect 16050 14656 16058 14720
rect 15738 14655 16058 14656
rect 17769 14650 17835 14653
rect 18321 14650 18387 14653
rect 17769 14648 18387 14650
rect 17769 14592 17774 14648
rect 17830 14592 18326 14648
rect 18382 14592 18387 14648
rect 17769 14590 18387 14592
rect 18462 14650 18522 14726
rect 19333 14784 24400 14786
rect 19333 14728 19338 14784
rect 19394 14728 24400 14784
rect 19333 14726 24400 14728
rect 19333 14723 19399 14726
rect 23920 14696 24400 14726
rect 20713 14650 20779 14653
rect 18462 14648 20779 14650
rect 18462 14592 20718 14648
rect 20774 14592 20779 14648
rect 18462 14590 20779 14592
rect 17769 14587 17835 14590
rect 18321 14587 18387 14590
rect 20713 14587 20779 14590
rect 3417 14514 3483 14517
rect 8569 14514 8635 14517
rect 3417 14512 8635 14514
rect 3417 14456 3422 14512
rect 3478 14456 8574 14512
rect 8630 14456 8635 14512
rect 3417 14454 8635 14456
rect 3417 14451 3483 14454
rect 8569 14451 8635 14454
rect 13445 14514 13511 14517
rect 15745 14514 15811 14517
rect 13445 14512 15811 14514
rect 13445 14456 13450 14512
rect 13506 14456 15750 14512
rect 15806 14456 15811 14512
rect 13445 14454 15811 14456
rect 13445 14451 13511 14454
rect 15745 14451 15811 14454
rect 17401 14514 17467 14517
rect 20437 14514 20503 14517
rect 17401 14512 20503 14514
rect 17401 14456 17406 14512
rect 17462 14456 20442 14512
rect 20498 14456 20503 14512
rect 17401 14454 20503 14456
rect 17401 14451 17467 14454
rect 20437 14451 20503 14454
rect 1853 14378 1919 14381
rect 8845 14378 8911 14381
rect 1853 14376 8911 14378
rect 1853 14320 1858 14376
rect 1914 14320 8850 14376
rect 8906 14320 8911 14376
rect 1853 14318 8911 14320
rect 1853 14315 1919 14318
rect 8845 14315 8911 14318
rect 10317 14378 10383 14381
rect 12341 14378 12407 14381
rect 10317 14376 12407 14378
rect 10317 14320 10322 14376
rect 10378 14320 12346 14376
rect 12402 14320 12407 14376
rect 10317 14318 12407 14320
rect 10317 14315 10383 14318
rect 12341 14315 12407 14318
rect 19333 14378 19399 14381
rect 19333 14376 23858 14378
rect 19333 14320 19338 14376
rect 19394 14320 23858 14376
rect 19333 14318 23858 14320
rect 19333 14315 19399 14318
rect 10412 14182 11944 14242
rect 4642 14176 4962 14177
rect 4642 14112 4650 14176
rect 4714 14112 4730 14176
rect 4794 14112 4810 14176
rect 4874 14112 4890 14176
rect 4954 14112 4962 14176
rect 4642 14111 4962 14112
rect 6821 14106 6887 14109
rect 5030 14104 6887 14106
rect 5030 14048 6826 14104
rect 6882 14048 6887 14104
rect 5030 14046 6887 14048
rect 4889 13970 4955 13973
rect 5030 13970 5090 14046
rect 6821 14043 6887 14046
rect 4889 13968 5090 13970
rect 4889 13912 4894 13968
rect 4950 13912 5090 13968
rect 4889 13910 5090 13912
rect 5901 13970 5967 13973
rect 10041 13970 10107 13973
rect 10412 13970 10472 14182
rect 5901 13968 6010 13970
rect 5901 13912 5906 13968
rect 5962 13912 6010 13968
rect 4889 13907 4955 13910
rect 5901 13907 6010 13912
rect 10041 13968 10472 13970
rect 10041 13912 10046 13968
rect 10102 13912 10472 13968
rect 10041 13910 10472 13912
rect 11884 13970 11944 14182
rect 13118 14180 13124 14244
rect 13188 14242 13194 14244
rect 16113 14242 16179 14245
rect 13188 14240 16179 14242
rect 13188 14184 16118 14240
rect 16174 14184 16179 14240
rect 13188 14182 16179 14184
rect 13188 14180 13194 14182
rect 16113 14179 16179 14182
rect 12040 14176 12360 14177
rect 12040 14112 12048 14176
rect 12112 14112 12128 14176
rect 12192 14112 12208 14176
rect 12272 14112 12288 14176
rect 12352 14112 12360 14176
rect 12040 14111 12360 14112
rect 19437 14176 19757 14177
rect 19437 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19605 14176
rect 19669 14112 19685 14176
rect 19749 14112 19757 14176
rect 19437 14111 19757 14112
rect 23798 14106 23858 14318
rect 23920 14106 24400 14136
rect 23798 14046 24400 14106
rect 23920 14016 24400 14046
rect 15101 13970 15167 13973
rect 11884 13968 15167 13970
rect 11884 13912 15106 13968
rect 15162 13912 15167 13968
rect 11884 13910 15167 13912
rect 10041 13907 10107 13910
rect 15101 13907 15167 13910
rect 4245 13834 4311 13837
rect 5165 13834 5231 13837
rect 4245 13832 5231 13834
rect 4245 13776 4250 13832
rect 4306 13776 5170 13832
rect 5226 13776 5231 13832
rect 4245 13774 5231 13776
rect 4245 13771 4311 13774
rect 5165 13771 5231 13774
rect 4245 13700 4311 13701
rect 5165 13700 5231 13701
rect 4245 13696 4292 13700
rect 4356 13698 4362 13700
rect 4245 13640 4250 13696
rect 4245 13636 4292 13640
rect 4356 13638 4402 13698
rect 5165 13696 5212 13700
rect 5276 13698 5282 13700
rect 5165 13640 5170 13696
rect 4356 13636 4362 13638
rect 5165 13636 5212 13640
rect 5276 13638 5322 13698
rect 5276 13636 5282 13638
rect 4245 13635 4311 13636
rect 5165 13635 5231 13636
rect 4153 13426 4219 13429
rect 4470 13426 4476 13428
rect 4153 13424 4476 13426
rect 4153 13368 4158 13424
rect 4214 13368 4476 13424
rect 4153 13366 4476 13368
rect 4153 13363 4219 13366
rect 4470 13364 4476 13366
rect 4540 13364 4546 13428
rect 5950 13290 6010 13907
rect 15326 13772 15332 13836
rect 15396 13834 15402 13836
rect 15653 13834 15719 13837
rect 15396 13832 15719 13834
rect 15396 13776 15658 13832
rect 15714 13776 15719 13832
rect 15396 13774 15719 13776
rect 15396 13772 15402 13774
rect 15653 13771 15719 13774
rect 8341 13632 8661 13633
rect 8341 13568 8349 13632
rect 8413 13568 8429 13632
rect 8493 13568 8509 13632
rect 8573 13568 8589 13632
rect 8653 13568 8661 13632
rect 8341 13567 8661 13568
rect 15738 13632 16058 13633
rect 15738 13568 15746 13632
rect 15810 13568 15826 13632
rect 15890 13568 15906 13632
rect 15970 13568 15986 13632
rect 16050 13568 16058 13632
rect 15738 13567 16058 13568
rect 18873 13562 18939 13565
rect 16208 13560 18939 13562
rect 16208 13504 18878 13560
rect 18934 13504 18939 13560
rect 16208 13502 18939 13504
rect 9581 13426 9647 13429
rect 13997 13426 14063 13429
rect 9581 13424 14063 13426
rect 9581 13368 9586 13424
rect 9642 13368 14002 13424
rect 14058 13368 14063 13424
rect 9581 13366 14063 13368
rect 9581 13363 9647 13366
rect 13997 13363 14063 13366
rect 14181 13426 14247 13429
rect 16208 13426 16268 13502
rect 18873 13499 18939 13502
rect 14181 13424 16268 13426
rect 14181 13368 14186 13424
rect 14242 13368 16268 13424
rect 14181 13366 16268 13368
rect 14181 13363 14247 13366
rect 17902 13364 17908 13428
rect 17972 13426 17978 13428
rect 23920 13426 24400 13456
rect 17972 13366 24400 13426
rect 17972 13364 17978 13366
rect 23920 13336 24400 13366
rect 6085 13290 6151 13293
rect 5950 13288 6151 13290
rect 5950 13232 6090 13288
rect 6146 13232 6151 13288
rect 5950 13230 6151 13232
rect 6085 13227 6151 13230
rect 11881 13290 11947 13293
rect 20345 13290 20411 13293
rect 11881 13288 20411 13290
rect 11881 13232 11886 13288
rect 11942 13232 20350 13288
rect 20406 13232 20411 13288
rect 11881 13230 20411 13232
rect 11881 13227 11947 13230
rect 20345 13227 20411 13230
rect 5349 13154 5415 13157
rect 5901 13154 5967 13157
rect 5349 13152 5967 13154
rect 5349 13096 5354 13152
rect 5410 13096 5906 13152
rect 5962 13096 5967 13152
rect 5349 13094 5967 13096
rect 5349 13091 5415 13094
rect 5901 13091 5967 13094
rect 4642 13088 4962 13089
rect 4642 13024 4650 13088
rect 4714 13024 4730 13088
rect 4794 13024 4810 13088
rect 4874 13024 4890 13088
rect 4954 13024 4962 13088
rect 4642 13023 4962 13024
rect 12040 13088 12360 13089
rect 12040 13024 12048 13088
rect 12112 13024 12128 13088
rect 12192 13024 12208 13088
rect 12272 13024 12288 13088
rect 12352 13024 12360 13088
rect 12040 13023 12360 13024
rect 19437 13088 19757 13089
rect 19437 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19605 13088
rect 19669 13024 19685 13088
rect 19749 13024 19757 13088
rect 19437 13023 19757 13024
rect 9121 13018 9187 13021
rect 17861 13018 17927 13021
rect 18689 13018 18755 13021
rect 9121 13016 9690 13018
rect 9121 12960 9126 13016
rect 9182 12960 9690 13016
rect 9121 12958 9690 12960
rect 9121 12955 9187 12958
rect 1669 12882 1735 12885
rect 8017 12882 8083 12885
rect 1669 12880 8083 12882
rect 1669 12824 1674 12880
rect 1730 12824 8022 12880
rect 8078 12824 8083 12880
rect 1669 12822 8083 12824
rect 1669 12819 1735 12822
rect 8017 12819 8083 12822
rect 5022 12684 5028 12748
rect 5092 12746 5098 12748
rect 5257 12746 5323 12749
rect 5092 12744 5323 12746
rect 5092 12688 5262 12744
rect 5318 12688 5323 12744
rect 5092 12686 5323 12688
rect 5092 12684 5098 12686
rect 5257 12683 5323 12686
rect 7230 12684 7236 12748
rect 7300 12746 7306 12748
rect 8753 12746 8819 12749
rect 7300 12744 8819 12746
rect 7300 12688 8758 12744
rect 8814 12688 8819 12744
rect 7300 12686 8819 12688
rect 7300 12684 7306 12686
rect 8753 12683 8819 12686
rect 9630 12610 9690 12958
rect 17861 13016 18755 13018
rect 17861 12960 17866 13016
rect 17922 12960 18694 13016
rect 18750 12960 18755 13016
rect 17861 12958 18755 12960
rect 17861 12955 17927 12958
rect 18689 12955 18755 12958
rect 10777 12882 10843 12885
rect 14457 12882 14523 12885
rect 20437 12882 20503 12885
rect 10777 12880 20503 12882
rect 10777 12824 10782 12880
rect 10838 12824 14462 12880
rect 14518 12824 20442 12880
rect 20498 12824 20503 12880
rect 10777 12822 20503 12824
rect 10777 12819 10843 12822
rect 14457 12819 14523 12822
rect 20437 12819 20503 12822
rect 11789 12746 11855 12749
rect 14733 12746 14799 12749
rect 11789 12744 14799 12746
rect 11789 12688 11794 12744
rect 11850 12688 14738 12744
rect 14794 12688 14799 12744
rect 11789 12686 14799 12688
rect 11789 12683 11855 12686
rect 14733 12683 14799 12686
rect 17534 12684 17540 12748
rect 17604 12746 17610 12748
rect 20069 12746 20135 12749
rect 17604 12744 20135 12746
rect 17604 12688 20074 12744
rect 20130 12688 20135 12744
rect 17604 12686 20135 12688
rect 17604 12684 17610 12686
rect 20069 12683 20135 12686
rect 21449 12746 21515 12749
rect 23920 12746 24400 12776
rect 21449 12744 24400 12746
rect 21449 12688 21454 12744
rect 21510 12688 24400 12744
rect 21449 12686 24400 12688
rect 21449 12683 21515 12686
rect 23920 12656 24400 12686
rect 11053 12610 11119 12613
rect 8848 12608 11119 12610
rect 8848 12552 11058 12608
rect 11114 12552 11119 12608
rect 8848 12550 11119 12552
rect 8341 12544 8661 12545
rect 8341 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8509 12544
rect 8573 12480 8589 12544
rect 8653 12480 8661 12544
rect 8341 12479 8661 12480
rect 8848 12341 8908 12550
rect 11053 12547 11119 12550
rect 13997 12610 14063 12613
rect 15561 12610 15627 12613
rect 13997 12608 15627 12610
rect 13997 12552 14002 12608
rect 14058 12552 15566 12608
rect 15622 12552 15627 12608
rect 13997 12550 15627 12552
rect 13997 12547 14063 12550
rect 15561 12547 15627 12550
rect 16757 12610 16823 12613
rect 19609 12610 19675 12613
rect 16757 12608 19675 12610
rect 16757 12552 16762 12608
rect 16818 12552 19614 12608
rect 19670 12552 19675 12608
rect 16757 12550 19675 12552
rect 16757 12547 16823 12550
rect 19609 12547 19675 12550
rect 20069 12610 20135 12613
rect 20253 12610 20319 12613
rect 20069 12608 20319 12610
rect 20069 12552 20074 12608
rect 20130 12552 20258 12608
rect 20314 12552 20319 12608
rect 20069 12550 20319 12552
rect 20069 12547 20135 12550
rect 20253 12547 20319 12550
rect 15738 12544 16058 12545
rect 15738 12480 15746 12544
rect 15810 12480 15826 12544
rect 15890 12480 15906 12544
rect 15970 12480 15986 12544
rect 16050 12480 16058 12544
rect 15738 12479 16058 12480
rect 9949 12474 10015 12477
rect 10174 12474 10180 12476
rect 9949 12472 10180 12474
rect 9949 12416 9954 12472
rect 10010 12416 10180 12472
rect 9949 12414 10180 12416
rect 9949 12411 10015 12414
rect 10174 12412 10180 12414
rect 10244 12412 10250 12476
rect 13169 12474 13235 12477
rect 13629 12474 13695 12477
rect 13169 12472 13695 12474
rect 13169 12416 13174 12472
rect 13230 12416 13634 12472
rect 13690 12416 13695 12472
rect 13169 12414 13695 12416
rect 13169 12411 13235 12414
rect 13629 12411 13695 12414
rect 13905 12472 13971 12477
rect 13905 12416 13910 12472
rect 13966 12416 13971 12472
rect 13905 12411 13971 12416
rect 18454 12412 18460 12476
rect 18524 12474 18530 12476
rect 18597 12474 18663 12477
rect 18524 12472 18663 12474
rect 18524 12416 18602 12472
rect 18658 12416 18663 12472
rect 18524 12414 18663 12416
rect 18524 12412 18530 12414
rect 18597 12411 18663 12414
rect 19190 12412 19196 12476
rect 19260 12474 19266 12476
rect 19885 12474 19951 12477
rect 19260 12472 19951 12474
rect 19260 12416 19890 12472
rect 19946 12416 19951 12472
rect 19260 12414 19951 12416
rect 19260 12412 19266 12414
rect 19885 12411 19951 12414
rect 6269 12340 6335 12341
rect 6269 12336 6316 12340
rect 6380 12338 6386 12340
rect 6269 12280 6274 12336
rect 6269 12276 6316 12280
rect 6380 12278 6426 12338
rect 8845 12336 8911 12341
rect 8845 12280 8850 12336
rect 8906 12280 8911 12336
rect 6380 12276 6386 12278
rect 6269 12275 6335 12276
rect 8845 12275 8911 12280
rect 9213 12340 9279 12341
rect 9213 12336 9260 12340
rect 9324 12338 9330 12340
rect 10593 12338 10659 12341
rect 11094 12338 11100 12340
rect 9213 12280 9218 12336
rect 9213 12276 9260 12280
rect 9324 12278 9370 12338
rect 10593 12336 11100 12338
rect 10593 12280 10598 12336
rect 10654 12280 11100 12336
rect 10593 12278 11100 12280
rect 9324 12276 9330 12278
rect 9213 12275 9279 12276
rect 10593 12275 10659 12278
rect 11094 12276 11100 12278
rect 11164 12276 11170 12340
rect 11237 12338 11303 12341
rect 13908 12338 13968 12411
rect 11237 12336 13968 12338
rect 11237 12280 11242 12336
rect 11298 12280 13968 12336
rect 11237 12278 13968 12280
rect 14273 12338 14339 12341
rect 14733 12338 14799 12341
rect 14273 12336 14799 12338
rect 14273 12280 14278 12336
rect 14334 12280 14738 12336
rect 14794 12280 14799 12336
rect 14273 12278 14799 12280
rect 11237 12275 11303 12278
rect 14273 12275 14339 12278
rect 14733 12275 14799 12278
rect 17902 12276 17908 12340
rect 17972 12338 17978 12340
rect 18045 12338 18111 12341
rect 17972 12336 18111 12338
rect 17972 12280 18050 12336
rect 18106 12280 18111 12336
rect 17972 12278 18111 12280
rect 17972 12276 17978 12278
rect 18045 12275 18111 12278
rect 2497 12202 2563 12205
rect 8845 12202 8911 12205
rect 9305 12204 9371 12205
rect 9254 12202 9260 12204
rect 2497 12200 8911 12202
rect 2497 12144 2502 12200
rect 2558 12144 8850 12200
rect 8906 12144 8911 12200
rect 2497 12142 8911 12144
rect 9214 12142 9260 12202
rect 9324 12200 9371 12204
rect 9366 12144 9371 12200
rect 2497 12139 2563 12142
rect 8845 12139 8911 12142
rect 9254 12140 9260 12142
rect 9324 12140 9371 12144
rect 9305 12139 9371 12140
rect 9857 12202 9923 12205
rect 11329 12202 11395 12205
rect 9857 12200 11395 12202
rect 9857 12144 9862 12200
rect 9918 12144 11334 12200
rect 11390 12144 11395 12200
rect 9857 12142 11395 12144
rect 9857 12139 9923 12142
rect 11329 12139 11395 12142
rect 13169 12202 13235 12205
rect 13813 12202 13879 12205
rect 13169 12200 13879 12202
rect 13169 12144 13174 12200
rect 13230 12144 13818 12200
rect 13874 12144 13879 12200
rect 13169 12142 13879 12144
rect 13169 12139 13235 12142
rect 13813 12139 13879 12142
rect 20529 12202 20595 12205
rect 20662 12202 20668 12204
rect 20529 12200 20668 12202
rect 20529 12144 20534 12200
rect 20590 12144 20668 12200
rect 20529 12142 20668 12144
rect 20529 12139 20595 12142
rect 20662 12140 20668 12142
rect 20732 12140 20738 12204
rect 23920 12202 24400 12232
rect 20854 12142 24400 12202
rect 12985 12068 13051 12069
rect 12934 12066 12940 12068
rect 12858 12006 12940 12066
rect 13004 12066 13051 12068
rect 14273 12066 14339 12069
rect 13004 12064 14339 12066
rect 13046 12008 14278 12064
rect 14334 12008 14339 12064
rect 12934 12004 12940 12006
rect 13004 12006 14339 12008
rect 13004 12004 13051 12006
rect 12985 12003 13051 12004
rect 14273 12003 14339 12006
rect 20161 12064 20227 12069
rect 20161 12008 20166 12064
rect 20222 12008 20227 12064
rect 20161 12003 20227 12008
rect 20437 12066 20503 12069
rect 20854 12066 20914 12142
rect 23920 12112 24400 12142
rect 20437 12064 20914 12066
rect 20437 12008 20442 12064
rect 20498 12008 20914 12064
rect 20437 12006 20914 12008
rect 20437 12003 20503 12006
rect 4642 12000 4962 12001
rect 4642 11936 4650 12000
rect 4714 11936 4730 12000
rect 4794 11936 4810 12000
rect 4874 11936 4890 12000
rect 4954 11936 4962 12000
rect 4642 11935 4962 11936
rect 12040 12000 12360 12001
rect 12040 11936 12048 12000
rect 12112 11936 12128 12000
rect 12192 11936 12208 12000
rect 12272 11936 12288 12000
rect 12352 11936 12360 12000
rect 12040 11935 12360 11936
rect 19437 12000 19757 12001
rect 19437 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19605 12000
rect 19669 11936 19685 12000
rect 19749 11936 19757 12000
rect 19437 11935 19757 11936
rect 7465 11930 7531 11933
rect 7833 11930 7899 11933
rect 7465 11928 7899 11930
rect 7465 11872 7470 11928
rect 7526 11872 7838 11928
rect 7894 11872 7899 11928
rect 7465 11870 7899 11872
rect 7465 11867 7531 11870
rect 7833 11867 7899 11870
rect 9949 11930 10015 11933
rect 11697 11930 11763 11933
rect 9949 11928 11763 11930
rect 9949 11872 9954 11928
rect 10010 11872 11702 11928
rect 11758 11872 11763 11928
rect 9949 11870 11763 11872
rect 9949 11867 10015 11870
rect 11697 11867 11763 11870
rect 13169 11930 13235 11933
rect 15653 11930 15719 11933
rect 13169 11928 15719 11930
rect 13169 11872 13174 11928
rect 13230 11872 15658 11928
rect 15714 11872 15719 11928
rect 13169 11870 15719 11872
rect 13169 11867 13235 11870
rect 15653 11867 15719 11870
rect 4797 11794 4863 11797
rect 8845 11794 8911 11797
rect 4797 11792 8911 11794
rect 4797 11736 4802 11792
rect 4858 11736 8850 11792
rect 8906 11736 8911 11792
rect 4797 11734 8911 11736
rect 4797 11731 4863 11734
rect 8845 11731 8911 11734
rect 10317 11794 10383 11797
rect 15009 11794 15075 11797
rect 10317 11792 15075 11794
rect 10317 11736 10322 11792
rect 10378 11736 15014 11792
rect 15070 11736 15075 11792
rect 10317 11734 15075 11736
rect 10317 11731 10383 11734
rect 15009 11731 15075 11734
rect 19006 11732 19012 11796
rect 19076 11794 19082 11796
rect 20164 11794 20224 12003
rect 19076 11734 20224 11794
rect 19076 11732 19082 11734
rect 2957 11658 3023 11661
rect 7557 11658 7623 11661
rect 2957 11656 7623 11658
rect 2957 11600 2962 11656
rect 3018 11600 7562 11656
rect 7618 11600 7623 11656
rect 2957 11598 7623 11600
rect 2957 11595 3023 11598
rect 7557 11595 7623 11598
rect 14549 11658 14615 11661
rect 15745 11658 15811 11661
rect 14549 11656 15811 11658
rect 14549 11600 14554 11656
rect 14610 11600 15750 11656
rect 15806 11600 15811 11656
rect 14549 11598 15811 11600
rect 14549 11595 14615 11598
rect 15745 11595 15811 11598
rect 16205 11658 16271 11661
rect 16389 11658 16455 11661
rect 16798 11658 16804 11660
rect 16205 11656 16314 11658
rect 16205 11600 16210 11656
rect 16266 11600 16314 11656
rect 16205 11595 16314 11600
rect 16389 11656 16804 11658
rect 16389 11600 16394 11656
rect 16450 11600 16804 11656
rect 16389 11598 16804 11600
rect 16389 11595 16455 11598
rect 16798 11596 16804 11598
rect 16868 11596 16874 11660
rect 19609 11658 19675 11661
rect 21541 11658 21607 11661
rect 19609 11656 21607 11658
rect 19609 11600 19614 11656
rect 19670 11600 21546 11656
rect 21602 11600 21607 11656
rect 19609 11598 21607 11600
rect 19609 11595 19675 11598
rect 21541 11595 21607 11598
rect 8845 11522 8911 11525
rect 13169 11522 13235 11525
rect 8845 11520 13235 11522
rect 8845 11464 8850 11520
rect 8906 11464 13174 11520
rect 13230 11464 13235 11520
rect 8845 11462 13235 11464
rect 8845 11459 8911 11462
rect 13169 11459 13235 11462
rect 8341 11456 8661 11457
rect 8341 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8509 11456
rect 8573 11392 8589 11456
rect 8653 11392 8661 11456
rect 8341 11391 8661 11392
rect 15738 11456 16058 11457
rect 15738 11392 15746 11456
rect 15810 11392 15826 11456
rect 15890 11392 15906 11456
rect 15970 11392 15986 11456
rect 16050 11392 16058 11456
rect 15738 11391 16058 11392
rect 15193 11252 15259 11253
rect 15142 11250 15148 11252
rect 15102 11190 15148 11250
rect 15212 11248 15259 11252
rect 15254 11192 15259 11248
rect 15142 11188 15148 11190
rect 15212 11188 15259 11192
rect 15193 11187 15259 11188
rect 16254 11117 16314 11595
rect 19333 11522 19399 11525
rect 23920 11522 24400 11552
rect 19333 11520 24400 11522
rect 19333 11464 19338 11520
rect 19394 11464 24400 11520
rect 19333 11462 24400 11464
rect 19333 11459 19399 11462
rect 23920 11432 24400 11462
rect 18229 11252 18295 11253
rect 18229 11248 18276 11252
rect 18340 11250 18346 11252
rect 18229 11192 18234 11248
rect 18229 11188 18276 11192
rect 18340 11190 18386 11250
rect 18340 11188 18346 11190
rect 18229 11187 18295 11188
rect 3325 11114 3391 11117
rect 3693 11114 3759 11117
rect 3325 11112 3759 11114
rect 3325 11056 3330 11112
rect 3386 11056 3698 11112
rect 3754 11056 3759 11112
rect 3325 11054 3759 11056
rect 3325 11051 3391 11054
rect 3693 11051 3759 11054
rect 4889 11114 4955 11117
rect 11329 11114 11395 11117
rect 12801 11114 12867 11117
rect 13169 11114 13235 11117
rect 4889 11112 5090 11114
rect 4889 11056 4894 11112
rect 4950 11056 5090 11112
rect 4889 11054 5090 11056
rect 4889 11051 4955 11054
rect 4642 10912 4962 10913
rect 4642 10848 4650 10912
rect 4714 10848 4730 10912
rect 4794 10848 4810 10912
rect 4874 10848 4890 10912
rect 4954 10848 4962 10912
rect 4642 10847 4962 10848
rect 4889 10706 4955 10709
rect 5030 10706 5090 11054
rect 11329 11112 12496 11114
rect 11329 11056 11334 11112
rect 11390 11056 12496 11112
rect 11329 11054 12496 11056
rect 11329 11051 11395 11054
rect 12436 10978 12496 11054
rect 12801 11112 13235 11114
rect 12801 11056 12806 11112
rect 12862 11056 13174 11112
rect 13230 11056 13235 11112
rect 12801 11054 13235 11056
rect 12801 11051 12867 11054
rect 13169 11051 13235 11054
rect 13537 11114 13603 11117
rect 14641 11114 14707 11117
rect 14774 11114 14780 11116
rect 13537 11112 14780 11114
rect 13537 11056 13542 11112
rect 13598 11056 14646 11112
rect 14702 11056 14780 11112
rect 13537 11054 14780 11056
rect 13537 11051 13603 11054
rect 14641 11051 14707 11054
rect 14774 11052 14780 11054
rect 14844 11052 14850 11116
rect 16254 11112 16363 11117
rect 16254 11056 16302 11112
rect 16358 11056 16363 11112
rect 16254 11054 16363 11056
rect 16297 11051 16363 11054
rect 17493 10978 17559 10981
rect 12436 10976 17559 10978
rect 12436 10920 17498 10976
rect 17554 10920 17559 10976
rect 12436 10918 17559 10920
rect 17493 10915 17559 10918
rect 12040 10912 12360 10913
rect 12040 10848 12048 10912
rect 12112 10848 12128 10912
rect 12192 10848 12208 10912
rect 12272 10848 12288 10912
rect 12352 10848 12360 10912
rect 12040 10847 12360 10848
rect 19437 10912 19757 10913
rect 19437 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19605 10912
rect 19669 10848 19685 10912
rect 19749 10848 19757 10912
rect 19437 10847 19757 10848
rect 15929 10842 15995 10845
rect 18229 10842 18295 10845
rect 15929 10840 18295 10842
rect 15929 10784 15934 10840
rect 15990 10784 18234 10840
rect 18290 10784 18295 10840
rect 15929 10782 18295 10784
rect 15929 10779 15995 10782
rect 18229 10779 18295 10782
rect 20897 10842 20963 10845
rect 23920 10842 24400 10872
rect 20897 10840 24400 10842
rect 20897 10784 20902 10840
rect 20958 10784 24400 10840
rect 20897 10782 24400 10784
rect 20897 10779 20963 10782
rect 23920 10752 24400 10782
rect 6361 10708 6427 10709
rect 4889 10704 5090 10706
rect 4889 10648 4894 10704
rect 4950 10648 5090 10704
rect 4889 10646 5090 10648
rect 4889 10643 4955 10646
rect 6310 10644 6316 10708
rect 6380 10706 6427 10708
rect 9673 10706 9739 10709
rect 19885 10706 19951 10709
rect 6380 10704 6472 10706
rect 6422 10648 6472 10704
rect 6380 10646 6472 10648
rect 9673 10704 19951 10706
rect 9673 10648 9678 10704
rect 9734 10648 19890 10704
rect 19946 10648 19951 10704
rect 9673 10646 19951 10648
rect 6380 10644 6427 10646
rect 6361 10643 6427 10644
rect 9673 10643 9739 10646
rect 19885 10643 19951 10646
rect 6821 10570 6887 10573
rect 21173 10570 21239 10573
rect 6821 10568 21239 10570
rect 6821 10512 6826 10568
rect 6882 10512 21178 10568
rect 21234 10512 21239 10568
rect 6821 10510 21239 10512
rect 6821 10507 6887 10510
rect 21173 10507 21239 10510
rect 12433 10434 12499 10437
rect 15009 10434 15075 10437
rect 12433 10432 15075 10434
rect 12433 10376 12438 10432
rect 12494 10376 15014 10432
rect 15070 10376 15075 10432
rect 12433 10374 15075 10376
rect 12433 10371 12499 10374
rect 15009 10371 15075 10374
rect 16481 10434 16547 10437
rect 16665 10434 16731 10437
rect 16481 10432 16731 10434
rect 16481 10376 16486 10432
rect 16542 10376 16670 10432
rect 16726 10376 16731 10432
rect 16481 10374 16731 10376
rect 16481 10371 16547 10374
rect 16665 10371 16731 10374
rect 17585 10434 17651 10437
rect 17718 10434 17724 10436
rect 17585 10432 17724 10434
rect 17585 10376 17590 10432
rect 17646 10376 17724 10432
rect 17585 10374 17724 10376
rect 17585 10371 17651 10374
rect 17718 10372 17724 10374
rect 17788 10372 17794 10436
rect 18045 10434 18111 10437
rect 18413 10434 18479 10437
rect 18045 10432 18479 10434
rect 18045 10376 18050 10432
rect 18106 10376 18418 10432
rect 18474 10376 18479 10432
rect 18045 10374 18479 10376
rect 18045 10371 18111 10374
rect 18413 10371 18479 10374
rect 8341 10368 8661 10369
rect 8341 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8509 10368
rect 8573 10304 8589 10368
rect 8653 10304 8661 10368
rect 8341 10303 8661 10304
rect 15738 10368 16058 10369
rect 15738 10304 15746 10368
rect 15810 10304 15826 10368
rect 15890 10304 15906 10368
rect 15970 10304 15986 10368
rect 16050 10304 16058 10368
rect 15738 10303 16058 10304
rect 12525 10298 12591 10301
rect 13353 10298 13419 10301
rect 13905 10298 13971 10301
rect 12525 10296 13971 10298
rect 12525 10240 12530 10296
rect 12586 10240 13358 10296
rect 13414 10240 13910 10296
rect 13966 10240 13971 10296
rect 12525 10238 13971 10240
rect 12525 10235 12591 10238
rect 13353 10235 13419 10238
rect 13905 10235 13971 10238
rect 17861 10298 17927 10301
rect 18413 10298 18479 10301
rect 17861 10296 18479 10298
rect 17861 10240 17866 10296
rect 17922 10240 18418 10296
rect 18474 10240 18479 10296
rect 17861 10238 18479 10240
rect 17861 10235 17927 10238
rect 18413 10235 18479 10238
rect 7414 10100 7420 10164
rect 7484 10162 7490 10164
rect 15561 10162 15627 10165
rect 7484 10160 15627 10162
rect 7484 10104 15566 10160
rect 15622 10104 15627 10160
rect 7484 10102 15627 10104
rect 7484 10100 7490 10102
rect 15561 10099 15627 10102
rect 17861 10162 17927 10165
rect 23920 10162 24400 10192
rect 17861 10160 24400 10162
rect 17861 10104 17866 10160
rect 17922 10104 24400 10160
rect 17861 10102 24400 10104
rect 17861 10099 17927 10102
rect 23920 10072 24400 10102
rect 2221 10026 2287 10029
rect 4429 10026 4495 10029
rect 2221 10024 4495 10026
rect 2221 9968 2226 10024
rect 2282 9968 4434 10024
rect 4490 9968 4495 10024
rect 2221 9966 4495 9968
rect 2221 9963 2287 9966
rect 4429 9963 4495 9966
rect 11329 10026 11395 10029
rect 19701 10026 19767 10029
rect 11329 10024 19767 10026
rect 11329 9968 11334 10024
rect 11390 9968 19706 10024
rect 19762 9968 19767 10024
rect 11329 9966 19767 9968
rect 11329 9963 11395 9966
rect 19701 9963 19767 9966
rect 4642 9824 4962 9825
rect 4642 9760 4650 9824
rect 4714 9760 4730 9824
rect 4794 9760 4810 9824
rect 4874 9760 4890 9824
rect 4954 9760 4962 9824
rect 4642 9759 4962 9760
rect 12040 9824 12360 9825
rect 12040 9760 12048 9824
rect 12112 9760 12128 9824
rect 12192 9760 12208 9824
rect 12272 9760 12288 9824
rect 12352 9760 12360 9824
rect 12040 9759 12360 9760
rect 19437 9824 19757 9825
rect 19437 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19605 9824
rect 19669 9760 19685 9824
rect 19749 9760 19757 9824
rect 19437 9759 19757 9760
rect 8385 9754 8451 9757
rect 9765 9754 9831 9757
rect 8385 9752 9831 9754
rect 8385 9696 8390 9752
rect 8446 9696 9770 9752
rect 9826 9696 9831 9752
rect 8385 9694 9831 9696
rect 8385 9691 8451 9694
rect 9765 9691 9831 9694
rect 14958 9692 14964 9756
rect 15028 9754 15034 9756
rect 15028 9694 19258 9754
rect 15028 9692 15034 9694
rect 9438 9556 9444 9620
rect 9508 9618 9514 9620
rect 9857 9618 9923 9621
rect 12617 9618 12683 9621
rect 9508 9616 9923 9618
rect 9508 9560 9862 9616
rect 9918 9560 9923 9616
rect 9508 9558 9923 9560
rect 9508 9556 9514 9558
rect 9857 9555 9923 9558
rect 10780 9616 12683 9618
rect 10780 9560 12622 9616
rect 12678 9560 12683 9616
rect 10780 9558 12683 9560
rect 9121 9482 9187 9485
rect 10780 9482 10840 9558
rect 12617 9555 12683 9558
rect 16941 9618 17007 9621
rect 18086 9618 18092 9620
rect 16941 9616 18092 9618
rect 16941 9560 16946 9616
rect 17002 9560 18092 9616
rect 16941 9558 18092 9560
rect 16941 9555 17007 9558
rect 18086 9556 18092 9558
rect 18156 9556 18162 9620
rect 18822 9556 18828 9620
rect 18892 9618 18898 9620
rect 18965 9618 19031 9621
rect 18892 9616 19031 9618
rect 18892 9560 18970 9616
rect 19026 9560 19031 9616
rect 18892 9558 19031 9560
rect 19198 9618 19258 9694
rect 19885 9618 19951 9621
rect 20437 9618 20503 9621
rect 19198 9616 20503 9618
rect 19198 9560 19890 9616
rect 19946 9560 20442 9616
rect 20498 9560 20503 9616
rect 19198 9558 20503 9560
rect 18892 9556 18898 9558
rect 18965 9555 19031 9558
rect 19885 9555 19951 9558
rect 20437 9555 20503 9558
rect 9121 9480 10840 9482
rect 9121 9424 9126 9480
rect 9182 9424 10840 9480
rect 9121 9422 10840 9424
rect 9121 9419 9187 9422
rect 10910 9420 10916 9484
rect 10980 9482 10986 9484
rect 11053 9482 11119 9485
rect 10980 9480 11119 9482
rect 10980 9424 11058 9480
rect 11114 9424 11119 9480
rect 10980 9422 11119 9424
rect 10980 9420 10986 9422
rect 11053 9419 11119 9422
rect 11830 9420 11836 9484
rect 11900 9482 11906 9484
rect 17861 9482 17927 9485
rect 11900 9480 17927 9482
rect 11900 9424 17866 9480
rect 17922 9424 17927 9480
rect 11900 9422 17927 9424
rect 11900 9420 11906 9422
rect 17861 9419 17927 9422
rect 18505 9482 18571 9485
rect 19425 9482 19491 9485
rect 23920 9482 24400 9512
rect 18505 9480 19491 9482
rect 18505 9424 18510 9480
rect 18566 9424 19430 9480
rect 19486 9424 19491 9480
rect 18505 9422 19491 9424
rect 18505 9419 18571 9422
rect 19425 9419 19491 9422
rect 23798 9422 24400 9482
rect 10225 9348 10291 9349
rect 10174 9346 10180 9348
rect 10134 9286 10180 9346
rect 10244 9344 10291 9348
rect 10286 9288 10291 9344
rect 10174 9284 10180 9286
rect 10244 9284 10291 9288
rect 10358 9284 10364 9348
rect 10428 9346 10434 9348
rect 11145 9346 11211 9349
rect 10428 9344 11211 9346
rect 10428 9288 11150 9344
rect 11206 9288 11211 9344
rect 10428 9286 11211 9288
rect 10428 9284 10434 9286
rect 10225 9283 10291 9284
rect 11145 9283 11211 9286
rect 13169 9346 13235 9349
rect 15561 9346 15627 9349
rect 13169 9344 15627 9346
rect 13169 9288 13174 9344
rect 13230 9288 15566 9344
rect 15622 9288 15627 9344
rect 13169 9286 15627 9288
rect 13169 9283 13235 9286
rect 15561 9283 15627 9286
rect 16941 9346 17007 9349
rect 18965 9346 19031 9349
rect 23798 9346 23858 9422
rect 23920 9392 24400 9422
rect 16941 9344 18890 9346
rect 16941 9288 16946 9344
rect 17002 9288 18890 9344
rect 16941 9286 18890 9288
rect 16941 9283 17007 9286
rect 8341 9280 8661 9281
rect 8341 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8509 9280
rect 8573 9216 8589 9280
rect 8653 9216 8661 9280
rect 8341 9215 8661 9216
rect 15738 9280 16058 9281
rect 15738 9216 15746 9280
rect 15810 9216 15826 9280
rect 15890 9216 15906 9280
rect 15970 9216 15986 9280
rect 16050 9216 16058 9280
rect 15738 9215 16058 9216
rect 11329 9210 11395 9213
rect 8756 9208 11395 9210
rect 8756 9152 11334 9208
rect 11390 9152 11395 9208
rect 8756 9150 11395 9152
rect 0 9074 480 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 480 9014
rect 1485 9011 1551 9014
rect 6821 9074 6887 9077
rect 8293 9074 8359 9077
rect 8756 9074 8816 9150
rect 11329 9147 11395 9150
rect 16205 9210 16271 9213
rect 16573 9210 16639 9213
rect 18229 9210 18295 9213
rect 18413 9210 18479 9213
rect 16205 9208 16639 9210
rect 16205 9152 16210 9208
rect 16266 9152 16578 9208
rect 16634 9152 16639 9208
rect 16205 9150 16639 9152
rect 16205 9147 16271 9150
rect 16573 9147 16639 9150
rect 16990 9208 18479 9210
rect 16990 9152 18234 9208
rect 18290 9152 18418 9208
rect 18474 9152 18479 9208
rect 16990 9150 18479 9152
rect 18830 9210 18890 9286
rect 18965 9344 23858 9346
rect 18965 9288 18970 9344
rect 19026 9288 23858 9344
rect 18965 9286 23858 9288
rect 18965 9283 19031 9286
rect 19149 9210 19215 9213
rect 18830 9208 19215 9210
rect 18830 9152 19154 9208
rect 19210 9152 19215 9208
rect 18830 9150 19215 9152
rect 9305 9076 9371 9077
rect 6821 9072 7850 9074
rect 6821 9016 6826 9072
rect 6882 9016 7850 9072
rect 6821 9014 7850 9016
rect 6821 9011 6887 9014
rect 7790 8940 7850 9014
rect 8293 9072 8816 9074
rect 8293 9016 8298 9072
rect 8354 9016 8816 9072
rect 8293 9014 8816 9016
rect 8293 9011 8359 9014
rect 9254 9012 9260 9076
rect 9324 9074 9371 9076
rect 10225 9074 10291 9077
rect 11237 9074 11303 9077
rect 14457 9074 14523 9077
rect 9324 9072 9416 9074
rect 9366 9016 9416 9072
rect 9324 9014 9416 9016
rect 10225 9072 14523 9074
rect 10225 9016 10230 9072
rect 10286 9016 11242 9072
rect 11298 9016 14462 9072
rect 14518 9016 14523 9072
rect 10225 9014 14523 9016
rect 9324 9012 9371 9014
rect 9305 9011 9371 9012
rect 10225 9011 10291 9014
rect 11237 9011 11303 9014
rect 14457 9011 14523 9014
rect 14917 9074 14983 9077
rect 16990 9074 17050 9150
rect 18229 9147 18295 9150
rect 18413 9147 18479 9150
rect 19149 9147 19215 9150
rect 14917 9072 17050 9074
rect 14917 9016 14922 9072
rect 14978 9016 17050 9072
rect 14917 9014 17050 9016
rect 17125 9074 17191 9077
rect 19333 9074 19399 9077
rect 17125 9072 19399 9074
rect 17125 9016 17130 9072
rect 17186 9016 19338 9072
rect 19394 9016 19399 9072
rect 17125 9014 19399 9016
rect 14917 9011 14983 9014
rect 17125 9011 17191 9014
rect 19333 9011 19399 9014
rect 20069 9074 20135 9077
rect 20662 9074 20668 9076
rect 20069 9072 20668 9074
rect 20069 9016 20074 9072
rect 20130 9016 20668 9072
rect 20069 9014 20668 9016
rect 20069 9011 20135 9014
rect 20662 9012 20668 9014
rect 20732 9012 20738 9076
rect 7782 8876 7788 8940
rect 7852 8938 7858 8940
rect 18137 8938 18203 8941
rect 18270 8938 18276 8940
rect 7852 8878 17234 8938
rect 7852 8876 7858 8878
rect 5349 8802 5415 8805
rect 8201 8802 8267 8805
rect 5349 8800 8267 8802
rect 5349 8744 5354 8800
rect 5410 8744 8206 8800
rect 8262 8744 8267 8800
rect 5349 8742 8267 8744
rect 5349 8739 5415 8742
rect 8201 8739 8267 8742
rect 8477 8802 8543 8805
rect 9806 8802 9812 8804
rect 8477 8800 9812 8802
rect 8477 8744 8482 8800
rect 8538 8744 9812 8800
rect 8477 8742 9812 8744
rect 8477 8739 8543 8742
rect 9806 8740 9812 8742
rect 9876 8740 9882 8804
rect 10041 8802 10107 8805
rect 11513 8802 11579 8805
rect 10041 8800 11579 8802
rect 10041 8744 10046 8800
rect 10102 8744 11518 8800
rect 11574 8744 11579 8800
rect 10041 8742 11579 8744
rect 10041 8739 10107 8742
rect 11513 8739 11579 8742
rect 4642 8736 4962 8737
rect 4642 8672 4650 8736
rect 4714 8672 4730 8736
rect 4794 8672 4810 8736
rect 4874 8672 4890 8736
rect 4954 8672 4962 8736
rect 4642 8671 4962 8672
rect 12040 8736 12360 8737
rect 12040 8672 12048 8736
rect 12112 8672 12128 8736
rect 12192 8672 12208 8736
rect 12272 8672 12288 8736
rect 12352 8672 12360 8736
rect 12040 8671 12360 8672
rect 7005 8668 7071 8669
rect 7005 8666 7052 8668
rect 6960 8664 7052 8666
rect 6960 8608 7010 8664
rect 6960 8606 7052 8608
rect 7005 8604 7052 8606
rect 7116 8604 7122 8668
rect 7414 8604 7420 8668
rect 7484 8666 7490 8668
rect 8017 8666 8083 8669
rect 7484 8664 8083 8666
rect 7484 8608 8022 8664
rect 8078 8608 8083 8664
rect 7484 8606 8083 8608
rect 7484 8604 7490 8606
rect 7005 8603 7071 8604
rect 8017 8603 8083 8606
rect 8201 8666 8267 8669
rect 10685 8666 10751 8669
rect 8201 8664 10751 8666
rect 8201 8608 8206 8664
rect 8262 8608 10690 8664
rect 10746 8608 10751 8664
rect 8201 8606 10751 8608
rect 8201 8603 8267 8606
rect 10685 8603 10751 8606
rect 5073 8532 5139 8533
rect 5022 8530 5028 8532
rect 4982 8470 5028 8530
rect 5092 8528 5139 8532
rect 5134 8472 5139 8528
rect 5022 8468 5028 8470
rect 5092 8468 5139 8472
rect 5073 8467 5139 8468
rect 6085 8530 6151 8533
rect 7966 8530 7972 8532
rect 6085 8528 7972 8530
rect 6085 8472 6090 8528
rect 6146 8472 7972 8528
rect 6085 8470 7972 8472
rect 6085 8467 6151 8470
rect 7966 8468 7972 8470
rect 8036 8468 8042 8532
rect 8385 8530 8451 8533
rect 13118 8530 13124 8532
rect 8385 8528 13124 8530
rect 8385 8472 8390 8528
rect 8446 8472 13124 8528
rect 8385 8470 13124 8472
rect 8385 8467 8451 8470
rect 13118 8468 13124 8470
rect 13188 8468 13194 8532
rect 13353 8530 13419 8533
rect 15561 8530 15627 8533
rect 13353 8528 15627 8530
rect 13353 8472 13358 8528
rect 13414 8472 15566 8528
rect 15622 8472 15627 8528
rect 13353 8470 15627 8472
rect 17174 8530 17234 8878
rect 18137 8936 18276 8938
rect 18137 8880 18142 8936
rect 18198 8880 18276 8936
rect 18137 8878 18276 8880
rect 18137 8875 18203 8878
rect 18270 8876 18276 8878
rect 18340 8876 18346 8940
rect 22001 8802 22067 8805
rect 23920 8802 24400 8832
rect 22001 8800 24400 8802
rect 22001 8744 22006 8800
rect 22062 8744 24400 8800
rect 22001 8742 24400 8744
rect 22001 8739 22067 8742
rect 19437 8736 19757 8737
rect 19437 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19605 8736
rect 19669 8672 19685 8736
rect 19749 8672 19757 8736
rect 23920 8712 24400 8742
rect 19437 8671 19757 8672
rect 22737 8530 22803 8533
rect 17174 8528 22803 8530
rect 17174 8472 22742 8528
rect 22798 8472 22803 8528
rect 17174 8470 22803 8472
rect 13353 8467 13419 8470
rect 15561 8467 15627 8470
rect 22737 8467 22803 8470
rect 9673 8394 9739 8397
rect 10174 8394 10180 8396
rect 8158 8334 8816 8394
rect 5901 8260 5967 8261
rect 5901 8256 5948 8260
rect 6012 8258 6018 8260
rect 6545 8258 6611 8261
rect 8158 8258 8218 8334
rect 5901 8200 5906 8256
rect 5901 8196 5948 8200
rect 6012 8198 6058 8258
rect 6545 8256 8218 8258
rect 6545 8200 6550 8256
rect 6606 8200 8218 8256
rect 6545 8198 8218 8200
rect 8756 8258 8816 8334
rect 9673 8392 10180 8394
rect 9673 8336 9678 8392
rect 9734 8336 10180 8392
rect 9673 8334 10180 8336
rect 9673 8331 9739 8334
rect 10174 8332 10180 8334
rect 10244 8332 10250 8396
rect 16297 8394 16363 8397
rect 18413 8394 18479 8397
rect 16297 8392 18479 8394
rect 16297 8336 16302 8392
rect 16358 8336 18418 8392
rect 18474 8336 18479 8392
rect 16297 8334 18479 8336
rect 16297 8331 16363 8334
rect 18413 8331 18479 8334
rect 13854 8258 13860 8260
rect 8756 8198 13860 8258
rect 6012 8196 6018 8198
rect 5901 8195 5967 8196
rect 6545 8195 6611 8198
rect 13854 8196 13860 8198
rect 13924 8196 13930 8260
rect 17493 8258 17559 8261
rect 20989 8258 21055 8261
rect 17493 8256 21055 8258
rect 17493 8200 17498 8256
rect 17554 8200 20994 8256
rect 21050 8200 21055 8256
rect 17493 8198 21055 8200
rect 17493 8195 17559 8198
rect 20989 8195 21055 8198
rect 21265 8258 21331 8261
rect 23920 8258 24400 8288
rect 21265 8256 24400 8258
rect 21265 8200 21270 8256
rect 21326 8200 24400 8256
rect 21265 8198 24400 8200
rect 21265 8195 21331 8198
rect 8341 8192 8661 8193
rect 8341 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8509 8192
rect 8573 8128 8589 8192
rect 8653 8128 8661 8192
rect 8341 8127 8661 8128
rect 15738 8192 16058 8193
rect 15738 8128 15746 8192
rect 15810 8128 15826 8192
rect 15890 8128 15906 8192
rect 15970 8128 15986 8192
rect 16050 8128 16058 8192
rect 23920 8168 24400 8198
rect 15738 8127 16058 8128
rect 8753 8122 8819 8125
rect 8886 8122 8892 8124
rect 8753 8120 8892 8122
rect 8753 8064 8758 8120
rect 8814 8064 8892 8120
rect 8753 8062 8892 8064
rect 8753 8059 8819 8062
rect 8886 8060 8892 8062
rect 8956 8060 8962 8124
rect 9029 8122 9095 8125
rect 10225 8122 10291 8125
rect 9029 8120 10291 8122
rect 9029 8064 9034 8120
rect 9090 8064 10230 8120
rect 10286 8064 10291 8120
rect 9029 8062 10291 8064
rect 9029 8059 9095 8062
rect 10225 8059 10291 8062
rect 10961 8122 11027 8125
rect 14825 8122 14891 8125
rect 10961 8120 14891 8122
rect 10961 8064 10966 8120
rect 11022 8064 14830 8120
rect 14886 8064 14891 8120
rect 10961 8062 14891 8064
rect 10961 8059 11027 8062
rect 14825 8059 14891 8062
rect 18086 8060 18092 8124
rect 18156 8122 18162 8124
rect 19149 8122 19215 8125
rect 18156 8120 19215 8122
rect 18156 8064 19154 8120
rect 19210 8064 19215 8120
rect 18156 8062 19215 8064
rect 18156 8060 18162 8062
rect 19149 8059 19215 8062
rect 20846 8060 20852 8124
rect 20916 8122 20922 8124
rect 21357 8122 21423 8125
rect 20916 8120 21423 8122
rect 20916 8064 21362 8120
rect 21418 8064 21423 8120
rect 20916 8062 21423 8064
rect 20916 8060 20922 8062
rect 21357 8059 21423 8062
rect 2497 7986 2563 7989
rect 8017 7986 8083 7989
rect 2497 7984 8083 7986
rect 2497 7928 2502 7984
rect 2558 7928 8022 7984
rect 8078 7928 8083 7984
rect 2497 7926 8083 7928
rect 2497 7923 2563 7926
rect 8017 7923 8083 7926
rect 8201 7986 8267 7989
rect 17309 7986 17375 7989
rect 8201 7984 17375 7986
rect 8201 7928 8206 7984
rect 8262 7928 17314 7984
rect 17370 7928 17375 7984
rect 8201 7926 17375 7928
rect 8201 7923 8267 7926
rect 17309 7923 17375 7926
rect 7557 7850 7623 7853
rect 14641 7850 14707 7853
rect 19885 7850 19951 7853
rect 7557 7848 12496 7850
rect 7557 7792 7562 7848
rect 7618 7792 12496 7848
rect 7557 7790 12496 7792
rect 7557 7787 7623 7790
rect 5533 7714 5599 7717
rect 7230 7714 7236 7716
rect 5533 7712 7236 7714
rect 5533 7656 5538 7712
rect 5594 7656 7236 7712
rect 5533 7654 7236 7656
rect 5533 7651 5599 7654
rect 7230 7652 7236 7654
rect 7300 7652 7306 7716
rect 8477 7714 8543 7717
rect 10910 7714 10916 7716
rect 8477 7712 10916 7714
rect 8477 7656 8482 7712
rect 8538 7656 10916 7712
rect 8477 7654 10916 7656
rect 8477 7651 8543 7654
rect 10910 7652 10916 7654
rect 10980 7652 10986 7716
rect 12436 7714 12496 7790
rect 14641 7848 19951 7850
rect 14641 7792 14646 7848
rect 14702 7792 19890 7848
rect 19946 7792 19951 7848
rect 14641 7790 19951 7792
rect 14641 7787 14707 7790
rect 19885 7787 19951 7790
rect 12436 7654 18660 7714
rect 4642 7648 4962 7649
rect 4642 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4890 7648
rect 4954 7584 4962 7648
rect 4642 7583 4962 7584
rect 12040 7648 12360 7649
rect 12040 7584 12048 7648
rect 12112 7584 12128 7648
rect 12192 7584 12208 7648
rect 12272 7584 12288 7648
rect 12352 7584 12360 7648
rect 12040 7583 12360 7584
rect 7557 7578 7623 7581
rect 7782 7578 7788 7580
rect 7557 7576 7788 7578
rect 7557 7520 7562 7576
rect 7618 7520 7788 7576
rect 7557 7518 7788 7520
rect 7557 7515 7623 7518
rect 7782 7516 7788 7518
rect 7852 7516 7858 7580
rect 8477 7578 8543 7581
rect 11605 7578 11671 7581
rect 8477 7576 11671 7578
rect 8477 7520 8482 7576
rect 8538 7520 11610 7576
rect 11666 7520 11671 7576
rect 8477 7518 11671 7520
rect 8477 7515 8543 7518
rect 11605 7515 11671 7518
rect 12709 7578 12775 7581
rect 13445 7578 13511 7581
rect 17534 7578 17540 7580
rect 12709 7576 17540 7578
rect 12709 7520 12714 7576
rect 12770 7520 13450 7576
rect 13506 7520 17540 7576
rect 12709 7518 17540 7520
rect 12709 7515 12775 7518
rect 13445 7515 13511 7518
rect 17534 7516 17540 7518
rect 17604 7516 17610 7580
rect 8017 7442 8083 7445
rect 8150 7442 8156 7444
rect 8017 7440 8156 7442
rect 8017 7384 8022 7440
rect 8078 7384 8156 7440
rect 8017 7382 8156 7384
rect 8017 7379 8083 7382
rect 8150 7380 8156 7382
rect 8220 7380 8226 7444
rect 8293 7442 8359 7445
rect 9070 7442 9076 7444
rect 8293 7440 9076 7442
rect 8293 7384 8298 7440
rect 8354 7384 9076 7440
rect 8293 7382 9076 7384
rect 8293 7379 8359 7382
rect 9070 7380 9076 7382
rect 9140 7380 9146 7444
rect 9581 7442 9647 7445
rect 18454 7442 18460 7444
rect 9581 7440 18460 7442
rect 9581 7384 9586 7440
rect 9642 7384 18460 7440
rect 9581 7382 18460 7384
rect 9581 7379 9647 7382
rect 18454 7380 18460 7382
rect 18524 7380 18530 7444
rect 18600 7442 18660 7654
rect 19437 7648 19757 7649
rect 19437 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19605 7648
rect 19669 7584 19685 7648
rect 19749 7584 19757 7648
rect 19437 7583 19757 7584
rect 20989 7578 21055 7581
rect 21449 7578 21515 7581
rect 23920 7578 24400 7608
rect 20989 7576 24400 7578
rect 20989 7520 20994 7576
rect 21050 7520 21454 7576
rect 21510 7520 24400 7576
rect 20989 7518 24400 7520
rect 20989 7515 21055 7518
rect 21449 7515 21515 7518
rect 23920 7488 24400 7518
rect 20294 7442 20300 7444
rect 18600 7382 20300 7442
rect 20294 7380 20300 7382
rect 20364 7380 20370 7444
rect 7005 7308 7071 7309
rect 7005 7304 7052 7308
rect 7116 7306 7122 7308
rect 7741 7306 7807 7309
rect 12893 7306 12959 7309
rect 13670 7306 13676 7308
rect 7005 7248 7010 7304
rect 7005 7244 7052 7248
rect 7116 7246 7162 7306
rect 7741 7304 12818 7306
rect 7741 7248 7746 7304
rect 7802 7248 12818 7304
rect 7741 7246 12818 7248
rect 7116 7244 7122 7246
rect 7005 7243 7071 7244
rect 7741 7243 7807 7246
rect 9806 7108 9812 7172
rect 9876 7170 9882 7172
rect 11513 7170 11579 7173
rect 9876 7168 11579 7170
rect 9876 7112 11518 7168
rect 11574 7112 11579 7168
rect 9876 7110 11579 7112
rect 12758 7170 12818 7246
rect 12893 7304 13676 7306
rect 12893 7248 12898 7304
rect 12954 7248 13676 7304
rect 12893 7246 13676 7248
rect 12893 7243 12959 7246
rect 13670 7244 13676 7246
rect 13740 7306 13746 7308
rect 14457 7306 14523 7309
rect 13740 7304 14523 7306
rect 13740 7248 14462 7304
rect 14518 7248 14523 7304
rect 13740 7246 14523 7248
rect 13740 7244 13746 7246
rect 14457 7243 14523 7246
rect 15193 7170 15259 7173
rect 12758 7168 15259 7170
rect 12758 7112 15198 7168
rect 15254 7112 15259 7168
rect 12758 7110 15259 7112
rect 9876 7108 9882 7110
rect 11513 7107 11579 7110
rect 15193 7107 15259 7110
rect 8341 7104 8661 7105
rect 8341 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8509 7104
rect 8573 7040 8589 7104
rect 8653 7040 8661 7104
rect 8341 7039 8661 7040
rect 15738 7104 16058 7105
rect 15738 7040 15746 7104
rect 15810 7040 15826 7104
rect 15890 7040 15906 7104
rect 15970 7040 15986 7104
rect 16050 7040 16058 7104
rect 15738 7039 16058 7040
rect 8886 6972 8892 7036
rect 8956 7034 8962 7036
rect 9213 7034 9279 7037
rect 8956 7032 9279 7034
rect 8956 6976 9218 7032
rect 9274 6976 9279 7032
rect 8956 6974 9279 6976
rect 8956 6972 8962 6974
rect 9213 6971 9279 6974
rect 9857 7034 9923 7037
rect 10961 7034 11027 7037
rect 9857 7032 11027 7034
rect 9857 6976 9862 7032
rect 9918 6976 10966 7032
rect 11022 6976 11027 7032
rect 9857 6974 11027 6976
rect 9857 6971 9923 6974
rect 10961 6971 11027 6974
rect 13353 7034 13419 7037
rect 14365 7034 14431 7037
rect 13353 7032 14431 7034
rect 13353 6976 13358 7032
rect 13414 6976 14370 7032
rect 14426 6976 14431 7032
rect 13353 6974 14431 6976
rect 13353 6971 13419 6974
rect 14365 6971 14431 6974
rect 8017 6898 8083 6901
rect 16757 6898 16823 6901
rect 8017 6896 16823 6898
rect 8017 6840 8022 6896
rect 8078 6840 16762 6896
rect 16818 6840 16823 6896
rect 8017 6838 16823 6840
rect 8017 6835 8083 6838
rect 16757 6835 16823 6838
rect 20805 6898 20871 6901
rect 21265 6898 21331 6901
rect 20805 6896 21331 6898
rect 20805 6840 20810 6896
rect 20866 6840 21270 6896
rect 21326 6840 21331 6896
rect 20805 6838 21331 6840
rect 20805 6835 20871 6838
rect 21265 6835 21331 6838
rect 22737 6898 22803 6901
rect 23920 6898 24400 6928
rect 22737 6896 24400 6898
rect 22737 6840 22742 6896
rect 22798 6840 24400 6896
rect 22737 6838 24400 6840
rect 22737 6835 22803 6838
rect 23920 6808 24400 6838
rect 9029 6762 9095 6765
rect 19241 6762 19307 6765
rect 9029 6760 19307 6762
rect 9029 6704 9034 6760
rect 9090 6704 19246 6760
rect 19302 6704 19307 6760
rect 9029 6702 19307 6704
rect 9029 6699 9095 6702
rect 19241 6699 19307 6702
rect 9673 6626 9739 6629
rect 11697 6626 11763 6629
rect 9673 6624 11763 6626
rect 9673 6568 9678 6624
rect 9734 6568 11702 6624
rect 11758 6568 11763 6624
rect 9673 6566 11763 6568
rect 9673 6563 9739 6566
rect 11697 6563 11763 6566
rect 13118 6564 13124 6628
rect 13188 6626 13194 6628
rect 19190 6626 19196 6628
rect 13188 6566 19196 6626
rect 13188 6564 13194 6566
rect 19190 6564 19196 6566
rect 19260 6564 19266 6628
rect 4642 6560 4962 6561
rect 4642 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4890 6560
rect 4954 6496 4962 6560
rect 4642 6495 4962 6496
rect 12040 6560 12360 6561
rect 12040 6496 12048 6560
rect 12112 6496 12128 6560
rect 12192 6496 12208 6560
rect 12272 6496 12288 6560
rect 12352 6496 12360 6560
rect 12040 6495 12360 6496
rect 19437 6560 19757 6561
rect 19437 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19605 6560
rect 19669 6496 19685 6560
rect 19749 6496 19757 6560
rect 19437 6495 19757 6496
rect 18873 6490 18939 6493
rect 12758 6488 18939 6490
rect 12758 6432 18878 6488
rect 18934 6432 18939 6488
rect 12758 6430 18939 6432
rect 8385 6354 8451 6357
rect 12758 6354 12818 6430
rect 18873 6427 18939 6430
rect 8385 6352 12818 6354
rect 8385 6296 8390 6352
rect 8446 6296 12818 6352
rect 8385 6294 12818 6296
rect 12893 6354 12959 6357
rect 16389 6354 16455 6357
rect 16941 6354 17007 6357
rect 12893 6352 17007 6354
rect 12893 6296 12898 6352
rect 12954 6296 16394 6352
rect 16450 6296 16946 6352
rect 17002 6296 17007 6352
rect 12893 6294 17007 6296
rect 8385 6291 8451 6294
rect 12893 6291 12959 6294
rect 16389 6291 16455 6294
rect 16941 6291 17007 6294
rect 18137 6354 18203 6357
rect 19977 6354 20043 6357
rect 22921 6354 22987 6357
rect 18137 6352 20043 6354
rect 18137 6296 18142 6352
rect 18198 6296 19982 6352
rect 20038 6296 20043 6352
rect 18137 6294 20043 6296
rect 18137 6291 18203 6294
rect 19977 6291 20043 6294
rect 21038 6352 22987 6354
rect 21038 6296 22926 6352
rect 22982 6296 22987 6352
rect 21038 6294 22987 6296
rect 9121 6218 9187 6221
rect 13118 6218 13124 6220
rect 9121 6216 13124 6218
rect 9121 6160 9126 6216
rect 9182 6160 13124 6216
rect 9121 6158 13124 6160
rect 9121 6155 9187 6158
rect 13118 6156 13124 6158
rect 13188 6156 13194 6220
rect 15285 6218 15351 6221
rect 21038 6218 21098 6294
rect 22921 6291 22987 6294
rect 15285 6216 21098 6218
rect 15285 6160 15290 6216
rect 15346 6160 21098 6216
rect 15285 6158 21098 6160
rect 22461 6218 22527 6221
rect 23920 6218 24400 6248
rect 22461 6216 24400 6218
rect 22461 6160 22466 6216
rect 22522 6160 24400 6216
rect 22461 6158 24400 6160
rect 15285 6155 15351 6158
rect 22461 6155 22527 6158
rect 23920 6128 24400 6158
rect 13077 6082 13143 6085
rect 15561 6082 15627 6085
rect 13077 6080 15627 6082
rect 13077 6024 13082 6080
rect 13138 6024 15566 6080
rect 15622 6024 15627 6080
rect 13077 6022 15627 6024
rect 13077 6019 13143 6022
rect 15561 6019 15627 6022
rect 16941 6082 17007 6085
rect 19977 6082 20043 6085
rect 16941 6080 20043 6082
rect 16941 6024 16946 6080
rect 17002 6024 19982 6080
rect 20038 6024 20043 6080
rect 16941 6022 20043 6024
rect 16941 6019 17007 6022
rect 19977 6019 20043 6022
rect 8341 6016 8661 6017
rect 8341 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8509 6016
rect 8573 5952 8589 6016
rect 8653 5952 8661 6016
rect 8341 5951 8661 5952
rect 15738 6016 16058 6017
rect 15738 5952 15746 6016
rect 15810 5952 15826 6016
rect 15890 5952 15906 6016
rect 15970 5952 15986 6016
rect 16050 5952 16058 6016
rect 15738 5951 16058 5952
rect 9305 5946 9371 5949
rect 9438 5946 9444 5948
rect 9305 5944 9444 5946
rect 9305 5888 9310 5944
rect 9366 5888 9444 5944
rect 9305 5886 9444 5888
rect 9305 5883 9371 5886
rect 9438 5884 9444 5886
rect 9508 5884 9514 5948
rect 15142 5946 15148 5948
rect 9998 5886 15148 5946
rect 7557 5810 7623 5813
rect 9998 5810 10058 5886
rect 15142 5884 15148 5886
rect 15212 5884 15218 5948
rect 19609 5946 19675 5949
rect 22737 5946 22803 5949
rect 19609 5944 22803 5946
rect 19609 5888 19614 5944
rect 19670 5888 22742 5944
rect 22798 5888 22803 5944
rect 19609 5886 22803 5888
rect 19609 5883 19675 5886
rect 22737 5883 22803 5886
rect 7557 5808 10058 5810
rect 7557 5752 7562 5808
rect 7618 5752 10058 5808
rect 7557 5750 10058 5752
rect 10225 5810 10291 5813
rect 11830 5810 11836 5812
rect 10225 5808 11836 5810
rect 10225 5752 10230 5808
rect 10286 5752 11836 5808
rect 10225 5750 11836 5752
rect 7557 5747 7623 5750
rect 10225 5747 10291 5750
rect 11830 5748 11836 5750
rect 11900 5748 11906 5812
rect 12157 5810 12223 5813
rect 21173 5810 21239 5813
rect 12157 5808 21239 5810
rect 12157 5752 12162 5808
rect 12218 5752 21178 5808
rect 21234 5752 21239 5808
rect 12157 5750 21239 5752
rect 12157 5747 12223 5750
rect 21173 5747 21239 5750
rect 13813 5674 13879 5677
rect 20253 5674 20319 5677
rect 13813 5672 20319 5674
rect 13813 5616 13818 5672
rect 13874 5616 20258 5672
rect 20314 5616 20319 5672
rect 13813 5614 20319 5616
rect 13813 5611 13879 5614
rect 20253 5611 20319 5614
rect 12893 5540 12959 5541
rect 13629 5540 13695 5541
rect 12893 5536 12940 5540
rect 13004 5538 13010 5540
rect 13629 5538 13676 5540
rect 12893 5480 12898 5536
rect 12893 5476 12940 5480
rect 13004 5478 13050 5538
rect 13584 5536 13676 5538
rect 13584 5480 13634 5536
rect 13584 5478 13676 5480
rect 13004 5476 13010 5478
rect 13629 5476 13676 5478
rect 13740 5476 13746 5540
rect 15653 5538 15719 5541
rect 17125 5538 17191 5541
rect 15653 5536 17191 5538
rect 15653 5480 15658 5536
rect 15714 5480 17130 5536
rect 17186 5480 17191 5536
rect 15653 5478 17191 5480
rect 12893 5475 12959 5476
rect 13629 5475 13695 5476
rect 15653 5475 15719 5478
rect 17125 5475 17191 5478
rect 19885 5538 19951 5541
rect 20713 5538 20779 5541
rect 19885 5536 20779 5538
rect 19885 5480 19890 5536
rect 19946 5480 20718 5536
rect 20774 5480 20779 5536
rect 19885 5478 20779 5480
rect 19885 5475 19951 5478
rect 20713 5475 20779 5478
rect 22829 5538 22895 5541
rect 23920 5538 24400 5568
rect 22829 5536 24400 5538
rect 22829 5480 22834 5536
rect 22890 5480 24400 5536
rect 22829 5478 24400 5480
rect 22829 5475 22895 5478
rect 4642 5472 4962 5473
rect 4642 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4890 5472
rect 4954 5408 4962 5472
rect 4642 5407 4962 5408
rect 12040 5472 12360 5473
rect 12040 5408 12048 5472
rect 12112 5408 12128 5472
rect 12192 5408 12208 5472
rect 12272 5408 12288 5472
rect 12352 5408 12360 5472
rect 12040 5407 12360 5408
rect 19437 5472 19757 5473
rect 19437 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19605 5472
rect 19669 5408 19685 5472
rect 19749 5408 19757 5472
rect 23920 5448 24400 5478
rect 19437 5407 19757 5408
rect 7465 5402 7531 5405
rect 7598 5402 7604 5404
rect 7465 5400 7604 5402
rect 7465 5344 7470 5400
rect 7526 5344 7604 5400
rect 7465 5342 7604 5344
rect 7465 5339 7531 5342
rect 7598 5340 7604 5342
rect 7668 5340 7674 5404
rect 12709 5402 12775 5405
rect 19057 5402 19123 5405
rect 12709 5400 19123 5402
rect 12709 5344 12714 5400
rect 12770 5344 19062 5400
rect 19118 5344 19123 5400
rect 12709 5342 19123 5344
rect 12709 5339 12775 5342
rect 19057 5339 19123 5342
rect 9397 5266 9463 5269
rect 12617 5266 12683 5269
rect 9397 5264 12683 5266
rect 9397 5208 9402 5264
rect 9458 5208 12622 5264
rect 12678 5208 12683 5264
rect 9397 5206 12683 5208
rect 9397 5203 9463 5206
rect 12617 5203 12683 5206
rect 16798 5204 16804 5268
rect 16868 5266 16874 5268
rect 16941 5266 17007 5269
rect 16868 5264 17007 5266
rect 16868 5208 16946 5264
rect 17002 5208 17007 5264
rect 16868 5206 17007 5208
rect 16868 5204 16874 5206
rect 16941 5203 17007 5206
rect 8341 4928 8661 4929
rect 8341 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8509 4928
rect 8573 4864 8589 4928
rect 8653 4864 8661 4928
rect 8341 4863 8661 4864
rect 15738 4928 16058 4929
rect 15738 4864 15746 4928
rect 15810 4864 15826 4928
rect 15890 4864 15906 4928
rect 15970 4864 15986 4928
rect 16050 4864 16058 4928
rect 15738 4863 16058 4864
rect 9857 4858 9923 4861
rect 10358 4858 10364 4860
rect 9857 4856 10364 4858
rect 9857 4800 9862 4856
rect 9918 4800 10364 4856
rect 9857 4798 10364 4800
rect 9857 4795 9923 4798
rect 10358 4796 10364 4798
rect 10428 4796 10434 4860
rect 20529 4858 20595 4861
rect 23920 4858 24400 4888
rect 20529 4856 24400 4858
rect 20529 4800 20534 4856
rect 20590 4800 24400 4856
rect 20529 4798 24400 4800
rect 20529 4795 20595 4798
rect 23920 4768 24400 4798
rect 15193 4722 15259 4725
rect 15469 4722 15535 4725
rect 19006 4722 19012 4724
rect 15193 4720 19012 4722
rect 15193 4664 15198 4720
rect 15254 4664 15474 4720
rect 15530 4664 19012 4720
rect 15193 4662 19012 4664
rect 15193 4659 15259 4662
rect 15469 4659 15535 4662
rect 19006 4660 19012 4662
rect 19076 4660 19082 4724
rect 14641 4586 14707 4589
rect 20662 4586 20668 4588
rect 14641 4584 20668 4586
rect 14641 4528 14646 4584
rect 14702 4528 20668 4584
rect 14641 4526 20668 4528
rect 14641 4523 14707 4526
rect 20662 4524 20668 4526
rect 20732 4524 20738 4588
rect 15009 4450 15075 4453
rect 15745 4450 15811 4453
rect 15009 4448 15811 4450
rect 15009 4392 15014 4448
rect 15070 4392 15750 4448
rect 15806 4392 15811 4448
rect 15009 4390 15811 4392
rect 15009 4387 15075 4390
rect 15745 4387 15811 4390
rect 16297 4450 16363 4453
rect 16614 4450 16620 4452
rect 16297 4448 16620 4450
rect 16297 4392 16302 4448
rect 16358 4392 16620 4448
rect 16297 4390 16620 4392
rect 16297 4387 16363 4390
rect 16614 4388 16620 4390
rect 16684 4388 16690 4452
rect 4642 4384 4962 4385
rect 4642 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4890 4384
rect 4954 4320 4962 4384
rect 4642 4319 4962 4320
rect 12040 4384 12360 4385
rect 12040 4320 12048 4384
rect 12112 4320 12128 4384
rect 12192 4320 12208 4384
rect 12272 4320 12288 4384
rect 12352 4320 12360 4384
rect 12040 4319 12360 4320
rect 19437 4384 19757 4385
rect 19437 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19605 4384
rect 19669 4320 19685 4384
rect 19749 4320 19757 4384
rect 19437 4319 19757 4320
rect 14457 4314 14523 4317
rect 17125 4314 17191 4317
rect 14457 4312 17191 4314
rect 14457 4256 14462 4312
rect 14518 4256 17130 4312
rect 17186 4256 17191 4312
rect 14457 4254 17191 4256
rect 14457 4251 14523 4254
rect 17125 4251 17191 4254
rect 20621 4314 20687 4317
rect 23920 4314 24400 4344
rect 20621 4312 24400 4314
rect 20621 4256 20626 4312
rect 20682 4256 24400 4312
rect 20621 4254 24400 4256
rect 20621 4251 20687 4254
rect 23920 4224 24400 4254
rect 13813 4178 13879 4181
rect 16573 4178 16639 4181
rect 13813 4176 16639 4178
rect 13813 4120 13818 4176
rect 13874 4120 16578 4176
rect 16634 4120 16639 4176
rect 13813 4118 16639 4120
rect 13813 4115 13879 4118
rect 16573 4115 16639 4118
rect 15561 4042 15627 4045
rect 18229 4042 18295 4045
rect 15561 4040 18295 4042
rect 15561 3984 15566 4040
rect 15622 3984 18234 4040
rect 18290 3984 18295 4040
rect 15561 3982 18295 3984
rect 15561 3979 15627 3982
rect 18229 3979 18295 3982
rect 16665 3906 16731 3909
rect 21817 3906 21883 3909
rect 16665 3904 21883 3906
rect 16665 3848 16670 3904
rect 16726 3848 21822 3904
rect 21878 3848 21883 3904
rect 16665 3846 21883 3848
rect 16665 3843 16731 3846
rect 21817 3843 21883 3846
rect 8341 3840 8661 3841
rect 8341 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8509 3840
rect 8573 3776 8589 3840
rect 8653 3776 8661 3840
rect 8341 3775 8661 3776
rect 15738 3840 16058 3841
rect 15738 3776 15746 3840
rect 15810 3776 15826 3840
rect 15890 3776 15906 3840
rect 15970 3776 15986 3840
rect 16050 3776 16058 3840
rect 15738 3775 16058 3776
rect 16941 3770 17007 3773
rect 20846 3770 20852 3772
rect 16941 3768 20852 3770
rect 16941 3712 16946 3768
rect 17002 3712 20852 3768
rect 16941 3710 20852 3712
rect 16941 3707 17007 3710
rect 20846 3708 20852 3710
rect 20916 3708 20922 3772
rect 12985 3634 13051 3637
rect 13997 3634 14063 3637
rect 15745 3634 15811 3637
rect 12985 3632 15811 3634
rect 12985 3576 12990 3632
rect 13046 3576 14002 3632
rect 14058 3576 15750 3632
rect 15806 3576 15811 3632
rect 12985 3574 15811 3576
rect 12985 3571 13051 3574
rect 13997 3571 14063 3574
rect 15745 3571 15811 3574
rect 15929 3634 15995 3637
rect 18822 3634 18828 3636
rect 15929 3632 18828 3634
rect 15929 3576 15934 3632
rect 15990 3576 18828 3632
rect 15929 3574 18828 3576
rect 15929 3571 15995 3574
rect 18822 3572 18828 3574
rect 18892 3572 18898 3636
rect 20161 3634 20227 3637
rect 23920 3634 24400 3664
rect 20161 3632 24400 3634
rect 20161 3576 20166 3632
rect 20222 3576 24400 3632
rect 20161 3574 24400 3576
rect 20161 3571 20227 3574
rect 23920 3544 24400 3574
rect 14549 3498 14615 3501
rect 16941 3498 17007 3501
rect 19926 3498 19932 3500
rect 14549 3496 17007 3498
rect 14549 3440 14554 3496
rect 14610 3440 16946 3496
rect 17002 3440 17007 3496
rect 14549 3438 17007 3440
rect 14549 3435 14615 3438
rect 16941 3435 17007 3438
rect 18094 3438 19932 3498
rect 13077 3362 13143 3365
rect 18094 3362 18154 3438
rect 19926 3436 19932 3438
rect 19996 3436 20002 3500
rect 13077 3360 18154 3362
rect 13077 3304 13082 3360
rect 13138 3304 18154 3360
rect 13077 3302 18154 3304
rect 13077 3299 13143 3302
rect 19926 3300 19932 3364
rect 19996 3362 20002 3364
rect 20478 3362 20484 3364
rect 19996 3302 20484 3362
rect 19996 3300 20002 3302
rect 20478 3300 20484 3302
rect 20548 3300 20554 3364
rect 4642 3296 4962 3297
rect 4642 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4890 3296
rect 4954 3232 4962 3296
rect 4642 3231 4962 3232
rect 12040 3296 12360 3297
rect 12040 3232 12048 3296
rect 12112 3232 12128 3296
rect 12192 3232 12208 3296
rect 12272 3232 12288 3296
rect 12352 3232 12360 3296
rect 12040 3231 12360 3232
rect 19437 3296 19757 3297
rect 19437 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19605 3296
rect 19669 3232 19685 3296
rect 19749 3232 19757 3296
rect 19437 3231 19757 3232
rect 14273 3226 14339 3229
rect 16982 3226 16988 3228
rect 14273 3224 16988 3226
rect 14273 3168 14278 3224
rect 14334 3168 16988 3224
rect 14273 3166 16988 3168
rect 14273 3163 14339 3166
rect 16982 3164 16988 3166
rect 17052 3164 17058 3228
rect 0 3090 480 3120
rect 1945 3090 2011 3093
rect 0 3088 2011 3090
rect 0 3032 1950 3088
rect 2006 3032 2011 3088
rect 0 3030 2011 3032
rect 0 3000 480 3030
rect 1945 3027 2011 3030
rect 14733 3090 14799 3093
rect 15510 3090 15516 3092
rect 14733 3088 15516 3090
rect 14733 3032 14738 3088
rect 14794 3032 15516 3088
rect 14733 3030 15516 3032
rect 14733 3027 14799 3030
rect 15510 3028 15516 3030
rect 15580 3028 15586 3092
rect 15745 3090 15811 3093
rect 21725 3090 21791 3093
rect 15745 3088 21791 3090
rect 15745 3032 15750 3088
rect 15806 3032 21730 3088
rect 21786 3032 21791 3088
rect 15745 3030 21791 3032
rect 15745 3027 15811 3030
rect 21725 3027 21791 3030
rect 14365 2954 14431 2957
rect 19926 2954 19932 2956
rect 14365 2952 19932 2954
rect 14365 2896 14370 2952
rect 14426 2896 19932 2952
rect 14365 2894 19932 2896
rect 14365 2891 14431 2894
rect 19926 2892 19932 2894
rect 19996 2892 20002 2956
rect 20345 2954 20411 2957
rect 23920 2954 24400 2984
rect 20345 2952 24400 2954
rect 20345 2896 20350 2952
rect 20406 2896 24400 2952
rect 20345 2894 24400 2896
rect 20345 2891 20411 2894
rect 23920 2864 24400 2894
rect 16205 2818 16271 2821
rect 20110 2818 20116 2820
rect 16205 2816 20116 2818
rect 16205 2760 16210 2816
rect 16266 2760 20116 2816
rect 16205 2758 20116 2760
rect 16205 2755 16271 2758
rect 20110 2756 20116 2758
rect 20180 2756 20186 2820
rect 8341 2752 8661 2753
rect 8341 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8509 2752
rect 8573 2688 8589 2752
rect 8653 2688 8661 2752
rect 8341 2687 8661 2688
rect 15738 2752 16058 2753
rect 15738 2688 15746 2752
rect 15810 2688 15826 2752
rect 15890 2688 15906 2752
rect 15970 2688 15986 2752
rect 16050 2688 16058 2752
rect 15738 2687 16058 2688
rect 13353 2682 13419 2685
rect 15326 2682 15332 2684
rect 13353 2680 15332 2682
rect 13353 2624 13358 2680
rect 13414 2624 15332 2680
rect 13353 2622 15332 2624
rect 13353 2619 13419 2622
rect 15326 2620 15332 2622
rect 15396 2620 15402 2684
rect 15653 2546 15719 2549
rect 18873 2546 18939 2549
rect 15653 2544 18939 2546
rect 15653 2488 15658 2544
rect 15714 2488 18878 2544
rect 18934 2488 18939 2544
rect 15653 2486 18939 2488
rect 15653 2483 15719 2486
rect 18873 2483 18939 2486
rect 8569 2410 8635 2413
rect 8886 2410 8892 2412
rect 8569 2408 8892 2410
rect 8569 2352 8574 2408
rect 8630 2352 8892 2408
rect 8569 2350 8892 2352
rect 8569 2347 8635 2350
rect 8886 2348 8892 2350
rect 8956 2348 8962 2412
rect 16614 2348 16620 2412
rect 16684 2410 16690 2412
rect 16684 2350 23122 2410
rect 16684 2348 16690 2350
rect 15009 2274 15075 2277
rect 16941 2274 17007 2277
rect 15009 2272 17007 2274
rect 15009 2216 15014 2272
rect 15070 2216 16946 2272
rect 17002 2216 17007 2272
rect 15009 2214 17007 2216
rect 23062 2274 23122 2350
rect 23920 2274 24400 2304
rect 23062 2214 24400 2274
rect 15009 2211 15075 2214
rect 16941 2211 17007 2214
rect 4642 2208 4962 2209
rect 4642 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4890 2208
rect 4954 2144 4962 2208
rect 4642 2143 4962 2144
rect 12040 2208 12360 2209
rect 12040 2144 12048 2208
rect 12112 2144 12128 2208
rect 12192 2144 12208 2208
rect 12272 2144 12288 2208
rect 12352 2144 12360 2208
rect 12040 2143 12360 2144
rect 19437 2208 19757 2209
rect 19437 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19605 2208
rect 19669 2144 19685 2208
rect 19749 2144 19757 2208
rect 23920 2184 24400 2214
rect 19437 2143 19757 2144
rect 22369 1594 22435 1597
rect 23920 1594 24400 1624
rect 22369 1592 24400 1594
rect 22369 1536 22374 1592
rect 22430 1536 24400 1592
rect 22369 1534 24400 1536
rect 22369 1531 22435 1534
rect 23920 1504 24400 1534
rect 19333 914 19399 917
rect 23920 914 24400 944
rect 19333 912 24400 914
rect 19333 856 19338 912
rect 19394 856 24400 912
rect 19333 854 24400 856
rect 19333 851 19399 854
rect 23920 824 24400 854
rect 23013 370 23079 373
rect 23920 370 24400 400
rect 23013 368 24400 370
rect 23013 312 23018 368
rect 23074 312 24400 368
rect 23013 310 24400 312
rect 23013 307 23079 310
rect 23920 280 24400 310
<< via3 >>
rect 4650 21788 4714 21792
rect 4650 21732 4654 21788
rect 4654 21732 4710 21788
rect 4710 21732 4714 21788
rect 4650 21728 4714 21732
rect 4730 21788 4794 21792
rect 4730 21732 4734 21788
rect 4734 21732 4790 21788
rect 4790 21732 4794 21788
rect 4730 21728 4794 21732
rect 4810 21788 4874 21792
rect 4810 21732 4814 21788
rect 4814 21732 4870 21788
rect 4870 21732 4874 21788
rect 4810 21728 4874 21732
rect 4890 21788 4954 21792
rect 4890 21732 4894 21788
rect 4894 21732 4950 21788
rect 4950 21732 4954 21788
rect 4890 21728 4954 21732
rect 12048 21788 12112 21792
rect 12048 21732 12052 21788
rect 12052 21732 12108 21788
rect 12108 21732 12112 21788
rect 12048 21728 12112 21732
rect 12128 21788 12192 21792
rect 12128 21732 12132 21788
rect 12132 21732 12188 21788
rect 12188 21732 12192 21788
rect 12128 21728 12192 21732
rect 12208 21788 12272 21792
rect 12208 21732 12212 21788
rect 12212 21732 12268 21788
rect 12268 21732 12272 21788
rect 12208 21728 12272 21732
rect 12288 21788 12352 21792
rect 12288 21732 12292 21788
rect 12292 21732 12348 21788
rect 12348 21732 12352 21788
rect 12288 21728 12352 21732
rect 19445 21788 19509 21792
rect 19445 21732 19449 21788
rect 19449 21732 19505 21788
rect 19505 21732 19509 21788
rect 19445 21728 19509 21732
rect 19525 21788 19589 21792
rect 19525 21732 19529 21788
rect 19529 21732 19585 21788
rect 19585 21732 19589 21788
rect 19525 21728 19589 21732
rect 19605 21788 19669 21792
rect 19605 21732 19609 21788
rect 19609 21732 19665 21788
rect 19665 21732 19669 21788
rect 19605 21728 19669 21732
rect 19685 21788 19749 21792
rect 19685 21732 19689 21788
rect 19689 21732 19745 21788
rect 19745 21732 19749 21788
rect 19685 21728 19749 21732
rect 8349 21244 8413 21248
rect 8349 21188 8353 21244
rect 8353 21188 8409 21244
rect 8409 21188 8413 21244
rect 8349 21184 8413 21188
rect 8429 21244 8493 21248
rect 8429 21188 8433 21244
rect 8433 21188 8489 21244
rect 8489 21188 8493 21244
rect 8429 21184 8493 21188
rect 8509 21244 8573 21248
rect 8509 21188 8513 21244
rect 8513 21188 8569 21244
rect 8569 21188 8573 21244
rect 8509 21184 8573 21188
rect 8589 21244 8653 21248
rect 8589 21188 8593 21244
rect 8593 21188 8649 21244
rect 8649 21188 8653 21244
rect 8589 21184 8653 21188
rect 15746 21244 15810 21248
rect 15746 21188 15750 21244
rect 15750 21188 15806 21244
rect 15806 21188 15810 21244
rect 15746 21184 15810 21188
rect 15826 21244 15890 21248
rect 15826 21188 15830 21244
rect 15830 21188 15886 21244
rect 15886 21188 15890 21244
rect 15826 21184 15890 21188
rect 15906 21244 15970 21248
rect 15906 21188 15910 21244
rect 15910 21188 15966 21244
rect 15966 21188 15970 21244
rect 15906 21184 15970 21188
rect 15986 21244 16050 21248
rect 15986 21188 15990 21244
rect 15990 21188 16046 21244
rect 16046 21188 16050 21244
rect 15986 21184 16050 21188
rect 7604 20980 7668 21044
rect 14964 20708 15028 20772
rect 16988 20768 17052 20772
rect 16988 20712 17002 20768
rect 17002 20712 17052 20768
rect 16988 20708 17052 20712
rect 20484 20768 20548 20772
rect 20484 20712 20534 20768
rect 20534 20712 20548 20768
rect 20484 20708 20548 20712
rect 4650 20700 4714 20704
rect 4650 20644 4654 20700
rect 4654 20644 4710 20700
rect 4710 20644 4714 20700
rect 4650 20640 4714 20644
rect 4730 20700 4794 20704
rect 4730 20644 4734 20700
rect 4734 20644 4790 20700
rect 4790 20644 4794 20700
rect 4730 20640 4794 20644
rect 4810 20700 4874 20704
rect 4810 20644 4814 20700
rect 4814 20644 4870 20700
rect 4870 20644 4874 20700
rect 4810 20640 4874 20644
rect 4890 20700 4954 20704
rect 4890 20644 4894 20700
rect 4894 20644 4950 20700
rect 4950 20644 4954 20700
rect 4890 20640 4954 20644
rect 12048 20700 12112 20704
rect 12048 20644 12052 20700
rect 12052 20644 12108 20700
rect 12108 20644 12112 20700
rect 12048 20640 12112 20644
rect 12128 20700 12192 20704
rect 12128 20644 12132 20700
rect 12132 20644 12188 20700
rect 12188 20644 12192 20700
rect 12128 20640 12192 20644
rect 12208 20700 12272 20704
rect 12208 20644 12212 20700
rect 12212 20644 12268 20700
rect 12268 20644 12272 20700
rect 12208 20640 12272 20644
rect 12288 20700 12352 20704
rect 12288 20644 12292 20700
rect 12292 20644 12348 20700
rect 12348 20644 12352 20700
rect 12288 20640 12352 20644
rect 19445 20700 19509 20704
rect 19445 20644 19449 20700
rect 19449 20644 19505 20700
rect 19505 20644 19509 20700
rect 19445 20640 19509 20644
rect 19525 20700 19589 20704
rect 19525 20644 19529 20700
rect 19529 20644 19585 20700
rect 19585 20644 19589 20700
rect 19525 20640 19589 20644
rect 19605 20700 19669 20704
rect 19605 20644 19609 20700
rect 19609 20644 19665 20700
rect 19665 20644 19669 20700
rect 19605 20640 19669 20644
rect 19685 20700 19749 20704
rect 19685 20644 19689 20700
rect 19689 20644 19745 20700
rect 19745 20644 19749 20700
rect 19685 20640 19749 20644
rect 7604 20300 7668 20364
rect 8349 20156 8413 20160
rect 8349 20100 8353 20156
rect 8353 20100 8409 20156
rect 8409 20100 8413 20156
rect 8349 20096 8413 20100
rect 8429 20156 8493 20160
rect 8429 20100 8433 20156
rect 8433 20100 8489 20156
rect 8489 20100 8493 20156
rect 8429 20096 8493 20100
rect 8509 20156 8573 20160
rect 8509 20100 8513 20156
rect 8513 20100 8569 20156
rect 8569 20100 8573 20156
rect 8509 20096 8573 20100
rect 8589 20156 8653 20160
rect 8589 20100 8593 20156
rect 8593 20100 8649 20156
rect 8649 20100 8653 20156
rect 8589 20096 8653 20100
rect 15746 20156 15810 20160
rect 15746 20100 15750 20156
rect 15750 20100 15806 20156
rect 15806 20100 15810 20156
rect 15746 20096 15810 20100
rect 15826 20156 15890 20160
rect 15826 20100 15830 20156
rect 15830 20100 15886 20156
rect 15886 20100 15890 20156
rect 15826 20096 15890 20100
rect 15906 20156 15970 20160
rect 15906 20100 15910 20156
rect 15910 20100 15966 20156
rect 15966 20100 15970 20156
rect 15906 20096 15970 20100
rect 15986 20156 16050 20160
rect 15986 20100 15990 20156
rect 15990 20100 16046 20156
rect 16046 20100 16050 20156
rect 15986 20096 16050 20100
rect 5948 19892 6012 19956
rect 20116 19756 20180 19820
rect 4650 19612 4714 19616
rect 4650 19556 4654 19612
rect 4654 19556 4710 19612
rect 4710 19556 4714 19612
rect 4650 19552 4714 19556
rect 4730 19612 4794 19616
rect 4730 19556 4734 19612
rect 4734 19556 4790 19612
rect 4790 19556 4794 19612
rect 4730 19552 4794 19556
rect 4810 19612 4874 19616
rect 4810 19556 4814 19612
rect 4814 19556 4870 19612
rect 4870 19556 4874 19612
rect 4810 19552 4874 19556
rect 4890 19612 4954 19616
rect 4890 19556 4894 19612
rect 4894 19556 4950 19612
rect 4950 19556 4954 19612
rect 4890 19552 4954 19556
rect 12048 19612 12112 19616
rect 12048 19556 12052 19612
rect 12052 19556 12108 19612
rect 12108 19556 12112 19612
rect 12048 19552 12112 19556
rect 12128 19612 12192 19616
rect 12128 19556 12132 19612
rect 12132 19556 12188 19612
rect 12188 19556 12192 19612
rect 12128 19552 12192 19556
rect 12208 19612 12272 19616
rect 12208 19556 12212 19612
rect 12212 19556 12268 19612
rect 12268 19556 12272 19612
rect 12208 19552 12272 19556
rect 12288 19612 12352 19616
rect 12288 19556 12292 19612
rect 12292 19556 12348 19612
rect 12348 19556 12352 19612
rect 12288 19552 12352 19556
rect 19445 19612 19509 19616
rect 19445 19556 19449 19612
rect 19449 19556 19505 19612
rect 19505 19556 19509 19612
rect 19445 19552 19509 19556
rect 19525 19612 19589 19616
rect 19525 19556 19529 19612
rect 19529 19556 19585 19612
rect 19585 19556 19589 19612
rect 19525 19552 19589 19556
rect 19605 19612 19669 19616
rect 19605 19556 19609 19612
rect 19609 19556 19665 19612
rect 19665 19556 19669 19612
rect 19605 19552 19669 19556
rect 19685 19612 19749 19616
rect 19685 19556 19689 19612
rect 19689 19556 19745 19612
rect 19745 19556 19749 19612
rect 19685 19552 19749 19556
rect 19932 19408 19996 19412
rect 19932 19352 19946 19408
rect 19946 19352 19996 19408
rect 19932 19348 19996 19352
rect 8892 19212 8956 19276
rect 8349 19068 8413 19072
rect 8349 19012 8353 19068
rect 8353 19012 8409 19068
rect 8409 19012 8413 19068
rect 8349 19008 8413 19012
rect 8429 19068 8493 19072
rect 8429 19012 8433 19068
rect 8433 19012 8489 19068
rect 8489 19012 8493 19068
rect 8429 19008 8493 19012
rect 8509 19068 8573 19072
rect 8509 19012 8513 19068
rect 8513 19012 8569 19068
rect 8569 19012 8573 19068
rect 8509 19008 8573 19012
rect 8589 19068 8653 19072
rect 8589 19012 8593 19068
rect 8593 19012 8649 19068
rect 8649 19012 8653 19068
rect 8589 19008 8653 19012
rect 15746 19068 15810 19072
rect 15746 19012 15750 19068
rect 15750 19012 15806 19068
rect 15806 19012 15810 19068
rect 15746 19008 15810 19012
rect 15826 19068 15890 19072
rect 15826 19012 15830 19068
rect 15830 19012 15886 19068
rect 15886 19012 15890 19068
rect 15826 19008 15890 19012
rect 15906 19068 15970 19072
rect 15906 19012 15910 19068
rect 15910 19012 15966 19068
rect 15966 19012 15970 19068
rect 15906 19008 15970 19012
rect 15986 19068 16050 19072
rect 15986 19012 15990 19068
rect 15990 19012 16046 19068
rect 16046 19012 16050 19068
rect 15986 19008 16050 19012
rect 4476 18864 4540 18868
rect 4476 18808 4490 18864
rect 4490 18808 4540 18864
rect 4476 18804 4540 18808
rect 5212 18532 5276 18596
rect 4650 18524 4714 18528
rect 4650 18468 4654 18524
rect 4654 18468 4710 18524
rect 4710 18468 4714 18524
rect 4650 18464 4714 18468
rect 4730 18524 4794 18528
rect 4730 18468 4734 18524
rect 4734 18468 4790 18524
rect 4790 18468 4794 18524
rect 4730 18464 4794 18468
rect 4810 18524 4874 18528
rect 4810 18468 4814 18524
rect 4814 18468 4870 18524
rect 4870 18468 4874 18524
rect 4810 18464 4874 18468
rect 4890 18524 4954 18528
rect 4890 18468 4894 18524
rect 4894 18468 4950 18524
rect 4950 18468 4954 18524
rect 4890 18464 4954 18468
rect 12048 18524 12112 18528
rect 12048 18468 12052 18524
rect 12052 18468 12108 18524
rect 12108 18468 12112 18524
rect 12048 18464 12112 18468
rect 12128 18524 12192 18528
rect 12128 18468 12132 18524
rect 12132 18468 12188 18524
rect 12188 18468 12192 18524
rect 12128 18464 12192 18468
rect 12208 18524 12272 18528
rect 12208 18468 12212 18524
rect 12212 18468 12268 18524
rect 12268 18468 12272 18524
rect 12208 18464 12272 18468
rect 12288 18524 12352 18528
rect 12288 18468 12292 18524
rect 12292 18468 12348 18524
rect 12348 18468 12352 18524
rect 12288 18464 12352 18468
rect 19445 18524 19509 18528
rect 19445 18468 19449 18524
rect 19449 18468 19505 18524
rect 19505 18468 19509 18524
rect 19445 18464 19509 18468
rect 19525 18524 19589 18528
rect 19525 18468 19529 18524
rect 19529 18468 19585 18524
rect 19585 18468 19589 18524
rect 19525 18464 19589 18468
rect 19605 18524 19669 18528
rect 19605 18468 19609 18524
rect 19609 18468 19665 18524
rect 19665 18468 19669 18524
rect 19605 18464 19669 18468
rect 19685 18524 19749 18528
rect 19685 18468 19689 18524
rect 19689 18468 19745 18524
rect 19745 18468 19749 18524
rect 19685 18464 19749 18468
rect 17724 18320 17788 18324
rect 17724 18264 17738 18320
rect 17738 18264 17788 18320
rect 17724 18260 17788 18264
rect 20668 18260 20732 18324
rect 9628 18124 9692 18188
rect 4292 17988 4356 18052
rect 9812 17988 9876 18052
rect 20300 17988 20364 18052
rect 8349 17980 8413 17984
rect 8349 17924 8353 17980
rect 8353 17924 8409 17980
rect 8409 17924 8413 17980
rect 8349 17920 8413 17924
rect 8429 17980 8493 17984
rect 8429 17924 8433 17980
rect 8433 17924 8489 17980
rect 8489 17924 8493 17980
rect 8429 17920 8493 17924
rect 8509 17980 8573 17984
rect 8509 17924 8513 17980
rect 8513 17924 8569 17980
rect 8569 17924 8573 17980
rect 8509 17920 8573 17924
rect 8589 17980 8653 17984
rect 8589 17924 8593 17980
rect 8593 17924 8649 17980
rect 8649 17924 8653 17980
rect 8589 17920 8653 17924
rect 15746 17980 15810 17984
rect 15746 17924 15750 17980
rect 15750 17924 15806 17980
rect 15806 17924 15810 17980
rect 15746 17920 15810 17924
rect 15826 17980 15890 17984
rect 15826 17924 15830 17980
rect 15830 17924 15886 17980
rect 15886 17924 15890 17980
rect 15826 17920 15890 17924
rect 15906 17980 15970 17984
rect 15906 17924 15910 17980
rect 15910 17924 15966 17980
rect 15966 17924 15970 17980
rect 15906 17920 15970 17924
rect 15986 17980 16050 17984
rect 15986 17924 15990 17980
rect 15990 17924 16046 17980
rect 16046 17924 16050 17980
rect 15986 17920 16050 17924
rect 4650 17436 4714 17440
rect 4650 17380 4654 17436
rect 4654 17380 4710 17436
rect 4710 17380 4714 17436
rect 4650 17376 4714 17380
rect 4730 17436 4794 17440
rect 4730 17380 4734 17436
rect 4734 17380 4790 17436
rect 4790 17380 4794 17436
rect 4730 17376 4794 17380
rect 4810 17436 4874 17440
rect 4810 17380 4814 17436
rect 4814 17380 4870 17436
rect 4870 17380 4874 17436
rect 4810 17376 4874 17380
rect 4890 17436 4954 17440
rect 4890 17380 4894 17436
rect 4894 17380 4950 17436
rect 4950 17380 4954 17436
rect 4890 17376 4954 17380
rect 12048 17436 12112 17440
rect 12048 17380 12052 17436
rect 12052 17380 12108 17436
rect 12108 17380 12112 17436
rect 12048 17376 12112 17380
rect 12128 17436 12192 17440
rect 12128 17380 12132 17436
rect 12132 17380 12188 17436
rect 12188 17380 12192 17436
rect 12128 17376 12192 17380
rect 12208 17436 12272 17440
rect 12208 17380 12212 17436
rect 12212 17380 12268 17436
rect 12268 17380 12272 17436
rect 12208 17376 12272 17380
rect 12288 17436 12352 17440
rect 12288 17380 12292 17436
rect 12292 17380 12348 17436
rect 12348 17380 12352 17436
rect 12288 17376 12352 17380
rect 19445 17436 19509 17440
rect 19445 17380 19449 17436
rect 19449 17380 19505 17436
rect 19505 17380 19509 17436
rect 19445 17376 19509 17380
rect 19525 17436 19589 17440
rect 19525 17380 19529 17436
rect 19529 17380 19585 17436
rect 19585 17380 19589 17436
rect 19525 17376 19589 17380
rect 19605 17436 19669 17440
rect 19605 17380 19609 17436
rect 19609 17380 19665 17436
rect 19665 17380 19669 17436
rect 19605 17376 19669 17380
rect 19685 17436 19749 17440
rect 19685 17380 19689 17436
rect 19689 17380 19745 17436
rect 19745 17380 19749 17436
rect 19685 17376 19749 17380
rect 4476 17036 4540 17100
rect 8349 16892 8413 16896
rect 8349 16836 8353 16892
rect 8353 16836 8409 16892
rect 8409 16836 8413 16892
rect 8349 16832 8413 16836
rect 8429 16892 8493 16896
rect 8429 16836 8433 16892
rect 8433 16836 8489 16892
rect 8489 16836 8493 16892
rect 8429 16832 8493 16836
rect 8509 16892 8573 16896
rect 8509 16836 8513 16892
rect 8513 16836 8569 16892
rect 8569 16836 8573 16892
rect 8509 16832 8573 16836
rect 8589 16892 8653 16896
rect 8589 16836 8593 16892
rect 8593 16836 8649 16892
rect 8649 16836 8653 16892
rect 8589 16832 8653 16836
rect 15746 16892 15810 16896
rect 15746 16836 15750 16892
rect 15750 16836 15806 16892
rect 15806 16836 15810 16892
rect 15746 16832 15810 16836
rect 15826 16892 15890 16896
rect 15826 16836 15830 16892
rect 15830 16836 15886 16892
rect 15886 16836 15890 16892
rect 15826 16832 15890 16836
rect 15906 16892 15970 16896
rect 15906 16836 15910 16892
rect 15910 16836 15966 16892
rect 15966 16836 15970 16892
rect 15906 16832 15970 16836
rect 15986 16892 16050 16896
rect 15986 16836 15990 16892
rect 15990 16836 16046 16892
rect 16046 16836 16050 16892
rect 15986 16832 16050 16836
rect 9260 16492 9324 16556
rect 9628 16492 9692 16556
rect 4650 16348 4714 16352
rect 4650 16292 4654 16348
rect 4654 16292 4710 16348
rect 4710 16292 4714 16348
rect 4650 16288 4714 16292
rect 4730 16348 4794 16352
rect 4730 16292 4734 16348
rect 4734 16292 4790 16348
rect 4790 16292 4794 16348
rect 4730 16288 4794 16292
rect 4810 16348 4874 16352
rect 4810 16292 4814 16348
rect 4814 16292 4870 16348
rect 4870 16292 4874 16348
rect 4810 16288 4874 16292
rect 4890 16348 4954 16352
rect 4890 16292 4894 16348
rect 4894 16292 4950 16348
rect 4950 16292 4954 16348
rect 4890 16288 4954 16292
rect 12048 16348 12112 16352
rect 12048 16292 12052 16348
rect 12052 16292 12108 16348
rect 12108 16292 12112 16348
rect 12048 16288 12112 16292
rect 12128 16348 12192 16352
rect 12128 16292 12132 16348
rect 12132 16292 12188 16348
rect 12188 16292 12192 16348
rect 12128 16288 12192 16292
rect 12208 16348 12272 16352
rect 12208 16292 12212 16348
rect 12212 16292 12268 16348
rect 12268 16292 12272 16348
rect 12208 16288 12272 16292
rect 12288 16348 12352 16352
rect 12288 16292 12292 16348
rect 12292 16292 12348 16348
rect 12348 16292 12352 16348
rect 12288 16288 12352 16292
rect 19445 16348 19509 16352
rect 19445 16292 19449 16348
rect 19449 16292 19505 16348
rect 19505 16292 19509 16348
rect 19445 16288 19509 16292
rect 19525 16348 19589 16352
rect 19525 16292 19529 16348
rect 19529 16292 19585 16348
rect 19585 16292 19589 16348
rect 19525 16288 19589 16292
rect 19605 16348 19669 16352
rect 19605 16292 19609 16348
rect 19609 16292 19665 16348
rect 19665 16292 19669 16348
rect 19605 16288 19669 16292
rect 19685 16348 19749 16352
rect 19685 16292 19689 16348
rect 19689 16292 19745 16348
rect 19745 16292 19749 16348
rect 19685 16288 19749 16292
rect 9812 16280 9876 16284
rect 9812 16224 9826 16280
rect 9826 16224 9876 16280
rect 9812 16220 9876 16224
rect 11100 16084 11164 16148
rect 8349 15804 8413 15808
rect 8349 15748 8353 15804
rect 8353 15748 8409 15804
rect 8409 15748 8413 15804
rect 8349 15744 8413 15748
rect 8429 15804 8493 15808
rect 8429 15748 8433 15804
rect 8433 15748 8489 15804
rect 8489 15748 8493 15804
rect 8429 15744 8493 15748
rect 8509 15804 8573 15808
rect 8509 15748 8513 15804
rect 8513 15748 8569 15804
rect 8569 15748 8573 15804
rect 8509 15744 8573 15748
rect 8589 15804 8653 15808
rect 8589 15748 8593 15804
rect 8593 15748 8649 15804
rect 8649 15748 8653 15804
rect 8589 15744 8653 15748
rect 15746 15804 15810 15808
rect 15746 15748 15750 15804
rect 15750 15748 15806 15804
rect 15806 15748 15810 15804
rect 15746 15744 15810 15748
rect 15826 15804 15890 15808
rect 15826 15748 15830 15804
rect 15830 15748 15886 15804
rect 15886 15748 15890 15804
rect 15826 15744 15890 15748
rect 15906 15804 15970 15808
rect 15906 15748 15910 15804
rect 15910 15748 15966 15804
rect 15966 15748 15970 15804
rect 15906 15744 15970 15748
rect 15986 15804 16050 15808
rect 15986 15748 15990 15804
rect 15990 15748 16046 15804
rect 16046 15748 16050 15804
rect 15986 15744 16050 15748
rect 7972 15540 8036 15604
rect 15516 15404 15580 15468
rect 9076 15268 9140 15332
rect 13860 15328 13924 15332
rect 13860 15272 13874 15328
rect 13874 15272 13924 15328
rect 13860 15268 13924 15272
rect 4650 15260 4714 15264
rect 4650 15204 4654 15260
rect 4654 15204 4710 15260
rect 4710 15204 4714 15260
rect 4650 15200 4714 15204
rect 4730 15260 4794 15264
rect 4730 15204 4734 15260
rect 4734 15204 4790 15260
rect 4790 15204 4794 15260
rect 4730 15200 4794 15204
rect 4810 15260 4874 15264
rect 4810 15204 4814 15260
rect 4814 15204 4870 15260
rect 4870 15204 4874 15260
rect 4810 15200 4874 15204
rect 4890 15260 4954 15264
rect 4890 15204 4894 15260
rect 4894 15204 4950 15260
rect 4950 15204 4954 15260
rect 4890 15200 4954 15204
rect 12048 15260 12112 15264
rect 12048 15204 12052 15260
rect 12052 15204 12108 15260
rect 12108 15204 12112 15260
rect 12048 15200 12112 15204
rect 12128 15260 12192 15264
rect 12128 15204 12132 15260
rect 12132 15204 12188 15260
rect 12188 15204 12192 15260
rect 12128 15200 12192 15204
rect 12208 15260 12272 15264
rect 12208 15204 12212 15260
rect 12212 15204 12268 15260
rect 12268 15204 12272 15260
rect 12208 15200 12272 15204
rect 12288 15260 12352 15264
rect 12288 15204 12292 15260
rect 12292 15204 12348 15260
rect 12348 15204 12352 15260
rect 12288 15200 12352 15204
rect 19445 15260 19509 15264
rect 19445 15204 19449 15260
rect 19449 15204 19505 15260
rect 19505 15204 19509 15260
rect 19445 15200 19509 15204
rect 19525 15260 19589 15264
rect 19525 15204 19529 15260
rect 19529 15204 19585 15260
rect 19585 15204 19589 15260
rect 19525 15200 19589 15204
rect 19605 15260 19669 15264
rect 19605 15204 19609 15260
rect 19609 15204 19665 15260
rect 19665 15204 19669 15260
rect 19605 15200 19669 15204
rect 19685 15260 19749 15264
rect 19685 15204 19689 15260
rect 19689 15204 19745 15260
rect 19745 15204 19749 15260
rect 19685 15200 19749 15204
rect 10180 15056 10244 15060
rect 10180 15000 10230 15056
rect 10230 15000 10244 15056
rect 10180 14996 10244 15000
rect 14780 14996 14844 15060
rect 8156 14860 8220 14924
rect 4476 14724 4540 14788
rect 8349 14716 8413 14720
rect 8349 14660 8353 14716
rect 8353 14660 8409 14716
rect 8409 14660 8413 14716
rect 8349 14656 8413 14660
rect 8429 14716 8493 14720
rect 8429 14660 8433 14716
rect 8433 14660 8489 14716
rect 8489 14660 8493 14716
rect 8429 14656 8493 14660
rect 8509 14716 8573 14720
rect 8509 14660 8513 14716
rect 8513 14660 8569 14716
rect 8569 14660 8573 14716
rect 8509 14656 8573 14660
rect 8589 14716 8653 14720
rect 8589 14660 8593 14716
rect 8593 14660 8649 14716
rect 8649 14660 8653 14716
rect 8589 14656 8653 14660
rect 15746 14716 15810 14720
rect 15746 14660 15750 14716
rect 15750 14660 15806 14716
rect 15806 14660 15810 14716
rect 15746 14656 15810 14660
rect 15826 14716 15890 14720
rect 15826 14660 15830 14716
rect 15830 14660 15886 14716
rect 15886 14660 15890 14716
rect 15826 14656 15890 14660
rect 15906 14716 15970 14720
rect 15906 14660 15910 14716
rect 15910 14660 15966 14716
rect 15966 14660 15970 14716
rect 15906 14656 15970 14660
rect 15986 14716 16050 14720
rect 15986 14660 15990 14716
rect 15990 14660 16046 14716
rect 16046 14660 16050 14716
rect 15986 14656 16050 14660
rect 4650 14172 4714 14176
rect 4650 14116 4654 14172
rect 4654 14116 4710 14172
rect 4710 14116 4714 14172
rect 4650 14112 4714 14116
rect 4730 14172 4794 14176
rect 4730 14116 4734 14172
rect 4734 14116 4790 14172
rect 4790 14116 4794 14172
rect 4730 14112 4794 14116
rect 4810 14172 4874 14176
rect 4810 14116 4814 14172
rect 4814 14116 4870 14172
rect 4870 14116 4874 14172
rect 4810 14112 4874 14116
rect 4890 14172 4954 14176
rect 4890 14116 4894 14172
rect 4894 14116 4950 14172
rect 4950 14116 4954 14172
rect 4890 14112 4954 14116
rect 13124 14180 13188 14244
rect 12048 14172 12112 14176
rect 12048 14116 12052 14172
rect 12052 14116 12108 14172
rect 12108 14116 12112 14172
rect 12048 14112 12112 14116
rect 12128 14172 12192 14176
rect 12128 14116 12132 14172
rect 12132 14116 12188 14172
rect 12188 14116 12192 14172
rect 12128 14112 12192 14116
rect 12208 14172 12272 14176
rect 12208 14116 12212 14172
rect 12212 14116 12268 14172
rect 12268 14116 12272 14172
rect 12208 14112 12272 14116
rect 12288 14172 12352 14176
rect 12288 14116 12292 14172
rect 12292 14116 12348 14172
rect 12348 14116 12352 14172
rect 12288 14112 12352 14116
rect 19445 14172 19509 14176
rect 19445 14116 19449 14172
rect 19449 14116 19505 14172
rect 19505 14116 19509 14172
rect 19445 14112 19509 14116
rect 19525 14172 19589 14176
rect 19525 14116 19529 14172
rect 19529 14116 19585 14172
rect 19585 14116 19589 14172
rect 19525 14112 19589 14116
rect 19605 14172 19669 14176
rect 19605 14116 19609 14172
rect 19609 14116 19665 14172
rect 19665 14116 19669 14172
rect 19605 14112 19669 14116
rect 19685 14172 19749 14176
rect 19685 14116 19689 14172
rect 19689 14116 19745 14172
rect 19745 14116 19749 14172
rect 19685 14112 19749 14116
rect 4292 13696 4356 13700
rect 4292 13640 4306 13696
rect 4306 13640 4356 13696
rect 4292 13636 4356 13640
rect 5212 13696 5276 13700
rect 5212 13640 5226 13696
rect 5226 13640 5276 13696
rect 5212 13636 5276 13640
rect 4476 13364 4540 13428
rect 15332 13772 15396 13836
rect 8349 13628 8413 13632
rect 8349 13572 8353 13628
rect 8353 13572 8409 13628
rect 8409 13572 8413 13628
rect 8349 13568 8413 13572
rect 8429 13628 8493 13632
rect 8429 13572 8433 13628
rect 8433 13572 8489 13628
rect 8489 13572 8493 13628
rect 8429 13568 8493 13572
rect 8509 13628 8573 13632
rect 8509 13572 8513 13628
rect 8513 13572 8569 13628
rect 8569 13572 8573 13628
rect 8509 13568 8573 13572
rect 8589 13628 8653 13632
rect 8589 13572 8593 13628
rect 8593 13572 8649 13628
rect 8649 13572 8653 13628
rect 8589 13568 8653 13572
rect 15746 13628 15810 13632
rect 15746 13572 15750 13628
rect 15750 13572 15806 13628
rect 15806 13572 15810 13628
rect 15746 13568 15810 13572
rect 15826 13628 15890 13632
rect 15826 13572 15830 13628
rect 15830 13572 15886 13628
rect 15886 13572 15890 13628
rect 15826 13568 15890 13572
rect 15906 13628 15970 13632
rect 15906 13572 15910 13628
rect 15910 13572 15966 13628
rect 15966 13572 15970 13628
rect 15906 13568 15970 13572
rect 15986 13628 16050 13632
rect 15986 13572 15990 13628
rect 15990 13572 16046 13628
rect 16046 13572 16050 13628
rect 15986 13568 16050 13572
rect 17908 13364 17972 13428
rect 4650 13084 4714 13088
rect 4650 13028 4654 13084
rect 4654 13028 4710 13084
rect 4710 13028 4714 13084
rect 4650 13024 4714 13028
rect 4730 13084 4794 13088
rect 4730 13028 4734 13084
rect 4734 13028 4790 13084
rect 4790 13028 4794 13084
rect 4730 13024 4794 13028
rect 4810 13084 4874 13088
rect 4810 13028 4814 13084
rect 4814 13028 4870 13084
rect 4870 13028 4874 13084
rect 4810 13024 4874 13028
rect 4890 13084 4954 13088
rect 4890 13028 4894 13084
rect 4894 13028 4950 13084
rect 4950 13028 4954 13084
rect 4890 13024 4954 13028
rect 12048 13084 12112 13088
rect 12048 13028 12052 13084
rect 12052 13028 12108 13084
rect 12108 13028 12112 13084
rect 12048 13024 12112 13028
rect 12128 13084 12192 13088
rect 12128 13028 12132 13084
rect 12132 13028 12188 13084
rect 12188 13028 12192 13084
rect 12128 13024 12192 13028
rect 12208 13084 12272 13088
rect 12208 13028 12212 13084
rect 12212 13028 12268 13084
rect 12268 13028 12272 13084
rect 12208 13024 12272 13028
rect 12288 13084 12352 13088
rect 12288 13028 12292 13084
rect 12292 13028 12348 13084
rect 12348 13028 12352 13084
rect 12288 13024 12352 13028
rect 19445 13084 19509 13088
rect 19445 13028 19449 13084
rect 19449 13028 19505 13084
rect 19505 13028 19509 13084
rect 19445 13024 19509 13028
rect 19525 13084 19589 13088
rect 19525 13028 19529 13084
rect 19529 13028 19585 13084
rect 19585 13028 19589 13084
rect 19525 13024 19589 13028
rect 19605 13084 19669 13088
rect 19605 13028 19609 13084
rect 19609 13028 19665 13084
rect 19665 13028 19669 13084
rect 19605 13024 19669 13028
rect 19685 13084 19749 13088
rect 19685 13028 19689 13084
rect 19689 13028 19745 13084
rect 19745 13028 19749 13084
rect 19685 13024 19749 13028
rect 5028 12684 5092 12748
rect 7236 12684 7300 12748
rect 17540 12684 17604 12748
rect 8349 12540 8413 12544
rect 8349 12484 8353 12540
rect 8353 12484 8409 12540
rect 8409 12484 8413 12540
rect 8349 12480 8413 12484
rect 8429 12540 8493 12544
rect 8429 12484 8433 12540
rect 8433 12484 8489 12540
rect 8489 12484 8493 12540
rect 8429 12480 8493 12484
rect 8509 12540 8573 12544
rect 8509 12484 8513 12540
rect 8513 12484 8569 12540
rect 8569 12484 8573 12540
rect 8509 12480 8573 12484
rect 8589 12540 8653 12544
rect 8589 12484 8593 12540
rect 8593 12484 8649 12540
rect 8649 12484 8653 12540
rect 8589 12480 8653 12484
rect 15746 12540 15810 12544
rect 15746 12484 15750 12540
rect 15750 12484 15806 12540
rect 15806 12484 15810 12540
rect 15746 12480 15810 12484
rect 15826 12540 15890 12544
rect 15826 12484 15830 12540
rect 15830 12484 15886 12540
rect 15886 12484 15890 12540
rect 15826 12480 15890 12484
rect 15906 12540 15970 12544
rect 15906 12484 15910 12540
rect 15910 12484 15966 12540
rect 15966 12484 15970 12540
rect 15906 12480 15970 12484
rect 15986 12540 16050 12544
rect 15986 12484 15990 12540
rect 15990 12484 16046 12540
rect 16046 12484 16050 12540
rect 15986 12480 16050 12484
rect 10180 12412 10244 12476
rect 18460 12412 18524 12476
rect 19196 12412 19260 12476
rect 6316 12336 6380 12340
rect 6316 12280 6330 12336
rect 6330 12280 6380 12336
rect 6316 12276 6380 12280
rect 9260 12336 9324 12340
rect 9260 12280 9274 12336
rect 9274 12280 9324 12336
rect 9260 12276 9324 12280
rect 11100 12276 11164 12340
rect 17908 12276 17972 12340
rect 9260 12200 9324 12204
rect 9260 12144 9310 12200
rect 9310 12144 9324 12200
rect 9260 12140 9324 12144
rect 20668 12140 20732 12204
rect 12940 12064 13004 12068
rect 12940 12008 12990 12064
rect 12990 12008 13004 12064
rect 12940 12004 13004 12008
rect 4650 11996 4714 12000
rect 4650 11940 4654 11996
rect 4654 11940 4710 11996
rect 4710 11940 4714 11996
rect 4650 11936 4714 11940
rect 4730 11996 4794 12000
rect 4730 11940 4734 11996
rect 4734 11940 4790 11996
rect 4790 11940 4794 11996
rect 4730 11936 4794 11940
rect 4810 11996 4874 12000
rect 4810 11940 4814 11996
rect 4814 11940 4870 11996
rect 4870 11940 4874 11996
rect 4810 11936 4874 11940
rect 4890 11996 4954 12000
rect 4890 11940 4894 11996
rect 4894 11940 4950 11996
rect 4950 11940 4954 11996
rect 4890 11936 4954 11940
rect 12048 11996 12112 12000
rect 12048 11940 12052 11996
rect 12052 11940 12108 11996
rect 12108 11940 12112 11996
rect 12048 11936 12112 11940
rect 12128 11996 12192 12000
rect 12128 11940 12132 11996
rect 12132 11940 12188 11996
rect 12188 11940 12192 11996
rect 12128 11936 12192 11940
rect 12208 11996 12272 12000
rect 12208 11940 12212 11996
rect 12212 11940 12268 11996
rect 12268 11940 12272 11996
rect 12208 11936 12272 11940
rect 12288 11996 12352 12000
rect 12288 11940 12292 11996
rect 12292 11940 12348 11996
rect 12348 11940 12352 11996
rect 12288 11936 12352 11940
rect 19445 11996 19509 12000
rect 19445 11940 19449 11996
rect 19449 11940 19505 11996
rect 19505 11940 19509 11996
rect 19445 11936 19509 11940
rect 19525 11996 19589 12000
rect 19525 11940 19529 11996
rect 19529 11940 19585 11996
rect 19585 11940 19589 11996
rect 19525 11936 19589 11940
rect 19605 11996 19669 12000
rect 19605 11940 19609 11996
rect 19609 11940 19665 11996
rect 19665 11940 19669 11996
rect 19605 11936 19669 11940
rect 19685 11996 19749 12000
rect 19685 11940 19689 11996
rect 19689 11940 19745 11996
rect 19745 11940 19749 11996
rect 19685 11936 19749 11940
rect 19012 11732 19076 11796
rect 16804 11596 16868 11660
rect 8349 11452 8413 11456
rect 8349 11396 8353 11452
rect 8353 11396 8409 11452
rect 8409 11396 8413 11452
rect 8349 11392 8413 11396
rect 8429 11452 8493 11456
rect 8429 11396 8433 11452
rect 8433 11396 8489 11452
rect 8489 11396 8493 11452
rect 8429 11392 8493 11396
rect 8509 11452 8573 11456
rect 8509 11396 8513 11452
rect 8513 11396 8569 11452
rect 8569 11396 8573 11452
rect 8509 11392 8573 11396
rect 8589 11452 8653 11456
rect 8589 11396 8593 11452
rect 8593 11396 8649 11452
rect 8649 11396 8653 11452
rect 8589 11392 8653 11396
rect 15746 11452 15810 11456
rect 15746 11396 15750 11452
rect 15750 11396 15806 11452
rect 15806 11396 15810 11452
rect 15746 11392 15810 11396
rect 15826 11452 15890 11456
rect 15826 11396 15830 11452
rect 15830 11396 15886 11452
rect 15886 11396 15890 11452
rect 15826 11392 15890 11396
rect 15906 11452 15970 11456
rect 15906 11396 15910 11452
rect 15910 11396 15966 11452
rect 15966 11396 15970 11452
rect 15906 11392 15970 11396
rect 15986 11452 16050 11456
rect 15986 11396 15990 11452
rect 15990 11396 16046 11452
rect 16046 11396 16050 11452
rect 15986 11392 16050 11396
rect 15148 11248 15212 11252
rect 15148 11192 15198 11248
rect 15198 11192 15212 11248
rect 15148 11188 15212 11192
rect 18276 11248 18340 11252
rect 18276 11192 18290 11248
rect 18290 11192 18340 11248
rect 18276 11188 18340 11192
rect 4650 10908 4714 10912
rect 4650 10852 4654 10908
rect 4654 10852 4710 10908
rect 4710 10852 4714 10908
rect 4650 10848 4714 10852
rect 4730 10908 4794 10912
rect 4730 10852 4734 10908
rect 4734 10852 4790 10908
rect 4790 10852 4794 10908
rect 4730 10848 4794 10852
rect 4810 10908 4874 10912
rect 4810 10852 4814 10908
rect 4814 10852 4870 10908
rect 4870 10852 4874 10908
rect 4810 10848 4874 10852
rect 4890 10908 4954 10912
rect 4890 10852 4894 10908
rect 4894 10852 4950 10908
rect 4950 10852 4954 10908
rect 4890 10848 4954 10852
rect 14780 11052 14844 11116
rect 12048 10908 12112 10912
rect 12048 10852 12052 10908
rect 12052 10852 12108 10908
rect 12108 10852 12112 10908
rect 12048 10848 12112 10852
rect 12128 10908 12192 10912
rect 12128 10852 12132 10908
rect 12132 10852 12188 10908
rect 12188 10852 12192 10908
rect 12128 10848 12192 10852
rect 12208 10908 12272 10912
rect 12208 10852 12212 10908
rect 12212 10852 12268 10908
rect 12268 10852 12272 10908
rect 12208 10848 12272 10852
rect 12288 10908 12352 10912
rect 12288 10852 12292 10908
rect 12292 10852 12348 10908
rect 12348 10852 12352 10908
rect 12288 10848 12352 10852
rect 19445 10908 19509 10912
rect 19445 10852 19449 10908
rect 19449 10852 19505 10908
rect 19505 10852 19509 10908
rect 19445 10848 19509 10852
rect 19525 10908 19589 10912
rect 19525 10852 19529 10908
rect 19529 10852 19585 10908
rect 19585 10852 19589 10908
rect 19525 10848 19589 10852
rect 19605 10908 19669 10912
rect 19605 10852 19609 10908
rect 19609 10852 19665 10908
rect 19665 10852 19669 10908
rect 19605 10848 19669 10852
rect 19685 10908 19749 10912
rect 19685 10852 19689 10908
rect 19689 10852 19745 10908
rect 19745 10852 19749 10908
rect 19685 10848 19749 10852
rect 6316 10704 6380 10708
rect 6316 10648 6366 10704
rect 6366 10648 6380 10704
rect 6316 10644 6380 10648
rect 17724 10372 17788 10436
rect 8349 10364 8413 10368
rect 8349 10308 8353 10364
rect 8353 10308 8409 10364
rect 8409 10308 8413 10364
rect 8349 10304 8413 10308
rect 8429 10364 8493 10368
rect 8429 10308 8433 10364
rect 8433 10308 8489 10364
rect 8489 10308 8493 10364
rect 8429 10304 8493 10308
rect 8509 10364 8573 10368
rect 8509 10308 8513 10364
rect 8513 10308 8569 10364
rect 8569 10308 8573 10364
rect 8509 10304 8573 10308
rect 8589 10364 8653 10368
rect 8589 10308 8593 10364
rect 8593 10308 8649 10364
rect 8649 10308 8653 10364
rect 8589 10304 8653 10308
rect 15746 10364 15810 10368
rect 15746 10308 15750 10364
rect 15750 10308 15806 10364
rect 15806 10308 15810 10364
rect 15746 10304 15810 10308
rect 15826 10364 15890 10368
rect 15826 10308 15830 10364
rect 15830 10308 15886 10364
rect 15886 10308 15890 10364
rect 15826 10304 15890 10308
rect 15906 10364 15970 10368
rect 15906 10308 15910 10364
rect 15910 10308 15966 10364
rect 15966 10308 15970 10364
rect 15906 10304 15970 10308
rect 15986 10364 16050 10368
rect 15986 10308 15990 10364
rect 15990 10308 16046 10364
rect 16046 10308 16050 10364
rect 15986 10304 16050 10308
rect 7420 10100 7484 10164
rect 4650 9820 4714 9824
rect 4650 9764 4654 9820
rect 4654 9764 4710 9820
rect 4710 9764 4714 9820
rect 4650 9760 4714 9764
rect 4730 9820 4794 9824
rect 4730 9764 4734 9820
rect 4734 9764 4790 9820
rect 4790 9764 4794 9820
rect 4730 9760 4794 9764
rect 4810 9820 4874 9824
rect 4810 9764 4814 9820
rect 4814 9764 4870 9820
rect 4870 9764 4874 9820
rect 4810 9760 4874 9764
rect 4890 9820 4954 9824
rect 4890 9764 4894 9820
rect 4894 9764 4950 9820
rect 4950 9764 4954 9820
rect 4890 9760 4954 9764
rect 12048 9820 12112 9824
rect 12048 9764 12052 9820
rect 12052 9764 12108 9820
rect 12108 9764 12112 9820
rect 12048 9760 12112 9764
rect 12128 9820 12192 9824
rect 12128 9764 12132 9820
rect 12132 9764 12188 9820
rect 12188 9764 12192 9820
rect 12128 9760 12192 9764
rect 12208 9820 12272 9824
rect 12208 9764 12212 9820
rect 12212 9764 12268 9820
rect 12268 9764 12272 9820
rect 12208 9760 12272 9764
rect 12288 9820 12352 9824
rect 12288 9764 12292 9820
rect 12292 9764 12348 9820
rect 12348 9764 12352 9820
rect 12288 9760 12352 9764
rect 19445 9820 19509 9824
rect 19445 9764 19449 9820
rect 19449 9764 19505 9820
rect 19505 9764 19509 9820
rect 19445 9760 19509 9764
rect 19525 9820 19589 9824
rect 19525 9764 19529 9820
rect 19529 9764 19585 9820
rect 19585 9764 19589 9820
rect 19525 9760 19589 9764
rect 19605 9820 19669 9824
rect 19605 9764 19609 9820
rect 19609 9764 19665 9820
rect 19665 9764 19669 9820
rect 19605 9760 19669 9764
rect 19685 9820 19749 9824
rect 19685 9764 19689 9820
rect 19689 9764 19745 9820
rect 19745 9764 19749 9820
rect 19685 9760 19749 9764
rect 14964 9692 15028 9756
rect 9444 9556 9508 9620
rect 18092 9556 18156 9620
rect 18828 9556 18892 9620
rect 10916 9420 10980 9484
rect 11836 9420 11900 9484
rect 10180 9344 10244 9348
rect 10180 9288 10230 9344
rect 10230 9288 10244 9344
rect 10180 9284 10244 9288
rect 10364 9284 10428 9348
rect 8349 9276 8413 9280
rect 8349 9220 8353 9276
rect 8353 9220 8409 9276
rect 8409 9220 8413 9276
rect 8349 9216 8413 9220
rect 8429 9276 8493 9280
rect 8429 9220 8433 9276
rect 8433 9220 8489 9276
rect 8489 9220 8493 9276
rect 8429 9216 8493 9220
rect 8509 9276 8573 9280
rect 8509 9220 8513 9276
rect 8513 9220 8569 9276
rect 8569 9220 8573 9276
rect 8509 9216 8573 9220
rect 8589 9276 8653 9280
rect 8589 9220 8593 9276
rect 8593 9220 8649 9276
rect 8649 9220 8653 9276
rect 8589 9216 8653 9220
rect 15746 9276 15810 9280
rect 15746 9220 15750 9276
rect 15750 9220 15806 9276
rect 15806 9220 15810 9276
rect 15746 9216 15810 9220
rect 15826 9276 15890 9280
rect 15826 9220 15830 9276
rect 15830 9220 15886 9276
rect 15886 9220 15890 9276
rect 15826 9216 15890 9220
rect 15906 9276 15970 9280
rect 15906 9220 15910 9276
rect 15910 9220 15966 9276
rect 15966 9220 15970 9276
rect 15906 9216 15970 9220
rect 15986 9276 16050 9280
rect 15986 9220 15990 9276
rect 15990 9220 16046 9276
rect 16046 9220 16050 9276
rect 15986 9216 16050 9220
rect 9260 9072 9324 9076
rect 9260 9016 9310 9072
rect 9310 9016 9324 9072
rect 9260 9012 9324 9016
rect 20668 9012 20732 9076
rect 7788 8876 7852 8940
rect 9812 8740 9876 8804
rect 4650 8732 4714 8736
rect 4650 8676 4654 8732
rect 4654 8676 4710 8732
rect 4710 8676 4714 8732
rect 4650 8672 4714 8676
rect 4730 8732 4794 8736
rect 4730 8676 4734 8732
rect 4734 8676 4790 8732
rect 4790 8676 4794 8732
rect 4730 8672 4794 8676
rect 4810 8732 4874 8736
rect 4810 8676 4814 8732
rect 4814 8676 4870 8732
rect 4870 8676 4874 8732
rect 4810 8672 4874 8676
rect 4890 8732 4954 8736
rect 4890 8676 4894 8732
rect 4894 8676 4950 8732
rect 4950 8676 4954 8732
rect 4890 8672 4954 8676
rect 12048 8732 12112 8736
rect 12048 8676 12052 8732
rect 12052 8676 12108 8732
rect 12108 8676 12112 8732
rect 12048 8672 12112 8676
rect 12128 8732 12192 8736
rect 12128 8676 12132 8732
rect 12132 8676 12188 8732
rect 12188 8676 12192 8732
rect 12128 8672 12192 8676
rect 12208 8732 12272 8736
rect 12208 8676 12212 8732
rect 12212 8676 12268 8732
rect 12268 8676 12272 8732
rect 12208 8672 12272 8676
rect 12288 8732 12352 8736
rect 12288 8676 12292 8732
rect 12292 8676 12348 8732
rect 12348 8676 12352 8732
rect 12288 8672 12352 8676
rect 7052 8664 7116 8668
rect 7052 8608 7066 8664
rect 7066 8608 7116 8664
rect 7052 8604 7116 8608
rect 7420 8604 7484 8668
rect 5028 8528 5092 8532
rect 5028 8472 5078 8528
rect 5078 8472 5092 8528
rect 5028 8468 5092 8472
rect 7972 8468 8036 8532
rect 13124 8468 13188 8532
rect 18276 8876 18340 8940
rect 19445 8732 19509 8736
rect 19445 8676 19449 8732
rect 19449 8676 19505 8732
rect 19505 8676 19509 8732
rect 19445 8672 19509 8676
rect 19525 8732 19589 8736
rect 19525 8676 19529 8732
rect 19529 8676 19585 8732
rect 19585 8676 19589 8732
rect 19525 8672 19589 8676
rect 19605 8732 19669 8736
rect 19605 8676 19609 8732
rect 19609 8676 19665 8732
rect 19665 8676 19669 8732
rect 19605 8672 19669 8676
rect 19685 8732 19749 8736
rect 19685 8676 19689 8732
rect 19689 8676 19745 8732
rect 19745 8676 19749 8732
rect 19685 8672 19749 8676
rect 5948 8256 6012 8260
rect 5948 8200 5962 8256
rect 5962 8200 6012 8256
rect 5948 8196 6012 8200
rect 10180 8332 10244 8396
rect 13860 8196 13924 8260
rect 8349 8188 8413 8192
rect 8349 8132 8353 8188
rect 8353 8132 8409 8188
rect 8409 8132 8413 8188
rect 8349 8128 8413 8132
rect 8429 8188 8493 8192
rect 8429 8132 8433 8188
rect 8433 8132 8489 8188
rect 8489 8132 8493 8188
rect 8429 8128 8493 8132
rect 8509 8188 8573 8192
rect 8509 8132 8513 8188
rect 8513 8132 8569 8188
rect 8569 8132 8573 8188
rect 8509 8128 8573 8132
rect 8589 8188 8653 8192
rect 8589 8132 8593 8188
rect 8593 8132 8649 8188
rect 8649 8132 8653 8188
rect 8589 8128 8653 8132
rect 15746 8188 15810 8192
rect 15746 8132 15750 8188
rect 15750 8132 15806 8188
rect 15806 8132 15810 8188
rect 15746 8128 15810 8132
rect 15826 8188 15890 8192
rect 15826 8132 15830 8188
rect 15830 8132 15886 8188
rect 15886 8132 15890 8188
rect 15826 8128 15890 8132
rect 15906 8188 15970 8192
rect 15906 8132 15910 8188
rect 15910 8132 15966 8188
rect 15966 8132 15970 8188
rect 15906 8128 15970 8132
rect 15986 8188 16050 8192
rect 15986 8132 15990 8188
rect 15990 8132 16046 8188
rect 16046 8132 16050 8188
rect 15986 8128 16050 8132
rect 8892 8060 8956 8124
rect 18092 8060 18156 8124
rect 20852 8060 20916 8124
rect 7236 7652 7300 7716
rect 10916 7652 10980 7716
rect 4650 7644 4714 7648
rect 4650 7588 4654 7644
rect 4654 7588 4710 7644
rect 4710 7588 4714 7644
rect 4650 7584 4714 7588
rect 4730 7644 4794 7648
rect 4730 7588 4734 7644
rect 4734 7588 4790 7644
rect 4790 7588 4794 7644
rect 4730 7584 4794 7588
rect 4810 7644 4874 7648
rect 4810 7588 4814 7644
rect 4814 7588 4870 7644
rect 4870 7588 4874 7644
rect 4810 7584 4874 7588
rect 4890 7644 4954 7648
rect 4890 7588 4894 7644
rect 4894 7588 4950 7644
rect 4950 7588 4954 7644
rect 4890 7584 4954 7588
rect 12048 7644 12112 7648
rect 12048 7588 12052 7644
rect 12052 7588 12108 7644
rect 12108 7588 12112 7644
rect 12048 7584 12112 7588
rect 12128 7644 12192 7648
rect 12128 7588 12132 7644
rect 12132 7588 12188 7644
rect 12188 7588 12192 7644
rect 12128 7584 12192 7588
rect 12208 7644 12272 7648
rect 12208 7588 12212 7644
rect 12212 7588 12268 7644
rect 12268 7588 12272 7644
rect 12208 7584 12272 7588
rect 12288 7644 12352 7648
rect 12288 7588 12292 7644
rect 12292 7588 12348 7644
rect 12348 7588 12352 7644
rect 12288 7584 12352 7588
rect 7788 7516 7852 7580
rect 17540 7516 17604 7580
rect 8156 7380 8220 7444
rect 9076 7380 9140 7444
rect 18460 7380 18524 7444
rect 19445 7644 19509 7648
rect 19445 7588 19449 7644
rect 19449 7588 19505 7644
rect 19505 7588 19509 7644
rect 19445 7584 19509 7588
rect 19525 7644 19589 7648
rect 19525 7588 19529 7644
rect 19529 7588 19585 7644
rect 19585 7588 19589 7644
rect 19525 7584 19589 7588
rect 19605 7644 19669 7648
rect 19605 7588 19609 7644
rect 19609 7588 19665 7644
rect 19665 7588 19669 7644
rect 19605 7584 19669 7588
rect 19685 7644 19749 7648
rect 19685 7588 19689 7644
rect 19689 7588 19745 7644
rect 19745 7588 19749 7644
rect 19685 7584 19749 7588
rect 20300 7380 20364 7444
rect 7052 7304 7116 7308
rect 7052 7248 7066 7304
rect 7066 7248 7116 7304
rect 7052 7244 7116 7248
rect 9812 7108 9876 7172
rect 13676 7244 13740 7308
rect 8349 7100 8413 7104
rect 8349 7044 8353 7100
rect 8353 7044 8409 7100
rect 8409 7044 8413 7100
rect 8349 7040 8413 7044
rect 8429 7100 8493 7104
rect 8429 7044 8433 7100
rect 8433 7044 8489 7100
rect 8489 7044 8493 7100
rect 8429 7040 8493 7044
rect 8509 7100 8573 7104
rect 8509 7044 8513 7100
rect 8513 7044 8569 7100
rect 8569 7044 8573 7100
rect 8509 7040 8573 7044
rect 8589 7100 8653 7104
rect 8589 7044 8593 7100
rect 8593 7044 8649 7100
rect 8649 7044 8653 7100
rect 8589 7040 8653 7044
rect 15746 7100 15810 7104
rect 15746 7044 15750 7100
rect 15750 7044 15806 7100
rect 15806 7044 15810 7100
rect 15746 7040 15810 7044
rect 15826 7100 15890 7104
rect 15826 7044 15830 7100
rect 15830 7044 15886 7100
rect 15886 7044 15890 7100
rect 15826 7040 15890 7044
rect 15906 7100 15970 7104
rect 15906 7044 15910 7100
rect 15910 7044 15966 7100
rect 15966 7044 15970 7100
rect 15906 7040 15970 7044
rect 15986 7100 16050 7104
rect 15986 7044 15990 7100
rect 15990 7044 16046 7100
rect 16046 7044 16050 7100
rect 15986 7040 16050 7044
rect 8892 6972 8956 7036
rect 13124 6564 13188 6628
rect 19196 6564 19260 6628
rect 4650 6556 4714 6560
rect 4650 6500 4654 6556
rect 4654 6500 4710 6556
rect 4710 6500 4714 6556
rect 4650 6496 4714 6500
rect 4730 6556 4794 6560
rect 4730 6500 4734 6556
rect 4734 6500 4790 6556
rect 4790 6500 4794 6556
rect 4730 6496 4794 6500
rect 4810 6556 4874 6560
rect 4810 6500 4814 6556
rect 4814 6500 4870 6556
rect 4870 6500 4874 6556
rect 4810 6496 4874 6500
rect 4890 6556 4954 6560
rect 4890 6500 4894 6556
rect 4894 6500 4950 6556
rect 4950 6500 4954 6556
rect 4890 6496 4954 6500
rect 12048 6556 12112 6560
rect 12048 6500 12052 6556
rect 12052 6500 12108 6556
rect 12108 6500 12112 6556
rect 12048 6496 12112 6500
rect 12128 6556 12192 6560
rect 12128 6500 12132 6556
rect 12132 6500 12188 6556
rect 12188 6500 12192 6556
rect 12128 6496 12192 6500
rect 12208 6556 12272 6560
rect 12208 6500 12212 6556
rect 12212 6500 12268 6556
rect 12268 6500 12272 6556
rect 12208 6496 12272 6500
rect 12288 6556 12352 6560
rect 12288 6500 12292 6556
rect 12292 6500 12348 6556
rect 12348 6500 12352 6556
rect 12288 6496 12352 6500
rect 19445 6556 19509 6560
rect 19445 6500 19449 6556
rect 19449 6500 19505 6556
rect 19505 6500 19509 6556
rect 19445 6496 19509 6500
rect 19525 6556 19589 6560
rect 19525 6500 19529 6556
rect 19529 6500 19585 6556
rect 19585 6500 19589 6556
rect 19525 6496 19589 6500
rect 19605 6556 19669 6560
rect 19605 6500 19609 6556
rect 19609 6500 19665 6556
rect 19665 6500 19669 6556
rect 19605 6496 19669 6500
rect 19685 6556 19749 6560
rect 19685 6500 19689 6556
rect 19689 6500 19745 6556
rect 19745 6500 19749 6556
rect 19685 6496 19749 6500
rect 13124 6156 13188 6220
rect 8349 6012 8413 6016
rect 8349 5956 8353 6012
rect 8353 5956 8409 6012
rect 8409 5956 8413 6012
rect 8349 5952 8413 5956
rect 8429 6012 8493 6016
rect 8429 5956 8433 6012
rect 8433 5956 8489 6012
rect 8489 5956 8493 6012
rect 8429 5952 8493 5956
rect 8509 6012 8573 6016
rect 8509 5956 8513 6012
rect 8513 5956 8569 6012
rect 8569 5956 8573 6012
rect 8509 5952 8573 5956
rect 8589 6012 8653 6016
rect 8589 5956 8593 6012
rect 8593 5956 8649 6012
rect 8649 5956 8653 6012
rect 8589 5952 8653 5956
rect 15746 6012 15810 6016
rect 15746 5956 15750 6012
rect 15750 5956 15806 6012
rect 15806 5956 15810 6012
rect 15746 5952 15810 5956
rect 15826 6012 15890 6016
rect 15826 5956 15830 6012
rect 15830 5956 15886 6012
rect 15886 5956 15890 6012
rect 15826 5952 15890 5956
rect 15906 6012 15970 6016
rect 15906 5956 15910 6012
rect 15910 5956 15966 6012
rect 15966 5956 15970 6012
rect 15906 5952 15970 5956
rect 15986 6012 16050 6016
rect 15986 5956 15990 6012
rect 15990 5956 16046 6012
rect 16046 5956 16050 6012
rect 15986 5952 16050 5956
rect 9444 5884 9508 5948
rect 15148 5884 15212 5948
rect 11836 5748 11900 5812
rect 12940 5536 13004 5540
rect 12940 5480 12954 5536
rect 12954 5480 13004 5536
rect 12940 5476 13004 5480
rect 13676 5536 13740 5540
rect 13676 5480 13690 5536
rect 13690 5480 13740 5536
rect 13676 5476 13740 5480
rect 4650 5468 4714 5472
rect 4650 5412 4654 5468
rect 4654 5412 4710 5468
rect 4710 5412 4714 5468
rect 4650 5408 4714 5412
rect 4730 5468 4794 5472
rect 4730 5412 4734 5468
rect 4734 5412 4790 5468
rect 4790 5412 4794 5468
rect 4730 5408 4794 5412
rect 4810 5468 4874 5472
rect 4810 5412 4814 5468
rect 4814 5412 4870 5468
rect 4870 5412 4874 5468
rect 4810 5408 4874 5412
rect 4890 5468 4954 5472
rect 4890 5412 4894 5468
rect 4894 5412 4950 5468
rect 4950 5412 4954 5468
rect 4890 5408 4954 5412
rect 12048 5468 12112 5472
rect 12048 5412 12052 5468
rect 12052 5412 12108 5468
rect 12108 5412 12112 5468
rect 12048 5408 12112 5412
rect 12128 5468 12192 5472
rect 12128 5412 12132 5468
rect 12132 5412 12188 5468
rect 12188 5412 12192 5468
rect 12128 5408 12192 5412
rect 12208 5468 12272 5472
rect 12208 5412 12212 5468
rect 12212 5412 12268 5468
rect 12268 5412 12272 5468
rect 12208 5408 12272 5412
rect 12288 5468 12352 5472
rect 12288 5412 12292 5468
rect 12292 5412 12348 5468
rect 12348 5412 12352 5468
rect 12288 5408 12352 5412
rect 19445 5468 19509 5472
rect 19445 5412 19449 5468
rect 19449 5412 19505 5468
rect 19505 5412 19509 5468
rect 19445 5408 19509 5412
rect 19525 5468 19589 5472
rect 19525 5412 19529 5468
rect 19529 5412 19585 5468
rect 19585 5412 19589 5468
rect 19525 5408 19589 5412
rect 19605 5468 19669 5472
rect 19605 5412 19609 5468
rect 19609 5412 19665 5468
rect 19665 5412 19669 5468
rect 19605 5408 19669 5412
rect 19685 5468 19749 5472
rect 19685 5412 19689 5468
rect 19689 5412 19745 5468
rect 19745 5412 19749 5468
rect 19685 5408 19749 5412
rect 7604 5340 7668 5404
rect 16804 5204 16868 5268
rect 8349 4924 8413 4928
rect 8349 4868 8353 4924
rect 8353 4868 8409 4924
rect 8409 4868 8413 4924
rect 8349 4864 8413 4868
rect 8429 4924 8493 4928
rect 8429 4868 8433 4924
rect 8433 4868 8489 4924
rect 8489 4868 8493 4924
rect 8429 4864 8493 4868
rect 8509 4924 8573 4928
rect 8509 4868 8513 4924
rect 8513 4868 8569 4924
rect 8569 4868 8573 4924
rect 8509 4864 8573 4868
rect 8589 4924 8653 4928
rect 8589 4868 8593 4924
rect 8593 4868 8649 4924
rect 8649 4868 8653 4924
rect 8589 4864 8653 4868
rect 15746 4924 15810 4928
rect 15746 4868 15750 4924
rect 15750 4868 15806 4924
rect 15806 4868 15810 4924
rect 15746 4864 15810 4868
rect 15826 4924 15890 4928
rect 15826 4868 15830 4924
rect 15830 4868 15886 4924
rect 15886 4868 15890 4924
rect 15826 4864 15890 4868
rect 15906 4924 15970 4928
rect 15906 4868 15910 4924
rect 15910 4868 15966 4924
rect 15966 4868 15970 4924
rect 15906 4864 15970 4868
rect 15986 4924 16050 4928
rect 15986 4868 15990 4924
rect 15990 4868 16046 4924
rect 16046 4868 16050 4924
rect 15986 4864 16050 4868
rect 10364 4796 10428 4860
rect 19012 4660 19076 4724
rect 20668 4524 20732 4588
rect 16620 4388 16684 4452
rect 4650 4380 4714 4384
rect 4650 4324 4654 4380
rect 4654 4324 4710 4380
rect 4710 4324 4714 4380
rect 4650 4320 4714 4324
rect 4730 4380 4794 4384
rect 4730 4324 4734 4380
rect 4734 4324 4790 4380
rect 4790 4324 4794 4380
rect 4730 4320 4794 4324
rect 4810 4380 4874 4384
rect 4810 4324 4814 4380
rect 4814 4324 4870 4380
rect 4870 4324 4874 4380
rect 4810 4320 4874 4324
rect 4890 4380 4954 4384
rect 4890 4324 4894 4380
rect 4894 4324 4950 4380
rect 4950 4324 4954 4380
rect 4890 4320 4954 4324
rect 12048 4380 12112 4384
rect 12048 4324 12052 4380
rect 12052 4324 12108 4380
rect 12108 4324 12112 4380
rect 12048 4320 12112 4324
rect 12128 4380 12192 4384
rect 12128 4324 12132 4380
rect 12132 4324 12188 4380
rect 12188 4324 12192 4380
rect 12128 4320 12192 4324
rect 12208 4380 12272 4384
rect 12208 4324 12212 4380
rect 12212 4324 12268 4380
rect 12268 4324 12272 4380
rect 12208 4320 12272 4324
rect 12288 4380 12352 4384
rect 12288 4324 12292 4380
rect 12292 4324 12348 4380
rect 12348 4324 12352 4380
rect 12288 4320 12352 4324
rect 19445 4380 19509 4384
rect 19445 4324 19449 4380
rect 19449 4324 19505 4380
rect 19505 4324 19509 4380
rect 19445 4320 19509 4324
rect 19525 4380 19589 4384
rect 19525 4324 19529 4380
rect 19529 4324 19585 4380
rect 19585 4324 19589 4380
rect 19525 4320 19589 4324
rect 19605 4380 19669 4384
rect 19605 4324 19609 4380
rect 19609 4324 19665 4380
rect 19665 4324 19669 4380
rect 19605 4320 19669 4324
rect 19685 4380 19749 4384
rect 19685 4324 19689 4380
rect 19689 4324 19745 4380
rect 19745 4324 19749 4380
rect 19685 4320 19749 4324
rect 8349 3836 8413 3840
rect 8349 3780 8353 3836
rect 8353 3780 8409 3836
rect 8409 3780 8413 3836
rect 8349 3776 8413 3780
rect 8429 3836 8493 3840
rect 8429 3780 8433 3836
rect 8433 3780 8489 3836
rect 8489 3780 8493 3836
rect 8429 3776 8493 3780
rect 8509 3836 8573 3840
rect 8509 3780 8513 3836
rect 8513 3780 8569 3836
rect 8569 3780 8573 3836
rect 8509 3776 8573 3780
rect 8589 3836 8653 3840
rect 8589 3780 8593 3836
rect 8593 3780 8649 3836
rect 8649 3780 8653 3836
rect 8589 3776 8653 3780
rect 15746 3836 15810 3840
rect 15746 3780 15750 3836
rect 15750 3780 15806 3836
rect 15806 3780 15810 3836
rect 15746 3776 15810 3780
rect 15826 3836 15890 3840
rect 15826 3780 15830 3836
rect 15830 3780 15886 3836
rect 15886 3780 15890 3836
rect 15826 3776 15890 3780
rect 15906 3836 15970 3840
rect 15906 3780 15910 3836
rect 15910 3780 15966 3836
rect 15966 3780 15970 3836
rect 15906 3776 15970 3780
rect 15986 3836 16050 3840
rect 15986 3780 15990 3836
rect 15990 3780 16046 3836
rect 16046 3780 16050 3836
rect 15986 3776 16050 3780
rect 20852 3708 20916 3772
rect 18828 3572 18892 3636
rect 19932 3436 19996 3500
rect 19932 3300 19996 3364
rect 20484 3300 20548 3364
rect 4650 3292 4714 3296
rect 4650 3236 4654 3292
rect 4654 3236 4710 3292
rect 4710 3236 4714 3292
rect 4650 3232 4714 3236
rect 4730 3292 4794 3296
rect 4730 3236 4734 3292
rect 4734 3236 4790 3292
rect 4790 3236 4794 3292
rect 4730 3232 4794 3236
rect 4810 3292 4874 3296
rect 4810 3236 4814 3292
rect 4814 3236 4870 3292
rect 4870 3236 4874 3292
rect 4810 3232 4874 3236
rect 4890 3292 4954 3296
rect 4890 3236 4894 3292
rect 4894 3236 4950 3292
rect 4950 3236 4954 3292
rect 4890 3232 4954 3236
rect 12048 3292 12112 3296
rect 12048 3236 12052 3292
rect 12052 3236 12108 3292
rect 12108 3236 12112 3292
rect 12048 3232 12112 3236
rect 12128 3292 12192 3296
rect 12128 3236 12132 3292
rect 12132 3236 12188 3292
rect 12188 3236 12192 3292
rect 12128 3232 12192 3236
rect 12208 3292 12272 3296
rect 12208 3236 12212 3292
rect 12212 3236 12268 3292
rect 12268 3236 12272 3292
rect 12208 3232 12272 3236
rect 12288 3292 12352 3296
rect 12288 3236 12292 3292
rect 12292 3236 12348 3292
rect 12348 3236 12352 3292
rect 12288 3232 12352 3236
rect 19445 3292 19509 3296
rect 19445 3236 19449 3292
rect 19449 3236 19505 3292
rect 19505 3236 19509 3292
rect 19445 3232 19509 3236
rect 19525 3292 19589 3296
rect 19525 3236 19529 3292
rect 19529 3236 19585 3292
rect 19585 3236 19589 3292
rect 19525 3232 19589 3236
rect 19605 3292 19669 3296
rect 19605 3236 19609 3292
rect 19609 3236 19665 3292
rect 19665 3236 19669 3292
rect 19605 3232 19669 3236
rect 19685 3292 19749 3296
rect 19685 3236 19689 3292
rect 19689 3236 19745 3292
rect 19745 3236 19749 3292
rect 19685 3232 19749 3236
rect 16988 3164 17052 3228
rect 15516 3028 15580 3092
rect 19932 2892 19996 2956
rect 20116 2756 20180 2820
rect 8349 2748 8413 2752
rect 8349 2692 8353 2748
rect 8353 2692 8409 2748
rect 8409 2692 8413 2748
rect 8349 2688 8413 2692
rect 8429 2748 8493 2752
rect 8429 2692 8433 2748
rect 8433 2692 8489 2748
rect 8489 2692 8493 2748
rect 8429 2688 8493 2692
rect 8509 2748 8573 2752
rect 8509 2692 8513 2748
rect 8513 2692 8569 2748
rect 8569 2692 8573 2748
rect 8509 2688 8573 2692
rect 8589 2748 8653 2752
rect 8589 2692 8593 2748
rect 8593 2692 8649 2748
rect 8649 2692 8653 2748
rect 8589 2688 8653 2692
rect 15746 2748 15810 2752
rect 15746 2692 15750 2748
rect 15750 2692 15806 2748
rect 15806 2692 15810 2748
rect 15746 2688 15810 2692
rect 15826 2748 15890 2752
rect 15826 2692 15830 2748
rect 15830 2692 15886 2748
rect 15886 2692 15890 2748
rect 15826 2688 15890 2692
rect 15906 2748 15970 2752
rect 15906 2692 15910 2748
rect 15910 2692 15966 2748
rect 15966 2692 15970 2748
rect 15906 2688 15970 2692
rect 15986 2748 16050 2752
rect 15986 2692 15990 2748
rect 15990 2692 16046 2748
rect 16046 2692 16050 2748
rect 15986 2688 16050 2692
rect 15332 2620 15396 2684
rect 8892 2348 8956 2412
rect 16620 2348 16684 2412
rect 4650 2204 4714 2208
rect 4650 2148 4654 2204
rect 4654 2148 4710 2204
rect 4710 2148 4714 2204
rect 4650 2144 4714 2148
rect 4730 2204 4794 2208
rect 4730 2148 4734 2204
rect 4734 2148 4790 2204
rect 4790 2148 4794 2204
rect 4730 2144 4794 2148
rect 4810 2204 4874 2208
rect 4810 2148 4814 2204
rect 4814 2148 4870 2204
rect 4870 2148 4874 2204
rect 4810 2144 4874 2148
rect 4890 2204 4954 2208
rect 4890 2148 4894 2204
rect 4894 2148 4950 2204
rect 4950 2148 4954 2204
rect 4890 2144 4954 2148
rect 12048 2204 12112 2208
rect 12048 2148 12052 2204
rect 12052 2148 12108 2204
rect 12108 2148 12112 2204
rect 12048 2144 12112 2148
rect 12128 2204 12192 2208
rect 12128 2148 12132 2204
rect 12132 2148 12188 2204
rect 12188 2148 12192 2204
rect 12128 2144 12192 2148
rect 12208 2204 12272 2208
rect 12208 2148 12212 2204
rect 12212 2148 12268 2204
rect 12268 2148 12272 2204
rect 12208 2144 12272 2148
rect 12288 2204 12352 2208
rect 12288 2148 12292 2204
rect 12292 2148 12348 2204
rect 12348 2148 12352 2204
rect 12288 2144 12352 2148
rect 19445 2204 19509 2208
rect 19445 2148 19449 2204
rect 19449 2148 19505 2204
rect 19505 2148 19509 2204
rect 19445 2144 19509 2148
rect 19525 2204 19589 2208
rect 19525 2148 19529 2204
rect 19529 2148 19585 2204
rect 19585 2148 19589 2204
rect 19525 2144 19589 2148
rect 19605 2204 19669 2208
rect 19605 2148 19609 2204
rect 19609 2148 19665 2204
rect 19665 2148 19669 2204
rect 19605 2144 19669 2148
rect 19685 2204 19749 2208
rect 19685 2148 19689 2204
rect 19689 2148 19745 2204
rect 19745 2148 19749 2204
rect 19685 2144 19749 2148
<< metal4 >>
rect 4642 21792 4963 21808
rect 4642 21728 4650 21792
rect 4714 21728 4730 21792
rect 4794 21728 4810 21792
rect 4874 21728 4890 21792
rect 4954 21728 4963 21792
rect 4642 20704 4963 21728
rect 8341 21248 8661 21808
rect 8341 21184 8349 21248
rect 8413 21184 8429 21248
rect 8493 21184 8509 21248
rect 8573 21184 8589 21248
rect 8653 21184 8661 21248
rect 7603 21044 7669 21045
rect 7603 20980 7604 21044
rect 7668 20980 7669 21044
rect 7603 20979 7669 20980
rect 4642 20640 4650 20704
rect 4714 20640 4730 20704
rect 4794 20640 4810 20704
rect 4874 20640 4890 20704
rect 4954 20640 4963 20704
rect 4642 19616 4963 20640
rect 7606 20365 7666 20979
rect 7603 20364 7669 20365
rect 7603 20300 7604 20364
rect 7668 20300 7669 20364
rect 7603 20299 7669 20300
rect 5947 19956 6013 19957
rect 5947 19892 5948 19956
rect 6012 19892 6013 19956
rect 5947 19891 6013 19892
rect 4642 19552 4650 19616
rect 4714 19552 4730 19616
rect 4794 19552 4810 19616
rect 4874 19552 4890 19616
rect 4954 19552 4963 19616
rect 4475 18868 4541 18869
rect 4475 18804 4476 18868
rect 4540 18804 4541 18868
rect 4475 18803 4541 18804
rect 4291 18052 4357 18053
rect 4291 17988 4292 18052
rect 4356 17988 4357 18052
rect 4291 17987 4357 17988
rect 4294 13701 4354 17987
rect 4478 17101 4538 18803
rect 4642 18528 4963 19552
rect 5211 18596 5277 18597
rect 5211 18532 5212 18596
rect 5276 18532 5277 18596
rect 5211 18531 5277 18532
rect 4642 18464 4650 18528
rect 4714 18464 4730 18528
rect 4794 18464 4810 18528
rect 4874 18464 4890 18528
rect 4954 18464 4963 18528
rect 4642 17440 4963 18464
rect 4642 17376 4650 17440
rect 4714 17376 4730 17440
rect 4794 17376 4810 17440
rect 4874 17376 4890 17440
rect 4954 17376 4963 17440
rect 4475 17100 4541 17101
rect 4475 17036 4476 17100
rect 4540 17036 4541 17100
rect 4475 17035 4541 17036
rect 4642 16352 4963 17376
rect 4642 16288 4650 16352
rect 4714 16288 4730 16352
rect 4794 16288 4810 16352
rect 4874 16288 4890 16352
rect 4954 16288 4963 16352
rect 4642 15264 4963 16288
rect 4642 15200 4650 15264
rect 4714 15200 4730 15264
rect 4794 15200 4810 15264
rect 4874 15200 4890 15264
rect 4954 15200 4963 15264
rect 4475 14788 4541 14789
rect 4475 14724 4476 14788
rect 4540 14724 4541 14788
rect 4475 14723 4541 14724
rect 4291 13700 4357 13701
rect 4291 13636 4292 13700
rect 4356 13636 4357 13700
rect 4291 13635 4357 13636
rect 4478 13429 4538 14723
rect 4642 14176 4963 15200
rect 4642 14112 4650 14176
rect 4714 14112 4730 14176
rect 4794 14112 4810 14176
rect 4874 14112 4890 14176
rect 4954 14112 4963 14176
rect 4475 13428 4541 13429
rect 4475 13364 4476 13428
rect 4540 13364 4541 13428
rect 4475 13363 4541 13364
rect 4642 13088 4963 14112
rect 5214 13701 5274 18531
rect 5211 13700 5277 13701
rect 5211 13636 5212 13700
rect 5276 13636 5277 13700
rect 5211 13635 5277 13636
rect 4642 13024 4650 13088
rect 4714 13024 4730 13088
rect 4794 13024 4810 13088
rect 4874 13024 4890 13088
rect 4954 13024 4963 13088
rect 4642 12000 4963 13024
rect 5027 12748 5093 12749
rect 5027 12684 5028 12748
rect 5092 12684 5093 12748
rect 5027 12683 5093 12684
rect 4642 11936 4650 12000
rect 4714 11936 4730 12000
rect 4794 11936 4810 12000
rect 4874 11936 4890 12000
rect 4954 11936 4963 12000
rect 4642 10912 4963 11936
rect 4642 10848 4650 10912
rect 4714 10848 4730 10912
rect 4794 10848 4810 10912
rect 4874 10848 4890 10912
rect 4954 10848 4963 10912
rect 4642 9824 4963 10848
rect 4642 9760 4650 9824
rect 4714 9760 4730 9824
rect 4794 9760 4810 9824
rect 4874 9760 4890 9824
rect 4954 9760 4963 9824
rect 4642 8736 4963 9760
rect 4642 8672 4650 8736
rect 4714 8672 4730 8736
rect 4794 8672 4810 8736
rect 4874 8672 4890 8736
rect 4954 8672 4963 8736
rect 4642 7648 4963 8672
rect 5030 8533 5090 12683
rect 5027 8532 5093 8533
rect 5027 8468 5028 8532
rect 5092 8468 5093 8532
rect 5027 8467 5093 8468
rect 5950 8261 6010 19891
rect 7235 12748 7301 12749
rect 7235 12684 7236 12748
rect 7300 12684 7301 12748
rect 7235 12683 7301 12684
rect 6315 12340 6381 12341
rect 6315 12276 6316 12340
rect 6380 12276 6381 12340
rect 6315 12275 6381 12276
rect 6318 10709 6378 12275
rect 6315 10708 6381 10709
rect 6315 10644 6316 10708
rect 6380 10644 6381 10708
rect 6315 10643 6381 10644
rect 7051 8668 7117 8669
rect 7051 8604 7052 8668
rect 7116 8604 7117 8668
rect 7051 8603 7117 8604
rect 5947 8260 6013 8261
rect 5947 8196 5948 8260
rect 6012 8196 6013 8260
rect 5947 8195 6013 8196
rect 4642 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4890 7648
rect 4954 7584 4963 7648
rect 4642 6560 4963 7584
rect 7054 7309 7114 8603
rect 7238 7717 7298 12683
rect 7419 10164 7485 10165
rect 7419 10100 7420 10164
rect 7484 10100 7485 10164
rect 7419 10099 7485 10100
rect 7422 8669 7482 10099
rect 7419 8668 7485 8669
rect 7419 8604 7420 8668
rect 7484 8604 7485 8668
rect 7419 8603 7485 8604
rect 7235 7716 7301 7717
rect 7235 7652 7236 7716
rect 7300 7652 7301 7716
rect 7235 7651 7301 7652
rect 7051 7308 7117 7309
rect 7051 7244 7052 7308
rect 7116 7244 7117 7308
rect 7051 7243 7117 7244
rect 4642 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4890 6560
rect 4954 6496 4963 6560
rect 4642 5472 4963 6496
rect 4642 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4890 5472
rect 4954 5408 4963 5472
rect 4642 4384 4963 5408
rect 7606 5405 7666 20299
rect 8341 20160 8661 21184
rect 8341 20096 8349 20160
rect 8413 20096 8429 20160
rect 8493 20096 8509 20160
rect 8573 20096 8589 20160
rect 8653 20096 8661 20160
rect 8341 19072 8661 20096
rect 12040 21792 12360 21808
rect 12040 21728 12048 21792
rect 12112 21728 12128 21792
rect 12192 21728 12208 21792
rect 12272 21728 12288 21792
rect 12352 21728 12360 21792
rect 12040 20704 12360 21728
rect 15738 21248 16058 21808
rect 15738 21184 15746 21248
rect 15810 21184 15826 21248
rect 15890 21184 15906 21248
rect 15970 21184 15986 21248
rect 16050 21184 16058 21248
rect 14963 20772 15029 20773
rect 14963 20708 14964 20772
rect 15028 20708 15029 20772
rect 14963 20707 15029 20708
rect 12040 20640 12048 20704
rect 12112 20640 12128 20704
rect 12192 20640 12208 20704
rect 12272 20640 12288 20704
rect 12352 20640 12360 20704
rect 12040 19616 12360 20640
rect 12040 19552 12048 19616
rect 12112 19552 12128 19616
rect 12192 19552 12208 19616
rect 12272 19552 12288 19616
rect 12352 19552 12360 19616
rect 8891 19276 8957 19277
rect 8891 19212 8892 19276
rect 8956 19212 8957 19276
rect 8891 19211 8957 19212
rect 8341 19008 8349 19072
rect 8413 19008 8429 19072
rect 8493 19008 8509 19072
rect 8573 19008 8589 19072
rect 8653 19008 8661 19072
rect 8341 17984 8661 19008
rect 8341 17920 8349 17984
rect 8413 17920 8429 17984
rect 8493 17920 8509 17984
rect 8573 17920 8589 17984
rect 8653 17920 8661 17984
rect 8341 16896 8661 17920
rect 8341 16832 8349 16896
rect 8413 16832 8429 16896
rect 8493 16832 8509 16896
rect 8573 16832 8589 16896
rect 8653 16832 8661 16896
rect 8341 15808 8661 16832
rect 8341 15744 8349 15808
rect 8413 15744 8429 15808
rect 8493 15744 8509 15808
rect 8573 15744 8589 15808
rect 8653 15744 8661 15808
rect 7971 15604 8037 15605
rect 7971 15540 7972 15604
rect 8036 15540 8037 15604
rect 7971 15539 8037 15540
rect 7787 8940 7853 8941
rect 7787 8876 7788 8940
rect 7852 8876 7853 8940
rect 7787 8875 7853 8876
rect 7790 7581 7850 8875
rect 7974 8533 8034 15539
rect 8155 14924 8221 14925
rect 8155 14860 8156 14924
rect 8220 14860 8221 14924
rect 8155 14859 8221 14860
rect 7971 8532 8037 8533
rect 7971 8468 7972 8532
rect 8036 8468 8037 8532
rect 7971 8467 8037 8468
rect 7787 7580 7853 7581
rect 7787 7516 7788 7580
rect 7852 7516 7853 7580
rect 7787 7515 7853 7516
rect 8158 7445 8218 14859
rect 8341 14720 8661 15744
rect 8341 14656 8349 14720
rect 8413 14656 8429 14720
rect 8493 14656 8509 14720
rect 8573 14656 8589 14720
rect 8653 14656 8661 14720
rect 8341 13632 8661 14656
rect 8341 13568 8349 13632
rect 8413 13568 8429 13632
rect 8493 13568 8509 13632
rect 8573 13568 8589 13632
rect 8653 13568 8661 13632
rect 8341 12544 8661 13568
rect 8341 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8509 12544
rect 8573 12480 8589 12544
rect 8653 12480 8661 12544
rect 8341 11456 8661 12480
rect 8341 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8509 11456
rect 8573 11392 8589 11456
rect 8653 11392 8661 11456
rect 8341 10368 8661 11392
rect 8341 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8509 10368
rect 8573 10304 8589 10368
rect 8653 10304 8661 10368
rect 8341 9280 8661 10304
rect 8341 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8509 9280
rect 8573 9216 8589 9280
rect 8653 9216 8661 9280
rect 8341 8192 8661 9216
rect 8341 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8509 8192
rect 8573 8128 8589 8192
rect 8653 8128 8661 8192
rect 8155 7444 8221 7445
rect 8155 7380 8156 7444
rect 8220 7380 8221 7444
rect 8155 7379 8221 7380
rect 8341 7104 8661 8128
rect 8894 8125 8954 19211
rect 12040 18528 12360 19552
rect 12040 18464 12048 18528
rect 12112 18464 12128 18528
rect 12192 18464 12208 18528
rect 12272 18464 12288 18528
rect 12352 18464 12360 18528
rect 9627 18188 9693 18189
rect 9627 18124 9628 18188
rect 9692 18124 9693 18188
rect 9627 18123 9693 18124
rect 9630 16557 9690 18123
rect 9811 18052 9877 18053
rect 9811 17988 9812 18052
rect 9876 17988 9877 18052
rect 9811 17987 9877 17988
rect 9259 16556 9325 16557
rect 9259 16492 9260 16556
rect 9324 16492 9325 16556
rect 9259 16491 9325 16492
rect 9627 16556 9693 16557
rect 9627 16492 9628 16556
rect 9692 16492 9693 16556
rect 9627 16491 9693 16492
rect 9075 15332 9141 15333
rect 9075 15268 9076 15332
rect 9140 15268 9141 15332
rect 9075 15267 9141 15268
rect 8891 8124 8957 8125
rect 8891 8060 8892 8124
rect 8956 8060 8957 8124
rect 8891 8059 8957 8060
rect 9078 7445 9138 15267
rect 9262 12341 9322 16491
rect 9814 16285 9874 17987
rect 12040 17440 12360 18464
rect 12040 17376 12048 17440
rect 12112 17376 12128 17440
rect 12192 17376 12208 17440
rect 12272 17376 12288 17440
rect 12352 17376 12360 17440
rect 12040 16352 12360 17376
rect 12040 16288 12048 16352
rect 12112 16288 12128 16352
rect 12192 16288 12208 16352
rect 12272 16288 12288 16352
rect 12352 16288 12360 16352
rect 9811 16284 9877 16285
rect 9811 16220 9812 16284
rect 9876 16220 9877 16284
rect 9811 16219 9877 16220
rect 11099 16148 11165 16149
rect 11099 16084 11100 16148
rect 11164 16084 11165 16148
rect 11099 16083 11165 16084
rect 10179 15060 10245 15061
rect 10179 14996 10180 15060
rect 10244 14996 10245 15060
rect 10179 14995 10245 14996
rect 10182 12477 10242 14995
rect 10179 12476 10245 12477
rect 10179 12412 10180 12476
rect 10244 12412 10245 12476
rect 10179 12411 10245 12412
rect 11102 12341 11162 16083
rect 12040 15264 12360 16288
rect 13859 15332 13925 15333
rect 13859 15268 13860 15332
rect 13924 15268 13925 15332
rect 13859 15267 13925 15268
rect 12040 15200 12048 15264
rect 12112 15200 12128 15264
rect 12192 15200 12208 15264
rect 12272 15200 12288 15264
rect 12352 15200 12360 15264
rect 12040 14176 12360 15200
rect 13123 14244 13189 14245
rect 13123 14180 13124 14244
rect 13188 14180 13189 14244
rect 13123 14179 13189 14180
rect 12040 14112 12048 14176
rect 12112 14112 12128 14176
rect 12192 14112 12208 14176
rect 12272 14112 12288 14176
rect 12352 14112 12360 14176
rect 12040 13088 12360 14112
rect 12040 13024 12048 13088
rect 12112 13024 12128 13088
rect 12192 13024 12208 13088
rect 12272 13024 12288 13088
rect 12352 13024 12360 13088
rect 9259 12340 9325 12341
rect 9259 12276 9260 12340
rect 9324 12276 9325 12340
rect 9259 12275 9325 12276
rect 11099 12340 11165 12341
rect 11099 12276 11100 12340
rect 11164 12276 11165 12340
rect 11099 12275 11165 12276
rect 9259 12204 9325 12205
rect 9259 12140 9260 12204
rect 9324 12140 9325 12204
rect 9259 12139 9325 12140
rect 9262 9077 9322 12139
rect 12040 12000 12360 13024
rect 12939 12068 13005 12069
rect 12939 12004 12940 12068
rect 13004 12004 13005 12068
rect 12939 12003 13005 12004
rect 12040 11936 12048 12000
rect 12112 11936 12128 12000
rect 12192 11936 12208 12000
rect 12272 11936 12288 12000
rect 12352 11936 12360 12000
rect 12040 10912 12360 11936
rect 12040 10848 12048 10912
rect 12112 10848 12128 10912
rect 12192 10848 12208 10912
rect 12272 10848 12288 10912
rect 12352 10848 12360 10912
rect 12040 9824 12360 10848
rect 12040 9760 12048 9824
rect 12112 9760 12128 9824
rect 12192 9760 12208 9824
rect 12272 9760 12288 9824
rect 12352 9760 12360 9824
rect 9443 9620 9509 9621
rect 9443 9556 9444 9620
rect 9508 9556 9509 9620
rect 9443 9555 9509 9556
rect 9259 9076 9325 9077
rect 9259 9012 9260 9076
rect 9324 9012 9325 9076
rect 9259 9011 9325 9012
rect 9075 7444 9141 7445
rect 9075 7380 9076 7444
rect 9140 7380 9141 7444
rect 9075 7379 9141 7380
rect 8341 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8509 7104
rect 8573 7040 8589 7104
rect 8653 7040 8661 7104
rect 8341 6016 8661 7040
rect 8891 7036 8957 7037
rect 8891 6972 8892 7036
rect 8956 6972 8957 7036
rect 8891 6971 8957 6972
rect 8341 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8509 6016
rect 8573 5952 8589 6016
rect 8653 5952 8661 6016
rect 7603 5404 7669 5405
rect 7603 5340 7604 5404
rect 7668 5340 7669 5404
rect 7603 5339 7669 5340
rect 4642 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4890 4384
rect 4954 4320 4963 4384
rect 4642 3296 4963 4320
rect 4642 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4890 3296
rect 4954 3232 4963 3296
rect 4642 2208 4963 3232
rect 4642 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4890 2208
rect 4954 2144 4963 2208
rect 4642 2128 4963 2144
rect 8341 4928 8661 5952
rect 8341 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8509 4928
rect 8573 4864 8589 4928
rect 8653 4864 8661 4928
rect 8341 3840 8661 4864
rect 8341 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8509 3840
rect 8573 3776 8589 3840
rect 8653 3776 8661 3840
rect 8341 2752 8661 3776
rect 8341 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8509 2752
rect 8573 2688 8589 2752
rect 8653 2688 8661 2752
rect 8341 2128 8661 2688
rect 8894 2413 8954 6971
rect 9446 5949 9506 9555
rect 10915 9484 10981 9485
rect 10915 9420 10916 9484
rect 10980 9420 10981 9484
rect 10915 9419 10981 9420
rect 11835 9484 11901 9485
rect 11835 9420 11836 9484
rect 11900 9420 11901 9484
rect 11835 9419 11901 9420
rect 10179 9348 10245 9349
rect 10179 9284 10180 9348
rect 10244 9284 10245 9348
rect 10179 9283 10245 9284
rect 10363 9348 10429 9349
rect 10363 9284 10364 9348
rect 10428 9284 10429 9348
rect 10363 9283 10429 9284
rect 9811 8804 9877 8805
rect 9811 8740 9812 8804
rect 9876 8740 9877 8804
rect 9811 8739 9877 8740
rect 9814 7173 9874 8739
rect 10182 8397 10242 9283
rect 10179 8396 10245 8397
rect 10179 8332 10180 8396
rect 10244 8332 10245 8396
rect 10179 8331 10245 8332
rect 9811 7172 9877 7173
rect 9811 7108 9812 7172
rect 9876 7108 9877 7172
rect 9811 7107 9877 7108
rect 9443 5948 9509 5949
rect 9443 5884 9444 5948
rect 9508 5884 9509 5948
rect 9443 5883 9509 5884
rect 10366 4861 10426 9283
rect 10918 7717 10978 9419
rect 10915 7716 10981 7717
rect 10915 7652 10916 7716
rect 10980 7652 10981 7716
rect 10915 7651 10981 7652
rect 11838 5813 11898 9419
rect 12040 8736 12360 9760
rect 12040 8672 12048 8736
rect 12112 8672 12128 8736
rect 12192 8672 12208 8736
rect 12272 8672 12288 8736
rect 12352 8672 12360 8736
rect 12040 7648 12360 8672
rect 12040 7584 12048 7648
rect 12112 7584 12128 7648
rect 12192 7584 12208 7648
rect 12272 7584 12288 7648
rect 12352 7584 12360 7648
rect 12040 6560 12360 7584
rect 12040 6496 12048 6560
rect 12112 6496 12128 6560
rect 12192 6496 12208 6560
rect 12272 6496 12288 6560
rect 12352 6496 12360 6560
rect 11835 5812 11901 5813
rect 11835 5748 11836 5812
rect 11900 5748 11901 5812
rect 11835 5747 11901 5748
rect 12040 5472 12360 6496
rect 12942 5541 13002 12003
rect 13126 8533 13186 14179
rect 13123 8532 13189 8533
rect 13123 8468 13124 8532
rect 13188 8468 13189 8532
rect 13123 8467 13189 8468
rect 13862 8261 13922 15267
rect 14779 15060 14845 15061
rect 14779 14996 14780 15060
rect 14844 14996 14845 15060
rect 14779 14995 14845 14996
rect 14782 11117 14842 14995
rect 14779 11116 14845 11117
rect 14779 11052 14780 11116
rect 14844 11052 14845 11116
rect 14779 11051 14845 11052
rect 14966 9757 15026 20707
rect 15738 20160 16058 21184
rect 19437 21792 19757 21808
rect 19437 21728 19445 21792
rect 19509 21728 19525 21792
rect 19589 21728 19605 21792
rect 19669 21728 19685 21792
rect 19749 21728 19757 21792
rect 16987 20772 17053 20773
rect 16987 20708 16988 20772
rect 17052 20708 17053 20772
rect 16987 20707 17053 20708
rect 15738 20096 15746 20160
rect 15810 20096 15826 20160
rect 15890 20096 15906 20160
rect 15970 20096 15986 20160
rect 16050 20096 16058 20160
rect 15738 19072 16058 20096
rect 15738 19008 15746 19072
rect 15810 19008 15826 19072
rect 15890 19008 15906 19072
rect 15970 19008 15986 19072
rect 16050 19008 16058 19072
rect 15738 17984 16058 19008
rect 15738 17920 15746 17984
rect 15810 17920 15826 17984
rect 15890 17920 15906 17984
rect 15970 17920 15986 17984
rect 16050 17920 16058 17984
rect 15738 16896 16058 17920
rect 15738 16832 15746 16896
rect 15810 16832 15826 16896
rect 15890 16832 15906 16896
rect 15970 16832 15986 16896
rect 16050 16832 16058 16896
rect 15738 15808 16058 16832
rect 15738 15744 15746 15808
rect 15810 15744 15826 15808
rect 15890 15744 15906 15808
rect 15970 15744 15986 15808
rect 16050 15744 16058 15808
rect 15515 15468 15581 15469
rect 15515 15404 15516 15468
rect 15580 15404 15581 15468
rect 15515 15403 15581 15404
rect 15331 13836 15397 13837
rect 15331 13772 15332 13836
rect 15396 13772 15397 13836
rect 15331 13771 15397 13772
rect 15147 11252 15213 11253
rect 15147 11188 15148 11252
rect 15212 11188 15213 11252
rect 15147 11187 15213 11188
rect 14963 9756 15029 9757
rect 14963 9692 14964 9756
rect 15028 9692 15029 9756
rect 14963 9691 15029 9692
rect 13859 8260 13925 8261
rect 13859 8196 13860 8260
rect 13924 8196 13925 8260
rect 13859 8195 13925 8196
rect 13675 7308 13741 7309
rect 13675 7244 13676 7308
rect 13740 7244 13741 7308
rect 13675 7243 13741 7244
rect 13123 6628 13189 6629
rect 13123 6564 13124 6628
rect 13188 6564 13189 6628
rect 13123 6563 13189 6564
rect 13126 6221 13186 6563
rect 13123 6220 13189 6221
rect 13123 6156 13124 6220
rect 13188 6156 13189 6220
rect 13123 6155 13189 6156
rect 13678 5541 13738 7243
rect 15150 5949 15210 11187
rect 15147 5948 15213 5949
rect 15147 5884 15148 5948
rect 15212 5884 15213 5948
rect 15147 5883 15213 5884
rect 12939 5540 13005 5541
rect 12939 5476 12940 5540
rect 13004 5476 13005 5540
rect 12939 5475 13005 5476
rect 13675 5540 13741 5541
rect 13675 5476 13676 5540
rect 13740 5476 13741 5540
rect 13675 5475 13741 5476
rect 12040 5408 12048 5472
rect 12112 5408 12128 5472
rect 12192 5408 12208 5472
rect 12272 5408 12288 5472
rect 12352 5408 12360 5472
rect 10363 4860 10429 4861
rect 10363 4796 10364 4860
rect 10428 4796 10429 4860
rect 10363 4795 10429 4796
rect 12040 4384 12360 5408
rect 12040 4320 12048 4384
rect 12112 4320 12128 4384
rect 12192 4320 12208 4384
rect 12272 4320 12288 4384
rect 12352 4320 12360 4384
rect 12040 3296 12360 4320
rect 12040 3232 12048 3296
rect 12112 3232 12128 3296
rect 12192 3232 12208 3296
rect 12272 3232 12288 3296
rect 12352 3232 12360 3296
rect 8891 2412 8957 2413
rect 8891 2348 8892 2412
rect 8956 2348 8957 2412
rect 8891 2347 8957 2348
rect 12040 2208 12360 3232
rect 15334 2685 15394 13771
rect 15518 3093 15578 15403
rect 15738 14720 16058 15744
rect 15738 14656 15746 14720
rect 15810 14656 15826 14720
rect 15890 14656 15906 14720
rect 15970 14656 15986 14720
rect 16050 14656 16058 14720
rect 15738 13632 16058 14656
rect 15738 13568 15746 13632
rect 15810 13568 15826 13632
rect 15890 13568 15906 13632
rect 15970 13568 15986 13632
rect 16050 13568 16058 13632
rect 15738 12544 16058 13568
rect 15738 12480 15746 12544
rect 15810 12480 15826 12544
rect 15890 12480 15906 12544
rect 15970 12480 15986 12544
rect 16050 12480 16058 12544
rect 15738 11456 16058 12480
rect 16803 11660 16869 11661
rect 16803 11596 16804 11660
rect 16868 11596 16869 11660
rect 16803 11595 16869 11596
rect 15738 11392 15746 11456
rect 15810 11392 15826 11456
rect 15890 11392 15906 11456
rect 15970 11392 15986 11456
rect 16050 11392 16058 11456
rect 15738 10368 16058 11392
rect 15738 10304 15746 10368
rect 15810 10304 15826 10368
rect 15890 10304 15906 10368
rect 15970 10304 15986 10368
rect 16050 10304 16058 10368
rect 15738 9280 16058 10304
rect 15738 9216 15746 9280
rect 15810 9216 15826 9280
rect 15890 9216 15906 9280
rect 15970 9216 15986 9280
rect 16050 9216 16058 9280
rect 15738 8192 16058 9216
rect 15738 8128 15746 8192
rect 15810 8128 15826 8192
rect 15890 8128 15906 8192
rect 15970 8128 15986 8192
rect 16050 8128 16058 8192
rect 15738 7104 16058 8128
rect 15738 7040 15746 7104
rect 15810 7040 15826 7104
rect 15890 7040 15906 7104
rect 15970 7040 15986 7104
rect 16050 7040 16058 7104
rect 15738 6016 16058 7040
rect 15738 5952 15746 6016
rect 15810 5952 15826 6016
rect 15890 5952 15906 6016
rect 15970 5952 15986 6016
rect 16050 5952 16058 6016
rect 15738 4928 16058 5952
rect 16806 5269 16866 11595
rect 16803 5268 16869 5269
rect 16803 5204 16804 5268
rect 16868 5204 16869 5268
rect 16803 5203 16869 5204
rect 15738 4864 15746 4928
rect 15810 4864 15826 4928
rect 15890 4864 15906 4928
rect 15970 4864 15986 4928
rect 16050 4864 16058 4928
rect 15738 3840 16058 4864
rect 16619 4452 16685 4453
rect 16619 4388 16620 4452
rect 16684 4388 16685 4452
rect 16619 4387 16685 4388
rect 15738 3776 15746 3840
rect 15810 3776 15826 3840
rect 15890 3776 15906 3840
rect 15970 3776 15986 3840
rect 16050 3776 16058 3840
rect 15515 3092 15581 3093
rect 15515 3028 15516 3092
rect 15580 3028 15581 3092
rect 15515 3027 15581 3028
rect 15738 2752 16058 3776
rect 15738 2688 15746 2752
rect 15810 2688 15826 2752
rect 15890 2688 15906 2752
rect 15970 2688 15986 2752
rect 16050 2688 16058 2752
rect 15331 2684 15397 2685
rect 15331 2620 15332 2684
rect 15396 2620 15397 2684
rect 15331 2619 15397 2620
rect 12040 2144 12048 2208
rect 12112 2144 12128 2208
rect 12192 2144 12208 2208
rect 12272 2144 12288 2208
rect 12352 2144 12360 2208
rect 12040 2128 12360 2144
rect 15738 2128 16058 2688
rect 16622 2413 16682 4387
rect 16990 3229 17050 20707
rect 19437 20704 19757 21728
rect 20483 20772 20549 20773
rect 20483 20708 20484 20772
rect 20548 20708 20549 20772
rect 20483 20707 20549 20708
rect 19437 20640 19445 20704
rect 19509 20640 19525 20704
rect 19589 20640 19605 20704
rect 19669 20640 19685 20704
rect 19749 20640 19757 20704
rect 19437 19616 19757 20640
rect 20115 19820 20181 19821
rect 20115 19756 20116 19820
rect 20180 19756 20181 19820
rect 20115 19755 20181 19756
rect 19437 19552 19445 19616
rect 19509 19552 19525 19616
rect 19589 19552 19605 19616
rect 19669 19552 19685 19616
rect 19749 19552 19757 19616
rect 19437 18528 19757 19552
rect 19931 19412 19997 19413
rect 19931 19348 19932 19412
rect 19996 19348 19997 19412
rect 19931 19347 19997 19348
rect 19437 18464 19445 18528
rect 19509 18464 19525 18528
rect 19589 18464 19605 18528
rect 19669 18464 19685 18528
rect 19749 18464 19757 18528
rect 17723 18324 17789 18325
rect 17723 18260 17724 18324
rect 17788 18260 17789 18324
rect 17723 18259 17789 18260
rect 17539 12748 17605 12749
rect 17539 12684 17540 12748
rect 17604 12684 17605 12748
rect 17539 12683 17605 12684
rect 17542 7581 17602 12683
rect 17726 10437 17786 18259
rect 19437 17440 19757 18464
rect 19437 17376 19445 17440
rect 19509 17376 19525 17440
rect 19589 17376 19605 17440
rect 19669 17376 19685 17440
rect 19749 17376 19757 17440
rect 19437 16352 19757 17376
rect 19437 16288 19445 16352
rect 19509 16288 19525 16352
rect 19589 16288 19605 16352
rect 19669 16288 19685 16352
rect 19749 16288 19757 16352
rect 19437 15264 19757 16288
rect 19437 15200 19445 15264
rect 19509 15200 19525 15264
rect 19589 15200 19605 15264
rect 19669 15200 19685 15264
rect 19749 15200 19757 15264
rect 19437 14176 19757 15200
rect 19437 14112 19445 14176
rect 19509 14112 19525 14176
rect 19589 14112 19605 14176
rect 19669 14112 19685 14176
rect 19749 14112 19757 14176
rect 17907 13428 17973 13429
rect 17907 13364 17908 13428
rect 17972 13364 17973 13428
rect 17907 13363 17973 13364
rect 17910 12341 17970 13363
rect 19437 13088 19757 14112
rect 19437 13024 19445 13088
rect 19509 13024 19525 13088
rect 19589 13024 19605 13088
rect 19669 13024 19685 13088
rect 19749 13024 19757 13088
rect 18459 12476 18525 12477
rect 18459 12412 18460 12476
rect 18524 12412 18525 12476
rect 18459 12411 18525 12412
rect 19195 12476 19261 12477
rect 19195 12412 19196 12476
rect 19260 12412 19261 12476
rect 19195 12411 19261 12412
rect 17907 12340 17973 12341
rect 17907 12276 17908 12340
rect 17972 12276 17973 12340
rect 17907 12275 17973 12276
rect 18275 11252 18341 11253
rect 18275 11188 18276 11252
rect 18340 11188 18341 11252
rect 18275 11187 18341 11188
rect 17723 10436 17789 10437
rect 17723 10372 17724 10436
rect 17788 10372 17789 10436
rect 17723 10371 17789 10372
rect 18091 9620 18157 9621
rect 18091 9556 18092 9620
rect 18156 9556 18157 9620
rect 18091 9555 18157 9556
rect 18094 8125 18154 9555
rect 18278 8941 18338 11187
rect 18275 8940 18341 8941
rect 18275 8876 18276 8940
rect 18340 8876 18341 8940
rect 18275 8875 18341 8876
rect 18091 8124 18157 8125
rect 18091 8060 18092 8124
rect 18156 8060 18157 8124
rect 18091 8059 18157 8060
rect 17539 7580 17605 7581
rect 17539 7516 17540 7580
rect 17604 7516 17605 7580
rect 17539 7515 17605 7516
rect 18462 7445 18522 12411
rect 19011 11796 19077 11797
rect 19011 11732 19012 11796
rect 19076 11732 19077 11796
rect 19011 11731 19077 11732
rect 18827 9620 18893 9621
rect 18827 9556 18828 9620
rect 18892 9556 18893 9620
rect 18827 9555 18893 9556
rect 18459 7444 18525 7445
rect 18459 7380 18460 7444
rect 18524 7380 18525 7444
rect 18459 7379 18525 7380
rect 18830 3637 18890 9555
rect 19014 4725 19074 11731
rect 19198 6629 19258 12411
rect 19437 12000 19757 13024
rect 19437 11936 19445 12000
rect 19509 11936 19525 12000
rect 19589 11936 19605 12000
rect 19669 11936 19685 12000
rect 19749 11936 19757 12000
rect 19437 10912 19757 11936
rect 19437 10848 19445 10912
rect 19509 10848 19525 10912
rect 19589 10848 19605 10912
rect 19669 10848 19685 10912
rect 19749 10848 19757 10912
rect 19437 9824 19757 10848
rect 19437 9760 19445 9824
rect 19509 9760 19525 9824
rect 19589 9760 19605 9824
rect 19669 9760 19685 9824
rect 19749 9760 19757 9824
rect 19437 8736 19757 9760
rect 19437 8672 19445 8736
rect 19509 8672 19525 8736
rect 19589 8672 19605 8736
rect 19669 8672 19685 8736
rect 19749 8672 19757 8736
rect 19437 7648 19757 8672
rect 19437 7584 19445 7648
rect 19509 7584 19525 7648
rect 19589 7584 19605 7648
rect 19669 7584 19685 7648
rect 19749 7584 19757 7648
rect 19195 6628 19261 6629
rect 19195 6564 19196 6628
rect 19260 6564 19261 6628
rect 19195 6563 19261 6564
rect 19437 6560 19757 7584
rect 19437 6496 19445 6560
rect 19509 6496 19525 6560
rect 19589 6496 19605 6560
rect 19669 6496 19685 6560
rect 19749 6496 19757 6560
rect 19437 5472 19757 6496
rect 19437 5408 19445 5472
rect 19509 5408 19525 5472
rect 19589 5408 19605 5472
rect 19669 5408 19685 5472
rect 19749 5408 19757 5472
rect 19011 4724 19077 4725
rect 19011 4660 19012 4724
rect 19076 4660 19077 4724
rect 19011 4659 19077 4660
rect 19437 4384 19757 5408
rect 19437 4320 19445 4384
rect 19509 4320 19525 4384
rect 19589 4320 19605 4384
rect 19669 4320 19685 4384
rect 19749 4320 19757 4384
rect 18827 3636 18893 3637
rect 18827 3572 18828 3636
rect 18892 3572 18893 3636
rect 18827 3571 18893 3572
rect 19437 3296 19757 4320
rect 19934 3501 19994 19347
rect 19931 3500 19997 3501
rect 19931 3436 19932 3500
rect 19996 3436 19997 3500
rect 19931 3435 19997 3436
rect 19931 3364 19997 3365
rect 19931 3300 19932 3364
rect 19996 3300 19997 3364
rect 19931 3299 19997 3300
rect 19437 3232 19445 3296
rect 19509 3232 19525 3296
rect 19589 3232 19605 3296
rect 19669 3232 19685 3296
rect 19749 3232 19757 3296
rect 16987 3228 17053 3229
rect 16987 3164 16988 3228
rect 17052 3164 17053 3228
rect 16987 3163 17053 3164
rect 16619 2412 16685 2413
rect 16619 2348 16620 2412
rect 16684 2348 16685 2412
rect 16619 2347 16685 2348
rect 19437 2208 19757 3232
rect 19934 2957 19994 3299
rect 19931 2956 19997 2957
rect 19931 2892 19932 2956
rect 19996 2892 19997 2956
rect 19931 2891 19997 2892
rect 20118 2821 20178 19755
rect 20299 18052 20365 18053
rect 20299 17988 20300 18052
rect 20364 17988 20365 18052
rect 20299 17987 20365 17988
rect 20302 7445 20362 17987
rect 20299 7444 20365 7445
rect 20299 7380 20300 7444
rect 20364 7380 20365 7444
rect 20299 7379 20365 7380
rect 20486 3365 20546 20707
rect 20667 18324 20733 18325
rect 20667 18260 20668 18324
rect 20732 18260 20733 18324
rect 20667 18259 20733 18260
rect 20670 12205 20730 18259
rect 20667 12204 20733 12205
rect 20667 12140 20668 12204
rect 20732 12140 20733 12204
rect 20667 12139 20733 12140
rect 20667 9076 20733 9077
rect 20667 9012 20668 9076
rect 20732 9012 20733 9076
rect 20667 9011 20733 9012
rect 20670 4589 20730 9011
rect 20851 8124 20917 8125
rect 20851 8060 20852 8124
rect 20916 8060 20917 8124
rect 20851 8059 20917 8060
rect 20667 4588 20733 4589
rect 20667 4524 20668 4588
rect 20732 4524 20733 4588
rect 20667 4523 20733 4524
rect 20854 3773 20914 8059
rect 20851 3772 20917 3773
rect 20851 3708 20852 3772
rect 20916 3708 20917 3772
rect 20851 3707 20917 3708
rect 20483 3364 20549 3365
rect 20483 3300 20484 3364
rect 20548 3300 20549 3364
rect 20483 3299 20549 3300
rect 20115 2820 20181 2821
rect 20115 2756 20116 2820
rect 20180 2756 20181 2820
rect 20115 2755 20181 2756
rect 19437 2144 19445 2208
rect 19509 2144 19525 2208
rect 19589 2144 19605 2208
rect 19669 2144 19685 2208
rect 19749 2144 19757 2208
rect 19437 2128 19757 2144
use sky130_fd_sc_hd__buf_2  _68_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1748 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_19
timestamp 1606821651
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _64_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4876 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_31 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1606821651
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1606821651
transform 1 0 5152 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1606821651
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606821651
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606821651
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606821651
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606821651
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606821651
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606821651
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606821651
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606821651
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_123
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_131
timestamp 1606821651
transform 1 0 13156 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14260 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 14352 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13248 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 13340 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1606821651
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_141
timestamp 1606821651
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_152
timestamp 1606821651
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_163
timestamp 1606821651
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1606821651
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606821651
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 15272 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1606821651
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 16192 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 16284 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 17204 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 18216 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606821651
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606821651
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 20700 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 20056 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1606821651
transform 1 0 19964 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_203
timestamp 1606821651
transform 1 0 19780 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606821651
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_202
timestamp 1606821651
transform 1 0 19688 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_211
timestamp 1606821651
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606821651
transform 1 0 22356 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 23276 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 23276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1606821651
transform 1 0 22632 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_229
timestamp 1606821651
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_235
timestamp 1606821651
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606821651
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606821651
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606821651
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606821651
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1606821651
transform 1 0 10764 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 12144 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1606821651
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1606821651
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1606821651
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1606821651
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606821651
transform 1 0 15548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 17112 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16100 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_161
timestamp 1606821651
transform 1 0 15916 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_172
timestamp 1606821651
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 18952 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_190
timestamp 1606821651
transform 1 0 18584 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1606821651
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1606821651
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 21344 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 23276 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_236
timestamp 1606821651
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606821651
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606821651
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606821651
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606821651
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606821651
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 10304 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1606821651
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1606821651
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12604 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1606821651
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 14628 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13616 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 1606821651
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 16284 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1606821651
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1606821651
transform 1 0 19044 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606821651
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1606821651
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 19504 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_198
timestamp 1606821651
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_216
timestamp 1606821651
transform 1 0 20976 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 21344 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1606821651
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606821651
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606821651
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606821651
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606821651
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606821651
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_104
timestamp 1606821651
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 11868 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_115
timestamp 1606821651
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1606821651
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 13892 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1606821651
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1606821651
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606821651
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 15732 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_157
timestamp 1606821651
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 18768 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 17756 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_175
timestamp 1606821651
transform 1 0 17204 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1606821651
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 19780 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 21068 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1606821651
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606821651
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 23276 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1606821651
transform 1 0 22540 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_237
timestamp 1606821651
transform 1 0 22908 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606821651
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606821651
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7452 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_68
timestamp 1606821651
transform 1 0 7360 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1606821651
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_89
timestamp 1606821651
transform 1 0 9292 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1606821651
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1606821651
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1606821651
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 13432 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1606821651
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_150
timestamp 1606821651
transform 1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16836 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15180 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1606821651
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 19044 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_180
timestamp 1606821651
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1606821651
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 20608 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 21160 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1606821651
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1606821651
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1606821651
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 23276 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_234
timestamp 1606821651
transform 1 0 22632 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606821651
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606821651
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606821651
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1606821651
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5888 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5612 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_44
timestamp 1606821651
transform 1 0 5152 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_61
timestamp 1606821651
transform 1 0 6716 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_47
timestamp 1606821651
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1606821651
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 7636 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8648 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_69
timestamp 1606821651
transform 1 0 7452 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1606821651
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_70
timestamp 1606821651
transform 1 0 7544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_80
timestamp 1606821651
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1606821651
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606821651
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9660 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 10028 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1606821651
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1606821651
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 10580 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 10672 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 12236 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 12696 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_119
timestamp 1606821651
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606821651
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14352 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 13892 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1606821651
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1606821651
transform 1 0 14720 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1606821651
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17112 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16008 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16100 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1606821651
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1606821651
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1606821651
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 18216 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18768 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18768 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1606821651
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1606821651
transform 1 0 17480 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_190
timestamp 1606821651
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 20700 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1606821651
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606821651
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1606821651
transform 1 0 20240 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_212
timestamp 1606821651
transform 1 0 20608 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_218
timestamp 1606821651
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 21436 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 22448 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 21344 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 23276 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_230
timestamp 1606821651
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_236
timestamp 1606821651
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1606821651
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606821651
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4508 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1606821651
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5520 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 6532 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1606821651
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 1606821651
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1606821651
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1606821651
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 9844 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606821651
transform 1 0 10396 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606821651
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_99
timestamp 1606821651
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1606821651
transform 1 0 12052 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1606821651
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_122
timestamp 1606821651
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 13524 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1606821651
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606821651
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15640 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1606821651
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1606821651
transform 1 0 17296 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17756 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1606821651
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19412 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1606821651
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_208
timestamp 1606821651
transform 1 0 20240 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1606821651
transform 1 0 22540 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 23276 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1606821651
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_236
timestamp 1606821651
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606821651
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1606821651
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1606821651
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1606821651
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606821651
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1606821651
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7452 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1606821651
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 10120 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1606821651
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 11776 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1606821651
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606821651
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 13432 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1606821651
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 15824 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_9_156
timestamp 1606821651
transform 1 0 15456 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 18400 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606821651
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 20516 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1606821651
transform 1 0 20332 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1606821651
transform 1 0 22172 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 23276 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_227
timestamp 1606821651
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_235
timestamp 1606821651
transform 1 0 22724 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1606821651
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  Test_en_FTB00
timestamp 1606821651
transform 1 0 4508 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1606821651
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1606821651
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606821651
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6532 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606821651
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_49
timestamp 1606821651
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_55
timestamp 1606821651
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1606821651
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1606821651
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606821651
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1606821651
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 12972 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1606821651
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1606821651
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606821651
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 15364 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15916 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_159
timestamp 1606821651
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1606821651
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17940 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1606821651
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19596 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01
timestamp 1606821651
transform 1 0 20976 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_199
timestamp 1606821651
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1606821651
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_215
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 21712 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 23276 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_222
timestamp 1606821651
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_233
timestamp 1606821651
transform 1 0 22540 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_237
timestamp 1606821651
transform 1 0 22908 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2852 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1606821651
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_28
timestamp 1606821651
transform 1 0 3680 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_36
timestamp 1606821651
transform 1 0 4416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 7084 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1606821651
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7636 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1606821651
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1606821651
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9660 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1606821651
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1606821651
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1606821651
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 14996 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 13340 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1606821651
transform 1 0 14812 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15548 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1606821651
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1606821651
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 19136 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1606821651
transform 1 0 17204 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1606821651
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1606821651
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 20792 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1606821651
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 22448 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 23276 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_230
timestamp 1606821651
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1606821651
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2852 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1606821651
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1606821651
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1606821651
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1606821651
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1606821651
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1606821651
transform 1 0 5888 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1606821651
transform 1 0 6256 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7544 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1606821651
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1606821651
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10672 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 12236 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_113
timestamp 1606821651
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_119
timestamp 1606821651
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1606821651
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606821651
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16468 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15456 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1606821651
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 18308 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_12_183
timestamp 1606821651
transform 1 0 17940 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 20424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_208
timestamp 1606821651
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1606821651
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 21252 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 23276 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_235
timestamp 1606821651
transform 1 0 22724 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1606821651
transform 1 0 1564 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2024 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 3036 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1606821651
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_8
timestamp 1606821651
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 4140 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_37
timestamp 1606821651
transform 1 0 4508 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_43
timestamp 1606821651
transform 1 0 5060 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1606821651
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1606821651
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606821651
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 5796 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1606821651
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606821651
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1606821651
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 7728 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_13_66
timestamp 1606821651
transform 1 0 7176 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1606821651
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_67
timestamp 1606821651
transform 1 0 7268 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_73
timestamp 1606821651
transform 1 0 7820 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 10396 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1606821651
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606821651
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1606821651
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_114
timestamp 1606821651
transform 1 0 11592 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_117
timestamp 1606821651
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 11316 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 11684 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1606821651
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 12696 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 12696 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606821651
transform 1 0 14628 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.clb_clk
timestamp 1606821651
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1606821651
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1606821651
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1606821651
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1606821651
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15456 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_170
timestamp 1606821651
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_172
timestamp 1606821651
transform 1 0 16928 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 19136 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18216 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 17204 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18124 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606821651
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_194
timestamp 1606821651
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_184
timestamp 1606821651
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 19872 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 20424 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_217
timestamp 1606821651
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_202
timestamp 1606821651
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_208
timestamp 1606821651
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1606821651
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 21252 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 21344 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 21804 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 23276 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1606821651
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_223
timestamp 1606821651
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_234
timestamp 1606821651
transform 1 0 22632 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 1656 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 3312 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606821651
transform 1 0 4968 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_22
timestamp 1606821651
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1606821651
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1606821651
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 7452 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 9108 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_66
timestamp 1606821651
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1606821651
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 9936 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 9384 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1606821651
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 12604 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_112
timestamp 1606821651
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606821651
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606821651
transform 1 0 14260 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1606821651
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15916 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1606821651
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18216 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 17572 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1606821651
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1606821651
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1606821651
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1606821651
transform 1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 19504 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1606821651
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1606821651
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 22356 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 21344 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_229
timestamp 1606821651
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_235
timestamp 1606821651
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 1472 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_20
timestamp 1606821651
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606821651
transform 1 0 3404 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 3128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1606821651
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1606821651
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1606821651
transform 1 0 6808 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 5152 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1606821651
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1606821651
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 7268 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_83
timestamp 1606821651
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 9936 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 10488 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_100
timestamp 1606821651
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 12236 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 12788 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_118
timestamp 1606821651
transform 1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1606821651
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_143
timestamp 1606821651
transform 1 0 14260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1606821651
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 15640 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1606821651
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 17296 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 17940 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_16_180
timestamp 1606821651
transform 1 0 17664 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_204
timestamp 1606821651
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1606821651
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 23276 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_235
timestamp 1606821651
transform 1 0 22724 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 1472 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1606821651
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 3128 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 4140 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 5060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1606821651
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_37
timestamp 1606821651
transform 1 0 4508 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606821651
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 8832 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606821651
transform 1 0 7176 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1606821651
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 9384 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 10396 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1606821651
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1606821651
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.clb_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 12604 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1606821651
transform 1 0 11868 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 14444 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15916 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 15272 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_158
timestamp 1606821651
transform 1 0 15640 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1606821651
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 19044 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606821651
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1606821651
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1606821651
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 21344 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1606821651
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 1564 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_21
timestamp 1606821651
transform 1 0 3036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 5060 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606821651
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1606821651
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 5336 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 6992 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_55
timestamp 1606821651
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_61
timestamp 1606821651
transform 1 0 6716 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1606821651
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1606821651
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 9844 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.clb_clk
timestamp 1606821651
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606821651
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1606821651
transform 1 0 10212 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_106
timestamp 1606821651
transform 1 0 10856 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 11408 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1606821651
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1606821651
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 16008 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 15456 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1606821651
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_171
timestamp 1606821651
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 18952 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17480 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_176
timestamp 1606821651
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19504 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1606821651
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1606821651
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1606821651
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1606821651
transform 1 0 22540 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 23276 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1606821651
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_236
timestamp 1606821651
transform 1 0 22816 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1606821651
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_8
timestamp 1606821651
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 1656 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 1472 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_21
timestamp 1606821651
transform 1 0 3036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 2024 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 3680 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 4508 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1606821651
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606821651
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_35
timestamp 1606821651
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 5336 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 6164 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6716 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_44
timestamp 1606821651
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_55
timestamp 1606821651
transform 1 0 6164 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_53
timestamp 1606821651
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_59
timestamp 1606821651
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8464 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 8372 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1606821651
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1606821651
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 10396 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 10672 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1606821651
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1606821651
transform 1 0 10304 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1606821651
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1606821651
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12144 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 12604 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1606821651
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 13616 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_19_141
timestamp 1606821651
transform 1 0 14076 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1606821651
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606821651
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 15180 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 16744 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1606821651
transform 1 0 16652 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18216 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18676 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606821651
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1606821651
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19688 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1606821651
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_213
timestamp 1606821651
transform 1 0 20700 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1606821651
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 20332 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_218
timestamp 1606821651
transform 1 0 21160 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_217
timestamp 1606821651
transform 1 0 21068 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 21160 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606821651
transform 1 0 22172 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 21344 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 23276 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_227
timestamp 1606821651
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1606821651
transform 1 0 22540 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_237
timestamp 1606821651
transform 1 0 22908 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_236
timestamp 1606821651
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1472 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1606821651
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606821651
transform 1 0 4232 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_31
timestamp 1606821651
transform 1 0 3956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1606821651
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1606821651
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1606821651
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8280 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1606821651
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_76
timestamp 1606821651
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1606821651
transform 1 0 10396 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 10672 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 9936 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_94
timestamp 1606821651
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_100
timestamp 1606821651
transform 1 0 10304 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606821651
transform 1 0 11684 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 12788 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1606821651
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1606821651
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_143
timestamp 1606821651
transform 1 0 14260 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_151
timestamp 1606821651
transform 1 0 14996 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1606821651
transform 1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1606821651
transform 1 0 15272 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 16284 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606821651
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_157
timestamp 1606821651
transform 1 0 15548 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606821651
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 19688 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1606821651
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 21804 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_223
timestamp 1606821651
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_234
timestamp 1606821651
transform 1 0 22632 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1656 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5060 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_22
timestamp 1606821651
transform 1 0 3128 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1606821651
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1606821651
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6624 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 6072 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1606821651
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1606821651
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 8280 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1606821651
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1606821651
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9844 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 11500 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 12420 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 1606821651
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1606821651
transform 1 0 12328 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13892 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1606821651
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 16100 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17756 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19412 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 21160 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 20424 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1606821651
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1606821651
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1606821651
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_215
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 23276 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1606821651
transform 1 0 22632 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1840 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_6
timestamp 1606821651
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 4140 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_24
timestamp 1606821651
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_31
timestamp 1606821651
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1606821651
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1606821651
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606821651
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1606821651
transform 1 0 8464 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8924 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1606821651
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_83
timestamp 1606821651
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10672 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_101
timestamp 1606821651
transform 1 0 10396 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606821651
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13432 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 14996 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1606821651
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_150
timestamp 1606821651
transform 1 0 14904 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1606821651
transform 1 0 16468 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 15272 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1606821651
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_170
timestamp 1606821651
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  clk_0_FTB00
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1606821651
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1606821651
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 19320 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 21436 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_219
timestamp 1606821651
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_230
timestamp 1606821651
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1606821651
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1472 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_20
timestamp 1606821651
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1606821651
transform 1 0 3128 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 4968 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 4416 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1606821651
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_40
timestamp 1606821651
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7084 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1606821651
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_81
timestamp 1606821651
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 11040 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 10764 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606821651
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_102
timestamp 1606821651
transform 1 0 10488 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13156 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1606821651
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1606821651
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606821651
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 17388 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17940 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_175
timestamp 1606821651
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_181
timestamp 1606821651
transform 1 0 17756 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19780 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_199
timestamp 1606821651
transform 1 0 19412 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606821651
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1606821651
transform 1 0 22540 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 23276 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_231
timestamp 1606821651
transform 1 0 22356 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_236
timestamp 1606821651
transform 1 0 22816 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606821651
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2024 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1606821651
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 3772 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_26
timestamp 1606821651
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1606821651
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 8924 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1606821651
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1606821651
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 13064 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1606821651
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606821651
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_127
timestamp 1606821651
transform 1 0 12788 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1606821651
transform 1 0 13340 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15548 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_154
timestamp 1606821651
transform 1 0 15272 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_173
timestamp 1606821651
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 17204 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1606821651
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19688 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1606821651
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_218
timestamp 1606821651
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 21344 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 23276 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1606821651
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1932 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2116 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1606821651
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606821651
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5060 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4784 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3772 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1606821651
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1606821651
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1606821651
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1606821651
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6256 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 5888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_52
timestamp 1606821651
transform 1 0 5888 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_49
timestamp 1606821651
transform 1 0 5612 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606821651
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8464 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7912 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1606821651
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_78
timestamp 1606821651
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10304 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606821651
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1606821651
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1606821651
transform 1 0 9936 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11684 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12604 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 11316 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_114
timestamp 1606821651
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_131
timestamp 1606821651
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_116
timestamp 1606821651
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1606821651
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13340 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_150
timestamp 1606821651
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606821651
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_146
timestamp 1606821651
transform 1 0 14536 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_142
timestamp 1606821651
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 14536 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 14628 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15088 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16744 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 16928 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1606821651
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_168
timestamp 1606821651
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18584 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 17204 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 17756 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_179
timestamp 1606821651
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1606821651
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1606821651
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19412 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 19688 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 20240 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1606821651
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1606821651
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_199
timestamp 1606821651
transform 1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_206
timestamp 1606821651
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1606821651
transform 1 0 22540 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 21896 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 23276 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_231
timestamp 1606821651
transform 1 0 22356 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_236
timestamp 1606821651
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_224
timestamp 1606821651
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_235
timestamp 1606821651
transform 1 0 22724 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2208 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1606821651
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1606821651
transform 1 0 4232 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4784 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1606821651
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_38
timestamp 1606821651
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6440 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1606821651
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1606821651
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8096 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1606821651
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1606821651
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606821651
transform 1 0 10304 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606821651
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_97
timestamp 1606821651
transform 1 0 10028 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 11960 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 12880 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1606821651
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_122
timestamp 1606821651
transform 1 0 12328 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606821651
transform 1 0 14628 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_144
timestamp 1606821651
transform 1 0 14352 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606821651
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606821651
transform 1 0 16928 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1606821651
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 19044 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 17388 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_175
timestamp 1606821651
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1606821651
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_204
timestamp 1606821651
transform 1 0 19872 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606821651
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_218
timestamp 1606821651
transform 1 0 21160 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 21344 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 23276 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_236
timestamp 1606821651
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2300 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1606821651
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 4048 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4600 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_29
timestamp 1606821651
transform 1 0 3772 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1606821651
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1606821651
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1606821651
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606821651
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1606821651
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8280 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1606821651
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 10212 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1606821651
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1606821651
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 12972 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_115
timestamp 1606821651
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606821651
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_127
timestamp 1606821651
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 14628 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 1606821651
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16652 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15640 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_156
timestamp 1606821651
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_167
timestamp 1606821651
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606821651
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_178
timestamp 1606821651
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 20056 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 20608 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_200
timestamp 1606821651
transform 1 0 19504 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1606821651
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 21804 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 23276 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_221
timestamp 1606821651
transform 1 0 21436 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_234
timestamp 1606821651
transform 1 0 22632 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2300 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1606821651
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 5060 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606821651
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1606821651
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 6808 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1606821651
transform 1 0 6256 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1606821651
transform 1 0 5888 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_60
timestamp 1606821651
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 7912 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_71
timestamp 1606821651
transform 1 0 7636 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 10212 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1606821651
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1606821651
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11868 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1606821651
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606821651
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13524 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1606821651
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_144
timestamp 1606821651
transform 1 0 14352 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1606821651
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15364 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_154
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_171
timestamp 1606821651
transform 1 0 16836 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 19044 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 17388 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_193
timestamp 1606821651
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1606821651
transform 1 0 20056 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_204
timestamp 1606821651
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1606821651
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 23276 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_235
timestamp 1606821651
transform 1 0 22724 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1606821651
transform 1 0 3036 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1606821651
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4692 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1606821651
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 6992 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_48
timestamp 1606821651
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606821651
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 7544 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 8556 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_68
timestamp 1606821651
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1606821651
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 10304 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_31_97
timestamp 1606821651
transform 1 0 10028 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1606821651
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606821651
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606821651
transform 1 0 13708 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 14260 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15088 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1606821651
transform 1 0 13248 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_136
timestamp 1606821651
transform 1 0 13616 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_141
timestamp 1606821651
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16284 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1606821651
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_161
timestamp 1606821651
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_174
timestamp 1606821651
transform 1 0 17112 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1606821651
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1606821651
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 20976 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1606821651
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1606821651
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_215
timestamp 1606821651
transform 1 0 20884 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_232
timestamp 1606821651
transform 1 0 22448 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606821651
transform 1 0 3036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_19
timestamp 1606821651
transform 1 0 2852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 4416 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_25
timestamp 1606821651
transform 1 0 3404 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1606821651
transform 1 0 6256 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_52
timestamp 1606821651
transform 1 0 5888 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_65
timestamp 1606821651
transform 1 0 7084 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 7912 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_72
timestamp 1606821651
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 10396 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1606821651
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1606821651
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_98
timestamp 1606821651
transform 1 0 10120 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 12052 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1606821651
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606821651
transform 1 0 14720 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 13524 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1606821651
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1606821651
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1606821651
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606821651
transform 1 0 17020 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1606821651
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1606821651
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1606821651
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1606821651
transform 1 0 17756 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_32_178
timestamp 1606821651
transform 1 0 17480 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1606821651
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1606821651
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_208
timestamp 1606821651
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_215
timestamp 1606821651
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1606821651
transform 1 0 21252 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1606821651
transform 1 0 22264 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 23276 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1606821651
transform 1 0 22080 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_235
timestamp 1606821651
transform 1 0 22724 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606821651
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1606821651
transform 1 0 1656 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1606821651
transform 1 0 1932 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606821651
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606821651
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1606821651
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_7
timestamp 1606821651
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606821651
transform 1 0 5060 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1606821651
transform 1 0 3404 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 5060 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1606821651
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_22
timestamp 1606821651
transform 1 0 3128 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_41
timestamp 1606821651
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_25
timestamp 1606821651
transform 1 0 3404 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1606821651
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 5888 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1606821651
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1606821651
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1606821651
transform 1 0 5428 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_51
timestamp 1606821651
transform 1 0 5796 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 7544 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 8464 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_78
timestamp 1606821651
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_68
timestamp 1606821651
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_86
timestamp 1606821651
transform 1 0 9016 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 11040 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 10396 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1606821651
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1606821651
transform 1 0 9936 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_100
timestamp 1606821651
transform 1 0 10304 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_102
timestamp 1606821651
transform 1 0 10488 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606821651
transform 1 0 12696 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 13064 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1606821651
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_117
timestamp 1606821651
transform 1 0 11868 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1606821651
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_123
timestamp 1606821651
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_130
timestamp 1606821651
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_124
timestamp 1606821651
transform 1 0 12512 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 13248 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1606821651
transform 1 0 14904 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1606821651
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_146
timestamp 1606821651
transform 1 0 14536 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1606821651
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606821651
transform 1 0 16928 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1606821651
transform 1 0 16560 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1606821651
transform 1 0 15272 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1606821651
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1606821651
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_170
timestamp 1606821651
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 17480 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1606821651
transform 1 0 19136 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1606821651
transform 1 0 18032 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1606821651
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1606821651
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_176
timestamp 1606821651
transform 1 0 17296 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1606821651
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 19688 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1606821651
transform 1 0 20884 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1606821651
transform 1 0 20792 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1606821651
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_200
timestamp 1606821651
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_211
timestamp 1606821651
transform 1 0 20516 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1606821651
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1606821651
transform 1 0 22540 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1606821651
transform 1 0 22448 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606821651
transform -1 0 23276 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606821651
transform -1 0 23276 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_230
timestamp 1606821651
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1606821651
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_231
timestamp 1606821651
transform 1 0 22356 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_236
timestamp 1606821651
transform 1 0 22816 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606821651
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1606821651
transform 1 0 2944 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 1932 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1606821651
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1606821651
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_18
timestamp 1606821651
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606821651
transform 1 0 5060 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1606821651
transform 1 0 4048 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1606821651
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_29
timestamp 1606821651
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1606821651
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 5796 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1606821651
transform 1 0 6900 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1606821651
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_47
timestamp 1606821651
transform 1 0 5428 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_60
timestamp 1606821651
transform 1 0 6624 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1606821651
transform 1 0 7912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_72
timestamp 1606821651
transform 1 0 7728 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_77
timestamp 1606821651
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606821651
transform 1 0 9752 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1606821651
transform 1 0 10672 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1606821651
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_88
timestamp 1606821651
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_92
timestamp 1606821651
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_98
timestamp 1606821651
transform 1 0 10120 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1606821651
transform 1 0 12604 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1606821651
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_120
timestamp 1606821651
transform 1 0 12144 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606821651
transform 1 0 14812 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 13616 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_134
timestamp 1606821651
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_145
timestamp 1606821651
transform 1 0 14444 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1606821651
transform 1 0 15456 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16468 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1606821651
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_153
timestamp 1606821651
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_165
timestamp 1606821651
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606821651
transform 1 0 17664 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606821651
transform 1 0 18308 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1606821651
transform 1 0 18860 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1606821651
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1606821651
transform 1 0 17296 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_184
timestamp 1606821651
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_191
timestamp 1606821651
transform 1 0 18676 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1606821651
transform 1 0 21160 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1606821651
transform 1 0 20516 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1606821651
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_209
timestamp 1606821651
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_215
timestamp 1606821651
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1606821651
transform 1 0 22172 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1606821651
transform -1 0 23276 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_227
timestamp 1606821651
transform 1 0 21988 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_233
timestamp 1606821651
transform 1 0 22540 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_237
timestamp 1606821651
transform 1 0 22908 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 8574 0 8630 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 16946 23920 17002 24400 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 12070 0 12126 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 17590 23920 17646 24400 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal3 s 23920 6808 24400 6928 6 Test_en_E_in
port 4 nsew default input
rlabel metal3 s 23920 6128 24400 6248 6 Test_en_E_out
port 5 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 Test_en_W_in
port 6 nsew default input
rlabel metal3 s 0 15104 480 15224 6 Test_en_W_out
port 7 nsew default tristate
rlabel metal2 s 1674 0 1730 480 6 bottom_width_0_height_0__pin_50_
port 8 nsew default tristate
rlabel metal2 s 5078 0 5134 480 6 bottom_width_0_height_0__pin_51_
port 9 nsew default tristate
rlabel metal3 s 0 8984 480 9104 6 ccff_head
port 10 nsew default input
rlabel metal3 s 23920 5448 24400 5568 6 ccff_tail
port 11 nsew default tristate
rlabel metal2 s 18234 23920 18290 24400 6 clk_0_N_in
port 12 nsew default input
rlabel metal2 s 15566 0 15622 480 6 clk_0_S_in
port 13 nsew default input
rlabel metal3 s 23920 8168 24400 8288 6 prog_clk_0_E_out
port 14 nsew default tristate
rlabel metal3 s 23920 7488 24400 7608 6 prog_clk_0_N_in
port 15 nsew default input
rlabel metal2 s 18878 23920 18934 24400 6 prog_clk_0_N_out
port 16 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 prog_clk_0_S_in
port 17 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_0_S_out
port 18 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 prog_clk_0_W_out
port 19 nsew default tristate
rlabel metal3 s 23920 8712 24400 8832 6 right_width_0_height_0__pin_16_
port 20 nsew default input
rlabel metal3 s 23920 9392 24400 9512 6 right_width_0_height_0__pin_17_
port 21 nsew default input
rlabel metal3 s 23920 10072 24400 10192 6 right_width_0_height_0__pin_18_
port 22 nsew default input
rlabel metal3 s 23920 10752 24400 10872 6 right_width_0_height_0__pin_19_
port 23 nsew default input
rlabel metal3 s 23920 11432 24400 11552 6 right_width_0_height_0__pin_20_
port 24 nsew default input
rlabel metal3 s 23920 12112 24400 12232 6 right_width_0_height_0__pin_21_
port 25 nsew default input
rlabel metal3 s 23920 12656 24400 12776 6 right_width_0_height_0__pin_22_
port 26 nsew default input
rlabel metal3 s 23920 13336 24400 13456 6 right_width_0_height_0__pin_23_
port 27 nsew default input
rlabel metal3 s 23920 14016 24400 14136 6 right_width_0_height_0__pin_24_
port 28 nsew default input
rlabel metal3 s 23920 14696 24400 14816 6 right_width_0_height_0__pin_25_
port 29 nsew default input
rlabel metal3 s 23920 15376 24400 15496 6 right_width_0_height_0__pin_26_
port 30 nsew default input
rlabel metal3 s 23920 16056 24400 16176 6 right_width_0_height_0__pin_27_
port 31 nsew default input
rlabel metal3 s 23920 16600 24400 16720 6 right_width_0_height_0__pin_28_
port 32 nsew default input
rlabel metal3 s 23920 17280 24400 17400 6 right_width_0_height_0__pin_29_
port 33 nsew default input
rlabel metal3 s 23920 17960 24400 18080 6 right_width_0_height_0__pin_30_
port 34 nsew default input
rlabel metal3 s 23920 18640 24400 18760 6 right_width_0_height_0__pin_31_
port 35 nsew default input
rlabel metal3 s 23920 280 24400 400 6 right_width_0_height_0__pin_42_lower
port 36 nsew default tristate
rlabel metal3 s 23920 19320 24400 19440 6 right_width_0_height_0__pin_42_upper
port 37 nsew default tristate
rlabel metal3 s 23920 824 24400 944 6 right_width_0_height_0__pin_43_lower
port 38 nsew default tristate
rlabel metal3 s 23920 20000 24400 20120 6 right_width_0_height_0__pin_43_upper
port 39 nsew default tristate
rlabel metal3 s 23920 1504 24400 1624 6 right_width_0_height_0__pin_44_lower
port 40 nsew default tristate
rlabel metal3 s 23920 20544 24400 20664 6 right_width_0_height_0__pin_44_upper
port 41 nsew default tristate
rlabel metal3 s 23920 2184 24400 2304 6 right_width_0_height_0__pin_45_lower
port 42 nsew default tristate
rlabel metal3 s 23920 21224 24400 21344 6 right_width_0_height_0__pin_45_upper
port 43 nsew default tristate
rlabel metal3 s 23920 2864 24400 2984 6 right_width_0_height_0__pin_46_lower
port 44 nsew default tristate
rlabel metal3 s 23920 21904 24400 22024 6 right_width_0_height_0__pin_46_upper
port 45 nsew default tristate
rlabel metal3 s 23920 3544 24400 3664 6 right_width_0_height_0__pin_47_lower
port 46 nsew default tristate
rlabel metal3 s 23920 22584 24400 22704 6 right_width_0_height_0__pin_47_upper
port 47 nsew default tristate
rlabel metal3 s 23920 4224 24400 4344 6 right_width_0_height_0__pin_48_lower
port 48 nsew default tristate
rlabel metal3 s 23920 23264 24400 23384 6 right_width_0_height_0__pin_48_upper
port 49 nsew default tristate
rlabel metal3 s 23920 4768 24400 4888 6 right_width_0_height_0__pin_49_lower
port 50 nsew default tristate
rlabel metal3 s 23920 23944 24400 24064 6 right_width_0_height_0__pin_49_upper
port 51 nsew default tristate
rlabel metal2 s 5354 23920 5410 24400 6 top_width_0_height_0__pin_0_
port 52 nsew default input
rlabel metal2 s 11794 23920 11850 24400 6 top_width_0_height_0__pin_10_
port 53 nsew default input
rlabel metal2 s 12438 23920 12494 24400 6 top_width_0_height_0__pin_11_
port 54 nsew default input
rlabel metal2 s 13082 23920 13138 24400 6 top_width_0_height_0__pin_12_
port 55 nsew default input
rlabel metal2 s 13726 23920 13782 24400 6 top_width_0_height_0__pin_13_
port 56 nsew default input
rlabel metal2 s 14370 23920 14426 24400 6 top_width_0_height_0__pin_14_
port 57 nsew default input
rlabel metal2 s 15014 23920 15070 24400 6 top_width_0_height_0__pin_15_
port 58 nsew default input
rlabel metal2 s 5998 23920 6054 24400 6 top_width_0_height_0__pin_1_
port 59 nsew default input
rlabel metal2 s 6642 23920 6698 24400 6 top_width_0_height_0__pin_2_
port 60 nsew default input
rlabel metal2 s 15658 23920 15714 24400 6 top_width_0_height_0__pin_32_
port 61 nsew default input
rlabel metal2 s 16302 23920 16358 24400 6 top_width_0_height_0__pin_33_
port 62 nsew default input
rlabel metal2 s 19522 23920 19578 24400 6 top_width_0_height_0__pin_34_lower
port 63 nsew default tristate
rlabel metal2 s 294 23920 350 24400 6 top_width_0_height_0__pin_34_upper
port 64 nsew default tristate
rlabel metal2 s 20166 23920 20222 24400 6 top_width_0_height_0__pin_35_lower
port 65 nsew default tristate
rlabel metal2 s 846 23920 902 24400 6 top_width_0_height_0__pin_35_upper
port 66 nsew default tristate
rlabel metal2 s 20810 23920 20866 24400 6 top_width_0_height_0__pin_36_lower
port 67 nsew default tristate
rlabel metal2 s 1490 23920 1546 24400 6 top_width_0_height_0__pin_36_upper
port 68 nsew default tristate
rlabel metal2 s 21454 23920 21510 24400 6 top_width_0_height_0__pin_37_lower
port 69 nsew default tristate
rlabel metal2 s 2134 23920 2190 24400 6 top_width_0_height_0__pin_37_upper
port 70 nsew default tristate
rlabel metal2 s 22098 23920 22154 24400 6 top_width_0_height_0__pin_38_lower
port 71 nsew default tristate
rlabel metal2 s 2778 23920 2834 24400 6 top_width_0_height_0__pin_38_upper
port 72 nsew default tristate
rlabel metal2 s 22742 23920 22798 24400 6 top_width_0_height_0__pin_39_lower
port 73 nsew default tristate
rlabel metal2 s 3422 23920 3478 24400 6 top_width_0_height_0__pin_39_upper
port 74 nsew default tristate
rlabel metal2 s 7286 23920 7342 24400 6 top_width_0_height_0__pin_3_
port 75 nsew default input
rlabel metal2 s 23386 23920 23442 24400 6 top_width_0_height_0__pin_40_lower
port 76 nsew default tristate
rlabel metal2 s 4066 23920 4122 24400 6 top_width_0_height_0__pin_40_upper
port 77 nsew default tristate
rlabel metal2 s 24030 23920 24086 24400 6 top_width_0_height_0__pin_41_lower
port 78 nsew default tristate
rlabel metal2 s 4710 23920 4766 24400 6 top_width_0_height_0__pin_41_upper
port 79 nsew default tristate
rlabel metal2 s 7930 23920 7986 24400 6 top_width_0_height_0__pin_4_
port 80 nsew default input
rlabel metal2 s 8574 23920 8630 24400 6 top_width_0_height_0__pin_5_
port 81 nsew default input
rlabel metal2 s 9218 23920 9274 24400 6 top_width_0_height_0__pin_6_
port 82 nsew default input
rlabel metal2 s 9862 23920 9918 24400 6 top_width_0_height_0__pin_7_
port 83 nsew default input
rlabel metal2 s 10506 23920 10562 24400 6 top_width_0_height_0__pin_8_
port 84 nsew default input
rlabel metal2 s 11150 23920 11206 24400 6 top_width_0_height_0__pin_9_
port 85 nsew default input
rlabel metal4 s 4643 2128 4963 21808 6 VPWR
port 86 nsew default input
rlabel metal4 s 8341 2128 8661 21808 6 VGND
port 87 nsew default input
<< properties >>
string FIXED_BBOX 0 0 24400 24400
<< end >>
