magic
tech sky130A
magscale 1 2
timestamp 1606236591
<< viali >>
rect 1777 8449 1811 8483
rect 1869 8313 1903 8347
rect 2789 8313 2823 8347
rect 2237 8041 2271 8075
rect 2053 7905 2087 7939
rect 2743 7497 2777 7531
rect 2672 7293 2706 7327
rect 2605 6341 2639 6375
rect 2973 6205 3007 6239
rect 3341 6137 3375 6171
rect 5825 5797 5859 5831
rect 5733 5661 5767 5695
rect 6745 5661 6779 5695
rect 2237 4029 2271 4063
rect 2504 3961 2538 3995
rect 3617 3893 3651 3927
<< metal1 >>
rect 1104 14714 7820 14736
rect 1104 14662 3246 14714
rect 3298 14662 3310 14714
rect 3362 14662 3374 14714
rect 3426 14662 3438 14714
rect 3490 14662 5510 14714
rect 5562 14662 5574 14714
rect 5626 14662 5638 14714
rect 5690 14662 5702 14714
rect 5754 14662 7820 14714
rect 1104 14640 7820 14662
rect 1104 14170 7820 14192
rect 1104 14118 2114 14170
rect 2166 14118 2178 14170
rect 2230 14118 2242 14170
rect 2294 14118 2306 14170
rect 2358 14118 4378 14170
rect 4430 14118 4442 14170
rect 4494 14118 4506 14170
rect 4558 14118 4570 14170
rect 4622 14118 6642 14170
rect 6694 14118 6706 14170
rect 6758 14118 6770 14170
rect 6822 14118 6834 14170
rect 6886 14118 7820 14170
rect 1104 14096 7820 14118
rect 1104 13626 7820 13648
rect 1104 13574 3246 13626
rect 3298 13574 3310 13626
rect 3362 13574 3374 13626
rect 3426 13574 3438 13626
rect 3490 13574 5510 13626
rect 5562 13574 5574 13626
rect 5626 13574 5638 13626
rect 5690 13574 5702 13626
rect 5754 13574 7820 13626
rect 1104 13552 7820 13574
rect 1104 13082 7820 13104
rect 1104 13030 2114 13082
rect 2166 13030 2178 13082
rect 2230 13030 2242 13082
rect 2294 13030 2306 13082
rect 2358 13030 4378 13082
rect 4430 13030 4442 13082
rect 4494 13030 4506 13082
rect 4558 13030 4570 13082
rect 4622 13030 6642 13082
rect 6694 13030 6706 13082
rect 6758 13030 6770 13082
rect 6822 13030 6834 13082
rect 6886 13030 7820 13082
rect 1104 13008 7820 13030
rect 1104 12538 7820 12560
rect 1104 12486 3246 12538
rect 3298 12486 3310 12538
rect 3362 12486 3374 12538
rect 3426 12486 3438 12538
rect 3490 12486 5510 12538
rect 5562 12486 5574 12538
rect 5626 12486 5638 12538
rect 5690 12486 5702 12538
rect 5754 12486 7820 12538
rect 1104 12464 7820 12486
rect 1104 11994 7820 12016
rect 1104 11942 2114 11994
rect 2166 11942 2178 11994
rect 2230 11942 2242 11994
rect 2294 11942 2306 11994
rect 2358 11942 4378 11994
rect 4430 11942 4442 11994
rect 4494 11942 4506 11994
rect 4558 11942 4570 11994
rect 4622 11942 6642 11994
rect 6694 11942 6706 11994
rect 6758 11942 6770 11994
rect 6822 11942 6834 11994
rect 6886 11942 7820 11994
rect 1104 11920 7820 11942
rect 1104 11450 7820 11472
rect 1104 11398 3246 11450
rect 3298 11398 3310 11450
rect 3362 11398 3374 11450
rect 3426 11398 3438 11450
rect 3490 11398 5510 11450
rect 5562 11398 5574 11450
rect 5626 11398 5638 11450
rect 5690 11398 5702 11450
rect 5754 11398 7820 11450
rect 1104 11376 7820 11398
rect 1104 10906 7820 10928
rect 1104 10854 2114 10906
rect 2166 10854 2178 10906
rect 2230 10854 2242 10906
rect 2294 10854 2306 10906
rect 2358 10854 4378 10906
rect 4430 10854 4442 10906
rect 4494 10854 4506 10906
rect 4558 10854 4570 10906
rect 4622 10854 6642 10906
rect 6694 10854 6706 10906
rect 6758 10854 6770 10906
rect 6822 10854 6834 10906
rect 6886 10854 7820 10906
rect 1104 10832 7820 10854
rect 1104 10362 7820 10384
rect 1104 10310 3246 10362
rect 3298 10310 3310 10362
rect 3362 10310 3374 10362
rect 3426 10310 3438 10362
rect 3490 10310 5510 10362
rect 5562 10310 5574 10362
rect 5626 10310 5638 10362
rect 5690 10310 5702 10362
rect 5754 10310 7820 10362
rect 1104 10288 7820 10310
rect 1104 9818 7820 9840
rect 1104 9766 2114 9818
rect 2166 9766 2178 9818
rect 2230 9766 2242 9818
rect 2294 9766 2306 9818
rect 2358 9766 4378 9818
rect 4430 9766 4442 9818
rect 4494 9766 4506 9818
rect 4558 9766 4570 9818
rect 4622 9766 6642 9818
rect 6694 9766 6706 9818
rect 6758 9766 6770 9818
rect 6822 9766 6834 9818
rect 6886 9766 7820 9818
rect 1104 9744 7820 9766
rect 1104 9274 7820 9296
rect 1104 9222 3246 9274
rect 3298 9222 3310 9274
rect 3362 9222 3374 9274
rect 3426 9222 3438 9274
rect 3490 9222 5510 9274
rect 5562 9222 5574 9274
rect 5626 9222 5638 9274
rect 5690 9222 5702 9274
rect 5754 9222 7820 9274
rect 1104 9200 7820 9222
rect 1104 8730 7820 8752
rect 1104 8678 2114 8730
rect 2166 8678 2178 8730
rect 2230 8678 2242 8730
rect 2294 8678 2306 8730
rect 2358 8678 4378 8730
rect 4430 8678 4442 8730
rect 4494 8678 4506 8730
rect 4558 8678 4570 8730
rect 4622 8678 6642 8730
rect 6694 8678 6706 8730
rect 6758 8678 6770 8730
rect 6822 8678 6834 8730
rect 6886 8678 7820 8730
rect 1104 8656 7820 8678
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 2774 8480 2780 8492
rect 1811 8452 2780 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 1854 8344 1860 8356
rect 1815 8316 1860 8344
rect 1854 8304 1860 8316
rect 1912 8304 1918 8356
rect 1946 8304 1952 8356
rect 2004 8344 2010 8356
rect 2777 8347 2835 8353
rect 2777 8344 2789 8347
rect 2004 8316 2789 8344
rect 2004 8304 2010 8316
rect 2777 8313 2789 8316
rect 2823 8313 2835 8347
rect 2777 8307 2835 8313
rect 1104 8186 7820 8208
rect 1104 8134 3246 8186
rect 3298 8134 3310 8186
rect 3362 8134 3374 8186
rect 3426 8134 3438 8186
rect 3490 8134 5510 8186
rect 5562 8134 5574 8186
rect 5626 8134 5638 8186
rect 5690 8134 5702 8186
rect 5754 8134 7820 8186
rect 1104 8112 7820 8134
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 1946 7896 1952 7948
rect 2004 7936 2010 7948
rect 2041 7939 2099 7945
rect 2041 7936 2053 7939
rect 2004 7908 2053 7936
rect 2004 7896 2010 7908
rect 2041 7905 2053 7908
rect 2087 7905 2099 7939
rect 2041 7899 2099 7905
rect 1104 7642 7820 7664
rect 1104 7590 2114 7642
rect 2166 7590 2178 7642
rect 2230 7590 2242 7642
rect 2294 7590 2306 7642
rect 2358 7590 4378 7642
rect 4430 7590 4442 7642
rect 4494 7590 4506 7642
rect 4558 7590 4570 7642
rect 4622 7590 6642 7642
rect 6694 7590 6706 7642
rect 6758 7590 6770 7642
rect 6822 7590 6834 7642
rect 6886 7590 7820 7642
rect 1104 7568 7820 7590
rect 1854 7488 1860 7540
rect 1912 7528 1918 7540
rect 2731 7531 2789 7537
rect 2731 7528 2743 7531
rect 1912 7500 2743 7528
rect 1912 7488 1918 7500
rect 2731 7497 2743 7500
rect 2777 7497 2789 7531
rect 2731 7491 2789 7497
rect 2660 7327 2718 7333
rect 2660 7293 2672 7327
rect 2706 7324 2718 7327
rect 5350 7324 5356 7336
rect 2706 7296 5356 7324
rect 2706 7293 2718 7296
rect 2660 7287 2718 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 1104 7098 7820 7120
rect 1104 7046 3246 7098
rect 3298 7046 3310 7098
rect 3362 7046 3374 7098
rect 3426 7046 3438 7098
rect 3490 7046 5510 7098
rect 5562 7046 5574 7098
rect 5626 7046 5638 7098
rect 5690 7046 5702 7098
rect 5754 7046 7820 7098
rect 1104 7024 7820 7046
rect 1104 6554 7820 6576
rect 1104 6502 2114 6554
rect 2166 6502 2178 6554
rect 2230 6502 2242 6554
rect 2294 6502 2306 6554
rect 2358 6502 4378 6554
rect 4430 6502 4442 6554
rect 4494 6502 4506 6554
rect 4558 6502 4570 6554
rect 4622 6502 6642 6554
rect 6694 6502 6706 6554
rect 6758 6502 6770 6554
rect 6822 6502 6834 6554
rect 6886 6502 7820 6554
rect 1104 6480 7820 6502
rect 2593 6375 2651 6381
rect 2593 6341 2605 6375
rect 2639 6372 2651 6375
rect 2866 6372 2872 6384
rect 2639 6344 2872 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 2958 6236 2964 6248
rect 2919 6208 2964 6236
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 3329 6171 3387 6177
rect 3329 6137 3341 6171
rect 3375 6168 3387 6171
rect 5350 6168 5356 6180
rect 3375 6140 5356 6168
rect 3375 6137 3387 6140
rect 3329 6131 3387 6137
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 1104 6010 7820 6032
rect 1104 5958 3246 6010
rect 3298 5958 3310 6010
rect 3362 5958 3374 6010
rect 3426 5958 3438 6010
rect 3490 5958 5510 6010
rect 5562 5958 5574 6010
rect 5626 5958 5638 6010
rect 5690 5958 5702 6010
rect 5754 5958 7820 6010
rect 1104 5936 7820 5958
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 5813 5831 5871 5837
rect 5813 5828 5825 5831
rect 5408 5800 5825 5828
rect 5408 5788 5414 5800
rect 5813 5797 5825 5800
rect 5859 5797 5871 5831
rect 5813 5791 5871 5797
rect 4154 5652 4160 5704
rect 4212 5692 4218 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 4212 5664 5733 5692
rect 4212 5652 4218 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 7834 5692 7840 5704
rect 6779 5664 7840 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 1104 5466 7820 5488
rect 1104 5414 2114 5466
rect 2166 5414 2178 5466
rect 2230 5414 2242 5466
rect 2294 5414 2306 5466
rect 2358 5414 4378 5466
rect 4430 5414 4442 5466
rect 4494 5414 4506 5466
rect 4558 5414 4570 5466
rect 4622 5414 6642 5466
rect 6694 5414 6706 5466
rect 6758 5414 6770 5466
rect 6822 5414 6834 5466
rect 6886 5414 7820 5466
rect 1104 5392 7820 5414
rect 1104 4922 7820 4944
rect 1104 4870 3246 4922
rect 3298 4870 3310 4922
rect 3362 4870 3374 4922
rect 3426 4870 3438 4922
rect 3490 4870 5510 4922
rect 5562 4870 5574 4922
rect 5626 4870 5638 4922
rect 5690 4870 5702 4922
rect 5754 4870 7820 4922
rect 1104 4848 7820 4870
rect 1104 4378 7820 4400
rect 1104 4326 2114 4378
rect 2166 4326 2178 4378
rect 2230 4326 2242 4378
rect 2294 4326 2306 4378
rect 2358 4326 4378 4378
rect 4430 4326 4442 4378
rect 4494 4326 4506 4378
rect 4558 4326 4570 4378
rect 4622 4326 6642 4378
rect 6694 4326 6706 4378
rect 6758 4326 6770 4378
rect 6822 4326 6834 4378
rect 6886 4326 7820 4378
rect 1104 4304 7820 4326
rect 1118 4020 1124 4072
rect 1176 4060 1182 4072
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 1176 4032 2237 4060
rect 1176 4020 1182 4032
rect 2225 4029 2237 4032
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 2492 3995 2550 4001
rect 2492 3961 2504 3995
rect 2538 3992 2550 3995
rect 3142 3992 3148 4004
rect 2538 3964 3148 3992
rect 2538 3961 2550 3964
rect 2492 3955 2550 3961
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 3605 3927 3663 3933
rect 3605 3924 3617 3927
rect 3016 3896 3617 3924
rect 3016 3884 3022 3896
rect 3605 3893 3617 3896
rect 3651 3924 3663 3927
rect 5810 3924 5816 3936
rect 3651 3896 5816 3924
rect 3651 3893 3663 3896
rect 3605 3887 3663 3893
rect 5810 3884 5816 3896
rect 5868 3884 5874 3936
rect 1104 3834 7820 3856
rect 1104 3782 3246 3834
rect 3298 3782 3310 3834
rect 3362 3782 3374 3834
rect 3426 3782 3438 3834
rect 3490 3782 5510 3834
rect 5562 3782 5574 3834
rect 5626 3782 5638 3834
rect 5690 3782 5702 3834
rect 5754 3782 7820 3834
rect 1104 3760 7820 3782
rect 1104 3290 7820 3312
rect 1104 3238 2114 3290
rect 2166 3238 2178 3290
rect 2230 3238 2242 3290
rect 2294 3238 2306 3290
rect 2358 3238 4378 3290
rect 4430 3238 4442 3290
rect 4494 3238 4506 3290
rect 4558 3238 4570 3290
rect 4622 3238 6642 3290
rect 6694 3238 6706 3290
rect 6758 3238 6770 3290
rect 6822 3238 6834 3290
rect 6886 3238 7820 3290
rect 1104 3216 7820 3238
rect 1104 2746 7820 2768
rect 1104 2694 3246 2746
rect 3298 2694 3310 2746
rect 3362 2694 3374 2746
rect 3426 2694 3438 2746
rect 3490 2694 5510 2746
rect 5562 2694 5574 2746
rect 5626 2694 5638 2746
rect 5690 2694 5702 2746
rect 5754 2694 7820 2746
rect 1104 2672 7820 2694
rect 1104 2202 7820 2224
rect 1104 2150 2114 2202
rect 2166 2150 2178 2202
rect 2230 2150 2242 2202
rect 2294 2150 2306 2202
rect 2358 2150 4378 2202
rect 4430 2150 4442 2202
rect 4494 2150 4506 2202
rect 4558 2150 4570 2202
rect 4622 2150 6642 2202
rect 6694 2150 6706 2202
rect 6758 2150 6770 2202
rect 6822 2150 6834 2202
rect 6886 2150 7820 2202
rect 1104 2128 7820 2150
<< via1 >>
rect 3246 14662 3298 14714
rect 3310 14662 3362 14714
rect 3374 14662 3426 14714
rect 3438 14662 3490 14714
rect 5510 14662 5562 14714
rect 5574 14662 5626 14714
rect 5638 14662 5690 14714
rect 5702 14662 5754 14714
rect 2114 14118 2166 14170
rect 2178 14118 2230 14170
rect 2242 14118 2294 14170
rect 2306 14118 2358 14170
rect 4378 14118 4430 14170
rect 4442 14118 4494 14170
rect 4506 14118 4558 14170
rect 4570 14118 4622 14170
rect 6642 14118 6694 14170
rect 6706 14118 6758 14170
rect 6770 14118 6822 14170
rect 6834 14118 6886 14170
rect 3246 13574 3298 13626
rect 3310 13574 3362 13626
rect 3374 13574 3426 13626
rect 3438 13574 3490 13626
rect 5510 13574 5562 13626
rect 5574 13574 5626 13626
rect 5638 13574 5690 13626
rect 5702 13574 5754 13626
rect 2114 13030 2166 13082
rect 2178 13030 2230 13082
rect 2242 13030 2294 13082
rect 2306 13030 2358 13082
rect 4378 13030 4430 13082
rect 4442 13030 4494 13082
rect 4506 13030 4558 13082
rect 4570 13030 4622 13082
rect 6642 13030 6694 13082
rect 6706 13030 6758 13082
rect 6770 13030 6822 13082
rect 6834 13030 6886 13082
rect 3246 12486 3298 12538
rect 3310 12486 3362 12538
rect 3374 12486 3426 12538
rect 3438 12486 3490 12538
rect 5510 12486 5562 12538
rect 5574 12486 5626 12538
rect 5638 12486 5690 12538
rect 5702 12486 5754 12538
rect 2114 11942 2166 11994
rect 2178 11942 2230 11994
rect 2242 11942 2294 11994
rect 2306 11942 2358 11994
rect 4378 11942 4430 11994
rect 4442 11942 4494 11994
rect 4506 11942 4558 11994
rect 4570 11942 4622 11994
rect 6642 11942 6694 11994
rect 6706 11942 6758 11994
rect 6770 11942 6822 11994
rect 6834 11942 6886 11994
rect 3246 11398 3298 11450
rect 3310 11398 3362 11450
rect 3374 11398 3426 11450
rect 3438 11398 3490 11450
rect 5510 11398 5562 11450
rect 5574 11398 5626 11450
rect 5638 11398 5690 11450
rect 5702 11398 5754 11450
rect 2114 10854 2166 10906
rect 2178 10854 2230 10906
rect 2242 10854 2294 10906
rect 2306 10854 2358 10906
rect 4378 10854 4430 10906
rect 4442 10854 4494 10906
rect 4506 10854 4558 10906
rect 4570 10854 4622 10906
rect 6642 10854 6694 10906
rect 6706 10854 6758 10906
rect 6770 10854 6822 10906
rect 6834 10854 6886 10906
rect 3246 10310 3298 10362
rect 3310 10310 3362 10362
rect 3374 10310 3426 10362
rect 3438 10310 3490 10362
rect 5510 10310 5562 10362
rect 5574 10310 5626 10362
rect 5638 10310 5690 10362
rect 5702 10310 5754 10362
rect 2114 9766 2166 9818
rect 2178 9766 2230 9818
rect 2242 9766 2294 9818
rect 2306 9766 2358 9818
rect 4378 9766 4430 9818
rect 4442 9766 4494 9818
rect 4506 9766 4558 9818
rect 4570 9766 4622 9818
rect 6642 9766 6694 9818
rect 6706 9766 6758 9818
rect 6770 9766 6822 9818
rect 6834 9766 6886 9818
rect 3246 9222 3298 9274
rect 3310 9222 3362 9274
rect 3374 9222 3426 9274
rect 3438 9222 3490 9274
rect 5510 9222 5562 9274
rect 5574 9222 5626 9274
rect 5638 9222 5690 9274
rect 5702 9222 5754 9274
rect 2114 8678 2166 8730
rect 2178 8678 2230 8730
rect 2242 8678 2294 8730
rect 2306 8678 2358 8730
rect 4378 8678 4430 8730
rect 4442 8678 4494 8730
rect 4506 8678 4558 8730
rect 4570 8678 4622 8730
rect 6642 8678 6694 8730
rect 6706 8678 6758 8730
rect 6770 8678 6822 8730
rect 6834 8678 6886 8730
rect 2780 8440 2832 8492
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 1952 8304 2004 8356
rect 3246 8134 3298 8186
rect 3310 8134 3362 8186
rect 3374 8134 3426 8186
rect 3438 8134 3490 8186
rect 5510 8134 5562 8186
rect 5574 8134 5626 8186
rect 5638 8134 5690 8186
rect 5702 8134 5754 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 1952 7896 2004 7948
rect 2114 7590 2166 7642
rect 2178 7590 2230 7642
rect 2242 7590 2294 7642
rect 2306 7590 2358 7642
rect 4378 7590 4430 7642
rect 4442 7590 4494 7642
rect 4506 7590 4558 7642
rect 4570 7590 4622 7642
rect 6642 7590 6694 7642
rect 6706 7590 6758 7642
rect 6770 7590 6822 7642
rect 6834 7590 6886 7642
rect 1860 7488 1912 7540
rect 5356 7284 5408 7336
rect 3246 7046 3298 7098
rect 3310 7046 3362 7098
rect 3374 7046 3426 7098
rect 3438 7046 3490 7098
rect 5510 7046 5562 7098
rect 5574 7046 5626 7098
rect 5638 7046 5690 7098
rect 5702 7046 5754 7098
rect 2114 6502 2166 6554
rect 2178 6502 2230 6554
rect 2242 6502 2294 6554
rect 2306 6502 2358 6554
rect 4378 6502 4430 6554
rect 4442 6502 4494 6554
rect 4506 6502 4558 6554
rect 4570 6502 4622 6554
rect 6642 6502 6694 6554
rect 6706 6502 6758 6554
rect 6770 6502 6822 6554
rect 6834 6502 6886 6554
rect 2872 6332 2924 6384
rect 2964 6239 3016 6248
rect 2964 6205 2973 6239
rect 2973 6205 3007 6239
rect 3007 6205 3016 6239
rect 2964 6196 3016 6205
rect 5356 6128 5408 6180
rect 3246 5958 3298 6010
rect 3310 5958 3362 6010
rect 3374 5958 3426 6010
rect 3438 5958 3490 6010
rect 5510 5958 5562 6010
rect 5574 5958 5626 6010
rect 5638 5958 5690 6010
rect 5702 5958 5754 6010
rect 5356 5788 5408 5840
rect 4160 5652 4212 5704
rect 7840 5652 7892 5704
rect 2114 5414 2166 5466
rect 2178 5414 2230 5466
rect 2242 5414 2294 5466
rect 2306 5414 2358 5466
rect 4378 5414 4430 5466
rect 4442 5414 4494 5466
rect 4506 5414 4558 5466
rect 4570 5414 4622 5466
rect 6642 5414 6694 5466
rect 6706 5414 6758 5466
rect 6770 5414 6822 5466
rect 6834 5414 6886 5466
rect 3246 4870 3298 4922
rect 3310 4870 3362 4922
rect 3374 4870 3426 4922
rect 3438 4870 3490 4922
rect 5510 4870 5562 4922
rect 5574 4870 5626 4922
rect 5638 4870 5690 4922
rect 5702 4870 5754 4922
rect 2114 4326 2166 4378
rect 2178 4326 2230 4378
rect 2242 4326 2294 4378
rect 2306 4326 2358 4378
rect 4378 4326 4430 4378
rect 4442 4326 4494 4378
rect 4506 4326 4558 4378
rect 4570 4326 4622 4378
rect 6642 4326 6694 4378
rect 6706 4326 6758 4378
rect 6770 4326 6822 4378
rect 6834 4326 6886 4378
rect 1124 4020 1176 4072
rect 3148 3952 3200 4004
rect 2964 3884 3016 3936
rect 5816 3884 5868 3936
rect 3246 3782 3298 3834
rect 3310 3782 3362 3834
rect 3374 3782 3426 3834
rect 3438 3782 3490 3834
rect 5510 3782 5562 3834
rect 5574 3782 5626 3834
rect 5638 3782 5690 3834
rect 5702 3782 5754 3834
rect 2114 3238 2166 3290
rect 2178 3238 2230 3290
rect 2242 3238 2294 3290
rect 2306 3238 2358 3290
rect 4378 3238 4430 3290
rect 4442 3238 4494 3290
rect 4506 3238 4558 3290
rect 4570 3238 4622 3290
rect 6642 3238 6694 3290
rect 6706 3238 6758 3290
rect 6770 3238 6822 3290
rect 6834 3238 6886 3290
rect 3246 2694 3298 2746
rect 3310 2694 3362 2746
rect 3374 2694 3426 2746
rect 3438 2694 3490 2746
rect 5510 2694 5562 2746
rect 5574 2694 5626 2746
rect 5638 2694 5690 2746
rect 5702 2694 5754 2746
rect 2114 2150 2166 2202
rect 2178 2150 2230 2202
rect 2242 2150 2294 2202
rect 2306 2150 2358 2202
rect 4378 2150 4430 2202
rect 4442 2150 4494 2202
rect 4506 2150 4558 2202
rect 4570 2150 4622 2202
rect 6642 2150 6694 2202
rect 6706 2150 6758 2202
rect 6770 2150 6822 2202
rect 6834 2150 6886 2202
<< metal2 >>
rect 2778 15328 2834 15337
rect 2778 15263 2834 15272
rect 2088 14172 2384 14192
rect 2144 14170 2168 14172
rect 2224 14170 2248 14172
rect 2304 14170 2328 14172
rect 2166 14118 2168 14170
rect 2230 14118 2242 14170
rect 2304 14118 2306 14170
rect 2144 14116 2168 14118
rect 2224 14116 2248 14118
rect 2304 14116 2328 14118
rect 2088 14096 2384 14116
rect 2088 13084 2384 13104
rect 2144 13082 2168 13084
rect 2224 13082 2248 13084
rect 2304 13082 2328 13084
rect 2166 13030 2168 13082
rect 2230 13030 2242 13082
rect 2304 13030 2306 13082
rect 2144 13028 2168 13030
rect 2224 13028 2248 13030
rect 2304 13028 2328 13030
rect 2088 13008 2384 13028
rect 2088 11996 2384 12016
rect 2144 11994 2168 11996
rect 2224 11994 2248 11996
rect 2304 11994 2328 11996
rect 2166 11942 2168 11994
rect 2230 11942 2242 11994
rect 2304 11942 2306 11994
rect 2144 11940 2168 11942
rect 2224 11940 2248 11942
rect 2304 11940 2328 11942
rect 2088 11920 2384 11940
rect 2088 10908 2384 10928
rect 2144 10906 2168 10908
rect 2224 10906 2248 10908
rect 2304 10906 2328 10908
rect 2166 10854 2168 10906
rect 2230 10854 2242 10906
rect 2304 10854 2306 10906
rect 2144 10852 2168 10854
rect 2224 10852 2248 10854
rect 2304 10852 2328 10854
rect 2088 10832 2384 10852
rect 2088 9820 2384 9840
rect 2144 9818 2168 9820
rect 2224 9818 2248 9820
rect 2304 9818 2328 9820
rect 2166 9766 2168 9818
rect 2230 9766 2242 9818
rect 2304 9766 2306 9818
rect 2144 9764 2168 9766
rect 2224 9764 2248 9766
rect 2304 9764 2328 9766
rect 2088 9744 2384 9764
rect 2088 8732 2384 8752
rect 2144 8730 2168 8732
rect 2224 8730 2248 8732
rect 2304 8730 2328 8732
rect 2166 8678 2168 8730
rect 2230 8678 2242 8730
rect 2304 8678 2306 8730
rect 2144 8676 2168 8678
rect 2224 8676 2248 8678
rect 2304 8676 2328 8678
rect 2088 8656 2384 8676
rect 2226 8528 2282 8537
rect 2792 8498 2820 15263
rect 3220 14716 3516 14736
rect 3276 14714 3300 14716
rect 3356 14714 3380 14716
rect 3436 14714 3460 14716
rect 3298 14662 3300 14714
rect 3362 14662 3374 14714
rect 3436 14662 3438 14714
rect 3276 14660 3300 14662
rect 3356 14660 3380 14662
rect 3436 14660 3460 14662
rect 3220 14640 3516 14660
rect 5484 14716 5780 14736
rect 5540 14714 5564 14716
rect 5620 14714 5644 14716
rect 5700 14714 5724 14716
rect 5562 14662 5564 14714
rect 5626 14662 5638 14714
rect 5700 14662 5702 14714
rect 5540 14660 5564 14662
rect 5620 14660 5644 14662
rect 5700 14660 5724 14662
rect 5484 14640 5780 14660
rect 4352 14172 4648 14192
rect 4408 14170 4432 14172
rect 4488 14170 4512 14172
rect 4568 14170 4592 14172
rect 4430 14118 4432 14170
rect 4494 14118 4506 14170
rect 4568 14118 4570 14170
rect 4408 14116 4432 14118
rect 4488 14116 4512 14118
rect 4568 14116 4592 14118
rect 4352 14096 4648 14116
rect 6616 14172 6912 14192
rect 6672 14170 6696 14172
rect 6752 14170 6776 14172
rect 6832 14170 6856 14172
rect 6694 14118 6696 14170
rect 6758 14118 6770 14170
rect 6832 14118 6834 14170
rect 6672 14116 6696 14118
rect 6752 14116 6776 14118
rect 6832 14116 6856 14118
rect 6616 14096 6912 14116
rect 3220 13628 3516 13648
rect 3276 13626 3300 13628
rect 3356 13626 3380 13628
rect 3436 13626 3460 13628
rect 3298 13574 3300 13626
rect 3362 13574 3374 13626
rect 3436 13574 3438 13626
rect 3276 13572 3300 13574
rect 3356 13572 3380 13574
rect 3436 13572 3460 13574
rect 3220 13552 3516 13572
rect 5484 13628 5780 13648
rect 5540 13626 5564 13628
rect 5620 13626 5644 13628
rect 5700 13626 5724 13628
rect 5562 13574 5564 13626
rect 5626 13574 5638 13626
rect 5700 13574 5702 13626
rect 5540 13572 5564 13574
rect 5620 13572 5644 13574
rect 5700 13572 5724 13574
rect 5484 13552 5780 13572
rect 4352 13084 4648 13104
rect 4408 13082 4432 13084
rect 4488 13082 4512 13084
rect 4568 13082 4592 13084
rect 4430 13030 4432 13082
rect 4494 13030 4506 13082
rect 4568 13030 4570 13082
rect 4408 13028 4432 13030
rect 4488 13028 4512 13030
rect 4568 13028 4592 13030
rect 4352 13008 4648 13028
rect 6616 13084 6912 13104
rect 6672 13082 6696 13084
rect 6752 13082 6776 13084
rect 6832 13082 6856 13084
rect 6694 13030 6696 13082
rect 6758 13030 6770 13082
rect 6832 13030 6834 13082
rect 6672 13028 6696 13030
rect 6752 13028 6776 13030
rect 6832 13028 6856 13030
rect 6616 13008 6912 13028
rect 3220 12540 3516 12560
rect 3276 12538 3300 12540
rect 3356 12538 3380 12540
rect 3436 12538 3460 12540
rect 3298 12486 3300 12538
rect 3362 12486 3374 12538
rect 3436 12486 3438 12538
rect 3276 12484 3300 12486
rect 3356 12484 3380 12486
rect 3436 12484 3460 12486
rect 3220 12464 3516 12484
rect 5484 12540 5780 12560
rect 5540 12538 5564 12540
rect 5620 12538 5644 12540
rect 5700 12538 5724 12540
rect 5562 12486 5564 12538
rect 5626 12486 5638 12538
rect 5700 12486 5702 12538
rect 5540 12484 5564 12486
rect 5620 12484 5644 12486
rect 5700 12484 5724 12486
rect 5484 12464 5780 12484
rect 4352 11996 4648 12016
rect 4408 11994 4432 11996
rect 4488 11994 4512 11996
rect 4568 11994 4592 11996
rect 4430 11942 4432 11994
rect 4494 11942 4506 11994
rect 4568 11942 4570 11994
rect 4408 11940 4432 11942
rect 4488 11940 4512 11942
rect 4568 11940 4592 11942
rect 4352 11920 4648 11940
rect 6616 11996 6912 12016
rect 6672 11994 6696 11996
rect 6752 11994 6776 11996
rect 6832 11994 6856 11996
rect 6694 11942 6696 11994
rect 6758 11942 6770 11994
rect 6832 11942 6834 11994
rect 6672 11940 6696 11942
rect 6752 11940 6776 11942
rect 6832 11940 6856 11942
rect 6616 11920 6912 11940
rect 2870 11792 2926 11801
rect 2870 11727 2926 11736
rect 2226 8463 2282 8472
rect 2780 8492 2832 8498
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1872 7546 1900 8298
rect 1964 7954 1992 8298
rect 2240 8090 2268 8463
rect 2780 8434 2832 8440
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1124 4072 1176 4078
rect 1124 4014 1176 4020
rect 1136 480 1164 4014
rect 1964 1737 1992 7890
rect 2088 7644 2384 7664
rect 2144 7642 2168 7644
rect 2224 7642 2248 7644
rect 2304 7642 2328 7644
rect 2166 7590 2168 7642
rect 2230 7590 2242 7642
rect 2304 7590 2306 7642
rect 2144 7588 2168 7590
rect 2224 7588 2248 7590
rect 2304 7588 2328 7590
rect 2088 7568 2384 7588
rect 2088 6556 2384 6576
rect 2144 6554 2168 6556
rect 2224 6554 2248 6556
rect 2304 6554 2328 6556
rect 2166 6502 2168 6554
rect 2230 6502 2242 6554
rect 2304 6502 2306 6554
rect 2144 6500 2168 6502
rect 2224 6500 2248 6502
rect 2304 6500 2328 6502
rect 2088 6480 2384 6500
rect 2884 6390 2912 11727
rect 3220 11452 3516 11472
rect 3276 11450 3300 11452
rect 3356 11450 3380 11452
rect 3436 11450 3460 11452
rect 3298 11398 3300 11450
rect 3362 11398 3374 11450
rect 3436 11398 3438 11450
rect 3276 11396 3300 11398
rect 3356 11396 3380 11398
rect 3436 11396 3460 11398
rect 3220 11376 3516 11396
rect 5484 11452 5780 11472
rect 5540 11450 5564 11452
rect 5620 11450 5644 11452
rect 5700 11450 5724 11452
rect 5562 11398 5564 11450
rect 5626 11398 5638 11450
rect 5700 11398 5702 11450
rect 5540 11396 5564 11398
rect 5620 11396 5644 11398
rect 5700 11396 5724 11398
rect 5484 11376 5780 11396
rect 4352 10908 4648 10928
rect 4408 10906 4432 10908
rect 4488 10906 4512 10908
rect 4568 10906 4592 10908
rect 4430 10854 4432 10906
rect 4494 10854 4506 10906
rect 4568 10854 4570 10906
rect 4408 10852 4432 10854
rect 4488 10852 4512 10854
rect 4568 10852 4592 10854
rect 4352 10832 4648 10852
rect 6616 10908 6912 10928
rect 6672 10906 6696 10908
rect 6752 10906 6776 10908
rect 6832 10906 6856 10908
rect 6694 10854 6696 10906
rect 6758 10854 6770 10906
rect 6832 10854 6834 10906
rect 6672 10852 6696 10854
rect 6752 10852 6776 10854
rect 6832 10852 6856 10854
rect 6616 10832 6912 10852
rect 3220 10364 3516 10384
rect 3276 10362 3300 10364
rect 3356 10362 3380 10364
rect 3436 10362 3460 10364
rect 3298 10310 3300 10362
rect 3362 10310 3374 10362
rect 3436 10310 3438 10362
rect 3276 10308 3300 10310
rect 3356 10308 3380 10310
rect 3436 10308 3460 10310
rect 3220 10288 3516 10308
rect 5484 10364 5780 10384
rect 5540 10362 5564 10364
rect 5620 10362 5644 10364
rect 5700 10362 5724 10364
rect 5562 10310 5564 10362
rect 5626 10310 5638 10362
rect 5700 10310 5702 10362
rect 5540 10308 5564 10310
rect 5620 10308 5644 10310
rect 5700 10308 5724 10310
rect 5484 10288 5780 10308
rect 4352 9820 4648 9840
rect 4408 9818 4432 9820
rect 4488 9818 4512 9820
rect 4568 9818 4592 9820
rect 4430 9766 4432 9818
rect 4494 9766 4506 9818
rect 4568 9766 4570 9818
rect 4408 9764 4432 9766
rect 4488 9764 4512 9766
rect 4568 9764 4592 9766
rect 4352 9744 4648 9764
rect 6616 9820 6912 9840
rect 6672 9818 6696 9820
rect 6752 9818 6776 9820
rect 6832 9818 6856 9820
rect 6694 9766 6696 9818
rect 6758 9766 6770 9818
rect 6832 9766 6834 9818
rect 6672 9764 6696 9766
rect 6752 9764 6776 9766
rect 6832 9764 6856 9766
rect 6616 9744 6912 9764
rect 3220 9276 3516 9296
rect 3276 9274 3300 9276
rect 3356 9274 3380 9276
rect 3436 9274 3460 9276
rect 3298 9222 3300 9274
rect 3362 9222 3374 9274
rect 3436 9222 3438 9274
rect 3276 9220 3300 9222
rect 3356 9220 3380 9222
rect 3436 9220 3460 9222
rect 3220 9200 3516 9220
rect 5484 9276 5780 9296
rect 5540 9274 5564 9276
rect 5620 9274 5644 9276
rect 5700 9274 5724 9276
rect 5562 9222 5564 9274
rect 5626 9222 5638 9274
rect 5700 9222 5702 9274
rect 5540 9220 5564 9222
rect 5620 9220 5644 9222
rect 5700 9220 5724 9222
rect 5484 9200 5780 9220
rect 4352 8732 4648 8752
rect 4408 8730 4432 8732
rect 4488 8730 4512 8732
rect 4568 8730 4592 8732
rect 4430 8678 4432 8730
rect 4494 8678 4506 8730
rect 4568 8678 4570 8730
rect 4408 8676 4432 8678
rect 4488 8676 4512 8678
rect 4568 8676 4592 8678
rect 4352 8656 4648 8676
rect 6616 8732 6912 8752
rect 6672 8730 6696 8732
rect 6752 8730 6776 8732
rect 6832 8730 6856 8732
rect 6694 8678 6696 8730
rect 6758 8678 6770 8730
rect 6832 8678 6834 8730
rect 6672 8676 6696 8678
rect 6752 8676 6776 8678
rect 6832 8676 6856 8678
rect 6616 8656 6912 8676
rect 5354 8528 5410 8537
rect 5354 8463 5410 8472
rect 3220 8188 3516 8208
rect 3276 8186 3300 8188
rect 3356 8186 3380 8188
rect 3436 8186 3460 8188
rect 3298 8134 3300 8186
rect 3362 8134 3374 8186
rect 3436 8134 3438 8186
rect 3276 8132 3300 8134
rect 3356 8132 3380 8134
rect 3436 8132 3460 8134
rect 3220 8112 3516 8132
rect 4352 7644 4648 7664
rect 4408 7642 4432 7644
rect 4488 7642 4512 7644
rect 4568 7642 4592 7644
rect 4430 7590 4432 7642
rect 4494 7590 4506 7642
rect 4568 7590 4570 7642
rect 4408 7588 4432 7590
rect 4488 7588 4512 7590
rect 4568 7588 4592 7590
rect 4352 7568 4648 7588
rect 5368 7342 5396 8463
rect 5484 8188 5780 8208
rect 5540 8186 5564 8188
rect 5620 8186 5644 8188
rect 5700 8186 5724 8188
rect 5562 8134 5564 8186
rect 5626 8134 5638 8186
rect 5700 8134 5702 8186
rect 5540 8132 5564 8134
rect 5620 8132 5644 8134
rect 5700 8132 5724 8134
rect 5484 8112 5780 8132
rect 6616 7644 6912 7664
rect 6672 7642 6696 7644
rect 6752 7642 6776 7644
rect 6832 7642 6856 7644
rect 6694 7590 6696 7642
rect 6758 7590 6770 7642
rect 6832 7590 6834 7642
rect 6672 7588 6696 7590
rect 6752 7588 6776 7590
rect 6832 7588 6856 7590
rect 6616 7568 6912 7588
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 3220 7100 3516 7120
rect 3276 7098 3300 7100
rect 3356 7098 3380 7100
rect 3436 7098 3460 7100
rect 3298 7046 3300 7098
rect 3362 7046 3374 7098
rect 3436 7046 3438 7098
rect 3276 7044 3300 7046
rect 3356 7044 3380 7046
rect 3436 7044 3460 7046
rect 3220 7024 3516 7044
rect 4352 6556 4648 6576
rect 4408 6554 4432 6556
rect 4488 6554 4512 6556
rect 4568 6554 4592 6556
rect 4430 6502 4432 6554
rect 4494 6502 4506 6554
rect 4568 6502 4570 6554
rect 4408 6500 4432 6502
rect 4488 6500 4512 6502
rect 4568 6500 4592 6502
rect 4352 6480 4648 6500
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2088 5468 2384 5488
rect 2144 5466 2168 5468
rect 2224 5466 2248 5468
rect 2304 5466 2328 5468
rect 2166 5414 2168 5466
rect 2230 5414 2242 5466
rect 2304 5414 2306 5466
rect 2144 5412 2168 5414
rect 2224 5412 2248 5414
rect 2304 5412 2328 5414
rect 2088 5392 2384 5412
rect 2088 4380 2384 4400
rect 2144 4378 2168 4380
rect 2224 4378 2248 4380
rect 2304 4378 2328 4380
rect 2166 4326 2168 4378
rect 2230 4326 2242 4378
rect 2304 4326 2306 4378
rect 2144 4324 2168 4326
rect 2224 4324 2248 4326
rect 2304 4324 2328 4326
rect 2088 4304 2384 4324
rect 2976 3942 3004 6190
rect 5368 6186 5396 7278
rect 5484 7100 5780 7120
rect 5540 7098 5564 7100
rect 5620 7098 5644 7100
rect 5700 7098 5724 7100
rect 5562 7046 5564 7098
rect 5626 7046 5638 7098
rect 5700 7046 5702 7098
rect 5540 7044 5564 7046
rect 5620 7044 5644 7046
rect 5700 7044 5724 7046
rect 5484 7024 5780 7044
rect 6616 6556 6912 6576
rect 6672 6554 6696 6556
rect 6752 6554 6776 6556
rect 6832 6554 6856 6556
rect 6694 6502 6696 6554
rect 6758 6502 6770 6554
rect 6832 6502 6834 6554
rect 6672 6500 6696 6502
rect 6752 6500 6776 6502
rect 6832 6500 6856 6502
rect 6616 6480 6912 6500
rect 5356 6180 5408 6186
rect 5356 6122 5408 6128
rect 3220 6012 3516 6032
rect 3276 6010 3300 6012
rect 3356 6010 3380 6012
rect 3436 6010 3460 6012
rect 3298 5958 3300 6010
rect 3362 5958 3374 6010
rect 3436 5958 3438 6010
rect 3276 5956 3300 5958
rect 3356 5956 3380 5958
rect 3436 5956 3460 5958
rect 3220 5936 3516 5956
rect 5368 5846 5396 6122
rect 5484 6012 5780 6032
rect 5540 6010 5564 6012
rect 5620 6010 5644 6012
rect 5700 6010 5724 6012
rect 5562 5958 5564 6010
rect 5626 5958 5638 6010
rect 5700 5958 5702 6010
rect 5540 5956 5564 5958
rect 5620 5956 5644 5958
rect 5700 5956 5724 5958
rect 5484 5936 5780 5956
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 4066 5128 4122 5137
rect 4172 5114 4200 5646
rect 4352 5468 4648 5488
rect 4408 5466 4432 5468
rect 4488 5466 4512 5468
rect 4568 5466 4592 5468
rect 4430 5414 4432 5466
rect 4494 5414 4506 5466
rect 4568 5414 4570 5466
rect 4408 5412 4432 5414
rect 4488 5412 4512 5414
rect 4568 5412 4592 5414
rect 4352 5392 4648 5412
rect 6616 5468 6912 5488
rect 6672 5466 6696 5468
rect 6752 5466 6776 5468
rect 6832 5466 6856 5468
rect 6694 5414 6696 5466
rect 6758 5414 6770 5466
rect 6832 5414 6834 5466
rect 6672 5412 6696 5414
rect 6752 5412 6776 5414
rect 6832 5412 6856 5414
rect 6616 5392 6912 5412
rect 4122 5086 4200 5114
rect 4066 5063 4122 5072
rect 3220 4924 3516 4944
rect 3276 4922 3300 4924
rect 3356 4922 3380 4924
rect 3436 4922 3460 4924
rect 3298 4870 3300 4922
rect 3362 4870 3374 4922
rect 3436 4870 3438 4922
rect 3276 4868 3300 4870
rect 3356 4868 3380 4870
rect 3436 4868 3460 4870
rect 3220 4848 3516 4868
rect 5484 4924 5780 4944
rect 5540 4922 5564 4924
rect 5620 4922 5644 4924
rect 5700 4922 5724 4924
rect 5562 4870 5564 4922
rect 5626 4870 5638 4922
rect 5700 4870 5702 4922
rect 5540 4868 5564 4870
rect 5620 4868 5644 4870
rect 5700 4868 5724 4870
rect 5484 4848 5780 4868
rect 4352 4380 4648 4400
rect 4408 4378 4432 4380
rect 4488 4378 4512 4380
rect 4568 4378 4592 4380
rect 4430 4326 4432 4378
rect 4494 4326 4506 4378
rect 4568 4326 4570 4378
rect 4408 4324 4432 4326
rect 4488 4324 4512 4326
rect 4568 4324 4592 4326
rect 4352 4304 4648 4324
rect 6616 4380 6912 4400
rect 6672 4378 6696 4380
rect 6752 4378 6776 4380
rect 6832 4378 6856 4380
rect 6694 4326 6696 4378
rect 6758 4326 6770 4378
rect 6832 4326 6834 4378
rect 6672 4324 6696 4326
rect 6752 4324 6776 4326
rect 6832 4324 6856 4326
rect 6616 4304 6912 4324
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2088 3292 2384 3312
rect 2144 3290 2168 3292
rect 2224 3290 2248 3292
rect 2304 3290 2328 3292
rect 2166 3238 2168 3290
rect 2230 3238 2242 3290
rect 2304 3238 2306 3290
rect 2144 3236 2168 3238
rect 2224 3236 2248 3238
rect 2304 3236 2328 3238
rect 2088 3216 2384 3236
rect 2088 2204 2384 2224
rect 2144 2202 2168 2204
rect 2224 2202 2248 2204
rect 2304 2202 2328 2204
rect 2166 2150 2168 2202
rect 2230 2150 2242 2202
rect 2304 2150 2306 2202
rect 2144 2148 2168 2150
rect 2224 2148 2248 2150
rect 2304 2148 2328 2150
rect 2088 2128 2384 2148
rect 3160 1986 3188 3946
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 3220 3836 3516 3856
rect 3276 3834 3300 3836
rect 3356 3834 3380 3836
rect 3436 3834 3460 3836
rect 3298 3782 3300 3834
rect 3362 3782 3374 3834
rect 3436 3782 3438 3834
rect 3276 3780 3300 3782
rect 3356 3780 3380 3782
rect 3436 3780 3460 3782
rect 3220 3760 3516 3780
rect 5484 3836 5780 3856
rect 5540 3834 5564 3836
rect 5620 3834 5644 3836
rect 5700 3834 5724 3836
rect 5562 3782 5564 3834
rect 5626 3782 5638 3834
rect 5700 3782 5702 3834
rect 5540 3780 5564 3782
rect 5620 3780 5644 3782
rect 5700 3780 5724 3782
rect 5484 3760 5780 3780
rect 4352 3292 4648 3312
rect 4408 3290 4432 3292
rect 4488 3290 4512 3292
rect 4568 3290 4592 3292
rect 4430 3238 4432 3290
rect 4494 3238 4506 3290
rect 4568 3238 4570 3290
rect 4408 3236 4432 3238
rect 4488 3236 4512 3238
rect 4568 3236 4592 3238
rect 4352 3216 4648 3236
rect 3220 2748 3516 2768
rect 3276 2746 3300 2748
rect 3356 2746 3380 2748
rect 3436 2746 3460 2748
rect 3298 2694 3300 2746
rect 3362 2694 3374 2746
rect 3436 2694 3438 2746
rect 3276 2692 3300 2694
rect 3356 2692 3380 2694
rect 3436 2692 3460 2694
rect 3220 2672 3516 2692
rect 5484 2748 5780 2768
rect 5540 2746 5564 2748
rect 5620 2746 5644 2748
rect 5700 2746 5724 2748
rect 5562 2694 5564 2746
rect 5626 2694 5638 2746
rect 5700 2694 5702 2746
rect 5540 2692 5564 2694
rect 5620 2692 5644 2694
rect 5700 2692 5724 2694
rect 5484 2672 5780 2692
rect 5828 2530 5856 3878
rect 6616 3292 6912 3312
rect 6672 3290 6696 3292
rect 6752 3290 6776 3292
rect 6832 3290 6856 3292
rect 6694 3238 6696 3290
rect 6758 3238 6770 3290
rect 6832 3238 6834 3290
rect 6672 3236 6696 3238
rect 6752 3236 6776 3238
rect 6832 3236 6856 3238
rect 6616 3216 6912 3236
rect 5644 2502 5856 2530
rect 4352 2204 4648 2224
rect 4408 2202 4432 2204
rect 4488 2202 4512 2204
rect 4568 2202 4592 2204
rect 4430 2150 4432 2202
rect 4494 2150 4506 2202
rect 4568 2150 4570 2202
rect 4408 2148 4432 2150
rect 4488 2148 4512 2150
rect 4568 2148 4592 2150
rect 4352 2128 4648 2148
rect 3160 1958 3372 1986
rect 1950 1728 2006 1737
rect 1950 1663 2006 1672
rect 3344 480 3372 1958
rect 5644 480 5672 2502
rect 6616 2204 6912 2224
rect 6672 2202 6696 2204
rect 6752 2202 6776 2204
rect 6832 2202 6856 2204
rect 6694 2150 6696 2202
rect 6758 2150 6770 2202
rect 6832 2150 6834 2202
rect 6672 2148 6696 2150
rect 6752 2148 6776 2150
rect 6832 2148 6856 2150
rect 6616 2128 6912 2148
rect 7852 480 7880 5646
rect 1122 0 1178 480
rect 3330 0 3386 480
rect 5630 0 5686 480
rect 7838 0 7894 480
<< via2 >>
rect 2778 15272 2834 15328
rect 2088 14170 2144 14172
rect 2168 14170 2224 14172
rect 2248 14170 2304 14172
rect 2328 14170 2384 14172
rect 2088 14118 2114 14170
rect 2114 14118 2144 14170
rect 2168 14118 2178 14170
rect 2178 14118 2224 14170
rect 2248 14118 2294 14170
rect 2294 14118 2304 14170
rect 2328 14118 2358 14170
rect 2358 14118 2384 14170
rect 2088 14116 2144 14118
rect 2168 14116 2224 14118
rect 2248 14116 2304 14118
rect 2328 14116 2384 14118
rect 2088 13082 2144 13084
rect 2168 13082 2224 13084
rect 2248 13082 2304 13084
rect 2328 13082 2384 13084
rect 2088 13030 2114 13082
rect 2114 13030 2144 13082
rect 2168 13030 2178 13082
rect 2178 13030 2224 13082
rect 2248 13030 2294 13082
rect 2294 13030 2304 13082
rect 2328 13030 2358 13082
rect 2358 13030 2384 13082
rect 2088 13028 2144 13030
rect 2168 13028 2224 13030
rect 2248 13028 2304 13030
rect 2328 13028 2384 13030
rect 2088 11994 2144 11996
rect 2168 11994 2224 11996
rect 2248 11994 2304 11996
rect 2328 11994 2384 11996
rect 2088 11942 2114 11994
rect 2114 11942 2144 11994
rect 2168 11942 2178 11994
rect 2178 11942 2224 11994
rect 2248 11942 2294 11994
rect 2294 11942 2304 11994
rect 2328 11942 2358 11994
rect 2358 11942 2384 11994
rect 2088 11940 2144 11942
rect 2168 11940 2224 11942
rect 2248 11940 2304 11942
rect 2328 11940 2384 11942
rect 2088 10906 2144 10908
rect 2168 10906 2224 10908
rect 2248 10906 2304 10908
rect 2328 10906 2384 10908
rect 2088 10854 2114 10906
rect 2114 10854 2144 10906
rect 2168 10854 2178 10906
rect 2178 10854 2224 10906
rect 2248 10854 2294 10906
rect 2294 10854 2304 10906
rect 2328 10854 2358 10906
rect 2358 10854 2384 10906
rect 2088 10852 2144 10854
rect 2168 10852 2224 10854
rect 2248 10852 2304 10854
rect 2328 10852 2384 10854
rect 2088 9818 2144 9820
rect 2168 9818 2224 9820
rect 2248 9818 2304 9820
rect 2328 9818 2384 9820
rect 2088 9766 2114 9818
rect 2114 9766 2144 9818
rect 2168 9766 2178 9818
rect 2178 9766 2224 9818
rect 2248 9766 2294 9818
rect 2294 9766 2304 9818
rect 2328 9766 2358 9818
rect 2358 9766 2384 9818
rect 2088 9764 2144 9766
rect 2168 9764 2224 9766
rect 2248 9764 2304 9766
rect 2328 9764 2384 9766
rect 2088 8730 2144 8732
rect 2168 8730 2224 8732
rect 2248 8730 2304 8732
rect 2328 8730 2384 8732
rect 2088 8678 2114 8730
rect 2114 8678 2144 8730
rect 2168 8678 2178 8730
rect 2178 8678 2224 8730
rect 2248 8678 2294 8730
rect 2294 8678 2304 8730
rect 2328 8678 2358 8730
rect 2358 8678 2384 8730
rect 2088 8676 2144 8678
rect 2168 8676 2224 8678
rect 2248 8676 2304 8678
rect 2328 8676 2384 8678
rect 2226 8472 2282 8528
rect 3220 14714 3276 14716
rect 3300 14714 3356 14716
rect 3380 14714 3436 14716
rect 3460 14714 3516 14716
rect 3220 14662 3246 14714
rect 3246 14662 3276 14714
rect 3300 14662 3310 14714
rect 3310 14662 3356 14714
rect 3380 14662 3426 14714
rect 3426 14662 3436 14714
rect 3460 14662 3490 14714
rect 3490 14662 3516 14714
rect 3220 14660 3276 14662
rect 3300 14660 3356 14662
rect 3380 14660 3436 14662
rect 3460 14660 3516 14662
rect 5484 14714 5540 14716
rect 5564 14714 5620 14716
rect 5644 14714 5700 14716
rect 5724 14714 5780 14716
rect 5484 14662 5510 14714
rect 5510 14662 5540 14714
rect 5564 14662 5574 14714
rect 5574 14662 5620 14714
rect 5644 14662 5690 14714
rect 5690 14662 5700 14714
rect 5724 14662 5754 14714
rect 5754 14662 5780 14714
rect 5484 14660 5540 14662
rect 5564 14660 5620 14662
rect 5644 14660 5700 14662
rect 5724 14660 5780 14662
rect 4352 14170 4408 14172
rect 4432 14170 4488 14172
rect 4512 14170 4568 14172
rect 4592 14170 4648 14172
rect 4352 14118 4378 14170
rect 4378 14118 4408 14170
rect 4432 14118 4442 14170
rect 4442 14118 4488 14170
rect 4512 14118 4558 14170
rect 4558 14118 4568 14170
rect 4592 14118 4622 14170
rect 4622 14118 4648 14170
rect 4352 14116 4408 14118
rect 4432 14116 4488 14118
rect 4512 14116 4568 14118
rect 4592 14116 4648 14118
rect 6616 14170 6672 14172
rect 6696 14170 6752 14172
rect 6776 14170 6832 14172
rect 6856 14170 6912 14172
rect 6616 14118 6642 14170
rect 6642 14118 6672 14170
rect 6696 14118 6706 14170
rect 6706 14118 6752 14170
rect 6776 14118 6822 14170
rect 6822 14118 6832 14170
rect 6856 14118 6886 14170
rect 6886 14118 6912 14170
rect 6616 14116 6672 14118
rect 6696 14116 6752 14118
rect 6776 14116 6832 14118
rect 6856 14116 6912 14118
rect 3220 13626 3276 13628
rect 3300 13626 3356 13628
rect 3380 13626 3436 13628
rect 3460 13626 3516 13628
rect 3220 13574 3246 13626
rect 3246 13574 3276 13626
rect 3300 13574 3310 13626
rect 3310 13574 3356 13626
rect 3380 13574 3426 13626
rect 3426 13574 3436 13626
rect 3460 13574 3490 13626
rect 3490 13574 3516 13626
rect 3220 13572 3276 13574
rect 3300 13572 3356 13574
rect 3380 13572 3436 13574
rect 3460 13572 3516 13574
rect 5484 13626 5540 13628
rect 5564 13626 5620 13628
rect 5644 13626 5700 13628
rect 5724 13626 5780 13628
rect 5484 13574 5510 13626
rect 5510 13574 5540 13626
rect 5564 13574 5574 13626
rect 5574 13574 5620 13626
rect 5644 13574 5690 13626
rect 5690 13574 5700 13626
rect 5724 13574 5754 13626
rect 5754 13574 5780 13626
rect 5484 13572 5540 13574
rect 5564 13572 5620 13574
rect 5644 13572 5700 13574
rect 5724 13572 5780 13574
rect 4352 13082 4408 13084
rect 4432 13082 4488 13084
rect 4512 13082 4568 13084
rect 4592 13082 4648 13084
rect 4352 13030 4378 13082
rect 4378 13030 4408 13082
rect 4432 13030 4442 13082
rect 4442 13030 4488 13082
rect 4512 13030 4558 13082
rect 4558 13030 4568 13082
rect 4592 13030 4622 13082
rect 4622 13030 4648 13082
rect 4352 13028 4408 13030
rect 4432 13028 4488 13030
rect 4512 13028 4568 13030
rect 4592 13028 4648 13030
rect 6616 13082 6672 13084
rect 6696 13082 6752 13084
rect 6776 13082 6832 13084
rect 6856 13082 6912 13084
rect 6616 13030 6642 13082
rect 6642 13030 6672 13082
rect 6696 13030 6706 13082
rect 6706 13030 6752 13082
rect 6776 13030 6822 13082
rect 6822 13030 6832 13082
rect 6856 13030 6886 13082
rect 6886 13030 6912 13082
rect 6616 13028 6672 13030
rect 6696 13028 6752 13030
rect 6776 13028 6832 13030
rect 6856 13028 6912 13030
rect 3220 12538 3276 12540
rect 3300 12538 3356 12540
rect 3380 12538 3436 12540
rect 3460 12538 3516 12540
rect 3220 12486 3246 12538
rect 3246 12486 3276 12538
rect 3300 12486 3310 12538
rect 3310 12486 3356 12538
rect 3380 12486 3426 12538
rect 3426 12486 3436 12538
rect 3460 12486 3490 12538
rect 3490 12486 3516 12538
rect 3220 12484 3276 12486
rect 3300 12484 3356 12486
rect 3380 12484 3436 12486
rect 3460 12484 3516 12486
rect 5484 12538 5540 12540
rect 5564 12538 5620 12540
rect 5644 12538 5700 12540
rect 5724 12538 5780 12540
rect 5484 12486 5510 12538
rect 5510 12486 5540 12538
rect 5564 12486 5574 12538
rect 5574 12486 5620 12538
rect 5644 12486 5690 12538
rect 5690 12486 5700 12538
rect 5724 12486 5754 12538
rect 5754 12486 5780 12538
rect 5484 12484 5540 12486
rect 5564 12484 5620 12486
rect 5644 12484 5700 12486
rect 5724 12484 5780 12486
rect 4352 11994 4408 11996
rect 4432 11994 4488 11996
rect 4512 11994 4568 11996
rect 4592 11994 4648 11996
rect 4352 11942 4378 11994
rect 4378 11942 4408 11994
rect 4432 11942 4442 11994
rect 4442 11942 4488 11994
rect 4512 11942 4558 11994
rect 4558 11942 4568 11994
rect 4592 11942 4622 11994
rect 4622 11942 4648 11994
rect 4352 11940 4408 11942
rect 4432 11940 4488 11942
rect 4512 11940 4568 11942
rect 4592 11940 4648 11942
rect 6616 11994 6672 11996
rect 6696 11994 6752 11996
rect 6776 11994 6832 11996
rect 6856 11994 6912 11996
rect 6616 11942 6642 11994
rect 6642 11942 6672 11994
rect 6696 11942 6706 11994
rect 6706 11942 6752 11994
rect 6776 11942 6822 11994
rect 6822 11942 6832 11994
rect 6856 11942 6886 11994
rect 6886 11942 6912 11994
rect 6616 11940 6672 11942
rect 6696 11940 6752 11942
rect 6776 11940 6832 11942
rect 6856 11940 6912 11942
rect 2870 11736 2926 11792
rect 2088 7642 2144 7644
rect 2168 7642 2224 7644
rect 2248 7642 2304 7644
rect 2328 7642 2384 7644
rect 2088 7590 2114 7642
rect 2114 7590 2144 7642
rect 2168 7590 2178 7642
rect 2178 7590 2224 7642
rect 2248 7590 2294 7642
rect 2294 7590 2304 7642
rect 2328 7590 2358 7642
rect 2358 7590 2384 7642
rect 2088 7588 2144 7590
rect 2168 7588 2224 7590
rect 2248 7588 2304 7590
rect 2328 7588 2384 7590
rect 2088 6554 2144 6556
rect 2168 6554 2224 6556
rect 2248 6554 2304 6556
rect 2328 6554 2384 6556
rect 2088 6502 2114 6554
rect 2114 6502 2144 6554
rect 2168 6502 2178 6554
rect 2178 6502 2224 6554
rect 2248 6502 2294 6554
rect 2294 6502 2304 6554
rect 2328 6502 2358 6554
rect 2358 6502 2384 6554
rect 2088 6500 2144 6502
rect 2168 6500 2224 6502
rect 2248 6500 2304 6502
rect 2328 6500 2384 6502
rect 3220 11450 3276 11452
rect 3300 11450 3356 11452
rect 3380 11450 3436 11452
rect 3460 11450 3516 11452
rect 3220 11398 3246 11450
rect 3246 11398 3276 11450
rect 3300 11398 3310 11450
rect 3310 11398 3356 11450
rect 3380 11398 3426 11450
rect 3426 11398 3436 11450
rect 3460 11398 3490 11450
rect 3490 11398 3516 11450
rect 3220 11396 3276 11398
rect 3300 11396 3356 11398
rect 3380 11396 3436 11398
rect 3460 11396 3516 11398
rect 5484 11450 5540 11452
rect 5564 11450 5620 11452
rect 5644 11450 5700 11452
rect 5724 11450 5780 11452
rect 5484 11398 5510 11450
rect 5510 11398 5540 11450
rect 5564 11398 5574 11450
rect 5574 11398 5620 11450
rect 5644 11398 5690 11450
rect 5690 11398 5700 11450
rect 5724 11398 5754 11450
rect 5754 11398 5780 11450
rect 5484 11396 5540 11398
rect 5564 11396 5620 11398
rect 5644 11396 5700 11398
rect 5724 11396 5780 11398
rect 4352 10906 4408 10908
rect 4432 10906 4488 10908
rect 4512 10906 4568 10908
rect 4592 10906 4648 10908
rect 4352 10854 4378 10906
rect 4378 10854 4408 10906
rect 4432 10854 4442 10906
rect 4442 10854 4488 10906
rect 4512 10854 4558 10906
rect 4558 10854 4568 10906
rect 4592 10854 4622 10906
rect 4622 10854 4648 10906
rect 4352 10852 4408 10854
rect 4432 10852 4488 10854
rect 4512 10852 4568 10854
rect 4592 10852 4648 10854
rect 6616 10906 6672 10908
rect 6696 10906 6752 10908
rect 6776 10906 6832 10908
rect 6856 10906 6912 10908
rect 6616 10854 6642 10906
rect 6642 10854 6672 10906
rect 6696 10854 6706 10906
rect 6706 10854 6752 10906
rect 6776 10854 6822 10906
rect 6822 10854 6832 10906
rect 6856 10854 6886 10906
rect 6886 10854 6912 10906
rect 6616 10852 6672 10854
rect 6696 10852 6752 10854
rect 6776 10852 6832 10854
rect 6856 10852 6912 10854
rect 3220 10362 3276 10364
rect 3300 10362 3356 10364
rect 3380 10362 3436 10364
rect 3460 10362 3516 10364
rect 3220 10310 3246 10362
rect 3246 10310 3276 10362
rect 3300 10310 3310 10362
rect 3310 10310 3356 10362
rect 3380 10310 3426 10362
rect 3426 10310 3436 10362
rect 3460 10310 3490 10362
rect 3490 10310 3516 10362
rect 3220 10308 3276 10310
rect 3300 10308 3356 10310
rect 3380 10308 3436 10310
rect 3460 10308 3516 10310
rect 5484 10362 5540 10364
rect 5564 10362 5620 10364
rect 5644 10362 5700 10364
rect 5724 10362 5780 10364
rect 5484 10310 5510 10362
rect 5510 10310 5540 10362
rect 5564 10310 5574 10362
rect 5574 10310 5620 10362
rect 5644 10310 5690 10362
rect 5690 10310 5700 10362
rect 5724 10310 5754 10362
rect 5754 10310 5780 10362
rect 5484 10308 5540 10310
rect 5564 10308 5620 10310
rect 5644 10308 5700 10310
rect 5724 10308 5780 10310
rect 4352 9818 4408 9820
rect 4432 9818 4488 9820
rect 4512 9818 4568 9820
rect 4592 9818 4648 9820
rect 4352 9766 4378 9818
rect 4378 9766 4408 9818
rect 4432 9766 4442 9818
rect 4442 9766 4488 9818
rect 4512 9766 4558 9818
rect 4558 9766 4568 9818
rect 4592 9766 4622 9818
rect 4622 9766 4648 9818
rect 4352 9764 4408 9766
rect 4432 9764 4488 9766
rect 4512 9764 4568 9766
rect 4592 9764 4648 9766
rect 6616 9818 6672 9820
rect 6696 9818 6752 9820
rect 6776 9818 6832 9820
rect 6856 9818 6912 9820
rect 6616 9766 6642 9818
rect 6642 9766 6672 9818
rect 6696 9766 6706 9818
rect 6706 9766 6752 9818
rect 6776 9766 6822 9818
rect 6822 9766 6832 9818
rect 6856 9766 6886 9818
rect 6886 9766 6912 9818
rect 6616 9764 6672 9766
rect 6696 9764 6752 9766
rect 6776 9764 6832 9766
rect 6856 9764 6912 9766
rect 3220 9274 3276 9276
rect 3300 9274 3356 9276
rect 3380 9274 3436 9276
rect 3460 9274 3516 9276
rect 3220 9222 3246 9274
rect 3246 9222 3276 9274
rect 3300 9222 3310 9274
rect 3310 9222 3356 9274
rect 3380 9222 3426 9274
rect 3426 9222 3436 9274
rect 3460 9222 3490 9274
rect 3490 9222 3516 9274
rect 3220 9220 3276 9222
rect 3300 9220 3356 9222
rect 3380 9220 3436 9222
rect 3460 9220 3516 9222
rect 5484 9274 5540 9276
rect 5564 9274 5620 9276
rect 5644 9274 5700 9276
rect 5724 9274 5780 9276
rect 5484 9222 5510 9274
rect 5510 9222 5540 9274
rect 5564 9222 5574 9274
rect 5574 9222 5620 9274
rect 5644 9222 5690 9274
rect 5690 9222 5700 9274
rect 5724 9222 5754 9274
rect 5754 9222 5780 9274
rect 5484 9220 5540 9222
rect 5564 9220 5620 9222
rect 5644 9220 5700 9222
rect 5724 9220 5780 9222
rect 4352 8730 4408 8732
rect 4432 8730 4488 8732
rect 4512 8730 4568 8732
rect 4592 8730 4648 8732
rect 4352 8678 4378 8730
rect 4378 8678 4408 8730
rect 4432 8678 4442 8730
rect 4442 8678 4488 8730
rect 4512 8678 4558 8730
rect 4558 8678 4568 8730
rect 4592 8678 4622 8730
rect 4622 8678 4648 8730
rect 4352 8676 4408 8678
rect 4432 8676 4488 8678
rect 4512 8676 4568 8678
rect 4592 8676 4648 8678
rect 6616 8730 6672 8732
rect 6696 8730 6752 8732
rect 6776 8730 6832 8732
rect 6856 8730 6912 8732
rect 6616 8678 6642 8730
rect 6642 8678 6672 8730
rect 6696 8678 6706 8730
rect 6706 8678 6752 8730
rect 6776 8678 6822 8730
rect 6822 8678 6832 8730
rect 6856 8678 6886 8730
rect 6886 8678 6912 8730
rect 6616 8676 6672 8678
rect 6696 8676 6752 8678
rect 6776 8676 6832 8678
rect 6856 8676 6912 8678
rect 5354 8472 5410 8528
rect 3220 8186 3276 8188
rect 3300 8186 3356 8188
rect 3380 8186 3436 8188
rect 3460 8186 3516 8188
rect 3220 8134 3246 8186
rect 3246 8134 3276 8186
rect 3300 8134 3310 8186
rect 3310 8134 3356 8186
rect 3380 8134 3426 8186
rect 3426 8134 3436 8186
rect 3460 8134 3490 8186
rect 3490 8134 3516 8186
rect 3220 8132 3276 8134
rect 3300 8132 3356 8134
rect 3380 8132 3436 8134
rect 3460 8132 3516 8134
rect 4352 7642 4408 7644
rect 4432 7642 4488 7644
rect 4512 7642 4568 7644
rect 4592 7642 4648 7644
rect 4352 7590 4378 7642
rect 4378 7590 4408 7642
rect 4432 7590 4442 7642
rect 4442 7590 4488 7642
rect 4512 7590 4558 7642
rect 4558 7590 4568 7642
rect 4592 7590 4622 7642
rect 4622 7590 4648 7642
rect 4352 7588 4408 7590
rect 4432 7588 4488 7590
rect 4512 7588 4568 7590
rect 4592 7588 4648 7590
rect 5484 8186 5540 8188
rect 5564 8186 5620 8188
rect 5644 8186 5700 8188
rect 5724 8186 5780 8188
rect 5484 8134 5510 8186
rect 5510 8134 5540 8186
rect 5564 8134 5574 8186
rect 5574 8134 5620 8186
rect 5644 8134 5690 8186
rect 5690 8134 5700 8186
rect 5724 8134 5754 8186
rect 5754 8134 5780 8186
rect 5484 8132 5540 8134
rect 5564 8132 5620 8134
rect 5644 8132 5700 8134
rect 5724 8132 5780 8134
rect 6616 7642 6672 7644
rect 6696 7642 6752 7644
rect 6776 7642 6832 7644
rect 6856 7642 6912 7644
rect 6616 7590 6642 7642
rect 6642 7590 6672 7642
rect 6696 7590 6706 7642
rect 6706 7590 6752 7642
rect 6776 7590 6822 7642
rect 6822 7590 6832 7642
rect 6856 7590 6886 7642
rect 6886 7590 6912 7642
rect 6616 7588 6672 7590
rect 6696 7588 6752 7590
rect 6776 7588 6832 7590
rect 6856 7588 6912 7590
rect 3220 7098 3276 7100
rect 3300 7098 3356 7100
rect 3380 7098 3436 7100
rect 3460 7098 3516 7100
rect 3220 7046 3246 7098
rect 3246 7046 3276 7098
rect 3300 7046 3310 7098
rect 3310 7046 3356 7098
rect 3380 7046 3426 7098
rect 3426 7046 3436 7098
rect 3460 7046 3490 7098
rect 3490 7046 3516 7098
rect 3220 7044 3276 7046
rect 3300 7044 3356 7046
rect 3380 7044 3436 7046
rect 3460 7044 3516 7046
rect 4352 6554 4408 6556
rect 4432 6554 4488 6556
rect 4512 6554 4568 6556
rect 4592 6554 4648 6556
rect 4352 6502 4378 6554
rect 4378 6502 4408 6554
rect 4432 6502 4442 6554
rect 4442 6502 4488 6554
rect 4512 6502 4558 6554
rect 4558 6502 4568 6554
rect 4592 6502 4622 6554
rect 4622 6502 4648 6554
rect 4352 6500 4408 6502
rect 4432 6500 4488 6502
rect 4512 6500 4568 6502
rect 4592 6500 4648 6502
rect 2088 5466 2144 5468
rect 2168 5466 2224 5468
rect 2248 5466 2304 5468
rect 2328 5466 2384 5468
rect 2088 5414 2114 5466
rect 2114 5414 2144 5466
rect 2168 5414 2178 5466
rect 2178 5414 2224 5466
rect 2248 5414 2294 5466
rect 2294 5414 2304 5466
rect 2328 5414 2358 5466
rect 2358 5414 2384 5466
rect 2088 5412 2144 5414
rect 2168 5412 2224 5414
rect 2248 5412 2304 5414
rect 2328 5412 2384 5414
rect 2088 4378 2144 4380
rect 2168 4378 2224 4380
rect 2248 4378 2304 4380
rect 2328 4378 2384 4380
rect 2088 4326 2114 4378
rect 2114 4326 2144 4378
rect 2168 4326 2178 4378
rect 2178 4326 2224 4378
rect 2248 4326 2294 4378
rect 2294 4326 2304 4378
rect 2328 4326 2358 4378
rect 2358 4326 2384 4378
rect 2088 4324 2144 4326
rect 2168 4324 2224 4326
rect 2248 4324 2304 4326
rect 2328 4324 2384 4326
rect 5484 7098 5540 7100
rect 5564 7098 5620 7100
rect 5644 7098 5700 7100
rect 5724 7098 5780 7100
rect 5484 7046 5510 7098
rect 5510 7046 5540 7098
rect 5564 7046 5574 7098
rect 5574 7046 5620 7098
rect 5644 7046 5690 7098
rect 5690 7046 5700 7098
rect 5724 7046 5754 7098
rect 5754 7046 5780 7098
rect 5484 7044 5540 7046
rect 5564 7044 5620 7046
rect 5644 7044 5700 7046
rect 5724 7044 5780 7046
rect 6616 6554 6672 6556
rect 6696 6554 6752 6556
rect 6776 6554 6832 6556
rect 6856 6554 6912 6556
rect 6616 6502 6642 6554
rect 6642 6502 6672 6554
rect 6696 6502 6706 6554
rect 6706 6502 6752 6554
rect 6776 6502 6822 6554
rect 6822 6502 6832 6554
rect 6856 6502 6886 6554
rect 6886 6502 6912 6554
rect 6616 6500 6672 6502
rect 6696 6500 6752 6502
rect 6776 6500 6832 6502
rect 6856 6500 6912 6502
rect 3220 6010 3276 6012
rect 3300 6010 3356 6012
rect 3380 6010 3436 6012
rect 3460 6010 3516 6012
rect 3220 5958 3246 6010
rect 3246 5958 3276 6010
rect 3300 5958 3310 6010
rect 3310 5958 3356 6010
rect 3380 5958 3426 6010
rect 3426 5958 3436 6010
rect 3460 5958 3490 6010
rect 3490 5958 3516 6010
rect 3220 5956 3276 5958
rect 3300 5956 3356 5958
rect 3380 5956 3436 5958
rect 3460 5956 3516 5958
rect 5484 6010 5540 6012
rect 5564 6010 5620 6012
rect 5644 6010 5700 6012
rect 5724 6010 5780 6012
rect 5484 5958 5510 6010
rect 5510 5958 5540 6010
rect 5564 5958 5574 6010
rect 5574 5958 5620 6010
rect 5644 5958 5690 6010
rect 5690 5958 5700 6010
rect 5724 5958 5754 6010
rect 5754 5958 5780 6010
rect 5484 5956 5540 5958
rect 5564 5956 5620 5958
rect 5644 5956 5700 5958
rect 5724 5956 5780 5958
rect 4066 5072 4122 5128
rect 4352 5466 4408 5468
rect 4432 5466 4488 5468
rect 4512 5466 4568 5468
rect 4592 5466 4648 5468
rect 4352 5414 4378 5466
rect 4378 5414 4408 5466
rect 4432 5414 4442 5466
rect 4442 5414 4488 5466
rect 4512 5414 4558 5466
rect 4558 5414 4568 5466
rect 4592 5414 4622 5466
rect 4622 5414 4648 5466
rect 4352 5412 4408 5414
rect 4432 5412 4488 5414
rect 4512 5412 4568 5414
rect 4592 5412 4648 5414
rect 6616 5466 6672 5468
rect 6696 5466 6752 5468
rect 6776 5466 6832 5468
rect 6856 5466 6912 5468
rect 6616 5414 6642 5466
rect 6642 5414 6672 5466
rect 6696 5414 6706 5466
rect 6706 5414 6752 5466
rect 6776 5414 6822 5466
rect 6822 5414 6832 5466
rect 6856 5414 6886 5466
rect 6886 5414 6912 5466
rect 6616 5412 6672 5414
rect 6696 5412 6752 5414
rect 6776 5412 6832 5414
rect 6856 5412 6912 5414
rect 3220 4922 3276 4924
rect 3300 4922 3356 4924
rect 3380 4922 3436 4924
rect 3460 4922 3516 4924
rect 3220 4870 3246 4922
rect 3246 4870 3276 4922
rect 3300 4870 3310 4922
rect 3310 4870 3356 4922
rect 3380 4870 3426 4922
rect 3426 4870 3436 4922
rect 3460 4870 3490 4922
rect 3490 4870 3516 4922
rect 3220 4868 3276 4870
rect 3300 4868 3356 4870
rect 3380 4868 3436 4870
rect 3460 4868 3516 4870
rect 5484 4922 5540 4924
rect 5564 4922 5620 4924
rect 5644 4922 5700 4924
rect 5724 4922 5780 4924
rect 5484 4870 5510 4922
rect 5510 4870 5540 4922
rect 5564 4870 5574 4922
rect 5574 4870 5620 4922
rect 5644 4870 5690 4922
rect 5690 4870 5700 4922
rect 5724 4870 5754 4922
rect 5754 4870 5780 4922
rect 5484 4868 5540 4870
rect 5564 4868 5620 4870
rect 5644 4868 5700 4870
rect 5724 4868 5780 4870
rect 4352 4378 4408 4380
rect 4432 4378 4488 4380
rect 4512 4378 4568 4380
rect 4592 4378 4648 4380
rect 4352 4326 4378 4378
rect 4378 4326 4408 4378
rect 4432 4326 4442 4378
rect 4442 4326 4488 4378
rect 4512 4326 4558 4378
rect 4558 4326 4568 4378
rect 4592 4326 4622 4378
rect 4622 4326 4648 4378
rect 4352 4324 4408 4326
rect 4432 4324 4488 4326
rect 4512 4324 4568 4326
rect 4592 4324 4648 4326
rect 6616 4378 6672 4380
rect 6696 4378 6752 4380
rect 6776 4378 6832 4380
rect 6856 4378 6912 4380
rect 6616 4326 6642 4378
rect 6642 4326 6672 4378
rect 6696 4326 6706 4378
rect 6706 4326 6752 4378
rect 6776 4326 6822 4378
rect 6822 4326 6832 4378
rect 6856 4326 6886 4378
rect 6886 4326 6912 4378
rect 6616 4324 6672 4326
rect 6696 4324 6752 4326
rect 6776 4324 6832 4326
rect 6856 4324 6912 4326
rect 2088 3290 2144 3292
rect 2168 3290 2224 3292
rect 2248 3290 2304 3292
rect 2328 3290 2384 3292
rect 2088 3238 2114 3290
rect 2114 3238 2144 3290
rect 2168 3238 2178 3290
rect 2178 3238 2224 3290
rect 2248 3238 2294 3290
rect 2294 3238 2304 3290
rect 2328 3238 2358 3290
rect 2358 3238 2384 3290
rect 2088 3236 2144 3238
rect 2168 3236 2224 3238
rect 2248 3236 2304 3238
rect 2328 3236 2384 3238
rect 2088 2202 2144 2204
rect 2168 2202 2224 2204
rect 2248 2202 2304 2204
rect 2328 2202 2384 2204
rect 2088 2150 2114 2202
rect 2114 2150 2144 2202
rect 2168 2150 2178 2202
rect 2178 2150 2224 2202
rect 2248 2150 2294 2202
rect 2294 2150 2304 2202
rect 2328 2150 2358 2202
rect 2358 2150 2384 2202
rect 2088 2148 2144 2150
rect 2168 2148 2224 2150
rect 2248 2148 2304 2150
rect 2328 2148 2384 2150
rect 3220 3834 3276 3836
rect 3300 3834 3356 3836
rect 3380 3834 3436 3836
rect 3460 3834 3516 3836
rect 3220 3782 3246 3834
rect 3246 3782 3276 3834
rect 3300 3782 3310 3834
rect 3310 3782 3356 3834
rect 3380 3782 3426 3834
rect 3426 3782 3436 3834
rect 3460 3782 3490 3834
rect 3490 3782 3516 3834
rect 3220 3780 3276 3782
rect 3300 3780 3356 3782
rect 3380 3780 3436 3782
rect 3460 3780 3516 3782
rect 5484 3834 5540 3836
rect 5564 3834 5620 3836
rect 5644 3834 5700 3836
rect 5724 3834 5780 3836
rect 5484 3782 5510 3834
rect 5510 3782 5540 3834
rect 5564 3782 5574 3834
rect 5574 3782 5620 3834
rect 5644 3782 5690 3834
rect 5690 3782 5700 3834
rect 5724 3782 5754 3834
rect 5754 3782 5780 3834
rect 5484 3780 5540 3782
rect 5564 3780 5620 3782
rect 5644 3780 5700 3782
rect 5724 3780 5780 3782
rect 4352 3290 4408 3292
rect 4432 3290 4488 3292
rect 4512 3290 4568 3292
rect 4592 3290 4648 3292
rect 4352 3238 4378 3290
rect 4378 3238 4408 3290
rect 4432 3238 4442 3290
rect 4442 3238 4488 3290
rect 4512 3238 4558 3290
rect 4558 3238 4568 3290
rect 4592 3238 4622 3290
rect 4622 3238 4648 3290
rect 4352 3236 4408 3238
rect 4432 3236 4488 3238
rect 4512 3236 4568 3238
rect 4592 3236 4648 3238
rect 3220 2746 3276 2748
rect 3300 2746 3356 2748
rect 3380 2746 3436 2748
rect 3460 2746 3516 2748
rect 3220 2694 3246 2746
rect 3246 2694 3276 2746
rect 3300 2694 3310 2746
rect 3310 2694 3356 2746
rect 3380 2694 3426 2746
rect 3426 2694 3436 2746
rect 3460 2694 3490 2746
rect 3490 2694 3516 2746
rect 3220 2692 3276 2694
rect 3300 2692 3356 2694
rect 3380 2692 3436 2694
rect 3460 2692 3516 2694
rect 5484 2746 5540 2748
rect 5564 2746 5620 2748
rect 5644 2746 5700 2748
rect 5724 2746 5780 2748
rect 5484 2694 5510 2746
rect 5510 2694 5540 2746
rect 5564 2694 5574 2746
rect 5574 2694 5620 2746
rect 5644 2694 5690 2746
rect 5690 2694 5700 2746
rect 5724 2694 5754 2746
rect 5754 2694 5780 2746
rect 5484 2692 5540 2694
rect 5564 2692 5620 2694
rect 5644 2692 5700 2694
rect 5724 2692 5780 2694
rect 6616 3290 6672 3292
rect 6696 3290 6752 3292
rect 6776 3290 6832 3292
rect 6856 3290 6912 3292
rect 6616 3238 6642 3290
rect 6642 3238 6672 3290
rect 6696 3238 6706 3290
rect 6706 3238 6752 3290
rect 6776 3238 6822 3290
rect 6822 3238 6832 3290
rect 6856 3238 6886 3290
rect 6886 3238 6912 3290
rect 6616 3236 6672 3238
rect 6696 3236 6752 3238
rect 6776 3236 6832 3238
rect 6856 3236 6912 3238
rect 4352 2202 4408 2204
rect 4432 2202 4488 2204
rect 4512 2202 4568 2204
rect 4592 2202 4648 2204
rect 4352 2150 4378 2202
rect 4378 2150 4408 2202
rect 4432 2150 4442 2202
rect 4442 2150 4488 2202
rect 4512 2150 4558 2202
rect 4558 2150 4568 2202
rect 4592 2150 4622 2202
rect 4622 2150 4648 2202
rect 4352 2148 4408 2150
rect 4432 2148 4488 2150
rect 4512 2148 4568 2150
rect 4592 2148 4648 2150
rect 1950 1672 2006 1728
rect 6616 2202 6672 2204
rect 6696 2202 6752 2204
rect 6776 2202 6832 2204
rect 6856 2202 6912 2204
rect 6616 2150 6642 2202
rect 6642 2150 6672 2202
rect 6696 2150 6706 2202
rect 6706 2150 6752 2202
rect 6776 2150 6822 2202
rect 6822 2150 6832 2202
rect 6856 2150 6886 2202
rect 6886 2150 6912 2202
rect 6616 2148 6672 2150
rect 6696 2148 6752 2150
rect 6776 2148 6832 2150
rect 6856 2148 6912 2150
<< metal3 >>
rect 0 15330 480 15360
rect 2773 15330 2839 15333
rect 0 15328 2839 15330
rect 0 15272 2778 15328
rect 2834 15272 2839 15328
rect 0 15270 2839 15272
rect 0 15240 480 15270
rect 2773 15267 2839 15270
rect 3208 14720 3528 14721
rect 3208 14656 3216 14720
rect 3280 14656 3296 14720
rect 3360 14656 3376 14720
rect 3440 14656 3456 14720
rect 3520 14656 3528 14720
rect 3208 14655 3528 14656
rect 5472 14720 5792 14721
rect 5472 14656 5480 14720
rect 5544 14656 5560 14720
rect 5624 14656 5640 14720
rect 5704 14656 5720 14720
rect 5784 14656 5792 14720
rect 5472 14655 5792 14656
rect 2076 14176 2396 14177
rect 2076 14112 2084 14176
rect 2148 14112 2164 14176
rect 2228 14112 2244 14176
rect 2308 14112 2324 14176
rect 2388 14112 2396 14176
rect 2076 14111 2396 14112
rect 4340 14176 4660 14177
rect 4340 14112 4348 14176
rect 4412 14112 4428 14176
rect 4492 14112 4508 14176
rect 4572 14112 4588 14176
rect 4652 14112 4660 14176
rect 4340 14111 4660 14112
rect 6604 14176 6924 14177
rect 6604 14112 6612 14176
rect 6676 14112 6692 14176
rect 6756 14112 6772 14176
rect 6836 14112 6852 14176
rect 6916 14112 6924 14176
rect 6604 14111 6924 14112
rect 3208 13632 3528 13633
rect 3208 13568 3216 13632
rect 3280 13568 3296 13632
rect 3360 13568 3376 13632
rect 3440 13568 3456 13632
rect 3520 13568 3528 13632
rect 3208 13567 3528 13568
rect 5472 13632 5792 13633
rect 5472 13568 5480 13632
rect 5544 13568 5560 13632
rect 5624 13568 5640 13632
rect 5704 13568 5720 13632
rect 5784 13568 5792 13632
rect 5472 13567 5792 13568
rect 2076 13088 2396 13089
rect 2076 13024 2084 13088
rect 2148 13024 2164 13088
rect 2228 13024 2244 13088
rect 2308 13024 2324 13088
rect 2388 13024 2396 13088
rect 2076 13023 2396 13024
rect 4340 13088 4660 13089
rect 4340 13024 4348 13088
rect 4412 13024 4428 13088
rect 4492 13024 4508 13088
rect 4572 13024 4588 13088
rect 4652 13024 4660 13088
rect 4340 13023 4660 13024
rect 6604 13088 6924 13089
rect 6604 13024 6612 13088
rect 6676 13024 6692 13088
rect 6756 13024 6772 13088
rect 6836 13024 6852 13088
rect 6916 13024 6924 13088
rect 6604 13023 6924 13024
rect 3208 12544 3528 12545
rect 3208 12480 3216 12544
rect 3280 12480 3296 12544
rect 3360 12480 3376 12544
rect 3440 12480 3456 12544
rect 3520 12480 3528 12544
rect 3208 12479 3528 12480
rect 5472 12544 5792 12545
rect 5472 12480 5480 12544
rect 5544 12480 5560 12544
rect 5624 12480 5640 12544
rect 5704 12480 5720 12544
rect 5784 12480 5792 12544
rect 5472 12479 5792 12480
rect 2076 12000 2396 12001
rect 0 11930 480 11960
rect 2076 11936 2084 12000
rect 2148 11936 2164 12000
rect 2228 11936 2244 12000
rect 2308 11936 2324 12000
rect 2388 11936 2396 12000
rect 2076 11935 2396 11936
rect 4340 12000 4660 12001
rect 4340 11936 4348 12000
rect 4412 11936 4428 12000
rect 4492 11936 4508 12000
rect 4572 11936 4588 12000
rect 4652 11936 4660 12000
rect 4340 11935 4660 11936
rect 6604 12000 6924 12001
rect 6604 11936 6612 12000
rect 6676 11936 6692 12000
rect 6756 11936 6772 12000
rect 6836 11936 6852 12000
rect 6916 11936 6924 12000
rect 6604 11935 6924 11936
rect 0 11870 1962 11930
rect 0 11840 480 11870
rect 1902 11794 1962 11870
rect 2865 11794 2931 11797
rect 1902 11792 2931 11794
rect 1902 11736 2870 11792
rect 2926 11736 2931 11792
rect 1902 11734 2931 11736
rect 2865 11731 2931 11734
rect 3208 11456 3528 11457
rect 3208 11392 3216 11456
rect 3280 11392 3296 11456
rect 3360 11392 3376 11456
rect 3440 11392 3456 11456
rect 3520 11392 3528 11456
rect 3208 11391 3528 11392
rect 5472 11456 5792 11457
rect 5472 11392 5480 11456
rect 5544 11392 5560 11456
rect 5624 11392 5640 11456
rect 5704 11392 5720 11456
rect 5784 11392 5792 11456
rect 5472 11391 5792 11392
rect 2076 10912 2396 10913
rect 2076 10848 2084 10912
rect 2148 10848 2164 10912
rect 2228 10848 2244 10912
rect 2308 10848 2324 10912
rect 2388 10848 2396 10912
rect 2076 10847 2396 10848
rect 4340 10912 4660 10913
rect 4340 10848 4348 10912
rect 4412 10848 4428 10912
rect 4492 10848 4508 10912
rect 4572 10848 4588 10912
rect 4652 10848 4660 10912
rect 4340 10847 4660 10848
rect 6604 10912 6924 10913
rect 6604 10848 6612 10912
rect 6676 10848 6692 10912
rect 6756 10848 6772 10912
rect 6836 10848 6852 10912
rect 6916 10848 6924 10912
rect 6604 10847 6924 10848
rect 3208 10368 3528 10369
rect 3208 10304 3216 10368
rect 3280 10304 3296 10368
rect 3360 10304 3376 10368
rect 3440 10304 3456 10368
rect 3520 10304 3528 10368
rect 3208 10303 3528 10304
rect 5472 10368 5792 10369
rect 5472 10304 5480 10368
rect 5544 10304 5560 10368
rect 5624 10304 5640 10368
rect 5704 10304 5720 10368
rect 5784 10304 5792 10368
rect 5472 10303 5792 10304
rect 2076 9824 2396 9825
rect 2076 9760 2084 9824
rect 2148 9760 2164 9824
rect 2228 9760 2244 9824
rect 2308 9760 2324 9824
rect 2388 9760 2396 9824
rect 2076 9759 2396 9760
rect 4340 9824 4660 9825
rect 4340 9760 4348 9824
rect 4412 9760 4428 9824
rect 4492 9760 4508 9824
rect 4572 9760 4588 9824
rect 4652 9760 4660 9824
rect 4340 9759 4660 9760
rect 6604 9824 6924 9825
rect 6604 9760 6612 9824
rect 6676 9760 6692 9824
rect 6756 9760 6772 9824
rect 6836 9760 6852 9824
rect 6916 9760 6924 9824
rect 6604 9759 6924 9760
rect 3208 9280 3528 9281
rect 3208 9216 3216 9280
rect 3280 9216 3296 9280
rect 3360 9216 3376 9280
rect 3440 9216 3456 9280
rect 3520 9216 3528 9280
rect 3208 9215 3528 9216
rect 5472 9280 5792 9281
rect 5472 9216 5480 9280
rect 5544 9216 5560 9280
rect 5624 9216 5640 9280
rect 5704 9216 5720 9280
rect 5784 9216 5792 9280
rect 5472 9215 5792 9216
rect 2076 8736 2396 8737
rect 2076 8672 2084 8736
rect 2148 8672 2164 8736
rect 2228 8672 2244 8736
rect 2308 8672 2324 8736
rect 2388 8672 2396 8736
rect 2076 8671 2396 8672
rect 4340 8736 4660 8737
rect 4340 8672 4348 8736
rect 4412 8672 4428 8736
rect 4492 8672 4508 8736
rect 4572 8672 4588 8736
rect 4652 8672 4660 8736
rect 4340 8671 4660 8672
rect 6604 8736 6924 8737
rect 6604 8672 6612 8736
rect 6676 8672 6692 8736
rect 6756 8672 6772 8736
rect 6836 8672 6852 8736
rect 6916 8672 6924 8736
rect 6604 8671 6924 8672
rect 0 8530 480 8560
rect 2221 8530 2287 8533
rect 0 8528 2287 8530
rect 0 8472 2226 8528
rect 2282 8472 2287 8528
rect 0 8470 2287 8472
rect 0 8440 480 8470
rect 2221 8467 2287 8470
rect 5349 8530 5415 8533
rect 8520 8530 9000 8560
rect 5349 8528 9000 8530
rect 5349 8472 5354 8528
rect 5410 8472 9000 8528
rect 5349 8470 9000 8472
rect 5349 8467 5415 8470
rect 8520 8440 9000 8470
rect 3208 8192 3528 8193
rect 3208 8128 3216 8192
rect 3280 8128 3296 8192
rect 3360 8128 3376 8192
rect 3440 8128 3456 8192
rect 3520 8128 3528 8192
rect 3208 8127 3528 8128
rect 5472 8192 5792 8193
rect 5472 8128 5480 8192
rect 5544 8128 5560 8192
rect 5624 8128 5640 8192
rect 5704 8128 5720 8192
rect 5784 8128 5792 8192
rect 5472 8127 5792 8128
rect 2076 7648 2396 7649
rect 2076 7584 2084 7648
rect 2148 7584 2164 7648
rect 2228 7584 2244 7648
rect 2308 7584 2324 7648
rect 2388 7584 2396 7648
rect 2076 7583 2396 7584
rect 4340 7648 4660 7649
rect 4340 7584 4348 7648
rect 4412 7584 4428 7648
rect 4492 7584 4508 7648
rect 4572 7584 4588 7648
rect 4652 7584 4660 7648
rect 4340 7583 4660 7584
rect 6604 7648 6924 7649
rect 6604 7584 6612 7648
rect 6676 7584 6692 7648
rect 6756 7584 6772 7648
rect 6836 7584 6852 7648
rect 6916 7584 6924 7648
rect 6604 7583 6924 7584
rect 3208 7104 3528 7105
rect 3208 7040 3216 7104
rect 3280 7040 3296 7104
rect 3360 7040 3376 7104
rect 3440 7040 3456 7104
rect 3520 7040 3528 7104
rect 3208 7039 3528 7040
rect 5472 7104 5792 7105
rect 5472 7040 5480 7104
rect 5544 7040 5560 7104
rect 5624 7040 5640 7104
rect 5704 7040 5720 7104
rect 5784 7040 5792 7104
rect 5472 7039 5792 7040
rect 2076 6560 2396 6561
rect 2076 6496 2084 6560
rect 2148 6496 2164 6560
rect 2228 6496 2244 6560
rect 2308 6496 2324 6560
rect 2388 6496 2396 6560
rect 2076 6495 2396 6496
rect 4340 6560 4660 6561
rect 4340 6496 4348 6560
rect 4412 6496 4428 6560
rect 4492 6496 4508 6560
rect 4572 6496 4588 6560
rect 4652 6496 4660 6560
rect 4340 6495 4660 6496
rect 6604 6560 6924 6561
rect 6604 6496 6612 6560
rect 6676 6496 6692 6560
rect 6756 6496 6772 6560
rect 6836 6496 6852 6560
rect 6916 6496 6924 6560
rect 6604 6495 6924 6496
rect 3208 6016 3528 6017
rect 3208 5952 3216 6016
rect 3280 5952 3296 6016
rect 3360 5952 3376 6016
rect 3440 5952 3456 6016
rect 3520 5952 3528 6016
rect 3208 5951 3528 5952
rect 5472 6016 5792 6017
rect 5472 5952 5480 6016
rect 5544 5952 5560 6016
rect 5624 5952 5640 6016
rect 5704 5952 5720 6016
rect 5784 5952 5792 6016
rect 5472 5951 5792 5952
rect 2076 5472 2396 5473
rect 2076 5408 2084 5472
rect 2148 5408 2164 5472
rect 2228 5408 2244 5472
rect 2308 5408 2324 5472
rect 2388 5408 2396 5472
rect 2076 5407 2396 5408
rect 4340 5472 4660 5473
rect 4340 5408 4348 5472
rect 4412 5408 4428 5472
rect 4492 5408 4508 5472
rect 4572 5408 4588 5472
rect 4652 5408 4660 5472
rect 4340 5407 4660 5408
rect 6604 5472 6924 5473
rect 6604 5408 6612 5472
rect 6676 5408 6692 5472
rect 6756 5408 6772 5472
rect 6836 5408 6852 5472
rect 6916 5408 6924 5472
rect 6604 5407 6924 5408
rect 0 5130 480 5160
rect 4061 5130 4127 5133
rect 0 5128 4127 5130
rect 0 5072 4066 5128
rect 4122 5072 4127 5128
rect 0 5070 4127 5072
rect 0 5040 480 5070
rect 4061 5067 4127 5070
rect 3208 4928 3528 4929
rect 3208 4864 3216 4928
rect 3280 4864 3296 4928
rect 3360 4864 3376 4928
rect 3440 4864 3456 4928
rect 3520 4864 3528 4928
rect 3208 4863 3528 4864
rect 5472 4928 5792 4929
rect 5472 4864 5480 4928
rect 5544 4864 5560 4928
rect 5624 4864 5640 4928
rect 5704 4864 5720 4928
rect 5784 4864 5792 4928
rect 5472 4863 5792 4864
rect 2076 4384 2396 4385
rect 2076 4320 2084 4384
rect 2148 4320 2164 4384
rect 2228 4320 2244 4384
rect 2308 4320 2324 4384
rect 2388 4320 2396 4384
rect 2076 4319 2396 4320
rect 4340 4384 4660 4385
rect 4340 4320 4348 4384
rect 4412 4320 4428 4384
rect 4492 4320 4508 4384
rect 4572 4320 4588 4384
rect 4652 4320 4660 4384
rect 4340 4319 4660 4320
rect 6604 4384 6924 4385
rect 6604 4320 6612 4384
rect 6676 4320 6692 4384
rect 6756 4320 6772 4384
rect 6836 4320 6852 4384
rect 6916 4320 6924 4384
rect 6604 4319 6924 4320
rect 3208 3840 3528 3841
rect 3208 3776 3216 3840
rect 3280 3776 3296 3840
rect 3360 3776 3376 3840
rect 3440 3776 3456 3840
rect 3520 3776 3528 3840
rect 3208 3775 3528 3776
rect 5472 3840 5792 3841
rect 5472 3776 5480 3840
rect 5544 3776 5560 3840
rect 5624 3776 5640 3840
rect 5704 3776 5720 3840
rect 5784 3776 5792 3840
rect 5472 3775 5792 3776
rect 2076 3296 2396 3297
rect 2076 3232 2084 3296
rect 2148 3232 2164 3296
rect 2228 3232 2244 3296
rect 2308 3232 2324 3296
rect 2388 3232 2396 3296
rect 2076 3231 2396 3232
rect 4340 3296 4660 3297
rect 4340 3232 4348 3296
rect 4412 3232 4428 3296
rect 4492 3232 4508 3296
rect 4572 3232 4588 3296
rect 4652 3232 4660 3296
rect 4340 3231 4660 3232
rect 6604 3296 6924 3297
rect 6604 3232 6612 3296
rect 6676 3232 6692 3296
rect 6756 3232 6772 3296
rect 6836 3232 6852 3296
rect 6916 3232 6924 3296
rect 6604 3231 6924 3232
rect 3208 2752 3528 2753
rect 3208 2688 3216 2752
rect 3280 2688 3296 2752
rect 3360 2688 3376 2752
rect 3440 2688 3456 2752
rect 3520 2688 3528 2752
rect 3208 2687 3528 2688
rect 5472 2752 5792 2753
rect 5472 2688 5480 2752
rect 5544 2688 5560 2752
rect 5624 2688 5640 2752
rect 5704 2688 5720 2752
rect 5784 2688 5792 2752
rect 5472 2687 5792 2688
rect 2076 2208 2396 2209
rect 2076 2144 2084 2208
rect 2148 2144 2164 2208
rect 2228 2144 2244 2208
rect 2308 2144 2324 2208
rect 2388 2144 2396 2208
rect 2076 2143 2396 2144
rect 4340 2208 4660 2209
rect 4340 2144 4348 2208
rect 4412 2144 4428 2208
rect 4492 2144 4508 2208
rect 4572 2144 4588 2208
rect 4652 2144 4660 2208
rect 4340 2143 4660 2144
rect 6604 2208 6924 2209
rect 6604 2144 6612 2208
rect 6676 2144 6692 2208
rect 6756 2144 6772 2208
rect 6836 2144 6852 2208
rect 6916 2144 6924 2208
rect 6604 2143 6924 2144
rect 0 1730 480 1760
rect 1945 1730 2011 1733
rect 0 1728 2011 1730
rect 0 1672 1950 1728
rect 2006 1672 2011 1728
rect 0 1670 2011 1672
rect 0 1640 480 1670
rect 1945 1667 2011 1670
<< via3 >>
rect 3216 14716 3280 14720
rect 3216 14660 3220 14716
rect 3220 14660 3276 14716
rect 3276 14660 3280 14716
rect 3216 14656 3280 14660
rect 3296 14716 3360 14720
rect 3296 14660 3300 14716
rect 3300 14660 3356 14716
rect 3356 14660 3360 14716
rect 3296 14656 3360 14660
rect 3376 14716 3440 14720
rect 3376 14660 3380 14716
rect 3380 14660 3436 14716
rect 3436 14660 3440 14716
rect 3376 14656 3440 14660
rect 3456 14716 3520 14720
rect 3456 14660 3460 14716
rect 3460 14660 3516 14716
rect 3516 14660 3520 14716
rect 3456 14656 3520 14660
rect 5480 14716 5544 14720
rect 5480 14660 5484 14716
rect 5484 14660 5540 14716
rect 5540 14660 5544 14716
rect 5480 14656 5544 14660
rect 5560 14716 5624 14720
rect 5560 14660 5564 14716
rect 5564 14660 5620 14716
rect 5620 14660 5624 14716
rect 5560 14656 5624 14660
rect 5640 14716 5704 14720
rect 5640 14660 5644 14716
rect 5644 14660 5700 14716
rect 5700 14660 5704 14716
rect 5640 14656 5704 14660
rect 5720 14716 5784 14720
rect 5720 14660 5724 14716
rect 5724 14660 5780 14716
rect 5780 14660 5784 14716
rect 5720 14656 5784 14660
rect 2084 14172 2148 14176
rect 2084 14116 2088 14172
rect 2088 14116 2144 14172
rect 2144 14116 2148 14172
rect 2084 14112 2148 14116
rect 2164 14172 2228 14176
rect 2164 14116 2168 14172
rect 2168 14116 2224 14172
rect 2224 14116 2228 14172
rect 2164 14112 2228 14116
rect 2244 14172 2308 14176
rect 2244 14116 2248 14172
rect 2248 14116 2304 14172
rect 2304 14116 2308 14172
rect 2244 14112 2308 14116
rect 2324 14172 2388 14176
rect 2324 14116 2328 14172
rect 2328 14116 2384 14172
rect 2384 14116 2388 14172
rect 2324 14112 2388 14116
rect 4348 14172 4412 14176
rect 4348 14116 4352 14172
rect 4352 14116 4408 14172
rect 4408 14116 4412 14172
rect 4348 14112 4412 14116
rect 4428 14172 4492 14176
rect 4428 14116 4432 14172
rect 4432 14116 4488 14172
rect 4488 14116 4492 14172
rect 4428 14112 4492 14116
rect 4508 14172 4572 14176
rect 4508 14116 4512 14172
rect 4512 14116 4568 14172
rect 4568 14116 4572 14172
rect 4508 14112 4572 14116
rect 4588 14172 4652 14176
rect 4588 14116 4592 14172
rect 4592 14116 4648 14172
rect 4648 14116 4652 14172
rect 4588 14112 4652 14116
rect 6612 14172 6676 14176
rect 6612 14116 6616 14172
rect 6616 14116 6672 14172
rect 6672 14116 6676 14172
rect 6612 14112 6676 14116
rect 6692 14172 6756 14176
rect 6692 14116 6696 14172
rect 6696 14116 6752 14172
rect 6752 14116 6756 14172
rect 6692 14112 6756 14116
rect 6772 14172 6836 14176
rect 6772 14116 6776 14172
rect 6776 14116 6832 14172
rect 6832 14116 6836 14172
rect 6772 14112 6836 14116
rect 6852 14172 6916 14176
rect 6852 14116 6856 14172
rect 6856 14116 6912 14172
rect 6912 14116 6916 14172
rect 6852 14112 6916 14116
rect 3216 13628 3280 13632
rect 3216 13572 3220 13628
rect 3220 13572 3276 13628
rect 3276 13572 3280 13628
rect 3216 13568 3280 13572
rect 3296 13628 3360 13632
rect 3296 13572 3300 13628
rect 3300 13572 3356 13628
rect 3356 13572 3360 13628
rect 3296 13568 3360 13572
rect 3376 13628 3440 13632
rect 3376 13572 3380 13628
rect 3380 13572 3436 13628
rect 3436 13572 3440 13628
rect 3376 13568 3440 13572
rect 3456 13628 3520 13632
rect 3456 13572 3460 13628
rect 3460 13572 3516 13628
rect 3516 13572 3520 13628
rect 3456 13568 3520 13572
rect 5480 13628 5544 13632
rect 5480 13572 5484 13628
rect 5484 13572 5540 13628
rect 5540 13572 5544 13628
rect 5480 13568 5544 13572
rect 5560 13628 5624 13632
rect 5560 13572 5564 13628
rect 5564 13572 5620 13628
rect 5620 13572 5624 13628
rect 5560 13568 5624 13572
rect 5640 13628 5704 13632
rect 5640 13572 5644 13628
rect 5644 13572 5700 13628
rect 5700 13572 5704 13628
rect 5640 13568 5704 13572
rect 5720 13628 5784 13632
rect 5720 13572 5724 13628
rect 5724 13572 5780 13628
rect 5780 13572 5784 13628
rect 5720 13568 5784 13572
rect 2084 13084 2148 13088
rect 2084 13028 2088 13084
rect 2088 13028 2144 13084
rect 2144 13028 2148 13084
rect 2084 13024 2148 13028
rect 2164 13084 2228 13088
rect 2164 13028 2168 13084
rect 2168 13028 2224 13084
rect 2224 13028 2228 13084
rect 2164 13024 2228 13028
rect 2244 13084 2308 13088
rect 2244 13028 2248 13084
rect 2248 13028 2304 13084
rect 2304 13028 2308 13084
rect 2244 13024 2308 13028
rect 2324 13084 2388 13088
rect 2324 13028 2328 13084
rect 2328 13028 2384 13084
rect 2384 13028 2388 13084
rect 2324 13024 2388 13028
rect 4348 13084 4412 13088
rect 4348 13028 4352 13084
rect 4352 13028 4408 13084
rect 4408 13028 4412 13084
rect 4348 13024 4412 13028
rect 4428 13084 4492 13088
rect 4428 13028 4432 13084
rect 4432 13028 4488 13084
rect 4488 13028 4492 13084
rect 4428 13024 4492 13028
rect 4508 13084 4572 13088
rect 4508 13028 4512 13084
rect 4512 13028 4568 13084
rect 4568 13028 4572 13084
rect 4508 13024 4572 13028
rect 4588 13084 4652 13088
rect 4588 13028 4592 13084
rect 4592 13028 4648 13084
rect 4648 13028 4652 13084
rect 4588 13024 4652 13028
rect 6612 13084 6676 13088
rect 6612 13028 6616 13084
rect 6616 13028 6672 13084
rect 6672 13028 6676 13084
rect 6612 13024 6676 13028
rect 6692 13084 6756 13088
rect 6692 13028 6696 13084
rect 6696 13028 6752 13084
rect 6752 13028 6756 13084
rect 6692 13024 6756 13028
rect 6772 13084 6836 13088
rect 6772 13028 6776 13084
rect 6776 13028 6832 13084
rect 6832 13028 6836 13084
rect 6772 13024 6836 13028
rect 6852 13084 6916 13088
rect 6852 13028 6856 13084
rect 6856 13028 6912 13084
rect 6912 13028 6916 13084
rect 6852 13024 6916 13028
rect 3216 12540 3280 12544
rect 3216 12484 3220 12540
rect 3220 12484 3276 12540
rect 3276 12484 3280 12540
rect 3216 12480 3280 12484
rect 3296 12540 3360 12544
rect 3296 12484 3300 12540
rect 3300 12484 3356 12540
rect 3356 12484 3360 12540
rect 3296 12480 3360 12484
rect 3376 12540 3440 12544
rect 3376 12484 3380 12540
rect 3380 12484 3436 12540
rect 3436 12484 3440 12540
rect 3376 12480 3440 12484
rect 3456 12540 3520 12544
rect 3456 12484 3460 12540
rect 3460 12484 3516 12540
rect 3516 12484 3520 12540
rect 3456 12480 3520 12484
rect 5480 12540 5544 12544
rect 5480 12484 5484 12540
rect 5484 12484 5540 12540
rect 5540 12484 5544 12540
rect 5480 12480 5544 12484
rect 5560 12540 5624 12544
rect 5560 12484 5564 12540
rect 5564 12484 5620 12540
rect 5620 12484 5624 12540
rect 5560 12480 5624 12484
rect 5640 12540 5704 12544
rect 5640 12484 5644 12540
rect 5644 12484 5700 12540
rect 5700 12484 5704 12540
rect 5640 12480 5704 12484
rect 5720 12540 5784 12544
rect 5720 12484 5724 12540
rect 5724 12484 5780 12540
rect 5780 12484 5784 12540
rect 5720 12480 5784 12484
rect 2084 11996 2148 12000
rect 2084 11940 2088 11996
rect 2088 11940 2144 11996
rect 2144 11940 2148 11996
rect 2084 11936 2148 11940
rect 2164 11996 2228 12000
rect 2164 11940 2168 11996
rect 2168 11940 2224 11996
rect 2224 11940 2228 11996
rect 2164 11936 2228 11940
rect 2244 11996 2308 12000
rect 2244 11940 2248 11996
rect 2248 11940 2304 11996
rect 2304 11940 2308 11996
rect 2244 11936 2308 11940
rect 2324 11996 2388 12000
rect 2324 11940 2328 11996
rect 2328 11940 2384 11996
rect 2384 11940 2388 11996
rect 2324 11936 2388 11940
rect 4348 11996 4412 12000
rect 4348 11940 4352 11996
rect 4352 11940 4408 11996
rect 4408 11940 4412 11996
rect 4348 11936 4412 11940
rect 4428 11996 4492 12000
rect 4428 11940 4432 11996
rect 4432 11940 4488 11996
rect 4488 11940 4492 11996
rect 4428 11936 4492 11940
rect 4508 11996 4572 12000
rect 4508 11940 4512 11996
rect 4512 11940 4568 11996
rect 4568 11940 4572 11996
rect 4508 11936 4572 11940
rect 4588 11996 4652 12000
rect 4588 11940 4592 11996
rect 4592 11940 4648 11996
rect 4648 11940 4652 11996
rect 4588 11936 4652 11940
rect 6612 11996 6676 12000
rect 6612 11940 6616 11996
rect 6616 11940 6672 11996
rect 6672 11940 6676 11996
rect 6612 11936 6676 11940
rect 6692 11996 6756 12000
rect 6692 11940 6696 11996
rect 6696 11940 6752 11996
rect 6752 11940 6756 11996
rect 6692 11936 6756 11940
rect 6772 11996 6836 12000
rect 6772 11940 6776 11996
rect 6776 11940 6832 11996
rect 6832 11940 6836 11996
rect 6772 11936 6836 11940
rect 6852 11996 6916 12000
rect 6852 11940 6856 11996
rect 6856 11940 6912 11996
rect 6912 11940 6916 11996
rect 6852 11936 6916 11940
rect 3216 11452 3280 11456
rect 3216 11396 3220 11452
rect 3220 11396 3276 11452
rect 3276 11396 3280 11452
rect 3216 11392 3280 11396
rect 3296 11452 3360 11456
rect 3296 11396 3300 11452
rect 3300 11396 3356 11452
rect 3356 11396 3360 11452
rect 3296 11392 3360 11396
rect 3376 11452 3440 11456
rect 3376 11396 3380 11452
rect 3380 11396 3436 11452
rect 3436 11396 3440 11452
rect 3376 11392 3440 11396
rect 3456 11452 3520 11456
rect 3456 11396 3460 11452
rect 3460 11396 3516 11452
rect 3516 11396 3520 11452
rect 3456 11392 3520 11396
rect 5480 11452 5544 11456
rect 5480 11396 5484 11452
rect 5484 11396 5540 11452
rect 5540 11396 5544 11452
rect 5480 11392 5544 11396
rect 5560 11452 5624 11456
rect 5560 11396 5564 11452
rect 5564 11396 5620 11452
rect 5620 11396 5624 11452
rect 5560 11392 5624 11396
rect 5640 11452 5704 11456
rect 5640 11396 5644 11452
rect 5644 11396 5700 11452
rect 5700 11396 5704 11452
rect 5640 11392 5704 11396
rect 5720 11452 5784 11456
rect 5720 11396 5724 11452
rect 5724 11396 5780 11452
rect 5780 11396 5784 11452
rect 5720 11392 5784 11396
rect 2084 10908 2148 10912
rect 2084 10852 2088 10908
rect 2088 10852 2144 10908
rect 2144 10852 2148 10908
rect 2084 10848 2148 10852
rect 2164 10908 2228 10912
rect 2164 10852 2168 10908
rect 2168 10852 2224 10908
rect 2224 10852 2228 10908
rect 2164 10848 2228 10852
rect 2244 10908 2308 10912
rect 2244 10852 2248 10908
rect 2248 10852 2304 10908
rect 2304 10852 2308 10908
rect 2244 10848 2308 10852
rect 2324 10908 2388 10912
rect 2324 10852 2328 10908
rect 2328 10852 2384 10908
rect 2384 10852 2388 10908
rect 2324 10848 2388 10852
rect 4348 10908 4412 10912
rect 4348 10852 4352 10908
rect 4352 10852 4408 10908
rect 4408 10852 4412 10908
rect 4348 10848 4412 10852
rect 4428 10908 4492 10912
rect 4428 10852 4432 10908
rect 4432 10852 4488 10908
rect 4488 10852 4492 10908
rect 4428 10848 4492 10852
rect 4508 10908 4572 10912
rect 4508 10852 4512 10908
rect 4512 10852 4568 10908
rect 4568 10852 4572 10908
rect 4508 10848 4572 10852
rect 4588 10908 4652 10912
rect 4588 10852 4592 10908
rect 4592 10852 4648 10908
rect 4648 10852 4652 10908
rect 4588 10848 4652 10852
rect 6612 10908 6676 10912
rect 6612 10852 6616 10908
rect 6616 10852 6672 10908
rect 6672 10852 6676 10908
rect 6612 10848 6676 10852
rect 6692 10908 6756 10912
rect 6692 10852 6696 10908
rect 6696 10852 6752 10908
rect 6752 10852 6756 10908
rect 6692 10848 6756 10852
rect 6772 10908 6836 10912
rect 6772 10852 6776 10908
rect 6776 10852 6832 10908
rect 6832 10852 6836 10908
rect 6772 10848 6836 10852
rect 6852 10908 6916 10912
rect 6852 10852 6856 10908
rect 6856 10852 6912 10908
rect 6912 10852 6916 10908
rect 6852 10848 6916 10852
rect 3216 10364 3280 10368
rect 3216 10308 3220 10364
rect 3220 10308 3276 10364
rect 3276 10308 3280 10364
rect 3216 10304 3280 10308
rect 3296 10364 3360 10368
rect 3296 10308 3300 10364
rect 3300 10308 3356 10364
rect 3356 10308 3360 10364
rect 3296 10304 3360 10308
rect 3376 10364 3440 10368
rect 3376 10308 3380 10364
rect 3380 10308 3436 10364
rect 3436 10308 3440 10364
rect 3376 10304 3440 10308
rect 3456 10364 3520 10368
rect 3456 10308 3460 10364
rect 3460 10308 3516 10364
rect 3516 10308 3520 10364
rect 3456 10304 3520 10308
rect 5480 10364 5544 10368
rect 5480 10308 5484 10364
rect 5484 10308 5540 10364
rect 5540 10308 5544 10364
rect 5480 10304 5544 10308
rect 5560 10364 5624 10368
rect 5560 10308 5564 10364
rect 5564 10308 5620 10364
rect 5620 10308 5624 10364
rect 5560 10304 5624 10308
rect 5640 10364 5704 10368
rect 5640 10308 5644 10364
rect 5644 10308 5700 10364
rect 5700 10308 5704 10364
rect 5640 10304 5704 10308
rect 5720 10364 5784 10368
rect 5720 10308 5724 10364
rect 5724 10308 5780 10364
rect 5780 10308 5784 10364
rect 5720 10304 5784 10308
rect 2084 9820 2148 9824
rect 2084 9764 2088 9820
rect 2088 9764 2144 9820
rect 2144 9764 2148 9820
rect 2084 9760 2148 9764
rect 2164 9820 2228 9824
rect 2164 9764 2168 9820
rect 2168 9764 2224 9820
rect 2224 9764 2228 9820
rect 2164 9760 2228 9764
rect 2244 9820 2308 9824
rect 2244 9764 2248 9820
rect 2248 9764 2304 9820
rect 2304 9764 2308 9820
rect 2244 9760 2308 9764
rect 2324 9820 2388 9824
rect 2324 9764 2328 9820
rect 2328 9764 2384 9820
rect 2384 9764 2388 9820
rect 2324 9760 2388 9764
rect 4348 9820 4412 9824
rect 4348 9764 4352 9820
rect 4352 9764 4408 9820
rect 4408 9764 4412 9820
rect 4348 9760 4412 9764
rect 4428 9820 4492 9824
rect 4428 9764 4432 9820
rect 4432 9764 4488 9820
rect 4488 9764 4492 9820
rect 4428 9760 4492 9764
rect 4508 9820 4572 9824
rect 4508 9764 4512 9820
rect 4512 9764 4568 9820
rect 4568 9764 4572 9820
rect 4508 9760 4572 9764
rect 4588 9820 4652 9824
rect 4588 9764 4592 9820
rect 4592 9764 4648 9820
rect 4648 9764 4652 9820
rect 4588 9760 4652 9764
rect 6612 9820 6676 9824
rect 6612 9764 6616 9820
rect 6616 9764 6672 9820
rect 6672 9764 6676 9820
rect 6612 9760 6676 9764
rect 6692 9820 6756 9824
rect 6692 9764 6696 9820
rect 6696 9764 6752 9820
rect 6752 9764 6756 9820
rect 6692 9760 6756 9764
rect 6772 9820 6836 9824
rect 6772 9764 6776 9820
rect 6776 9764 6832 9820
rect 6832 9764 6836 9820
rect 6772 9760 6836 9764
rect 6852 9820 6916 9824
rect 6852 9764 6856 9820
rect 6856 9764 6912 9820
rect 6912 9764 6916 9820
rect 6852 9760 6916 9764
rect 3216 9276 3280 9280
rect 3216 9220 3220 9276
rect 3220 9220 3276 9276
rect 3276 9220 3280 9276
rect 3216 9216 3280 9220
rect 3296 9276 3360 9280
rect 3296 9220 3300 9276
rect 3300 9220 3356 9276
rect 3356 9220 3360 9276
rect 3296 9216 3360 9220
rect 3376 9276 3440 9280
rect 3376 9220 3380 9276
rect 3380 9220 3436 9276
rect 3436 9220 3440 9276
rect 3376 9216 3440 9220
rect 3456 9276 3520 9280
rect 3456 9220 3460 9276
rect 3460 9220 3516 9276
rect 3516 9220 3520 9276
rect 3456 9216 3520 9220
rect 5480 9276 5544 9280
rect 5480 9220 5484 9276
rect 5484 9220 5540 9276
rect 5540 9220 5544 9276
rect 5480 9216 5544 9220
rect 5560 9276 5624 9280
rect 5560 9220 5564 9276
rect 5564 9220 5620 9276
rect 5620 9220 5624 9276
rect 5560 9216 5624 9220
rect 5640 9276 5704 9280
rect 5640 9220 5644 9276
rect 5644 9220 5700 9276
rect 5700 9220 5704 9276
rect 5640 9216 5704 9220
rect 5720 9276 5784 9280
rect 5720 9220 5724 9276
rect 5724 9220 5780 9276
rect 5780 9220 5784 9276
rect 5720 9216 5784 9220
rect 2084 8732 2148 8736
rect 2084 8676 2088 8732
rect 2088 8676 2144 8732
rect 2144 8676 2148 8732
rect 2084 8672 2148 8676
rect 2164 8732 2228 8736
rect 2164 8676 2168 8732
rect 2168 8676 2224 8732
rect 2224 8676 2228 8732
rect 2164 8672 2228 8676
rect 2244 8732 2308 8736
rect 2244 8676 2248 8732
rect 2248 8676 2304 8732
rect 2304 8676 2308 8732
rect 2244 8672 2308 8676
rect 2324 8732 2388 8736
rect 2324 8676 2328 8732
rect 2328 8676 2384 8732
rect 2384 8676 2388 8732
rect 2324 8672 2388 8676
rect 4348 8732 4412 8736
rect 4348 8676 4352 8732
rect 4352 8676 4408 8732
rect 4408 8676 4412 8732
rect 4348 8672 4412 8676
rect 4428 8732 4492 8736
rect 4428 8676 4432 8732
rect 4432 8676 4488 8732
rect 4488 8676 4492 8732
rect 4428 8672 4492 8676
rect 4508 8732 4572 8736
rect 4508 8676 4512 8732
rect 4512 8676 4568 8732
rect 4568 8676 4572 8732
rect 4508 8672 4572 8676
rect 4588 8732 4652 8736
rect 4588 8676 4592 8732
rect 4592 8676 4648 8732
rect 4648 8676 4652 8732
rect 4588 8672 4652 8676
rect 6612 8732 6676 8736
rect 6612 8676 6616 8732
rect 6616 8676 6672 8732
rect 6672 8676 6676 8732
rect 6612 8672 6676 8676
rect 6692 8732 6756 8736
rect 6692 8676 6696 8732
rect 6696 8676 6752 8732
rect 6752 8676 6756 8732
rect 6692 8672 6756 8676
rect 6772 8732 6836 8736
rect 6772 8676 6776 8732
rect 6776 8676 6832 8732
rect 6832 8676 6836 8732
rect 6772 8672 6836 8676
rect 6852 8732 6916 8736
rect 6852 8676 6856 8732
rect 6856 8676 6912 8732
rect 6912 8676 6916 8732
rect 6852 8672 6916 8676
rect 3216 8188 3280 8192
rect 3216 8132 3220 8188
rect 3220 8132 3276 8188
rect 3276 8132 3280 8188
rect 3216 8128 3280 8132
rect 3296 8188 3360 8192
rect 3296 8132 3300 8188
rect 3300 8132 3356 8188
rect 3356 8132 3360 8188
rect 3296 8128 3360 8132
rect 3376 8188 3440 8192
rect 3376 8132 3380 8188
rect 3380 8132 3436 8188
rect 3436 8132 3440 8188
rect 3376 8128 3440 8132
rect 3456 8188 3520 8192
rect 3456 8132 3460 8188
rect 3460 8132 3516 8188
rect 3516 8132 3520 8188
rect 3456 8128 3520 8132
rect 5480 8188 5544 8192
rect 5480 8132 5484 8188
rect 5484 8132 5540 8188
rect 5540 8132 5544 8188
rect 5480 8128 5544 8132
rect 5560 8188 5624 8192
rect 5560 8132 5564 8188
rect 5564 8132 5620 8188
rect 5620 8132 5624 8188
rect 5560 8128 5624 8132
rect 5640 8188 5704 8192
rect 5640 8132 5644 8188
rect 5644 8132 5700 8188
rect 5700 8132 5704 8188
rect 5640 8128 5704 8132
rect 5720 8188 5784 8192
rect 5720 8132 5724 8188
rect 5724 8132 5780 8188
rect 5780 8132 5784 8188
rect 5720 8128 5784 8132
rect 2084 7644 2148 7648
rect 2084 7588 2088 7644
rect 2088 7588 2144 7644
rect 2144 7588 2148 7644
rect 2084 7584 2148 7588
rect 2164 7644 2228 7648
rect 2164 7588 2168 7644
rect 2168 7588 2224 7644
rect 2224 7588 2228 7644
rect 2164 7584 2228 7588
rect 2244 7644 2308 7648
rect 2244 7588 2248 7644
rect 2248 7588 2304 7644
rect 2304 7588 2308 7644
rect 2244 7584 2308 7588
rect 2324 7644 2388 7648
rect 2324 7588 2328 7644
rect 2328 7588 2384 7644
rect 2384 7588 2388 7644
rect 2324 7584 2388 7588
rect 4348 7644 4412 7648
rect 4348 7588 4352 7644
rect 4352 7588 4408 7644
rect 4408 7588 4412 7644
rect 4348 7584 4412 7588
rect 4428 7644 4492 7648
rect 4428 7588 4432 7644
rect 4432 7588 4488 7644
rect 4488 7588 4492 7644
rect 4428 7584 4492 7588
rect 4508 7644 4572 7648
rect 4508 7588 4512 7644
rect 4512 7588 4568 7644
rect 4568 7588 4572 7644
rect 4508 7584 4572 7588
rect 4588 7644 4652 7648
rect 4588 7588 4592 7644
rect 4592 7588 4648 7644
rect 4648 7588 4652 7644
rect 4588 7584 4652 7588
rect 6612 7644 6676 7648
rect 6612 7588 6616 7644
rect 6616 7588 6672 7644
rect 6672 7588 6676 7644
rect 6612 7584 6676 7588
rect 6692 7644 6756 7648
rect 6692 7588 6696 7644
rect 6696 7588 6752 7644
rect 6752 7588 6756 7644
rect 6692 7584 6756 7588
rect 6772 7644 6836 7648
rect 6772 7588 6776 7644
rect 6776 7588 6832 7644
rect 6832 7588 6836 7644
rect 6772 7584 6836 7588
rect 6852 7644 6916 7648
rect 6852 7588 6856 7644
rect 6856 7588 6912 7644
rect 6912 7588 6916 7644
rect 6852 7584 6916 7588
rect 3216 7100 3280 7104
rect 3216 7044 3220 7100
rect 3220 7044 3276 7100
rect 3276 7044 3280 7100
rect 3216 7040 3280 7044
rect 3296 7100 3360 7104
rect 3296 7044 3300 7100
rect 3300 7044 3356 7100
rect 3356 7044 3360 7100
rect 3296 7040 3360 7044
rect 3376 7100 3440 7104
rect 3376 7044 3380 7100
rect 3380 7044 3436 7100
rect 3436 7044 3440 7100
rect 3376 7040 3440 7044
rect 3456 7100 3520 7104
rect 3456 7044 3460 7100
rect 3460 7044 3516 7100
rect 3516 7044 3520 7100
rect 3456 7040 3520 7044
rect 5480 7100 5544 7104
rect 5480 7044 5484 7100
rect 5484 7044 5540 7100
rect 5540 7044 5544 7100
rect 5480 7040 5544 7044
rect 5560 7100 5624 7104
rect 5560 7044 5564 7100
rect 5564 7044 5620 7100
rect 5620 7044 5624 7100
rect 5560 7040 5624 7044
rect 5640 7100 5704 7104
rect 5640 7044 5644 7100
rect 5644 7044 5700 7100
rect 5700 7044 5704 7100
rect 5640 7040 5704 7044
rect 5720 7100 5784 7104
rect 5720 7044 5724 7100
rect 5724 7044 5780 7100
rect 5780 7044 5784 7100
rect 5720 7040 5784 7044
rect 2084 6556 2148 6560
rect 2084 6500 2088 6556
rect 2088 6500 2144 6556
rect 2144 6500 2148 6556
rect 2084 6496 2148 6500
rect 2164 6556 2228 6560
rect 2164 6500 2168 6556
rect 2168 6500 2224 6556
rect 2224 6500 2228 6556
rect 2164 6496 2228 6500
rect 2244 6556 2308 6560
rect 2244 6500 2248 6556
rect 2248 6500 2304 6556
rect 2304 6500 2308 6556
rect 2244 6496 2308 6500
rect 2324 6556 2388 6560
rect 2324 6500 2328 6556
rect 2328 6500 2384 6556
rect 2384 6500 2388 6556
rect 2324 6496 2388 6500
rect 4348 6556 4412 6560
rect 4348 6500 4352 6556
rect 4352 6500 4408 6556
rect 4408 6500 4412 6556
rect 4348 6496 4412 6500
rect 4428 6556 4492 6560
rect 4428 6500 4432 6556
rect 4432 6500 4488 6556
rect 4488 6500 4492 6556
rect 4428 6496 4492 6500
rect 4508 6556 4572 6560
rect 4508 6500 4512 6556
rect 4512 6500 4568 6556
rect 4568 6500 4572 6556
rect 4508 6496 4572 6500
rect 4588 6556 4652 6560
rect 4588 6500 4592 6556
rect 4592 6500 4648 6556
rect 4648 6500 4652 6556
rect 4588 6496 4652 6500
rect 6612 6556 6676 6560
rect 6612 6500 6616 6556
rect 6616 6500 6672 6556
rect 6672 6500 6676 6556
rect 6612 6496 6676 6500
rect 6692 6556 6756 6560
rect 6692 6500 6696 6556
rect 6696 6500 6752 6556
rect 6752 6500 6756 6556
rect 6692 6496 6756 6500
rect 6772 6556 6836 6560
rect 6772 6500 6776 6556
rect 6776 6500 6832 6556
rect 6832 6500 6836 6556
rect 6772 6496 6836 6500
rect 6852 6556 6916 6560
rect 6852 6500 6856 6556
rect 6856 6500 6912 6556
rect 6912 6500 6916 6556
rect 6852 6496 6916 6500
rect 3216 6012 3280 6016
rect 3216 5956 3220 6012
rect 3220 5956 3276 6012
rect 3276 5956 3280 6012
rect 3216 5952 3280 5956
rect 3296 6012 3360 6016
rect 3296 5956 3300 6012
rect 3300 5956 3356 6012
rect 3356 5956 3360 6012
rect 3296 5952 3360 5956
rect 3376 6012 3440 6016
rect 3376 5956 3380 6012
rect 3380 5956 3436 6012
rect 3436 5956 3440 6012
rect 3376 5952 3440 5956
rect 3456 6012 3520 6016
rect 3456 5956 3460 6012
rect 3460 5956 3516 6012
rect 3516 5956 3520 6012
rect 3456 5952 3520 5956
rect 5480 6012 5544 6016
rect 5480 5956 5484 6012
rect 5484 5956 5540 6012
rect 5540 5956 5544 6012
rect 5480 5952 5544 5956
rect 5560 6012 5624 6016
rect 5560 5956 5564 6012
rect 5564 5956 5620 6012
rect 5620 5956 5624 6012
rect 5560 5952 5624 5956
rect 5640 6012 5704 6016
rect 5640 5956 5644 6012
rect 5644 5956 5700 6012
rect 5700 5956 5704 6012
rect 5640 5952 5704 5956
rect 5720 6012 5784 6016
rect 5720 5956 5724 6012
rect 5724 5956 5780 6012
rect 5780 5956 5784 6012
rect 5720 5952 5784 5956
rect 2084 5468 2148 5472
rect 2084 5412 2088 5468
rect 2088 5412 2144 5468
rect 2144 5412 2148 5468
rect 2084 5408 2148 5412
rect 2164 5468 2228 5472
rect 2164 5412 2168 5468
rect 2168 5412 2224 5468
rect 2224 5412 2228 5468
rect 2164 5408 2228 5412
rect 2244 5468 2308 5472
rect 2244 5412 2248 5468
rect 2248 5412 2304 5468
rect 2304 5412 2308 5468
rect 2244 5408 2308 5412
rect 2324 5468 2388 5472
rect 2324 5412 2328 5468
rect 2328 5412 2384 5468
rect 2384 5412 2388 5468
rect 2324 5408 2388 5412
rect 4348 5468 4412 5472
rect 4348 5412 4352 5468
rect 4352 5412 4408 5468
rect 4408 5412 4412 5468
rect 4348 5408 4412 5412
rect 4428 5468 4492 5472
rect 4428 5412 4432 5468
rect 4432 5412 4488 5468
rect 4488 5412 4492 5468
rect 4428 5408 4492 5412
rect 4508 5468 4572 5472
rect 4508 5412 4512 5468
rect 4512 5412 4568 5468
rect 4568 5412 4572 5468
rect 4508 5408 4572 5412
rect 4588 5468 4652 5472
rect 4588 5412 4592 5468
rect 4592 5412 4648 5468
rect 4648 5412 4652 5468
rect 4588 5408 4652 5412
rect 6612 5468 6676 5472
rect 6612 5412 6616 5468
rect 6616 5412 6672 5468
rect 6672 5412 6676 5468
rect 6612 5408 6676 5412
rect 6692 5468 6756 5472
rect 6692 5412 6696 5468
rect 6696 5412 6752 5468
rect 6752 5412 6756 5468
rect 6692 5408 6756 5412
rect 6772 5468 6836 5472
rect 6772 5412 6776 5468
rect 6776 5412 6832 5468
rect 6832 5412 6836 5468
rect 6772 5408 6836 5412
rect 6852 5468 6916 5472
rect 6852 5412 6856 5468
rect 6856 5412 6912 5468
rect 6912 5412 6916 5468
rect 6852 5408 6916 5412
rect 3216 4924 3280 4928
rect 3216 4868 3220 4924
rect 3220 4868 3276 4924
rect 3276 4868 3280 4924
rect 3216 4864 3280 4868
rect 3296 4924 3360 4928
rect 3296 4868 3300 4924
rect 3300 4868 3356 4924
rect 3356 4868 3360 4924
rect 3296 4864 3360 4868
rect 3376 4924 3440 4928
rect 3376 4868 3380 4924
rect 3380 4868 3436 4924
rect 3436 4868 3440 4924
rect 3376 4864 3440 4868
rect 3456 4924 3520 4928
rect 3456 4868 3460 4924
rect 3460 4868 3516 4924
rect 3516 4868 3520 4924
rect 3456 4864 3520 4868
rect 5480 4924 5544 4928
rect 5480 4868 5484 4924
rect 5484 4868 5540 4924
rect 5540 4868 5544 4924
rect 5480 4864 5544 4868
rect 5560 4924 5624 4928
rect 5560 4868 5564 4924
rect 5564 4868 5620 4924
rect 5620 4868 5624 4924
rect 5560 4864 5624 4868
rect 5640 4924 5704 4928
rect 5640 4868 5644 4924
rect 5644 4868 5700 4924
rect 5700 4868 5704 4924
rect 5640 4864 5704 4868
rect 5720 4924 5784 4928
rect 5720 4868 5724 4924
rect 5724 4868 5780 4924
rect 5780 4868 5784 4924
rect 5720 4864 5784 4868
rect 2084 4380 2148 4384
rect 2084 4324 2088 4380
rect 2088 4324 2144 4380
rect 2144 4324 2148 4380
rect 2084 4320 2148 4324
rect 2164 4380 2228 4384
rect 2164 4324 2168 4380
rect 2168 4324 2224 4380
rect 2224 4324 2228 4380
rect 2164 4320 2228 4324
rect 2244 4380 2308 4384
rect 2244 4324 2248 4380
rect 2248 4324 2304 4380
rect 2304 4324 2308 4380
rect 2244 4320 2308 4324
rect 2324 4380 2388 4384
rect 2324 4324 2328 4380
rect 2328 4324 2384 4380
rect 2384 4324 2388 4380
rect 2324 4320 2388 4324
rect 4348 4380 4412 4384
rect 4348 4324 4352 4380
rect 4352 4324 4408 4380
rect 4408 4324 4412 4380
rect 4348 4320 4412 4324
rect 4428 4380 4492 4384
rect 4428 4324 4432 4380
rect 4432 4324 4488 4380
rect 4488 4324 4492 4380
rect 4428 4320 4492 4324
rect 4508 4380 4572 4384
rect 4508 4324 4512 4380
rect 4512 4324 4568 4380
rect 4568 4324 4572 4380
rect 4508 4320 4572 4324
rect 4588 4380 4652 4384
rect 4588 4324 4592 4380
rect 4592 4324 4648 4380
rect 4648 4324 4652 4380
rect 4588 4320 4652 4324
rect 6612 4380 6676 4384
rect 6612 4324 6616 4380
rect 6616 4324 6672 4380
rect 6672 4324 6676 4380
rect 6612 4320 6676 4324
rect 6692 4380 6756 4384
rect 6692 4324 6696 4380
rect 6696 4324 6752 4380
rect 6752 4324 6756 4380
rect 6692 4320 6756 4324
rect 6772 4380 6836 4384
rect 6772 4324 6776 4380
rect 6776 4324 6832 4380
rect 6832 4324 6836 4380
rect 6772 4320 6836 4324
rect 6852 4380 6916 4384
rect 6852 4324 6856 4380
rect 6856 4324 6912 4380
rect 6912 4324 6916 4380
rect 6852 4320 6916 4324
rect 3216 3836 3280 3840
rect 3216 3780 3220 3836
rect 3220 3780 3276 3836
rect 3276 3780 3280 3836
rect 3216 3776 3280 3780
rect 3296 3836 3360 3840
rect 3296 3780 3300 3836
rect 3300 3780 3356 3836
rect 3356 3780 3360 3836
rect 3296 3776 3360 3780
rect 3376 3836 3440 3840
rect 3376 3780 3380 3836
rect 3380 3780 3436 3836
rect 3436 3780 3440 3836
rect 3376 3776 3440 3780
rect 3456 3836 3520 3840
rect 3456 3780 3460 3836
rect 3460 3780 3516 3836
rect 3516 3780 3520 3836
rect 3456 3776 3520 3780
rect 5480 3836 5544 3840
rect 5480 3780 5484 3836
rect 5484 3780 5540 3836
rect 5540 3780 5544 3836
rect 5480 3776 5544 3780
rect 5560 3836 5624 3840
rect 5560 3780 5564 3836
rect 5564 3780 5620 3836
rect 5620 3780 5624 3836
rect 5560 3776 5624 3780
rect 5640 3836 5704 3840
rect 5640 3780 5644 3836
rect 5644 3780 5700 3836
rect 5700 3780 5704 3836
rect 5640 3776 5704 3780
rect 5720 3836 5784 3840
rect 5720 3780 5724 3836
rect 5724 3780 5780 3836
rect 5780 3780 5784 3836
rect 5720 3776 5784 3780
rect 2084 3292 2148 3296
rect 2084 3236 2088 3292
rect 2088 3236 2144 3292
rect 2144 3236 2148 3292
rect 2084 3232 2148 3236
rect 2164 3292 2228 3296
rect 2164 3236 2168 3292
rect 2168 3236 2224 3292
rect 2224 3236 2228 3292
rect 2164 3232 2228 3236
rect 2244 3292 2308 3296
rect 2244 3236 2248 3292
rect 2248 3236 2304 3292
rect 2304 3236 2308 3292
rect 2244 3232 2308 3236
rect 2324 3292 2388 3296
rect 2324 3236 2328 3292
rect 2328 3236 2384 3292
rect 2384 3236 2388 3292
rect 2324 3232 2388 3236
rect 4348 3292 4412 3296
rect 4348 3236 4352 3292
rect 4352 3236 4408 3292
rect 4408 3236 4412 3292
rect 4348 3232 4412 3236
rect 4428 3292 4492 3296
rect 4428 3236 4432 3292
rect 4432 3236 4488 3292
rect 4488 3236 4492 3292
rect 4428 3232 4492 3236
rect 4508 3292 4572 3296
rect 4508 3236 4512 3292
rect 4512 3236 4568 3292
rect 4568 3236 4572 3292
rect 4508 3232 4572 3236
rect 4588 3292 4652 3296
rect 4588 3236 4592 3292
rect 4592 3236 4648 3292
rect 4648 3236 4652 3292
rect 4588 3232 4652 3236
rect 6612 3292 6676 3296
rect 6612 3236 6616 3292
rect 6616 3236 6672 3292
rect 6672 3236 6676 3292
rect 6612 3232 6676 3236
rect 6692 3292 6756 3296
rect 6692 3236 6696 3292
rect 6696 3236 6752 3292
rect 6752 3236 6756 3292
rect 6692 3232 6756 3236
rect 6772 3292 6836 3296
rect 6772 3236 6776 3292
rect 6776 3236 6832 3292
rect 6832 3236 6836 3292
rect 6772 3232 6836 3236
rect 6852 3292 6916 3296
rect 6852 3236 6856 3292
rect 6856 3236 6912 3292
rect 6912 3236 6916 3292
rect 6852 3232 6916 3236
rect 3216 2748 3280 2752
rect 3216 2692 3220 2748
rect 3220 2692 3276 2748
rect 3276 2692 3280 2748
rect 3216 2688 3280 2692
rect 3296 2748 3360 2752
rect 3296 2692 3300 2748
rect 3300 2692 3356 2748
rect 3356 2692 3360 2748
rect 3296 2688 3360 2692
rect 3376 2748 3440 2752
rect 3376 2692 3380 2748
rect 3380 2692 3436 2748
rect 3436 2692 3440 2748
rect 3376 2688 3440 2692
rect 3456 2748 3520 2752
rect 3456 2692 3460 2748
rect 3460 2692 3516 2748
rect 3516 2692 3520 2748
rect 3456 2688 3520 2692
rect 5480 2748 5544 2752
rect 5480 2692 5484 2748
rect 5484 2692 5540 2748
rect 5540 2692 5544 2748
rect 5480 2688 5544 2692
rect 5560 2748 5624 2752
rect 5560 2692 5564 2748
rect 5564 2692 5620 2748
rect 5620 2692 5624 2748
rect 5560 2688 5624 2692
rect 5640 2748 5704 2752
rect 5640 2692 5644 2748
rect 5644 2692 5700 2748
rect 5700 2692 5704 2748
rect 5640 2688 5704 2692
rect 5720 2748 5784 2752
rect 5720 2692 5724 2748
rect 5724 2692 5780 2748
rect 5780 2692 5784 2748
rect 5720 2688 5784 2692
rect 2084 2204 2148 2208
rect 2084 2148 2088 2204
rect 2088 2148 2144 2204
rect 2144 2148 2148 2204
rect 2084 2144 2148 2148
rect 2164 2204 2228 2208
rect 2164 2148 2168 2204
rect 2168 2148 2224 2204
rect 2224 2148 2228 2204
rect 2164 2144 2228 2148
rect 2244 2204 2308 2208
rect 2244 2148 2248 2204
rect 2248 2148 2304 2204
rect 2304 2148 2308 2204
rect 2244 2144 2308 2148
rect 2324 2204 2388 2208
rect 2324 2148 2328 2204
rect 2328 2148 2384 2204
rect 2384 2148 2388 2204
rect 2324 2144 2388 2148
rect 4348 2204 4412 2208
rect 4348 2148 4352 2204
rect 4352 2148 4408 2204
rect 4408 2148 4412 2204
rect 4348 2144 4412 2148
rect 4428 2204 4492 2208
rect 4428 2148 4432 2204
rect 4432 2148 4488 2204
rect 4488 2148 4492 2204
rect 4428 2144 4492 2148
rect 4508 2204 4572 2208
rect 4508 2148 4512 2204
rect 4512 2148 4568 2204
rect 4568 2148 4572 2204
rect 4508 2144 4572 2148
rect 4588 2204 4652 2208
rect 4588 2148 4592 2204
rect 4592 2148 4648 2204
rect 4648 2148 4652 2204
rect 4588 2144 4652 2148
rect 6612 2204 6676 2208
rect 6612 2148 6616 2204
rect 6616 2148 6672 2204
rect 6672 2148 6676 2204
rect 6612 2144 6676 2148
rect 6692 2204 6756 2208
rect 6692 2148 6696 2204
rect 6696 2148 6752 2204
rect 6752 2148 6756 2204
rect 6692 2144 6756 2148
rect 6772 2204 6836 2208
rect 6772 2148 6776 2204
rect 6776 2148 6832 2204
rect 6832 2148 6836 2204
rect 6772 2144 6836 2148
rect 6852 2204 6916 2208
rect 6852 2148 6856 2204
rect 6856 2148 6912 2204
rect 6912 2148 6916 2204
rect 6852 2144 6916 2148
<< metal4 >>
rect 2076 14176 2396 14736
rect 2076 14112 2084 14176
rect 2148 14112 2164 14176
rect 2228 14112 2244 14176
rect 2308 14112 2324 14176
rect 2388 14112 2396 14176
rect 2076 13088 2396 14112
rect 2076 13024 2084 13088
rect 2148 13024 2164 13088
rect 2228 13024 2244 13088
rect 2308 13024 2324 13088
rect 2388 13024 2396 13088
rect 2076 12000 2396 13024
rect 2076 11936 2084 12000
rect 2148 11936 2164 12000
rect 2228 11936 2244 12000
rect 2308 11936 2324 12000
rect 2388 11936 2396 12000
rect 2076 10912 2396 11936
rect 2076 10848 2084 10912
rect 2148 10848 2164 10912
rect 2228 10848 2244 10912
rect 2308 10848 2324 10912
rect 2388 10848 2396 10912
rect 2076 9824 2396 10848
rect 2076 9760 2084 9824
rect 2148 9760 2164 9824
rect 2228 9760 2244 9824
rect 2308 9760 2324 9824
rect 2388 9760 2396 9824
rect 2076 8736 2396 9760
rect 2076 8672 2084 8736
rect 2148 8672 2164 8736
rect 2228 8672 2244 8736
rect 2308 8672 2324 8736
rect 2388 8672 2396 8736
rect 2076 7648 2396 8672
rect 2076 7584 2084 7648
rect 2148 7584 2164 7648
rect 2228 7584 2244 7648
rect 2308 7584 2324 7648
rect 2388 7584 2396 7648
rect 2076 6560 2396 7584
rect 2076 6496 2084 6560
rect 2148 6496 2164 6560
rect 2228 6496 2244 6560
rect 2308 6496 2324 6560
rect 2388 6496 2396 6560
rect 2076 5472 2396 6496
rect 2076 5408 2084 5472
rect 2148 5408 2164 5472
rect 2228 5408 2244 5472
rect 2308 5408 2324 5472
rect 2388 5408 2396 5472
rect 2076 4384 2396 5408
rect 2076 4320 2084 4384
rect 2148 4320 2164 4384
rect 2228 4320 2244 4384
rect 2308 4320 2324 4384
rect 2388 4320 2396 4384
rect 2076 3296 2396 4320
rect 2076 3232 2084 3296
rect 2148 3232 2164 3296
rect 2228 3232 2244 3296
rect 2308 3232 2324 3296
rect 2388 3232 2396 3296
rect 2076 2208 2396 3232
rect 2076 2144 2084 2208
rect 2148 2144 2164 2208
rect 2228 2144 2244 2208
rect 2308 2144 2324 2208
rect 2388 2144 2396 2208
rect 2076 2128 2396 2144
rect 3208 14720 3528 14736
rect 3208 14656 3216 14720
rect 3280 14656 3296 14720
rect 3360 14656 3376 14720
rect 3440 14656 3456 14720
rect 3520 14656 3528 14720
rect 3208 13632 3528 14656
rect 3208 13568 3216 13632
rect 3280 13568 3296 13632
rect 3360 13568 3376 13632
rect 3440 13568 3456 13632
rect 3520 13568 3528 13632
rect 3208 12544 3528 13568
rect 3208 12480 3216 12544
rect 3280 12480 3296 12544
rect 3360 12480 3376 12544
rect 3440 12480 3456 12544
rect 3520 12480 3528 12544
rect 3208 11456 3528 12480
rect 3208 11392 3216 11456
rect 3280 11392 3296 11456
rect 3360 11392 3376 11456
rect 3440 11392 3456 11456
rect 3520 11392 3528 11456
rect 3208 10368 3528 11392
rect 3208 10304 3216 10368
rect 3280 10304 3296 10368
rect 3360 10304 3376 10368
rect 3440 10304 3456 10368
rect 3520 10304 3528 10368
rect 3208 9280 3528 10304
rect 3208 9216 3216 9280
rect 3280 9216 3296 9280
rect 3360 9216 3376 9280
rect 3440 9216 3456 9280
rect 3520 9216 3528 9280
rect 3208 8192 3528 9216
rect 3208 8128 3216 8192
rect 3280 8128 3296 8192
rect 3360 8128 3376 8192
rect 3440 8128 3456 8192
rect 3520 8128 3528 8192
rect 3208 7104 3528 8128
rect 3208 7040 3216 7104
rect 3280 7040 3296 7104
rect 3360 7040 3376 7104
rect 3440 7040 3456 7104
rect 3520 7040 3528 7104
rect 3208 6016 3528 7040
rect 3208 5952 3216 6016
rect 3280 5952 3296 6016
rect 3360 5952 3376 6016
rect 3440 5952 3456 6016
rect 3520 5952 3528 6016
rect 3208 4928 3528 5952
rect 3208 4864 3216 4928
rect 3280 4864 3296 4928
rect 3360 4864 3376 4928
rect 3440 4864 3456 4928
rect 3520 4864 3528 4928
rect 3208 3840 3528 4864
rect 3208 3776 3216 3840
rect 3280 3776 3296 3840
rect 3360 3776 3376 3840
rect 3440 3776 3456 3840
rect 3520 3776 3528 3840
rect 3208 2752 3528 3776
rect 3208 2688 3216 2752
rect 3280 2688 3296 2752
rect 3360 2688 3376 2752
rect 3440 2688 3456 2752
rect 3520 2688 3528 2752
rect 3208 2128 3528 2688
rect 4340 14176 4660 14736
rect 4340 14112 4348 14176
rect 4412 14112 4428 14176
rect 4492 14112 4508 14176
rect 4572 14112 4588 14176
rect 4652 14112 4660 14176
rect 4340 13088 4660 14112
rect 4340 13024 4348 13088
rect 4412 13024 4428 13088
rect 4492 13024 4508 13088
rect 4572 13024 4588 13088
rect 4652 13024 4660 13088
rect 4340 12000 4660 13024
rect 4340 11936 4348 12000
rect 4412 11936 4428 12000
rect 4492 11936 4508 12000
rect 4572 11936 4588 12000
rect 4652 11936 4660 12000
rect 4340 10912 4660 11936
rect 4340 10848 4348 10912
rect 4412 10848 4428 10912
rect 4492 10848 4508 10912
rect 4572 10848 4588 10912
rect 4652 10848 4660 10912
rect 4340 9824 4660 10848
rect 4340 9760 4348 9824
rect 4412 9760 4428 9824
rect 4492 9760 4508 9824
rect 4572 9760 4588 9824
rect 4652 9760 4660 9824
rect 4340 8736 4660 9760
rect 4340 8672 4348 8736
rect 4412 8672 4428 8736
rect 4492 8672 4508 8736
rect 4572 8672 4588 8736
rect 4652 8672 4660 8736
rect 4340 7648 4660 8672
rect 4340 7584 4348 7648
rect 4412 7584 4428 7648
rect 4492 7584 4508 7648
rect 4572 7584 4588 7648
rect 4652 7584 4660 7648
rect 4340 6560 4660 7584
rect 4340 6496 4348 6560
rect 4412 6496 4428 6560
rect 4492 6496 4508 6560
rect 4572 6496 4588 6560
rect 4652 6496 4660 6560
rect 4340 5472 4660 6496
rect 4340 5408 4348 5472
rect 4412 5408 4428 5472
rect 4492 5408 4508 5472
rect 4572 5408 4588 5472
rect 4652 5408 4660 5472
rect 4340 4384 4660 5408
rect 4340 4320 4348 4384
rect 4412 4320 4428 4384
rect 4492 4320 4508 4384
rect 4572 4320 4588 4384
rect 4652 4320 4660 4384
rect 4340 3296 4660 4320
rect 4340 3232 4348 3296
rect 4412 3232 4428 3296
rect 4492 3232 4508 3296
rect 4572 3232 4588 3296
rect 4652 3232 4660 3296
rect 4340 2208 4660 3232
rect 4340 2144 4348 2208
rect 4412 2144 4428 2208
rect 4492 2144 4508 2208
rect 4572 2144 4588 2208
rect 4652 2144 4660 2208
rect 4340 2128 4660 2144
rect 5472 14720 5792 14736
rect 5472 14656 5480 14720
rect 5544 14656 5560 14720
rect 5624 14656 5640 14720
rect 5704 14656 5720 14720
rect 5784 14656 5792 14720
rect 5472 13632 5792 14656
rect 5472 13568 5480 13632
rect 5544 13568 5560 13632
rect 5624 13568 5640 13632
rect 5704 13568 5720 13632
rect 5784 13568 5792 13632
rect 5472 12544 5792 13568
rect 5472 12480 5480 12544
rect 5544 12480 5560 12544
rect 5624 12480 5640 12544
rect 5704 12480 5720 12544
rect 5784 12480 5792 12544
rect 5472 11456 5792 12480
rect 5472 11392 5480 11456
rect 5544 11392 5560 11456
rect 5624 11392 5640 11456
rect 5704 11392 5720 11456
rect 5784 11392 5792 11456
rect 5472 10368 5792 11392
rect 5472 10304 5480 10368
rect 5544 10304 5560 10368
rect 5624 10304 5640 10368
rect 5704 10304 5720 10368
rect 5784 10304 5792 10368
rect 5472 9280 5792 10304
rect 5472 9216 5480 9280
rect 5544 9216 5560 9280
rect 5624 9216 5640 9280
rect 5704 9216 5720 9280
rect 5784 9216 5792 9280
rect 5472 8192 5792 9216
rect 5472 8128 5480 8192
rect 5544 8128 5560 8192
rect 5624 8128 5640 8192
rect 5704 8128 5720 8192
rect 5784 8128 5792 8192
rect 5472 7104 5792 8128
rect 5472 7040 5480 7104
rect 5544 7040 5560 7104
rect 5624 7040 5640 7104
rect 5704 7040 5720 7104
rect 5784 7040 5792 7104
rect 5472 6016 5792 7040
rect 5472 5952 5480 6016
rect 5544 5952 5560 6016
rect 5624 5952 5640 6016
rect 5704 5952 5720 6016
rect 5784 5952 5792 6016
rect 5472 4928 5792 5952
rect 5472 4864 5480 4928
rect 5544 4864 5560 4928
rect 5624 4864 5640 4928
rect 5704 4864 5720 4928
rect 5784 4864 5792 4928
rect 5472 3840 5792 4864
rect 5472 3776 5480 3840
rect 5544 3776 5560 3840
rect 5624 3776 5640 3840
rect 5704 3776 5720 3840
rect 5784 3776 5792 3840
rect 5472 2752 5792 3776
rect 5472 2688 5480 2752
rect 5544 2688 5560 2752
rect 5624 2688 5640 2752
rect 5704 2688 5720 2752
rect 5784 2688 5792 2752
rect 5472 2128 5792 2688
rect 6604 14176 6924 14736
rect 6604 14112 6612 14176
rect 6676 14112 6692 14176
rect 6756 14112 6772 14176
rect 6836 14112 6852 14176
rect 6916 14112 6924 14176
rect 6604 13088 6924 14112
rect 6604 13024 6612 13088
rect 6676 13024 6692 13088
rect 6756 13024 6772 13088
rect 6836 13024 6852 13088
rect 6916 13024 6924 13088
rect 6604 12000 6924 13024
rect 6604 11936 6612 12000
rect 6676 11936 6692 12000
rect 6756 11936 6772 12000
rect 6836 11936 6852 12000
rect 6916 11936 6924 12000
rect 6604 10912 6924 11936
rect 6604 10848 6612 10912
rect 6676 10848 6692 10912
rect 6756 10848 6772 10912
rect 6836 10848 6852 10912
rect 6916 10848 6924 10912
rect 6604 9824 6924 10848
rect 6604 9760 6612 9824
rect 6676 9760 6692 9824
rect 6756 9760 6772 9824
rect 6836 9760 6852 9824
rect 6916 9760 6924 9824
rect 6604 8736 6924 9760
rect 6604 8672 6612 8736
rect 6676 8672 6692 8736
rect 6756 8672 6772 8736
rect 6836 8672 6852 8736
rect 6916 8672 6924 8736
rect 6604 7648 6924 8672
rect 6604 7584 6612 7648
rect 6676 7584 6692 7648
rect 6756 7584 6772 7648
rect 6836 7584 6852 7648
rect 6916 7584 6924 7648
rect 6604 6560 6924 7584
rect 6604 6496 6612 6560
rect 6676 6496 6692 6560
rect 6756 6496 6772 6560
rect 6836 6496 6852 6560
rect 6916 6496 6924 6560
rect 6604 5472 6924 6496
rect 6604 5408 6612 5472
rect 6676 5408 6692 5472
rect 6756 5408 6772 5472
rect 6836 5408 6852 5472
rect 6916 5408 6924 5472
rect 6604 4384 6924 5408
rect 6604 4320 6612 4384
rect 6676 4320 6692 4384
rect 6756 4320 6772 4384
rect 6836 4320 6852 4384
rect 6916 4320 6924 4384
rect 6604 3296 6924 4320
rect 6604 3232 6612 3296
rect 6676 3232 6692 3296
rect 6756 3232 6772 3296
rect 6836 3232 6852 3296
rect 6916 3232 6924 3296
rect 6604 2208 6924 3232
rect 6604 2144 6612 2208
rect 6676 2144 6692 2208
rect 6756 2144 6772 2208
rect 6836 2144 6852 2208
rect 6916 2144 6924 2208
rect 6604 2128 6924 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 7820 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 7820 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 7820 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2208 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1605641404
transform 1 0 2116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_28
timestamp 1605641404
transform 1 0 3680 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_40
timestamp 1605641404
transform 1 0 4784 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_52
timestamp 1605641404
transform 1 0 5888 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1605641404
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 7820 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1605641404
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 7820 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_62
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 7820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2576 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_25
timestamp 1605641404
transform 1 0 3404 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5612 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_48
timestamp 1605641404
transform 1 0 5520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_37
timestamp 1605641404
transform 1 0 4508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_49
timestamp 1605641404
transform 1 0 5612 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_62
timestamp 1605641404
transform 1 0 6808 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 7820 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 7820 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1605641404
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1605641404
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 7820 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1605641404
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2576 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_19
timestamp 1605641404
transform 1 0 2852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1605641404
transform 1 0 3956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1605641404
transform 1 0 5060 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_55
timestamp 1605641404
transform 1 0 6164 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 7820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2024 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_9
timestamp 1605641404
transform 1 0 1932 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_14
timestamp 1605641404
transform 1 0 2392 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_26
timestamp 1605641404
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1605641404
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1605641404
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1605641404
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 7820 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1605641404
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1605641404
transform 1 0 1656 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_19
timestamp 1605641404
transform 1 0 2852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1605641404
transform 1 0 3956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1605641404
transform 1 0 5060 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_55
timestamp 1605641404
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 7820 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1605641404
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1605641404
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1605641404
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1605641404
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 7820 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1605641404
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1605641404
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1605641404
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1605641404
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1605641404
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1605641404
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1605641404
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1605641404
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 7820 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 7820 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1605641404
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1605641404
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1605641404
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1605641404
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1605641404
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 7820 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1605641404
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1605641404
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1605641404
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 7820 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1605641404
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1605641404
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1605641404
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1605641404
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1605641404
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 7820 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1605641404
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1605641404
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1605641404
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1605641404
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 7820 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1605641404
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1605641404
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1605641404
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1605641404
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1605641404
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1605641404
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 7820 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 7820 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_68
timestamp 1605641404
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1605641404
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1605641404
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1605641404
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1605641404
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1605641404
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_63
timestamp 1605641404
transform 1 0 6900 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 7820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1605641404
transform 1 0 7452 0 -1 14688
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 11840 480 11960 6 IO_ISOL_N
port 0 nsew default input
rlabel metal2 s 3330 0 3386 480 6 ccff_head
port 1 nsew default input
rlabel metal2 s 5630 0 5686 480 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 8520 8440 9000 8560 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 3 nsew default tristate
rlabel metal3 s 0 15240 480 15360 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 4 nsew default input
rlabel metal2 s 7838 0 7894 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 5 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 left_width_0_height_0__pin_0_
port 6 nsew default input
rlabel metal3 s 0 1640 480 1760 6 left_width_0_height_0__pin_1_lower
port 7 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 left_width_0_height_0__pin_1_upper
port 8 nsew default tristate
rlabel metal2 s 1122 0 1178 480 6 prog_clk
port 9 nsew default input
rlabel metal4 s 2076 2128 2396 14736 6 VPWR
port 10 nsew default input
rlabel metal4 s 3208 2128 3528 14736 6 VGND
port 11 nsew default input
<< properties >>
string FIXED_BBOX 0 0 9000 15360
<< end >>
