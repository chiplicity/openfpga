magic
tech sky130A
magscale 1 2
timestamp 1604668711
<< locali >>
rect 10241 25347 10275 25449
rect 12173 25143 12207 25313
rect 14197 25279 14231 25449
rect 22201 25347 22235 25449
rect 9505 23579 9539 23749
rect 4445 23103 4479 23205
rect 17693 22423 17727 22593
rect 3341 20791 3375 20893
rect 23305 16983 23339 17085
<< viali >>
rect 1409 25449 1443 25483
rect 2789 25449 2823 25483
rect 4261 25449 4295 25483
rect 5641 25449 5675 25483
rect 7573 25449 7607 25483
rect 8033 25449 8067 25483
rect 10241 25449 10275 25483
rect 10517 25449 10551 25483
rect 12633 25449 12667 25483
rect 14197 25449 14231 25483
rect 14473 25449 14507 25483
rect 17325 25449 17359 25483
rect 20177 25449 20211 25483
rect 22201 25449 22235 25483
rect 22385 25449 22419 25483
rect 23029 25449 23063 25483
rect 4077 25313 4111 25347
rect 6285 25313 6319 25347
rect 7113 25313 7147 25347
rect 8493 25313 8527 25347
rect 9965 25313 9999 25347
rect 10241 25313 10275 25347
rect 11345 25313 11379 25347
rect 12173 25313 12207 25347
rect 12449 25313 12483 25347
rect 13001 25313 13035 25347
rect 2881 25245 2915 25279
rect 3065 25245 3099 25279
rect 5733 25245 5767 25279
rect 5825 25245 5859 25279
rect 8585 25245 8619 25279
rect 8677 25245 8711 25279
rect 11437 25245 11471 25279
rect 11621 25245 11655 25279
rect 3801 25177 3835 25211
rect 5273 25177 5307 25211
rect 7297 25177 7331 25211
rect 10977 25177 11011 25211
rect 21557 25381 21591 25415
rect 23765 25381 23799 25415
rect 24409 25381 24443 25415
rect 14289 25313 14323 25347
rect 15853 25313 15887 25347
rect 15945 25313 15979 25347
rect 17141 25313 17175 25347
rect 18429 25313 18463 25347
rect 19993 25313 20027 25347
rect 21741 25313 21775 25347
rect 22201 25313 22235 25347
rect 22845 25313 22879 25347
rect 24501 25313 24535 25347
rect 25605 25313 25639 25347
rect 13093 25245 13127 25279
rect 13277 25245 13311 25279
rect 14197 25245 14231 25279
rect 16129 25245 16163 25279
rect 24685 25245 24719 25279
rect 15485 25177 15519 25211
rect 18613 25177 18647 25211
rect 21925 25177 21959 25211
rect 25789 25177 25823 25211
rect 1961 25109 1995 25143
rect 2329 25109 2363 25143
rect 2421 25109 2455 25143
rect 3433 25109 3467 25143
rect 4629 25109 4663 25143
rect 5089 25109 5123 25143
rect 6653 25109 6687 25143
rect 8125 25109 8159 25143
rect 9137 25109 9171 25143
rect 10149 25109 10183 25143
rect 11989 25109 12023 25143
rect 12173 25109 12207 25143
rect 15117 25109 15151 25143
rect 16589 25109 16623 25143
rect 18153 25109 18187 25143
rect 22661 25109 22695 25143
rect 24041 25109 24075 25143
rect 25237 25109 25271 25143
rect 10701 24905 10735 24939
rect 13001 24905 13035 24939
rect 16129 24905 16163 24939
rect 17509 24905 17543 24939
rect 18521 24905 18555 24939
rect 24777 24905 24811 24939
rect 21465 24837 21499 24871
rect 2145 24769 2179 24803
rect 2697 24769 2731 24803
rect 7297 24769 7331 24803
rect 7481 24769 7515 24803
rect 11897 24769 11931 24803
rect 13645 24769 13679 24803
rect 14381 24769 14415 24803
rect 15669 24769 15703 24803
rect 19993 24769 20027 24803
rect 21097 24769 21131 24803
rect 22569 24769 22603 24803
rect 24133 24769 24167 24803
rect 24225 24769 24259 24803
rect 25053 24769 25087 24803
rect 1961 24701 1995 24735
rect 3157 24701 3191 24735
rect 3424 24701 3458 24735
rect 5273 24701 5307 24735
rect 5641 24701 5675 24735
rect 6285 24701 6319 24735
rect 8217 24701 8251 24735
rect 8493 24701 8527 24735
rect 11345 24701 11379 24735
rect 12265 24701 12299 24735
rect 14933 24701 14967 24735
rect 16405 24701 16439 24735
rect 16589 24701 16623 24735
rect 18061 24701 18095 24735
rect 19073 24701 19107 24735
rect 22385 24701 22419 24735
rect 25237 24701 25271 24735
rect 6653 24633 6687 24667
rect 8760 24633 8794 24667
rect 11069 24633 11103 24667
rect 12909 24633 12943 24667
rect 15393 24633 15427 24667
rect 20913 24633 20947 24667
rect 21925 24633 21959 24667
rect 22477 24633 22511 24667
rect 23489 24633 23523 24667
rect 24041 24633 24075 24667
rect 25789 24633 25823 24667
rect 1593 24565 1627 24599
rect 2053 24565 2087 24599
rect 3065 24565 3099 24599
rect 4537 24565 4571 24599
rect 5825 24565 5859 24599
rect 6837 24565 6871 24599
rect 7205 24565 7239 24599
rect 9873 24565 9907 24599
rect 11529 24565 11563 24599
rect 13369 24565 13403 24599
rect 13461 24565 13495 24599
rect 14013 24565 14047 24599
rect 15025 24565 15059 24599
rect 15485 24565 15519 24599
rect 16773 24565 16807 24599
rect 17141 24565 17175 24599
rect 18245 24565 18279 24599
rect 18889 24565 18923 24599
rect 19257 24565 19291 24599
rect 20269 24565 20303 24599
rect 20453 24565 20487 24599
rect 20821 24565 20855 24599
rect 22017 24565 22051 24599
rect 23121 24565 23155 24599
rect 23673 24565 23707 24599
rect 25421 24565 25455 24599
rect 1869 24361 1903 24395
rect 2329 24361 2363 24395
rect 3893 24361 3927 24395
rect 4537 24361 4571 24395
rect 7665 24361 7699 24395
rect 8125 24361 8159 24395
rect 8769 24361 8803 24395
rect 10149 24361 10183 24395
rect 10701 24361 10735 24395
rect 11161 24361 11195 24395
rect 11805 24361 11839 24395
rect 14289 24361 14323 24395
rect 18337 24361 18371 24395
rect 19349 24361 19383 24395
rect 20085 24361 20119 24395
rect 23121 24361 23155 24395
rect 24317 24361 24351 24395
rect 25237 24361 25271 24395
rect 2789 24293 2823 24327
rect 2881 24293 2915 24327
rect 11069 24293 11103 24327
rect 12633 24293 12667 24327
rect 17785 24293 17819 24327
rect 22845 24293 22879 24327
rect 1409 24225 1443 24259
rect 6000 24225 6034 24259
rect 8217 24225 8251 24259
rect 12725 24225 12759 24259
rect 14105 24225 14139 24259
rect 16129 24225 16163 24259
rect 17693 24225 17727 24259
rect 19165 24225 19199 24259
rect 21281 24225 21315 24259
rect 22109 24225 22143 24259
rect 23673 24225 23707 24259
rect 25329 24225 25363 24259
rect 3065 24157 3099 24191
rect 4629 24157 4663 24191
rect 4813 24157 4847 24191
rect 5733 24157 5767 24191
rect 9689 24157 9723 24191
rect 11345 24157 11379 24191
rect 12173 24157 12207 24191
rect 12817 24157 12851 24191
rect 15577 24157 15611 24191
rect 16221 24157 16255 24191
rect 16313 24157 16347 24191
rect 17233 24157 17267 24191
rect 17877 24157 17911 24191
rect 22201 24157 22235 24191
rect 22293 24157 22327 24191
rect 23765 24157 23799 24191
rect 23857 24157 23891 24191
rect 25421 24157 25455 24191
rect 5549 24089 5583 24123
rect 7113 24089 7147 24123
rect 21649 24089 21683 24123
rect 1593 24021 1627 24055
rect 2421 24021 2455 24055
rect 3525 24021 3559 24055
rect 4169 24021 4203 24055
rect 5273 24021 5307 24055
rect 8401 24021 8435 24055
rect 9137 24021 9171 24055
rect 12265 24021 12299 24055
rect 13277 24021 13311 24055
rect 14657 24021 14691 24055
rect 15025 24021 15059 24055
rect 15761 24021 15795 24055
rect 17325 24021 17359 24055
rect 19073 24021 19107 24055
rect 20545 24021 20579 24055
rect 21741 24021 21775 24055
rect 23305 24021 23339 24055
rect 24869 24021 24903 24055
rect 1593 23817 1627 23851
rect 1961 23817 1995 23851
rect 9321 23817 9355 23851
rect 11805 23817 11839 23851
rect 12633 23817 12667 23851
rect 14381 23817 14415 23851
rect 14933 23817 14967 23851
rect 16865 23817 16899 23851
rect 17417 23817 17451 23851
rect 17785 23817 17819 23851
rect 20085 23817 20119 23851
rect 23673 23817 23707 23851
rect 24961 23817 24995 23851
rect 25421 23817 25455 23851
rect 25789 23817 25823 23851
rect 5365 23749 5399 23783
rect 9505 23749 9539 23783
rect 9597 23749 9631 23783
rect 12173 23749 12207 23783
rect 18337 23749 18371 23783
rect 19349 23749 19383 23783
rect 19809 23749 19843 23783
rect 2329 23681 2363 23715
rect 2881 23681 2915 23715
rect 3065 23681 3099 23715
rect 3985 23681 4019 23715
rect 6377 23681 6411 23715
rect 8861 23681 8895 23715
rect 1409 23613 1443 23647
rect 2789 23613 2823 23647
rect 3801 23613 3835 23647
rect 4241 23613 4275 23647
rect 6837 23613 6871 23647
rect 8585 23613 8619 23647
rect 13001 23681 13035 23715
rect 18797 23681 18831 23715
rect 18981 23681 19015 23715
rect 20361 23681 20395 23715
rect 24133 23681 24167 23715
rect 24317 23681 24351 23715
rect 9781 23613 9815 23647
rect 10037 23613 10071 23647
rect 15485 23613 15519 23647
rect 15752 23613 15786 23647
rect 18705 23613 18739 23647
rect 19901 23613 19935 23647
rect 20913 23613 20947 23647
rect 21180 23613 21214 23647
rect 24041 23613 24075 23647
rect 25237 23613 25271 23647
rect 3525 23545 3559 23579
rect 8125 23545 8159 23579
rect 9505 23545 9539 23579
rect 13268 23545 13302 23579
rect 23029 23545 23063 23579
rect 2421 23477 2455 23511
rect 6009 23477 6043 23511
rect 7021 23477 7055 23511
rect 7389 23477 7423 23511
rect 8217 23477 8251 23511
rect 8677 23477 8711 23511
rect 11161 23477 11195 23511
rect 15301 23477 15335 23511
rect 20821 23477 20855 23511
rect 22293 23477 22327 23511
rect 23305 23477 23339 23511
rect 2881 23273 2915 23307
rect 4353 23273 4387 23307
rect 4721 23273 4755 23307
rect 6285 23273 6319 23307
rect 7573 23273 7607 23307
rect 8401 23273 8435 23307
rect 8493 23273 8527 23307
rect 9689 23273 9723 23307
rect 10793 23273 10827 23307
rect 11069 23273 11103 23307
rect 12909 23273 12943 23307
rect 18337 23273 18371 23307
rect 18797 23273 18831 23307
rect 19717 23273 19751 23307
rect 21465 23273 21499 23307
rect 22937 23273 22971 23307
rect 24409 23273 24443 23307
rect 24501 23273 24535 23307
rect 25145 23273 25179 23307
rect 4445 23205 4479 23239
rect 7849 23205 7883 23239
rect 9413 23205 9447 23239
rect 10149 23205 10183 23239
rect 11796 23205 11830 23239
rect 16396 23205 16430 23239
rect 19625 23205 19659 23239
rect 21802 23205 21836 23239
rect 1409 23137 1443 23171
rect 2789 23137 2823 23171
rect 3433 23137 3467 23171
rect 5172 23137 5206 23171
rect 10057 23137 10091 23171
rect 11529 23137 11563 23171
rect 14105 23137 14139 23171
rect 3065 23069 3099 23103
rect 4445 23069 4479 23103
rect 4905 23069 4939 23103
rect 8677 23069 8711 23103
rect 10241 23069 10275 23103
rect 15117 23069 15151 23103
rect 16129 23069 16163 23103
rect 19165 23069 19199 23103
rect 19901 23069 19935 23103
rect 21557 23069 21591 23103
rect 24593 23069 24627 23103
rect 1961 23001 1995 23035
rect 8033 23001 8067 23035
rect 9137 23001 9171 23035
rect 17509 23001 17543 23035
rect 19257 23001 19291 23035
rect 23949 23001 23983 23035
rect 2329 22933 2363 22967
rect 2421 22933 2455 22967
rect 3801 22933 3835 22967
rect 6929 22933 6963 22967
rect 13553 22933 13587 22967
rect 14289 22933 14323 22967
rect 14657 22933 14691 22967
rect 15485 22933 15519 22967
rect 15945 22933 15979 22967
rect 20269 22933 20303 22967
rect 23489 22933 23523 22967
rect 24041 22933 24075 22967
rect 25513 22933 25547 22967
rect 3157 22729 3191 22763
rect 3341 22729 3375 22763
rect 4445 22729 4479 22763
rect 6561 22729 6595 22763
rect 7941 22729 7975 22763
rect 9413 22729 9447 22763
rect 11529 22729 11563 22763
rect 11897 22729 11931 22763
rect 13093 22729 13127 22763
rect 16405 22729 16439 22763
rect 19073 22729 19107 22763
rect 21005 22729 21039 22763
rect 22661 22729 22695 22763
rect 25053 22729 25087 22763
rect 25421 22729 25455 22763
rect 1777 22661 1811 22695
rect 2881 22661 2915 22695
rect 4905 22661 4939 22695
rect 5917 22661 5951 22695
rect 10517 22661 10551 22695
rect 15301 22661 15335 22695
rect 23673 22661 23707 22695
rect 2421 22593 2455 22627
rect 3893 22593 3927 22627
rect 5365 22593 5399 22627
rect 5457 22593 5491 22627
rect 7573 22593 7607 22627
rect 8033 22593 8067 22627
rect 9965 22593 9999 22627
rect 10977 22593 11011 22627
rect 11069 22593 11103 22627
rect 16957 22593 16991 22627
rect 17693 22593 17727 22627
rect 18613 22593 18647 22627
rect 22017 22593 22051 22627
rect 23489 22593 23523 22627
rect 24225 22593 24259 22627
rect 2237 22525 2271 22559
rect 3709 22525 3743 22559
rect 3801 22525 3835 22559
rect 5273 22525 5307 22559
rect 6837 22525 6871 22559
rect 12909 22525 12943 22559
rect 13921 22525 13955 22559
rect 16129 22525 16163 22559
rect 16865 22525 16899 22559
rect 1685 22457 1719 22491
rect 2145 22457 2179 22491
rect 8278 22457 8312 22491
rect 14166 22457 14200 22491
rect 16773 22457 16807 22491
rect 17509 22457 17543 22491
rect 18429 22525 18463 22559
rect 19625 22525 19659 22559
rect 21557 22525 21591 22559
rect 22477 22525 22511 22559
rect 24133 22525 24167 22559
rect 25237 22525 25271 22559
rect 25789 22525 25823 22559
rect 19870 22457 19904 22491
rect 24041 22457 24075 22491
rect 4813 22389 4847 22423
rect 7021 22389 7055 22423
rect 10333 22389 10367 22423
rect 10885 22389 10919 22423
rect 12725 22389 12759 22423
rect 13461 22389 13495 22423
rect 13737 22389 13771 22423
rect 17693 22389 17727 22423
rect 17785 22389 17819 22423
rect 18061 22389 18095 22423
rect 18521 22389 18555 22423
rect 19441 22389 19475 22423
rect 22293 22389 22327 22423
rect 23121 22389 23155 22423
rect 24685 22389 24719 22423
rect 1961 22185 1995 22219
rect 3065 22185 3099 22219
rect 3433 22185 3467 22219
rect 5181 22185 5215 22219
rect 5457 22185 5491 22219
rect 8585 22185 8619 22219
rect 9505 22185 9539 22219
rect 10333 22185 10367 22219
rect 10977 22185 11011 22219
rect 16221 22185 16255 22219
rect 16773 22185 16807 22219
rect 22201 22185 22235 22219
rect 23397 22185 23431 22219
rect 24777 22185 24811 22219
rect 4445 22117 4479 22151
rect 6460 22117 6494 22151
rect 9137 22117 9171 22151
rect 10241 22117 10275 22151
rect 11704 22117 11738 22151
rect 17141 22117 17175 22151
rect 23857 22117 23891 22151
rect 2053 22049 2087 22083
rect 5917 22049 5951 22083
rect 11345 22049 11379 22083
rect 14105 22049 14139 22083
rect 15669 22049 15703 22083
rect 17785 22049 17819 22083
rect 18593 22049 18627 22083
rect 23305 22049 23339 22083
rect 23765 22049 23799 22083
rect 24961 22049 24995 22083
rect 2145 21981 2179 22015
rect 4537 21981 4571 22015
rect 4721 21981 4755 22015
rect 6193 21981 6227 22015
rect 10517 21981 10551 22015
rect 11437 21981 11471 22015
rect 14657 21981 14691 22015
rect 17233 21981 17267 22015
rect 17417 21981 17451 22015
rect 18337 21981 18371 22015
rect 22293 21981 22327 22015
rect 22477 21981 22511 22015
rect 24041 21981 24075 22015
rect 4077 21913 4111 21947
rect 13369 21913 13403 21947
rect 14289 21913 14323 21947
rect 15117 21913 15151 21947
rect 15853 21913 15887 21947
rect 19717 21913 19751 21947
rect 21557 21913 21591 21947
rect 25145 21913 25179 21947
rect 1593 21845 1627 21879
rect 2605 21845 2639 21879
rect 3709 21845 3743 21879
rect 7573 21845 7607 21879
rect 8125 21845 8159 21879
rect 9873 21845 9907 21879
rect 12817 21845 12851 21879
rect 13921 21845 13955 21879
rect 15485 21845 15519 21879
rect 16681 21845 16715 21879
rect 18245 21845 18279 21879
rect 20269 21845 20303 21879
rect 21833 21845 21867 21879
rect 24501 21845 24535 21879
rect 2605 21641 2639 21675
rect 4721 21641 4755 21675
rect 5273 21641 5307 21675
rect 5917 21641 5951 21675
rect 8309 21641 8343 21675
rect 10241 21641 10275 21675
rect 10609 21641 10643 21675
rect 11805 21641 11839 21675
rect 12265 21641 12299 21675
rect 13093 21641 13127 21675
rect 16405 21641 16439 21675
rect 17877 21641 17911 21675
rect 21465 21641 21499 21675
rect 22569 21641 22603 21675
rect 24777 21641 24811 21675
rect 25513 21641 25547 21675
rect 23765 21573 23799 21607
rect 2053 21505 2087 21539
rect 2145 21505 2179 21539
rect 7481 21505 7515 21539
rect 7849 21505 7883 21539
rect 9689 21505 9723 21539
rect 9873 21505 9907 21539
rect 11345 21505 11379 21539
rect 13277 21505 13311 21539
rect 15577 21505 15611 21539
rect 17049 21505 17083 21539
rect 20913 21505 20947 21539
rect 22017 21505 22051 21539
rect 24317 21505 24351 21539
rect 1961 21437 1995 21471
rect 3341 21437 3375 21471
rect 6653 21437 6687 21471
rect 7205 21437 7239 21471
rect 7297 21437 7331 21471
rect 8769 21437 8803 21471
rect 11253 21437 11287 21471
rect 12633 21437 12667 21471
rect 13533 21437 13567 21471
rect 15945 21437 15979 21471
rect 18981 21437 19015 21471
rect 24133 21437 24167 21471
rect 25329 21437 25363 21471
rect 25881 21437 25915 21471
rect 3608 21369 3642 21403
rect 9137 21369 9171 21403
rect 9597 21369 9631 21403
rect 11161 21369 11195 21403
rect 16865 21369 16899 21403
rect 19226 21369 19260 21403
rect 23121 21369 23155 21403
rect 25145 21369 25179 21403
rect 1593 21301 1627 21335
rect 3249 21301 3283 21335
rect 6285 21301 6319 21335
rect 6837 21301 6871 21335
rect 9229 21301 9263 21335
rect 10793 21301 10827 21335
rect 14657 21301 14691 21335
rect 16313 21301 16347 21335
rect 16773 21301 16807 21335
rect 17417 21301 17451 21335
rect 18337 21301 18371 21335
rect 18797 21301 18831 21335
rect 20361 21301 20395 21335
rect 21373 21301 21407 21335
rect 21833 21301 21867 21335
rect 21925 21301 21959 21335
rect 23397 21301 23431 21335
rect 24225 21301 24259 21335
rect 1409 21097 1443 21131
rect 1869 21097 1903 21131
rect 2237 21097 2271 21131
rect 2421 21097 2455 21131
rect 7389 21097 7423 21131
rect 7941 21097 7975 21131
rect 9321 21097 9355 21131
rect 9965 21097 9999 21131
rect 10241 21097 10275 21131
rect 10517 21097 10551 21131
rect 11897 21097 11931 21131
rect 12081 21097 12115 21131
rect 13369 21097 13403 21131
rect 13645 21097 13679 21131
rect 15853 21097 15887 21131
rect 16405 21097 16439 21131
rect 19073 21097 19107 21131
rect 19257 21097 19291 21131
rect 21281 21097 21315 21131
rect 22017 21097 22051 21131
rect 22293 21097 22327 21131
rect 24317 21097 24351 21131
rect 2789 21029 2823 21063
rect 6009 21029 6043 21063
rect 14013 21029 14047 21063
rect 15577 21029 15611 21063
rect 17040 21029 17074 21063
rect 18705 21029 18739 21063
rect 21373 21029 21407 21063
rect 4333 20961 4367 20995
rect 7297 20961 7331 20995
rect 8493 20961 8527 20995
rect 10885 20961 10919 20995
rect 12449 20961 12483 20995
rect 14105 20961 14139 20995
rect 15669 20961 15703 20995
rect 19625 20961 19659 20995
rect 20637 20961 20671 20995
rect 22753 20961 22787 20995
rect 24225 20961 24259 20995
rect 2881 20893 2915 20927
rect 2973 20893 3007 20927
rect 3341 20893 3375 20927
rect 4077 20893 4111 20927
rect 7573 20893 7607 20927
rect 10977 20893 11011 20927
rect 11069 20893 11103 20927
rect 12541 20893 12575 20927
rect 12725 20893 12759 20927
rect 14197 20893 14231 20927
rect 16773 20893 16807 20927
rect 19717 20893 19751 20927
rect 19809 20893 19843 20927
rect 21465 20893 21499 20927
rect 24409 20893 24443 20927
rect 25421 20893 25455 20927
rect 3801 20825 3835 20859
rect 6469 20825 6503 20859
rect 6929 20825 6963 20859
rect 8677 20825 8711 20859
rect 15117 20825 15151 20859
rect 18153 20825 18187 20859
rect 20269 20825 20303 20859
rect 22937 20825 22971 20859
rect 23489 20825 23523 20859
rect 3341 20757 3375 20791
rect 3525 20757 3559 20791
rect 5457 20757 5491 20791
rect 6745 20757 6779 20791
rect 8309 20757 8343 20791
rect 11529 20757 11563 20791
rect 14657 20757 14691 20791
rect 20913 20757 20947 20791
rect 23857 20757 23891 20791
rect 24961 20757 24995 20791
rect 25329 20757 25363 20791
rect 2053 20553 2087 20587
rect 4445 20553 4479 20587
rect 5825 20553 5859 20587
rect 6285 20553 6319 20587
rect 6837 20553 6871 20587
rect 9965 20553 9999 20587
rect 10609 20553 10643 20587
rect 11713 20553 11747 20587
rect 14381 20553 14415 20587
rect 18245 20553 18279 20587
rect 19165 20553 19199 20587
rect 20545 20553 20579 20587
rect 22385 20553 22419 20587
rect 23029 20553 23063 20587
rect 23489 20553 23523 20587
rect 25421 20553 25455 20587
rect 3433 20417 3467 20451
rect 5089 20417 5123 20451
rect 7297 20417 7331 20451
rect 7389 20417 7423 20451
rect 12449 20417 12483 20451
rect 19717 20417 19751 20451
rect 24133 20417 24167 20451
rect 24317 20417 24351 20451
rect 1434 20349 1468 20383
rect 3249 20349 3283 20383
rect 4905 20349 4939 20383
rect 8125 20349 8159 20383
rect 8585 20349 8619 20383
rect 10885 20349 10919 20383
rect 15393 20349 15427 20383
rect 17325 20349 17359 20383
rect 18061 20349 18095 20383
rect 18705 20349 18739 20383
rect 19533 20349 19567 20383
rect 21005 20349 21039 20383
rect 25053 20349 25087 20383
rect 25237 20349 25271 20383
rect 25789 20349 25823 20383
rect 3341 20281 3375 20315
rect 4169 20281 4203 20315
rect 8830 20281 8864 20315
rect 12694 20281 12728 20315
rect 15660 20281 15694 20315
rect 21272 20281 21306 20315
rect 24041 20281 24075 20315
rect 1593 20213 1627 20247
rect 2329 20213 2363 20247
rect 2789 20213 2823 20247
rect 2881 20213 2915 20247
rect 4813 20213 4847 20247
rect 5457 20213 5491 20247
rect 6653 20213 6687 20247
rect 7205 20213 7239 20247
rect 8493 20213 8527 20247
rect 11069 20213 11103 20247
rect 12081 20213 12115 20247
rect 13829 20213 13863 20247
rect 14841 20213 14875 20247
rect 15209 20213 15243 20247
rect 16773 20213 16807 20247
rect 17785 20213 17819 20247
rect 18981 20213 19015 20247
rect 19625 20213 19659 20247
rect 20913 20213 20947 20247
rect 23673 20213 23707 20247
rect 24685 20213 24719 20247
rect 2421 20009 2455 20043
rect 2881 20009 2915 20043
rect 4077 20009 4111 20043
rect 8125 20009 8159 20043
rect 11069 20009 11103 20043
rect 12173 20009 12207 20043
rect 13553 20009 13587 20043
rect 13645 20009 13679 20043
rect 14657 20009 14691 20043
rect 16865 20009 16899 20043
rect 17417 20009 17451 20043
rect 19717 20009 19751 20043
rect 21097 20009 21131 20043
rect 21557 20009 21591 20043
rect 24869 20009 24903 20043
rect 24961 20009 24995 20043
rect 4445 19941 4479 19975
rect 6092 19941 6126 19975
rect 7849 19941 7883 19975
rect 9934 19941 9968 19975
rect 20729 19941 20763 19975
rect 25513 19941 25547 19975
rect 1409 19873 1443 19907
rect 2789 19873 2823 19907
rect 5181 19873 5215 19907
rect 5825 19873 5859 19907
rect 8309 19873 8343 19907
rect 12449 19873 12483 19907
rect 14013 19873 14047 19907
rect 14105 19873 14139 19907
rect 15025 19873 15059 19907
rect 15669 19873 15703 19907
rect 17233 19873 17267 19907
rect 18604 19873 18638 19907
rect 20913 19873 20947 19907
rect 22284 19873 22318 19907
rect 3065 19805 3099 19839
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 9689 19805 9723 19839
rect 11621 19805 11655 19839
rect 12633 19805 12667 19839
rect 14289 19805 14323 19839
rect 15761 19805 15795 19839
rect 15945 19805 15979 19839
rect 18337 19805 18371 19839
rect 22017 19805 22051 19839
rect 24409 19805 24443 19839
rect 25145 19805 25179 19839
rect 1593 19737 1627 19771
rect 8861 19737 8895 19771
rect 23397 19737 23431 19771
rect 24501 19737 24535 19771
rect 1869 19669 1903 19703
rect 2237 19669 2271 19703
rect 3709 19669 3743 19703
rect 5549 19669 5583 19703
rect 7205 19669 7239 19703
rect 8493 19669 8527 19703
rect 9321 19669 9355 19703
rect 13185 19669 13219 19703
rect 15301 19669 15335 19703
rect 16405 19669 16439 19703
rect 18061 19669 18095 19703
rect 20269 19669 20303 19703
rect 21925 19669 21959 19703
rect 23949 19669 23983 19703
rect 2973 19465 3007 19499
rect 5181 19465 5215 19499
rect 6285 19465 6319 19499
rect 10241 19465 10275 19499
rect 14381 19465 14415 19499
rect 16497 19465 16531 19499
rect 16865 19465 16899 19499
rect 17233 19465 17267 19499
rect 17785 19465 17819 19499
rect 25973 19465 26007 19499
rect 25605 19397 25639 19431
rect 1685 19329 1719 19363
rect 2421 19329 2455 19363
rect 4261 19329 4295 19363
rect 5733 19329 5767 19363
rect 7481 19329 7515 19363
rect 9689 19329 9723 19363
rect 9781 19329 9815 19363
rect 11437 19329 11471 19363
rect 13645 19329 13679 19363
rect 14565 19329 14599 19363
rect 18061 19329 18095 19363
rect 2329 19261 2363 19295
rect 4077 19261 4111 19295
rect 5549 19261 5583 19295
rect 6653 19261 6687 19295
rect 7849 19261 7883 19295
rect 9137 19261 9171 19295
rect 10701 19261 10735 19295
rect 11805 19261 11839 19295
rect 12265 19261 12299 19295
rect 12909 19261 12943 19295
rect 13461 19261 13495 19295
rect 14832 19261 14866 19295
rect 20361 19261 20395 19295
rect 20913 19261 20947 19295
rect 23673 19261 23707 19295
rect 23940 19261 23974 19295
rect 2237 19193 2271 19227
rect 3525 19193 3559 19227
rect 3985 19193 4019 19227
rect 5641 19193 5675 19227
rect 8677 19193 8711 19227
rect 11253 19193 11287 19227
rect 14105 19193 14139 19227
rect 18328 19193 18362 19227
rect 20085 19193 20119 19227
rect 21180 19193 21214 19227
rect 1869 19125 1903 19159
rect 3617 19125 3651 19159
rect 4629 19125 4663 19159
rect 5089 19125 5123 19159
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 7297 19125 7331 19159
rect 8401 19125 8435 19159
rect 9229 19125 9263 19159
rect 9597 19125 9631 19159
rect 10793 19125 10827 19159
rect 11161 19125 11195 19159
rect 13001 19125 13035 19159
rect 13369 19125 13403 19159
rect 15945 19125 15979 19159
rect 19441 19125 19475 19159
rect 20821 19125 20855 19159
rect 22293 19125 22327 19159
rect 22937 19125 22971 19159
rect 23397 19125 23431 19159
rect 25053 19125 25087 19159
rect 1869 18921 1903 18955
rect 2881 18921 2915 18955
rect 2973 18921 3007 18955
rect 5181 18921 5215 18955
rect 5825 18921 5859 18955
rect 7389 18921 7423 18955
rect 7849 18921 7883 18955
rect 9873 18921 9907 18955
rect 13369 18921 13403 18955
rect 14749 18921 14783 18955
rect 15025 18921 15059 18955
rect 17509 18921 17543 18955
rect 17877 18921 17911 18955
rect 18613 18921 18647 18955
rect 19073 18921 19107 18955
rect 22109 18921 22143 18955
rect 24777 18921 24811 18955
rect 25237 18921 25271 18955
rect 3709 18853 3743 18887
rect 4445 18853 4479 18887
rect 7297 18853 7331 18887
rect 8769 18853 8803 18887
rect 10885 18853 10919 18887
rect 14197 18853 14231 18887
rect 23581 18853 23615 18887
rect 25789 18853 25823 18887
rect 1777 18785 1811 18819
rect 2513 18785 2547 18819
rect 6193 18785 6227 18819
rect 6285 18785 6319 18819
rect 7757 18785 7791 18819
rect 10241 18785 10275 18819
rect 10333 18785 10367 18819
rect 11693 18785 11727 18819
rect 16313 18785 16347 18819
rect 17417 18785 17451 18819
rect 19441 18785 19475 18819
rect 21465 18785 21499 18819
rect 22017 18785 22051 18819
rect 23121 18785 23155 18819
rect 25145 18785 25179 18819
rect 2053 18717 2087 18751
rect 4537 18717 4571 18751
rect 4721 18717 4755 18751
rect 6469 18717 6503 18751
rect 7941 18717 7975 18751
rect 10425 18717 10459 18751
rect 11253 18717 11287 18751
rect 11437 18717 11471 18751
rect 16405 18717 16439 18751
rect 16497 18717 16531 18751
rect 17049 18717 17083 18751
rect 17969 18717 18003 18751
rect 18153 18717 18187 18751
rect 19533 18717 19567 18751
rect 19625 18717 19659 18751
rect 21189 18717 21223 18751
rect 22293 18717 22327 18751
rect 23673 18717 23707 18751
rect 23857 18717 23891 18751
rect 25421 18717 25455 18751
rect 4077 18649 4111 18683
rect 5733 18649 5767 18683
rect 9505 18649 9539 18683
rect 15945 18649 15979 18683
rect 20729 18649 20763 18683
rect 21649 18649 21683 18683
rect 23213 18649 23247 18683
rect 24685 18649 24719 18683
rect 1409 18581 1443 18615
rect 6929 18581 6963 18615
rect 8493 18581 8527 18615
rect 12817 18581 12851 18615
rect 13829 18581 13863 18615
rect 15485 18581 15519 18615
rect 18889 18581 18923 18615
rect 20177 18581 20211 18615
rect 22661 18581 22695 18615
rect 24225 18581 24259 18615
rect 4537 18377 4571 18411
rect 7849 18377 7883 18411
rect 12449 18377 12483 18411
rect 14105 18377 14139 18411
rect 17417 18377 17451 18411
rect 18061 18377 18095 18411
rect 21741 18377 21775 18411
rect 23489 18377 23523 18411
rect 24869 18377 24903 18411
rect 25421 18377 25455 18411
rect 25789 18377 25823 18411
rect 26249 18377 26283 18411
rect 5549 18309 5583 18343
rect 12265 18309 12299 18343
rect 19993 18309 20027 18343
rect 21373 18309 21407 18343
rect 1961 18241 1995 18275
rect 2145 18241 2179 18275
rect 2605 18241 2639 18275
rect 5089 18241 5123 18275
rect 6653 18241 6687 18275
rect 8493 18241 8527 18275
rect 13093 18241 13127 18275
rect 13461 18241 13495 18275
rect 14289 18241 14323 18275
rect 16957 18241 16991 18275
rect 18613 18241 18647 18275
rect 20545 18241 20579 18275
rect 20637 18241 20671 18275
rect 22385 18241 22419 18275
rect 22569 18241 22603 18275
rect 24133 18241 24167 18275
rect 24225 18241 24259 18275
rect 3157 18173 3191 18207
rect 3413 18173 3447 18207
rect 5641 18173 5675 18207
rect 8309 18173 8343 18207
rect 8861 18173 8895 18207
rect 9413 18173 9447 18207
rect 9669 18173 9703 18207
rect 12817 18173 12851 18207
rect 14556 18173 14590 18207
rect 18429 18173 18463 18207
rect 22293 18173 22327 18207
rect 25237 18173 25271 18207
rect 11805 18105 11839 18139
rect 16589 18105 16623 18139
rect 19073 18105 19107 18139
rect 23029 18105 23063 18139
rect 24041 18105 24075 18139
rect 1501 18037 1535 18071
rect 1869 18037 1903 18071
rect 2973 18037 3007 18071
rect 5825 18037 5859 18071
rect 6285 18037 6319 18071
rect 6837 18037 6871 18071
rect 7481 18037 7515 18071
rect 8217 18037 8251 18071
rect 9229 18037 9263 18071
rect 10793 18037 10827 18071
rect 11529 18037 11563 18071
rect 12909 18037 12943 18071
rect 15669 18037 15703 18071
rect 16313 18037 16347 18071
rect 17785 18037 17819 18071
rect 18521 18037 18555 18071
rect 19533 18037 19567 18071
rect 20085 18037 20119 18071
rect 20453 18037 20487 18071
rect 21925 18037 21959 18071
rect 23673 18037 23707 18071
rect 3433 17833 3467 17867
rect 3893 17833 3927 17867
rect 4629 17833 4663 17867
rect 6745 17833 6779 17867
rect 7113 17833 7147 17867
rect 8309 17833 8343 17867
rect 9137 17833 9171 17867
rect 10793 17833 10827 17867
rect 12817 17833 12851 17867
rect 13829 17833 13863 17867
rect 14657 17833 14691 17867
rect 16773 17833 16807 17867
rect 18337 17833 18371 17867
rect 18889 17833 18923 17867
rect 19349 17833 19383 17867
rect 19901 17833 19935 17867
rect 22293 17833 22327 17867
rect 22845 17833 22879 17867
rect 23305 17833 23339 17867
rect 7757 17765 7791 17799
rect 11682 17765 11716 17799
rect 13369 17765 13403 17799
rect 16497 17765 16531 17799
rect 17202 17765 17236 17799
rect 20729 17765 20763 17799
rect 21180 17765 21214 17799
rect 1768 17697 1802 17731
rect 5080 17697 5114 17731
rect 7665 17697 7699 17731
rect 10057 17697 10091 17731
rect 11437 17697 11471 17731
rect 15761 17697 15795 17731
rect 15853 17697 15887 17731
rect 19717 17697 19751 17731
rect 23765 17697 23799 17731
rect 24961 17697 24995 17731
rect 1501 17629 1535 17663
rect 4813 17629 4847 17663
rect 7849 17629 7883 17663
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 14197 17629 14231 17663
rect 15117 17629 15151 17663
rect 16037 17629 16071 17663
rect 16957 17629 16991 17663
rect 20913 17629 20947 17663
rect 23857 17629 23891 17663
rect 24041 17629 24075 17663
rect 2881 17493 2915 17527
rect 4353 17493 4387 17527
rect 6193 17493 6227 17527
rect 7297 17493 7331 17527
rect 8677 17493 8711 17527
rect 9413 17493 9447 17527
rect 9689 17493 9723 17527
rect 11253 17493 11287 17527
rect 15393 17493 15427 17527
rect 20361 17493 20395 17527
rect 23397 17493 23431 17527
rect 24409 17493 24443 17527
rect 24869 17493 24903 17527
rect 25145 17493 25179 17527
rect 25605 17493 25639 17527
rect 1869 17289 1903 17323
rect 3433 17289 3467 17323
rect 4721 17289 4755 17323
rect 6653 17289 6687 17323
rect 7021 17289 7055 17323
rect 7389 17289 7423 17323
rect 11805 17289 11839 17323
rect 12173 17289 12207 17323
rect 12633 17289 12667 17323
rect 13553 17289 13587 17323
rect 16405 17289 16439 17323
rect 17417 17289 17451 17323
rect 18429 17289 18463 17323
rect 19993 17289 20027 17323
rect 22477 17289 22511 17323
rect 4353 17221 4387 17255
rect 20545 17221 20579 17255
rect 20913 17221 20947 17255
rect 2053 17153 2087 17187
rect 5365 17153 5399 17187
rect 5457 17153 5491 17187
rect 11437 17153 11471 17187
rect 13737 17153 13771 17187
rect 16865 17153 16899 17187
rect 17049 17153 17083 17187
rect 17785 17153 17819 17187
rect 18613 17153 18647 17187
rect 21097 17153 21131 17187
rect 2320 17085 2354 17119
rect 5273 17085 5307 17119
rect 6837 17085 6871 17119
rect 8033 17085 8067 17119
rect 10609 17085 10643 17119
rect 11161 17085 11195 17119
rect 12449 17085 12483 17119
rect 12909 17085 12943 17119
rect 14004 17085 14038 17119
rect 16773 17085 16807 17119
rect 18869 17085 18903 17119
rect 21364 17085 21398 17119
rect 23305 17085 23339 17119
rect 23673 17085 23707 17119
rect 4077 17017 4111 17051
rect 7757 17017 7791 17051
rect 8300 17017 8334 17051
rect 11253 17017 11287 17051
rect 15669 17017 15703 17051
rect 23121 17017 23155 17051
rect 23940 17017 23974 17051
rect 4905 16949 4939 16983
rect 5917 16949 5951 16983
rect 9413 16949 9447 16983
rect 9965 16949 9999 16983
rect 10793 16949 10827 16983
rect 15117 16949 15151 16983
rect 16129 16949 16163 16983
rect 23305 16949 23339 16983
rect 23397 16949 23431 16983
rect 25053 16949 25087 16983
rect 25605 16949 25639 16983
rect 1409 16745 1443 16779
rect 1961 16745 1995 16779
rect 3433 16745 3467 16779
rect 4261 16745 4295 16779
rect 4905 16745 4939 16779
rect 6837 16745 6871 16779
rect 7481 16745 7515 16779
rect 7941 16745 7975 16779
rect 8309 16745 8343 16779
rect 9137 16745 9171 16779
rect 10977 16745 11011 16779
rect 15117 16745 15151 16779
rect 17693 16745 17727 16779
rect 18705 16745 18739 16779
rect 18797 16745 18831 16779
rect 19165 16745 19199 16779
rect 19809 16745 19843 16779
rect 20913 16745 20947 16779
rect 21281 16745 21315 16779
rect 22569 16745 22603 16779
rect 22937 16745 22971 16779
rect 24409 16745 24443 16779
rect 5365 16677 5399 16711
rect 5702 16677 5736 16711
rect 7849 16677 7883 16711
rect 10241 16677 10275 16711
rect 21373 16677 21407 16711
rect 23296 16677 23330 16711
rect 2789 16609 2823 16643
rect 3893 16609 3927 16643
rect 4077 16609 4111 16643
rect 9413 16609 9447 16643
rect 11253 16609 11287 16643
rect 11704 16609 11738 16643
rect 13921 16609 13955 16643
rect 15301 16609 15335 16643
rect 16313 16609 16347 16643
rect 16580 16609 16614 16643
rect 19257 16609 19291 16643
rect 20361 16609 20395 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 5457 16541 5491 16575
rect 8401 16541 8435 16575
rect 8585 16541 8619 16575
rect 10333 16541 10367 16575
rect 10517 16541 10551 16575
rect 11437 16541 11471 16575
rect 19441 16541 19475 16575
rect 21465 16541 21499 16575
rect 23029 16541 23063 16575
rect 9873 16473 9907 16507
rect 20729 16473 20763 16507
rect 21925 16473 21959 16507
rect 2237 16405 2271 16439
rect 2421 16405 2455 16439
rect 12817 16405 12851 16439
rect 13829 16405 13863 16439
rect 14381 16405 14415 16439
rect 15853 16405 15887 16439
rect 16221 16405 16255 16439
rect 18337 16405 18371 16439
rect 2421 16201 2455 16235
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 8769 16201 8803 16235
rect 9781 16201 9815 16235
rect 12449 16201 12483 16235
rect 13921 16201 13955 16235
rect 14013 16201 14047 16235
rect 15853 16201 15887 16235
rect 16405 16201 16439 16235
rect 19165 16201 19199 16235
rect 19901 16201 19935 16235
rect 21281 16201 21315 16235
rect 23029 16201 23063 16235
rect 23397 16201 23431 16235
rect 9321 16133 9355 16167
rect 19809 16133 19843 16167
rect 22753 16133 22787 16167
rect 2605 16065 2639 16099
rect 5089 16065 5123 16099
rect 5733 16065 5767 16099
rect 6837 16065 6871 16099
rect 13001 16065 13035 16099
rect 13461 16065 13495 16099
rect 14565 16065 14599 16099
rect 17049 16065 17083 16099
rect 18613 16065 18647 16099
rect 20361 16065 20395 16099
rect 20545 16065 20579 16099
rect 22017 16065 22051 16099
rect 23673 16065 23707 16099
rect 1409 15997 1443 16031
rect 9873 15997 9907 16031
rect 11805 15997 11839 16031
rect 17785 15997 17819 16031
rect 18521 15997 18555 16031
rect 21925 15997 21959 16031
rect 2053 15929 2087 15963
rect 2872 15929 2906 15963
rect 4721 15929 4755 15963
rect 5641 15929 5675 15963
rect 7104 15929 7138 15963
rect 10140 15929 10174 15963
rect 12265 15929 12299 15963
rect 12817 15929 12851 15963
rect 16773 15929 16807 15963
rect 18429 15929 18463 15963
rect 20269 15929 20303 15963
rect 21833 15929 21867 15963
rect 23918 15929 23952 15963
rect 1593 15861 1627 15895
rect 3985 15861 4019 15895
rect 5181 15861 5215 15895
rect 5549 15861 5583 15895
rect 8217 15861 8251 15895
rect 11253 15861 11287 15895
rect 12909 15861 12943 15895
rect 14381 15861 14415 15895
rect 14473 15861 14507 15895
rect 15485 15861 15519 15895
rect 16313 15861 16347 15895
rect 16865 15861 16899 15895
rect 17417 15861 17451 15895
rect 18061 15861 18095 15895
rect 21005 15861 21039 15895
rect 21465 15861 21499 15895
rect 25053 15861 25087 15895
rect 2053 15657 2087 15691
rect 3801 15657 3835 15691
rect 5549 15657 5583 15691
rect 8033 15657 8067 15691
rect 8769 15657 8803 15691
rect 9505 15657 9539 15691
rect 9873 15657 9907 15691
rect 10977 15657 11011 15691
rect 11345 15657 11379 15691
rect 12817 15657 12851 15691
rect 14105 15657 14139 15691
rect 15669 15657 15703 15691
rect 16405 15657 16439 15691
rect 17877 15657 17911 15691
rect 19165 15657 19199 15691
rect 19257 15657 19291 15691
rect 20729 15657 20763 15691
rect 21189 15657 21223 15691
rect 22937 15657 22971 15691
rect 23489 15657 23523 15691
rect 2421 15589 2455 15623
rect 3157 15589 3191 15623
rect 4813 15589 4847 15623
rect 6184 15589 6218 15623
rect 10241 15589 10275 15623
rect 3525 15521 3559 15555
rect 4721 15521 4755 15555
rect 5917 15521 5951 15555
rect 8585 15521 8619 15555
rect 9137 15521 9171 15555
rect 11437 15521 11471 15555
rect 11704 15521 11738 15555
rect 13921 15521 13955 15555
rect 15485 15521 15519 15555
rect 16497 15521 16531 15555
rect 16764 15521 16798 15555
rect 18797 15521 18831 15555
rect 19625 15521 19659 15555
rect 21813 15521 21847 15555
rect 24409 15521 24443 15555
rect 24501 15521 24535 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 4997 15453 5031 15487
rect 8309 15453 8343 15487
rect 10333 15453 10367 15487
rect 10425 15453 10459 15487
rect 19717 15453 19751 15487
rect 19809 15453 19843 15487
rect 21557 15453 21591 15487
rect 24685 15453 24719 15487
rect 4353 15385 4387 15419
rect 14381 15385 14415 15419
rect 23949 15385 23983 15419
rect 1593 15317 1627 15351
rect 7297 15317 7331 15351
rect 13369 15317 13403 15351
rect 20269 15317 20303 15351
rect 24041 15317 24075 15351
rect 1593 15113 1627 15147
rect 2145 15113 2179 15147
rect 4077 15113 4111 15147
rect 4445 15113 4479 15147
rect 6561 15113 6595 15147
rect 9965 15113 9999 15147
rect 10793 15113 10827 15147
rect 11805 15113 11839 15147
rect 14565 15113 14599 15147
rect 16589 15113 16623 15147
rect 16957 15113 16991 15147
rect 17509 15113 17543 15147
rect 21005 15113 21039 15147
rect 21925 15113 21959 15147
rect 23489 15113 23523 15147
rect 23857 15113 23891 15147
rect 25605 15113 25639 15147
rect 2697 15045 2731 15079
rect 4721 15045 4755 15079
rect 12725 15045 12759 15079
rect 17785 15045 17819 15079
rect 22661 15045 22695 15079
rect 24869 15045 24903 15079
rect 25237 15045 25271 15079
rect 3341 14977 3375 15011
rect 5825 14977 5859 15011
rect 6285 14977 6319 15011
rect 7573 14977 7607 15011
rect 7757 14977 7791 15011
rect 11437 14977 11471 15011
rect 13277 14977 13311 15011
rect 14657 14977 14691 15011
rect 18613 14977 18647 15011
rect 24317 14977 24351 15011
rect 24409 14977 24443 15011
rect 1409 14909 1443 14943
rect 3157 14909 3191 14943
rect 5549 14909 5583 14943
rect 12265 14909 12299 14943
rect 13185 14909 13219 14943
rect 18429 14909 18463 14943
rect 19625 14909 19659 14943
rect 22477 14909 22511 14943
rect 23029 14909 23063 14943
rect 25421 14909 25455 14943
rect 25973 14909 26007 14943
rect 7021 14841 7055 14875
rect 8002 14841 8036 14875
rect 10609 14841 10643 14875
rect 11161 14841 11195 14875
rect 14902 14841 14936 14875
rect 19892 14841 19926 14875
rect 2605 14773 2639 14807
rect 3065 14773 3099 14807
rect 5181 14773 5215 14807
rect 5641 14773 5675 14807
rect 9137 14773 9171 14807
rect 10241 14773 10275 14807
rect 11253 14773 11287 14807
rect 13093 14773 13127 14807
rect 13921 14773 13955 14807
rect 16037 14773 16071 14807
rect 18061 14773 18095 14807
rect 18521 14773 18555 14807
rect 19349 14773 19383 14807
rect 21557 14773 21591 14807
rect 24225 14773 24259 14807
rect 2145 14569 2179 14603
rect 3525 14569 3559 14603
rect 3893 14569 3927 14603
rect 4261 14569 4295 14603
rect 6285 14569 6319 14603
rect 9505 14569 9539 14603
rect 11621 14569 11655 14603
rect 11989 14569 12023 14603
rect 13185 14569 13219 14603
rect 13553 14569 13587 14603
rect 13645 14569 13679 14603
rect 17601 14569 17635 14603
rect 18245 14569 18279 14603
rect 18705 14569 18739 14603
rect 20545 14569 20579 14603
rect 22293 14569 22327 14603
rect 23857 14569 23891 14603
rect 24869 14569 24903 14603
rect 25605 14569 25639 14603
rect 2881 14501 2915 14535
rect 5917 14501 5951 14535
rect 6644 14501 6678 14535
rect 19073 14501 19107 14535
rect 20177 14501 20211 14535
rect 24317 14501 24351 14535
rect 1409 14433 1443 14467
rect 2789 14433 2823 14467
rect 5181 14433 5215 14467
rect 5273 14433 5307 14467
rect 6377 14433 6411 14467
rect 9956 14433 9990 14467
rect 12173 14433 12207 14467
rect 14013 14433 14047 14467
rect 16221 14433 16255 14467
rect 16477 14433 16511 14467
rect 21180 14433 21214 14467
rect 23397 14433 23431 14467
rect 24225 14433 24259 14467
rect 25421 14433 25455 14467
rect 2973 14365 3007 14399
rect 5365 14365 5399 14399
rect 9689 14365 9723 14399
rect 14105 14365 14139 14399
rect 14197 14365 14231 14399
rect 19165 14365 19199 14399
rect 19257 14365 19291 14399
rect 19809 14365 19843 14399
rect 20913 14365 20947 14399
rect 24409 14365 24443 14399
rect 4813 14297 4847 14331
rect 7757 14297 7791 14331
rect 8309 14297 8343 14331
rect 12357 14297 12391 14331
rect 1593 14229 1627 14263
rect 2421 14229 2455 14263
rect 4721 14229 4755 14263
rect 8769 14229 8803 14263
rect 9137 14229 9171 14263
rect 11069 14229 11103 14263
rect 12725 14229 12759 14263
rect 14657 14229 14691 14263
rect 15485 14229 15519 14263
rect 16037 14229 16071 14263
rect 18613 14229 18647 14263
rect 23029 14229 23063 14263
rect 23765 14229 23799 14263
rect 1593 14025 1627 14059
rect 1961 14025 1995 14059
rect 2697 14025 2731 14059
rect 4997 14025 5031 14059
rect 6377 14025 6411 14059
rect 7481 14025 7515 14059
rect 9045 14025 9079 14059
rect 9413 14025 9447 14059
rect 11529 14025 11563 14059
rect 12909 14025 12943 14059
rect 15853 14025 15887 14059
rect 17877 14025 17911 14059
rect 21281 14025 21315 14059
rect 21465 14025 21499 14059
rect 25421 14025 25455 14059
rect 2421 13957 2455 13991
rect 5181 13957 5215 13991
rect 8033 13957 8067 13991
rect 13369 13957 13403 13991
rect 14841 13957 14875 13991
rect 16957 13957 16991 13991
rect 18429 13957 18463 13991
rect 19993 13957 20027 13991
rect 23121 13957 23155 13991
rect 3525 13889 3559 13923
rect 4169 13889 4203 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 8677 13889 8711 13923
rect 16497 13889 16531 13923
rect 22017 13889 22051 13923
rect 24225 13889 24259 13923
rect 26157 13889 26191 13923
rect 1409 13821 1443 13855
rect 2513 13821 2547 13855
rect 3065 13821 3099 13855
rect 4721 13821 4755 13855
rect 7849 13821 7883 13855
rect 9597 13821 9631 13855
rect 9853 13821 9887 13855
rect 13461 13821 13495 13855
rect 15393 13821 15427 13855
rect 16405 13821 16439 13855
rect 18613 13821 18647 13855
rect 20637 13821 20671 13855
rect 21925 13821 21959 13855
rect 23489 13821 23523 13855
rect 24133 13821 24167 13855
rect 25053 13821 25087 13855
rect 25237 13821 25271 13855
rect 25789 13821 25823 13855
rect 4077 13753 4111 13787
rect 5549 13753 5583 13787
rect 6837 13753 6871 13787
rect 8401 13753 8435 13787
rect 8493 13753 8527 13787
rect 13706 13753 13740 13787
rect 18858 13753 18892 13787
rect 21833 13753 21867 13787
rect 24041 13753 24075 13787
rect 3617 13685 3651 13719
rect 3985 13685 4019 13719
rect 10977 13685 11011 13719
rect 12265 13685 12299 13719
rect 12449 13685 12483 13719
rect 15945 13685 15979 13719
rect 16313 13685 16347 13719
rect 21005 13685 21039 13719
rect 22477 13685 22511 13719
rect 23673 13685 23707 13719
rect 24685 13685 24719 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 2329 13481 2363 13515
rect 2697 13481 2731 13515
rect 3617 13481 3651 13515
rect 4261 13481 4295 13515
rect 4445 13481 4479 13515
rect 4905 13481 4939 13515
rect 5457 13481 5491 13515
rect 6009 13481 6043 13515
rect 6469 13481 6503 13515
rect 7021 13481 7055 13515
rect 7941 13481 7975 13515
rect 8401 13481 8435 13515
rect 9413 13481 9447 13515
rect 13829 13481 13863 13515
rect 14381 13481 14415 13515
rect 18705 13481 18739 13515
rect 19165 13481 19199 13515
rect 21189 13481 21223 13515
rect 22661 13481 22695 13515
rect 23673 13481 23707 13515
rect 24133 13481 24167 13515
rect 5825 13413 5859 13447
rect 7389 13413 7423 13447
rect 17018 13413 17052 13447
rect 19717 13413 19751 13447
rect 24225 13413 24259 13447
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 4813 13345 4847 13379
rect 6377 13345 6411 13379
rect 8493 13345 8527 13379
rect 10232 13345 10266 13379
rect 12716 13345 12750 13379
rect 15761 13345 15795 13379
rect 16773 13345 16807 13379
rect 19625 13345 19659 13379
rect 21548 13345 21582 13379
rect 25329 13345 25363 13379
rect 5089 13277 5123 13311
rect 6653 13277 6687 13311
rect 8677 13277 8711 13311
rect 9965 13277 9999 13311
rect 12449 13277 12483 13311
rect 19901 13277 19935 13311
rect 21281 13277 21315 13311
rect 24317 13277 24351 13311
rect 8033 13209 8067 13243
rect 18153 13209 18187 13243
rect 3157 13141 3191 13175
rect 11345 13141 11379 13175
rect 12173 13141 12207 13175
rect 15485 13141 15519 13175
rect 16313 13141 16347 13175
rect 19257 13141 19291 13175
rect 20269 13141 20303 13175
rect 20729 13141 20763 13175
rect 23305 13141 23339 13175
rect 23765 13141 23799 13175
rect 25513 13141 25547 13175
rect 1593 12937 1627 12971
rect 3525 12937 3559 12971
rect 5181 12937 5215 12971
rect 6285 12937 6319 12971
rect 6837 12937 6871 12971
rect 8125 12937 8159 12971
rect 8493 12937 8527 12971
rect 8769 12937 8803 12971
rect 9321 12937 9355 12971
rect 10333 12937 10367 12971
rect 10793 12937 10827 12971
rect 13001 12937 13035 12971
rect 13553 12937 13587 12971
rect 15025 12937 15059 12971
rect 16405 12937 16439 12971
rect 16773 12937 16807 12971
rect 17141 12937 17175 12971
rect 18061 12937 18095 12971
rect 19349 12937 19383 12971
rect 20637 12937 20671 12971
rect 21925 12937 21959 12971
rect 23673 12937 23707 12971
rect 24685 12937 24719 12971
rect 25053 12937 25087 12971
rect 26157 12937 26191 12971
rect 2697 12869 2731 12903
rect 3157 12869 3191 12903
rect 4997 12869 5031 12903
rect 15117 12869 15151 12903
rect 23029 12869 23063 12903
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 6561 12801 6595 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 9873 12801 9907 12835
rect 12541 12801 12575 12835
rect 14105 12801 14139 12835
rect 14657 12801 14691 12835
rect 15669 12801 15703 12835
rect 17509 12801 17543 12835
rect 18613 12801 18647 12835
rect 20269 12801 20303 12835
rect 21833 12801 21867 12835
rect 22385 12801 22419 12835
rect 22569 12801 22603 12835
rect 24133 12801 24167 12835
rect 24317 12801 24351 12835
rect 1409 12733 1443 12767
rect 2513 12733 2547 12767
rect 3617 12733 3651 12767
rect 4353 12733 4387 12767
rect 5549 12733 5583 12767
rect 7205 12733 7239 12767
rect 9689 12733 9723 12767
rect 13461 12733 13495 12767
rect 14013 12733 14047 12767
rect 15485 12733 15519 12767
rect 15577 12733 15611 12767
rect 16957 12733 16991 12767
rect 20085 12733 20119 12767
rect 25237 12733 25271 12767
rect 25789 12733 25823 12767
rect 2053 12665 2087 12699
rect 4721 12665 4755 12699
rect 9137 12665 9171 12699
rect 10977 12665 11011 12699
rect 18429 12665 18463 12699
rect 19993 12665 20027 12699
rect 22293 12665 22327 12699
rect 23397 12665 23431 12699
rect 24041 12665 24075 12699
rect 2329 12597 2363 12631
rect 3801 12597 3835 12631
rect 9781 12597 9815 12631
rect 12173 12597 12207 12631
rect 13921 12597 13955 12631
rect 17785 12597 17819 12631
rect 18521 12597 18555 12631
rect 19625 12597 19659 12631
rect 21373 12597 21407 12631
rect 25421 12597 25455 12631
rect 1777 12393 1811 12427
rect 2145 12393 2179 12427
rect 2881 12393 2915 12427
rect 3249 12393 3283 12427
rect 3893 12393 3927 12427
rect 4813 12393 4847 12427
rect 5641 12393 5675 12427
rect 7205 12393 7239 12427
rect 8953 12393 8987 12427
rect 9413 12393 9447 12427
rect 12909 12393 12943 12427
rect 18061 12393 18095 12427
rect 19717 12393 19751 12427
rect 21465 12393 21499 12427
rect 23765 12393 23799 12427
rect 24317 12393 24351 12427
rect 25329 12393 25363 12427
rect 2513 12325 2547 12359
rect 4537 12325 4571 12359
rect 10149 12325 10183 12359
rect 22652 12325 22686 12359
rect 1593 12257 1627 12291
rect 2697 12257 2731 12291
rect 5273 12257 5307 12291
rect 6009 12257 6043 12291
rect 6101 12257 6135 12291
rect 7573 12257 7607 12291
rect 10057 12257 10091 12291
rect 11529 12257 11563 12291
rect 11796 12257 11830 12291
rect 14013 12257 14047 12291
rect 15301 12257 15335 12291
rect 15568 12257 15602 12291
rect 18604 12257 18638 12291
rect 20729 12257 20763 12291
rect 21281 12257 21315 12291
rect 25237 12257 25271 12291
rect 6285 12189 6319 12223
rect 7665 12189 7699 12223
rect 7757 12189 7791 12223
rect 10241 12189 10275 12223
rect 14197 12189 14231 12223
rect 18337 12189 18371 12223
rect 21189 12189 21223 12223
rect 21925 12189 21959 12223
rect 22385 12189 22419 12223
rect 25421 12189 25455 12223
rect 8677 12121 8711 12155
rect 9689 12121 9723 12155
rect 10885 12121 10919 12155
rect 24869 12121 24903 12155
rect 6929 12053 6963 12087
rect 8309 12053 8343 12087
rect 11253 12053 11287 12087
rect 13645 12053 13679 12087
rect 15117 12053 15151 12087
rect 16681 12053 16715 12087
rect 17325 12053 17359 12087
rect 20361 12053 20395 12087
rect 1593 11849 1627 11883
rect 2789 11849 2823 11883
rect 4997 11849 5031 11883
rect 6101 11849 6135 11883
rect 6653 11849 6687 11883
rect 7205 11849 7239 11883
rect 9229 11849 9263 11883
rect 10241 11849 10275 11883
rect 10793 11849 10827 11883
rect 11805 11849 11839 11883
rect 13093 11849 13127 11883
rect 14657 11849 14691 11883
rect 15761 11849 15795 11883
rect 22661 11849 22695 11883
rect 23489 11849 23523 11883
rect 23673 11849 23707 11883
rect 24961 11849 24995 11883
rect 25421 11849 25455 11883
rect 1869 11781 1903 11815
rect 2237 11781 2271 11815
rect 4629 11781 4663 11815
rect 5733 11781 5767 11815
rect 7665 11781 7699 11815
rect 18061 11781 18095 11815
rect 5273 11713 5307 11747
rect 7573 11713 7607 11747
rect 8125 11713 8159 11747
rect 8309 11713 8343 11747
rect 8769 11713 8803 11747
rect 9781 11713 9815 11747
rect 11253 11713 11287 11747
rect 11437 11713 11471 11747
rect 13277 11713 13311 11747
rect 16221 11713 16255 11747
rect 16405 11713 16439 11747
rect 16865 11713 16899 11747
rect 17509 11713 17543 11747
rect 18613 11713 18647 11747
rect 22017 11713 22051 11747
rect 24133 11713 24167 11747
rect 24317 11713 24351 11747
rect 26157 11713 26191 11747
rect 1409 11645 1443 11679
rect 8033 11645 8067 11679
rect 9137 11645 9171 11679
rect 9597 11645 9631 11679
rect 10701 11645 10735 11679
rect 11161 11645 11195 11679
rect 15301 11645 15335 11679
rect 16129 11645 16163 11679
rect 18429 11645 18463 11679
rect 19901 11645 19935 11679
rect 22477 11645 22511 11679
rect 23029 11645 23063 11679
rect 24041 11645 24075 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 9689 11577 9723 11611
rect 12173 11577 12207 11611
rect 12817 11577 12851 11611
rect 13544 11577 13578 11611
rect 19073 11577 19107 11611
rect 19717 11577 19751 11611
rect 20168 11577 20202 11611
rect 17785 11509 17819 11543
rect 18521 11509 18555 11543
rect 21281 11509 21315 11543
rect 22293 11509 22327 11543
rect 6101 11305 6135 11339
rect 7297 11305 7331 11339
rect 7757 11305 7791 11339
rect 8401 11305 8435 11339
rect 9321 11305 9355 11339
rect 10149 11305 10183 11339
rect 10977 11305 11011 11339
rect 14197 11305 14231 11339
rect 16681 11305 16715 11339
rect 17785 11305 17819 11339
rect 18061 11305 18095 11339
rect 21557 11305 21591 11339
rect 23489 11305 23523 11339
rect 24041 11305 24075 11339
rect 24409 11305 24443 11339
rect 24961 11305 24995 11339
rect 9689 11237 9723 11271
rect 15117 11237 15151 11271
rect 15568 11237 15602 11271
rect 18604 11237 18638 11271
rect 25605 11237 25639 11271
rect 8493 11169 8527 11203
rect 10793 11169 10827 11203
rect 11345 11169 11379 11203
rect 12909 11169 12943 11203
rect 13553 11169 13587 11203
rect 15301 11169 15335 11203
rect 22365 11169 22399 11203
rect 8585 11101 8619 11135
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 12081 11101 12115 11135
rect 13001 11101 13035 11135
rect 13185 11101 13219 11135
rect 18337 11101 18371 11135
rect 21097 11101 21131 11135
rect 22109 11101 22143 11135
rect 25053 11101 25087 11135
rect 25145 11101 25179 11135
rect 5733 11033 5767 11067
rect 8033 11033 8067 11067
rect 12449 11033 12483 11067
rect 17417 11033 17451 11067
rect 19717 11033 19751 11067
rect 20269 11033 20303 11067
rect 22017 11033 22051 11067
rect 24593 11033 24627 11067
rect 12541 10965 12575 10999
rect 7757 10761 7791 10795
rect 8493 10761 8527 10795
rect 9229 10761 9263 10795
rect 10793 10761 10827 10795
rect 13829 10761 13863 10795
rect 15945 10761 15979 10795
rect 16313 10761 16347 10795
rect 17049 10761 17083 10795
rect 18245 10761 18279 10795
rect 19625 10761 19659 10795
rect 20085 10761 20119 10795
rect 23029 10761 23063 10795
rect 23489 10761 23523 10795
rect 23673 10761 23707 10795
rect 25145 10761 25179 10795
rect 25421 10761 25455 10795
rect 25881 10761 25915 10795
rect 12173 10693 12207 10727
rect 14933 10693 14967 10727
rect 17509 10693 17543 10727
rect 8125 10625 8159 10659
rect 9781 10625 9815 10659
rect 11253 10625 11287 10659
rect 11437 10625 11471 10659
rect 12449 10625 12483 10659
rect 15485 10625 15519 10659
rect 18705 10625 18739 10659
rect 18797 10625 18831 10659
rect 24225 10625 24259 10659
rect 9137 10557 9171 10591
rect 9597 10557 9631 10591
rect 16865 10557 16899 10591
rect 18613 10557 18647 10591
rect 19901 10557 19935 10591
rect 21005 10557 21039 10591
rect 21097 10557 21131 10591
rect 24685 10557 24719 10591
rect 25237 10557 25271 10591
rect 10609 10489 10643 10523
rect 11161 10489 11195 10523
rect 12716 10489 12750 10523
rect 15393 10489 15427 10523
rect 17877 10489 17911 10523
rect 21364 10489 21398 10523
rect 24041 10489 24075 10523
rect 9689 10421 9723 10455
rect 10333 10421 10367 10455
rect 11805 10421 11839 10455
rect 14381 10421 14415 10455
rect 14841 10421 14875 10455
rect 15301 10421 15335 10455
rect 16681 10421 16715 10455
rect 19349 10421 19383 10455
rect 20637 10421 20671 10455
rect 22477 10421 22511 10455
rect 24133 10421 24167 10455
rect 9321 10217 9355 10251
rect 10609 10217 10643 10251
rect 11621 10217 11655 10251
rect 15025 10217 15059 10251
rect 15577 10217 15611 10251
rect 18797 10217 18831 10251
rect 19165 10217 19199 10251
rect 19809 10217 19843 10251
rect 20913 10217 20947 10251
rect 24225 10217 24259 10251
rect 10149 10149 10183 10183
rect 16304 10149 16338 10183
rect 19257 10149 19291 10183
rect 21741 10149 21775 10183
rect 22192 10149 22226 10183
rect 8953 10081 8987 10115
rect 10977 10081 11011 10115
rect 12173 10081 12207 10115
rect 12440 10081 12474 10115
rect 16037 10081 16071 10115
rect 21925 10081 21959 10115
rect 24593 10081 24627 10115
rect 10517 10013 10551 10047
rect 11069 10013 11103 10047
rect 11161 10013 11195 10047
rect 11989 10013 12023 10047
rect 19349 10013 19383 10047
rect 18061 9945 18095 9979
rect 24777 9945 24811 9979
rect 13553 9877 13587 9911
rect 17417 9877 17451 9911
rect 18337 9877 18371 9911
rect 20269 9877 20303 9911
rect 23305 9877 23339 9911
rect 23857 9877 23891 9911
rect 25145 9877 25179 9911
rect 11161 9673 11195 9707
rect 12173 9673 12207 9707
rect 15117 9673 15151 9707
rect 22661 9673 22695 9707
rect 24409 9673 24443 9707
rect 10057 9605 10091 9639
rect 16221 9605 16255 9639
rect 17233 9605 17267 9639
rect 20269 9605 20303 9639
rect 24777 9605 24811 9639
rect 10701 9537 10735 9571
rect 13553 9537 13587 9571
rect 13737 9537 13771 9571
rect 16865 9537 16899 9571
rect 22293 9537 22327 9571
rect 10517 9469 10551 9503
rect 11897 9469 11931 9503
rect 18337 9469 18371 9503
rect 21189 9469 21223 9503
rect 22109 9469 22143 9503
rect 24593 9469 24627 9503
rect 25145 9469 25179 9503
rect 13277 9401 13311 9435
rect 14004 9401 14038 9435
rect 16129 9401 16163 9435
rect 16681 9401 16715 9435
rect 18582 9401 18616 9435
rect 21557 9401 21591 9435
rect 22017 9401 22051 9435
rect 9873 9333 9907 9367
rect 10425 9333 10459 9367
rect 11529 9333 11563 9367
rect 12541 9333 12575 9367
rect 15761 9333 15795 9367
rect 16589 9333 16623 9367
rect 17785 9333 17819 9367
rect 19717 9333 19751 9367
rect 21649 9333 21683 9367
rect 10057 9129 10091 9163
rect 10701 9129 10735 9163
rect 11897 9129 11931 9163
rect 13461 9129 13495 9163
rect 13921 9129 13955 9163
rect 14565 9129 14599 9163
rect 15577 9129 15611 9163
rect 16957 9129 16991 9163
rect 19441 9129 19475 9163
rect 19993 9129 20027 9163
rect 20913 9129 20947 9163
rect 22845 9129 22879 9163
rect 24777 9129 24811 9163
rect 13829 9061 13863 9095
rect 16589 9061 16623 9095
rect 22017 9061 22051 9095
rect 12265 8993 12299 9027
rect 13001 8993 13035 9027
rect 15945 8993 15979 9027
rect 17141 8993 17175 9027
rect 17408 8993 17442 9027
rect 19809 8993 19843 9027
rect 21281 8993 21315 9027
rect 22937 8993 22971 9027
rect 24593 8993 24627 9027
rect 12357 8925 12391 8959
rect 12541 8925 12575 8959
rect 14105 8925 14139 8959
rect 15117 8925 15151 8959
rect 16037 8925 16071 8959
rect 16129 8925 16163 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 23121 8925 23155 8959
rect 18521 8857 18555 8891
rect 22477 8857 22511 8891
rect 20729 8789 20763 8823
rect 11621 8585 11655 8619
rect 12909 8585 12943 8619
rect 14013 8585 14047 8619
rect 15669 8585 15703 8619
rect 17509 8585 17543 8619
rect 18889 8585 18923 8619
rect 19349 8585 19383 8619
rect 21281 8585 21315 8619
rect 22845 8585 22879 8619
rect 23213 8585 23247 8619
rect 25237 8585 25271 8619
rect 12817 8517 12851 8551
rect 14473 8517 14507 8551
rect 20913 8517 20947 8551
rect 13369 8449 13403 8483
rect 13553 8449 13587 8483
rect 15025 8449 15059 8483
rect 16313 8449 16347 8483
rect 16957 8449 16991 8483
rect 17877 8449 17911 8483
rect 19809 8449 19843 8483
rect 19901 8449 19935 8483
rect 21741 8449 21775 8483
rect 21833 8449 21867 8483
rect 24041 8449 24075 8483
rect 11253 8381 11287 8415
rect 13277 8381 13311 8415
rect 16865 8381 16899 8415
rect 19257 8381 19291 8415
rect 19717 8381 19751 8415
rect 20545 8381 20579 8415
rect 21649 8381 21683 8415
rect 25053 8381 25087 8415
rect 25513 8381 25547 8415
rect 11897 8313 11931 8347
rect 14381 8313 14415 8347
rect 14841 8313 14875 8347
rect 16773 8313 16807 8347
rect 18061 8313 18095 8347
rect 14933 8245 14967 8279
rect 16405 8245 16439 8279
rect 22477 8245 22511 8279
rect 24593 8245 24627 8279
rect 11897 8041 11931 8075
rect 13277 8041 13311 8075
rect 13645 8041 13679 8075
rect 15117 8041 15151 8075
rect 15669 8041 15703 8075
rect 16037 8041 16071 8075
rect 17877 8041 17911 8075
rect 20085 8041 20119 8075
rect 21557 8041 21591 8075
rect 22109 8041 22143 8075
rect 22845 8041 22879 8075
rect 23857 8041 23891 8075
rect 24869 8041 24903 8075
rect 12357 7973 12391 8007
rect 13001 7973 13035 8007
rect 20729 7973 20763 8007
rect 12265 7905 12299 7939
rect 13461 7905 13495 7939
rect 15485 7905 15519 7939
rect 16497 7905 16531 7939
rect 16764 7905 16798 7939
rect 19349 7905 19383 7939
rect 21373 7905 21407 7939
rect 22661 7905 22695 7939
rect 23673 7905 23707 7939
rect 24685 7905 24719 7939
rect 12449 7837 12483 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 14013 7701 14047 7735
rect 14565 7701 14599 7735
rect 16405 7701 16439 7735
rect 18981 7701 19015 7735
rect 11621 7497 11655 7531
rect 13461 7497 13495 7531
rect 15025 7497 15059 7531
rect 16405 7497 16439 7531
rect 18061 7497 18095 7531
rect 19165 7497 19199 7531
rect 19625 7497 19659 7531
rect 20637 7497 20671 7531
rect 23029 7497 23063 7531
rect 23857 7497 23891 7531
rect 24133 7497 24167 7531
rect 25513 7497 25547 7531
rect 15945 7429 15979 7463
rect 24869 7429 24903 7463
rect 15117 7361 15151 7395
rect 16313 7361 16347 7395
rect 16865 7361 16899 7395
rect 16957 7361 16991 7395
rect 17509 7361 17543 7395
rect 18705 7361 18739 7395
rect 20269 7361 20303 7395
rect 21189 7361 21223 7395
rect 22569 7361 22603 7395
rect 12725 7293 12759 7327
rect 16773 7293 16807 7327
rect 20085 7293 20119 7327
rect 23673 7293 23707 7327
rect 24501 7293 24535 7327
rect 24685 7293 24719 7327
rect 25145 7293 25179 7327
rect 17877 7225 17911 7259
rect 19533 7225 19567 7259
rect 11897 7157 11931 7191
rect 18429 7157 18463 7191
rect 18521 7157 18555 7191
rect 19993 7157 20027 7191
rect 15485 6953 15519 6987
rect 16865 6953 16899 6987
rect 17417 6953 17451 6987
rect 19073 6953 19107 6987
rect 19625 6953 19659 6987
rect 20085 6953 20119 6987
rect 16129 6817 16163 6851
rect 23765 6817 23799 6851
rect 24777 6817 24811 6851
rect 17509 6749 17543 6783
rect 17601 6749 17635 6783
rect 17049 6681 17083 6715
rect 23949 6681 23983 6715
rect 16497 6613 16531 6647
rect 18153 6613 18187 6647
rect 16221 6409 16255 6443
rect 16405 6409 16439 6443
rect 17877 6409 17911 6443
rect 23857 6409 23891 6443
rect 16957 6273 16991 6307
rect 16865 6205 16899 6239
rect 16773 6069 16807 6103
rect 17417 6069 17451 6103
rect 16405 5865 16439 5899
rect 17049 5865 17083 5899
rect 14289 2601 14323 2635
rect 12449 2465 12483 2499
rect 13176 2465 13210 2499
rect 11989 2397 12023 2431
rect 12909 2397 12943 2431
<< metal1 >>
rect 10042 25984 10048 26036
rect 10100 26024 10106 26036
rect 14826 26024 14832 26036
rect 10100 25996 14832 26024
rect 10100 25984 10106 25996
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 8018 25916 8024 25968
rect 8076 25956 8082 25968
rect 18598 25956 18604 25968
rect 8076 25928 18604 25956
rect 8076 25916 8082 25928
rect 18598 25916 18604 25928
rect 18656 25916 18662 25968
rect 13262 25848 13268 25900
rect 13320 25888 13326 25900
rect 21542 25888 21548 25900
rect 13320 25860 21548 25888
rect 13320 25848 13326 25860
rect 21542 25848 21548 25860
rect 21600 25848 21606 25900
rect 9582 25780 9588 25832
rect 9640 25820 9646 25832
rect 18046 25820 18052 25832
rect 9640 25792 18052 25820
rect 9640 25780 9646 25792
rect 18046 25780 18052 25792
rect 18104 25780 18110 25832
rect 10962 25712 10968 25764
rect 11020 25752 11026 25764
rect 16298 25752 16304 25764
rect 11020 25724 16304 25752
rect 11020 25712 11026 25724
rect 16298 25712 16304 25724
rect 16356 25712 16362 25764
rect 1394 25644 1400 25696
rect 1452 25684 1458 25696
rect 11698 25684 11704 25696
rect 1452 25656 11704 25684
rect 1452 25644 1458 25656
rect 11698 25644 11704 25656
rect 11756 25644 11762 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1394 25480 1400 25492
rect 1355 25452 1400 25480
rect 1394 25440 1400 25452
rect 1452 25440 1458 25492
rect 2777 25483 2835 25489
rect 2777 25449 2789 25483
rect 2823 25480 2835 25483
rect 2866 25480 2872 25492
rect 2823 25452 2872 25480
rect 2823 25449 2835 25452
rect 2777 25443 2835 25449
rect 2866 25440 2872 25452
rect 2924 25440 2930 25492
rect 2958 25440 2964 25492
rect 3016 25480 3022 25492
rect 4249 25483 4307 25489
rect 4249 25480 4261 25483
rect 3016 25452 4261 25480
rect 3016 25440 3022 25452
rect 4249 25449 4261 25452
rect 4295 25449 4307 25483
rect 4249 25443 4307 25449
rect 5074 25440 5080 25492
rect 5132 25480 5138 25492
rect 5629 25483 5687 25489
rect 5629 25480 5641 25483
rect 5132 25452 5641 25480
rect 5132 25440 5138 25452
rect 5629 25449 5641 25452
rect 5675 25449 5687 25483
rect 5629 25443 5687 25449
rect 7282 25440 7288 25492
rect 7340 25480 7346 25492
rect 7561 25483 7619 25489
rect 7561 25480 7573 25483
rect 7340 25452 7573 25480
rect 7340 25440 7346 25452
rect 7561 25449 7573 25452
rect 7607 25449 7619 25483
rect 8018 25480 8024 25492
rect 7979 25452 8024 25480
rect 7561 25443 7619 25449
rect 8018 25440 8024 25452
rect 8076 25440 8082 25492
rect 10229 25483 10287 25489
rect 10229 25449 10241 25483
rect 10275 25480 10287 25483
rect 10505 25483 10563 25489
rect 10505 25480 10517 25483
rect 10275 25452 10517 25480
rect 10275 25449 10287 25452
rect 10229 25443 10287 25449
rect 10505 25449 10517 25452
rect 10551 25480 10563 25483
rect 10962 25480 10968 25492
rect 10551 25452 10968 25480
rect 10551 25449 10563 25452
rect 10505 25443 10563 25449
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 12621 25483 12679 25489
rect 12621 25480 12633 25483
rect 11256 25452 12633 25480
rect 3970 25304 3976 25356
rect 4028 25344 4034 25356
rect 4065 25347 4123 25353
rect 4065 25344 4077 25347
rect 4028 25316 4077 25344
rect 4028 25304 4034 25316
rect 4065 25313 4077 25316
rect 4111 25344 4123 25347
rect 6273 25347 6331 25353
rect 6273 25344 6285 25347
rect 4111 25316 6285 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 6273 25313 6285 25316
rect 6319 25313 6331 25347
rect 6273 25307 6331 25313
rect 7101 25347 7159 25353
rect 7101 25313 7113 25347
rect 7147 25344 7159 25347
rect 8036 25344 8064 25440
rect 7147 25316 8064 25344
rect 8481 25347 8539 25353
rect 7147 25313 7159 25316
rect 7101 25307 7159 25313
rect 8481 25313 8493 25347
rect 8527 25344 8539 25347
rect 8754 25344 8760 25356
rect 8527 25316 8760 25344
rect 8527 25313 8539 25316
rect 8481 25307 8539 25313
rect 8754 25304 8760 25316
rect 8812 25344 8818 25356
rect 9582 25344 9588 25356
rect 8812 25316 9588 25344
rect 8812 25304 8818 25316
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 9953 25347 10011 25353
rect 9953 25313 9965 25347
rect 9999 25344 10011 25347
rect 10229 25347 10287 25353
rect 10229 25344 10241 25347
rect 9999 25316 10241 25344
rect 9999 25313 10011 25316
rect 9953 25307 10011 25313
rect 10229 25313 10241 25316
rect 10275 25313 10287 25347
rect 10229 25307 10287 25313
rect 10686 25304 10692 25356
rect 10744 25344 10750 25356
rect 11256 25344 11284 25452
rect 12621 25449 12633 25452
rect 12667 25449 12679 25483
rect 14185 25483 14243 25489
rect 14185 25480 14197 25483
rect 12621 25443 12679 25449
rect 13188 25452 14197 25480
rect 13188 25412 13216 25452
rect 14185 25449 14197 25452
rect 14231 25449 14243 25483
rect 14185 25443 14243 25449
rect 14461 25483 14519 25489
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 17126 25480 17132 25492
rect 14507 25452 17132 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 17126 25440 17132 25452
rect 17184 25440 17190 25492
rect 17313 25483 17371 25489
rect 17313 25449 17325 25483
rect 17359 25480 17371 25483
rect 20070 25480 20076 25492
rect 17359 25452 20076 25480
rect 17359 25449 17371 25452
rect 17313 25443 17371 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 20165 25483 20223 25489
rect 20165 25449 20177 25483
rect 20211 25480 20223 25483
rect 21818 25480 21824 25492
rect 20211 25452 21824 25480
rect 20211 25449 20223 25452
rect 20165 25443 20223 25449
rect 21818 25440 21824 25452
rect 21876 25440 21882 25492
rect 22189 25483 22247 25489
rect 22189 25449 22201 25483
rect 22235 25480 22247 25483
rect 22373 25483 22431 25489
rect 22373 25480 22385 25483
rect 22235 25452 22385 25480
rect 22235 25449 22247 25452
rect 22189 25443 22247 25449
rect 22373 25449 22385 25452
rect 22419 25480 22431 25483
rect 22830 25480 22836 25492
rect 22419 25452 22836 25480
rect 22419 25449 22431 25452
rect 22373 25443 22431 25449
rect 22830 25440 22836 25452
rect 22888 25440 22894 25492
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25480 23075 25483
rect 24762 25480 24768 25492
rect 23063 25452 24768 25480
rect 23063 25449 23075 25452
rect 23017 25443 23075 25449
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 16114 25412 16120 25424
rect 12360 25384 13216 25412
rect 13280 25384 16120 25412
rect 10744 25316 11284 25344
rect 10744 25304 10750 25316
rect 2866 25276 2872 25288
rect 2827 25248 2872 25276
rect 2866 25236 2872 25248
rect 2924 25236 2930 25288
rect 3050 25276 3056 25288
rect 3011 25248 3056 25276
rect 3050 25236 3056 25248
rect 3108 25236 3114 25288
rect 5534 25236 5540 25288
rect 5592 25276 5598 25288
rect 5721 25279 5779 25285
rect 5721 25276 5733 25279
rect 5592 25248 5733 25276
rect 5592 25236 5598 25248
rect 5721 25245 5733 25248
rect 5767 25245 5779 25279
rect 5721 25239 5779 25245
rect 5813 25279 5871 25285
rect 5813 25245 5825 25279
rect 5859 25245 5871 25279
rect 5813 25239 5871 25245
rect 3789 25211 3847 25217
rect 3789 25208 3801 25211
rect 2424 25180 3801 25208
rect 2424 25152 2452 25180
rect 3789 25177 3801 25180
rect 3835 25177 3847 25211
rect 3789 25171 3847 25177
rect 4062 25168 4068 25220
rect 4120 25208 4126 25220
rect 5261 25211 5319 25217
rect 5261 25208 5273 25211
rect 4120 25180 5273 25208
rect 4120 25168 4126 25180
rect 5261 25177 5273 25180
rect 5307 25177 5319 25211
rect 5261 25171 5319 25177
rect 5442 25168 5448 25220
rect 5500 25208 5506 25220
rect 5828 25208 5856 25239
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 8573 25279 8631 25285
rect 8573 25276 8585 25279
rect 8352 25248 8585 25276
rect 8352 25236 8358 25248
rect 8573 25245 8585 25248
rect 8619 25245 8631 25279
rect 8573 25239 8631 25245
rect 8665 25279 8723 25285
rect 8665 25245 8677 25279
rect 8711 25276 8723 25279
rect 9122 25276 9128 25288
rect 8711 25248 9128 25276
rect 8711 25245 8723 25248
rect 8665 25239 8723 25245
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 11256 25276 11284 25316
rect 11333 25347 11391 25353
rect 11333 25313 11345 25347
rect 11379 25344 11391 25347
rect 11790 25344 11796 25356
rect 11379 25316 11796 25344
rect 11379 25313 11391 25316
rect 11333 25307 11391 25313
rect 11790 25304 11796 25316
rect 11848 25344 11854 25356
rect 12161 25347 12219 25353
rect 12161 25344 12173 25347
rect 11848 25316 12173 25344
rect 11848 25304 11854 25316
rect 12161 25313 12173 25316
rect 12207 25313 12219 25347
rect 12161 25307 12219 25313
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 11256 25248 11437 25276
rect 11425 25245 11437 25248
rect 11471 25245 11483 25279
rect 11606 25276 11612 25288
rect 11567 25248 11612 25276
rect 11425 25239 11483 25245
rect 11606 25236 11612 25248
rect 11664 25236 11670 25288
rect 12360 25276 12388 25384
rect 12437 25347 12495 25353
rect 12437 25313 12449 25347
rect 12483 25344 12495 25347
rect 12986 25344 12992 25356
rect 12483 25316 12992 25344
rect 12483 25313 12495 25316
rect 12437 25307 12495 25313
rect 12986 25304 12992 25316
rect 13044 25304 13050 25356
rect 11716 25248 12388 25276
rect 5500 25180 5856 25208
rect 7285 25211 7343 25217
rect 5500 25168 5506 25180
rect 7285 25177 7297 25211
rect 7331 25208 7343 25211
rect 10594 25208 10600 25220
rect 7331 25180 10600 25208
rect 7331 25177 7343 25180
rect 7285 25171 7343 25177
rect 10594 25168 10600 25180
rect 10652 25168 10658 25220
rect 10962 25208 10968 25220
rect 10923 25180 10968 25208
rect 10962 25168 10968 25180
rect 11020 25168 11026 25220
rect 1946 25140 1952 25152
rect 1907 25112 1952 25140
rect 1946 25100 1952 25112
rect 2004 25100 2010 25152
rect 2314 25140 2320 25152
rect 2275 25112 2320 25140
rect 2314 25100 2320 25112
rect 2372 25100 2378 25152
rect 2406 25100 2412 25152
rect 2464 25140 2470 25152
rect 3418 25140 3424 25152
rect 2464 25112 2509 25140
rect 3379 25112 3424 25140
rect 2464 25100 2470 25112
rect 3418 25100 3424 25112
rect 3476 25100 3482 25152
rect 3510 25100 3516 25152
rect 3568 25140 3574 25152
rect 4617 25143 4675 25149
rect 4617 25140 4629 25143
rect 3568 25112 4629 25140
rect 3568 25100 3574 25112
rect 4617 25109 4629 25112
rect 4663 25109 4675 25143
rect 5074 25140 5080 25152
rect 5035 25112 5080 25140
rect 4617 25103 4675 25109
rect 5074 25100 5080 25112
rect 5132 25100 5138 25152
rect 6638 25140 6644 25152
rect 6599 25112 6644 25140
rect 6638 25100 6644 25112
rect 6696 25100 6702 25152
rect 8113 25143 8171 25149
rect 8113 25109 8125 25143
rect 8159 25140 8171 25143
rect 8938 25140 8944 25152
rect 8159 25112 8944 25140
rect 8159 25109 8171 25112
rect 8113 25103 8171 25109
rect 8938 25100 8944 25112
rect 8996 25100 9002 25152
rect 9122 25140 9128 25152
rect 9083 25112 9128 25140
rect 9122 25100 9128 25112
rect 9180 25100 9186 25152
rect 10137 25143 10195 25149
rect 10137 25109 10149 25143
rect 10183 25140 10195 25143
rect 11716 25140 11744 25248
rect 12710 25236 12716 25288
rect 12768 25276 12774 25288
rect 13081 25279 13139 25285
rect 13081 25276 13093 25279
rect 12768 25248 13093 25276
rect 12768 25236 12774 25248
rect 13081 25245 13093 25248
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 13170 25236 13176 25288
rect 13228 25276 13234 25288
rect 13280 25285 13308 25384
rect 16114 25372 16120 25384
rect 16172 25372 16178 25424
rect 21542 25412 21548 25424
rect 21503 25384 21548 25412
rect 21542 25372 21548 25384
rect 21600 25412 21606 25424
rect 23750 25412 23756 25424
rect 21600 25384 22876 25412
rect 23711 25384 23756 25412
rect 21600 25372 21606 25384
rect 14277 25347 14335 25353
rect 14277 25313 14289 25347
rect 14323 25344 14335 25347
rect 14458 25344 14464 25356
rect 14323 25316 14464 25344
rect 14323 25313 14335 25316
rect 14277 25307 14335 25313
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 15562 25304 15568 25356
rect 15620 25344 15626 25356
rect 15841 25347 15899 25353
rect 15841 25344 15853 25347
rect 15620 25316 15853 25344
rect 15620 25304 15626 25316
rect 15841 25313 15853 25316
rect 15887 25313 15899 25347
rect 15841 25307 15899 25313
rect 15933 25347 15991 25353
rect 15933 25313 15945 25347
rect 15979 25344 15991 25347
rect 16206 25344 16212 25356
rect 15979 25316 16212 25344
rect 15979 25313 15991 25316
rect 15933 25307 15991 25313
rect 16206 25304 16212 25316
rect 16264 25304 16270 25356
rect 17034 25304 17040 25356
rect 17092 25344 17098 25356
rect 22848 25353 22876 25384
rect 23750 25372 23756 25384
rect 23808 25372 23814 25424
rect 24394 25412 24400 25424
rect 24355 25384 24400 25412
rect 24394 25372 24400 25384
rect 24452 25372 24458 25424
rect 17129 25347 17187 25353
rect 17129 25344 17141 25347
rect 17092 25316 17141 25344
rect 17092 25304 17098 25316
rect 17129 25313 17141 25316
rect 17175 25313 17187 25347
rect 17129 25307 17187 25313
rect 18417 25347 18475 25353
rect 18417 25313 18429 25347
rect 18463 25313 18475 25347
rect 18417 25307 18475 25313
rect 19981 25347 20039 25353
rect 19981 25313 19993 25347
rect 20027 25313 20039 25347
rect 19981 25307 20039 25313
rect 21729 25347 21787 25353
rect 21729 25313 21741 25347
rect 21775 25344 21787 25347
rect 22189 25347 22247 25353
rect 22189 25344 22201 25347
rect 21775 25316 22201 25344
rect 21775 25313 21787 25316
rect 21729 25307 21787 25313
rect 22189 25313 22201 25316
rect 22235 25313 22247 25347
rect 22189 25307 22247 25313
rect 22833 25347 22891 25353
rect 22833 25313 22845 25347
rect 22879 25313 22891 25347
rect 24486 25344 24492 25356
rect 24447 25316 24492 25344
rect 22833 25307 22891 25313
rect 13265 25279 13323 25285
rect 13265 25276 13277 25279
rect 13228 25248 13277 25276
rect 13228 25236 13234 25248
rect 13265 25245 13277 25248
rect 13311 25245 13323 25279
rect 13265 25239 13323 25245
rect 14185 25279 14243 25285
rect 14185 25245 14197 25279
rect 14231 25276 14243 25279
rect 16114 25276 16120 25288
rect 14231 25248 15976 25276
rect 16075 25248 16120 25276
rect 14231 25245 14243 25248
rect 14185 25239 14243 25245
rect 15473 25211 15531 25217
rect 15473 25208 15485 25211
rect 13271 25180 15485 25208
rect 11974 25140 11980 25152
rect 10183 25112 11744 25140
rect 11935 25112 11980 25140
rect 10183 25109 10195 25112
rect 10137 25103 10195 25109
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12161 25143 12219 25149
rect 12161 25109 12173 25143
rect 12207 25140 12219 25143
rect 13271 25140 13299 25180
rect 15473 25177 15485 25180
rect 15519 25177 15531 25211
rect 15948 25208 15976 25248
rect 16114 25236 16120 25248
rect 16172 25236 16178 25288
rect 18432 25208 18460 25307
rect 19996 25276 20024 25307
rect 24486 25304 24492 25316
rect 24544 25304 24550 25356
rect 25590 25344 25596 25356
rect 25551 25316 25596 25344
rect 25590 25304 25596 25316
rect 25648 25304 25654 25356
rect 20070 25276 20076 25288
rect 19983 25248 20076 25276
rect 20070 25236 20076 25248
rect 20128 25276 20134 25288
rect 24673 25279 24731 25285
rect 20128 25248 24256 25276
rect 20128 25236 20134 25248
rect 18506 25208 18512 25220
rect 15948 25180 18512 25208
rect 15473 25171 15531 25177
rect 18506 25168 18512 25180
rect 18564 25168 18570 25220
rect 18601 25211 18659 25217
rect 18601 25177 18613 25211
rect 18647 25208 18659 25211
rect 20622 25208 20628 25220
rect 18647 25180 20628 25208
rect 18647 25177 18659 25180
rect 18601 25171 18659 25177
rect 20622 25168 20628 25180
rect 20680 25168 20686 25220
rect 21913 25211 21971 25217
rect 21913 25177 21925 25211
rect 21959 25208 21971 25211
rect 24118 25208 24124 25220
rect 21959 25180 24124 25208
rect 21959 25177 21971 25180
rect 21913 25171 21971 25177
rect 24118 25168 24124 25180
rect 24176 25168 24182 25220
rect 24228 25208 24256 25248
rect 24673 25245 24685 25279
rect 24719 25276 24731 25279
rect 24854 25276 24860 25288
rect 24719 25248 24860 25276
rect 24719 25245 24731 25248
rect 24673 25239 24731 25245
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 25777 25211 25835 25217
rect 25777 25208 25789 25211
rect 24228 25180 25789 25208
rect 25777 25177 25789 25180
rect 25823 25177 25835 25211
rect 25777 25171 25835 25177
rect 12207 25112 13299 25140
rect 15105 25143 15163 25149
rect 12207 25109 12219 25112
rect 12161 25103 12219 25109
rect 15105 25109 15117 25143
rect 15151 25140 15163 25143
rect 15286 25140 15292 25152
rect 15151 25112 15292 25140
rect 15151 25109 15163 25112
rect 15105 25103 15163 25109
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 16574 25140 16580 25152
rect 16535 25112 16580 25140
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 18138 25140 18144 25152
rect 18099 25112 18144 25140
rect 18138 25100 18144 25112
rect 18196 25100 18202 25152
rect 22554 25100 22560 25152
rect 22612 25140 22618 25152
rect 22649 25143 22707 25149
rect 22649 25140 22661 25143
rect 22612 25112 22661 25140
rect 22612 25100 22618 25112
rect 22649 25109 22661 25112
rect 22695 25109 22707 25143
rect 24026 25140 24032 25152
rect 23987 25112 24032 25140
rect 22649 25103 22707 25109
rect 24026 25100 24032 25112
rect 24084 25100 24090 25152
rect 25222 25140 25228 25152
rect 25183 25112 25228 25140
rect 25222 25100 25228 25112
rect 25280 25100 25286 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1394 24896 1400 24948
rect 1452 24936 1458 24948
rect 3510 24936 3516 24948
rect 1452 24908 3516 24936
rect 1452 24896 1458 24908
rect 3510 24896 3516 24908
rect 3568 24896 3574 24948
rect 4338 24896 4344 24948
rect 4396 24936 4402 24948
rect 8846 24936 8852 24948
rect 4396 24908 8852 24936
rect 4396 24896 4402 24908
rect 8846 24896 8852 24908
rect 8904 24896 8910 24948
rect 10686 24936 10692 24948
rect 10647 24908 10692 24936
rect 10686 24896 10692 24908
rect 10744 24896 10750 24948
rect 12986 24936 12992 24948
rect 12947 24908 12992 24936
rect 12986 24896 12992 24908
rect 13044 24896 13050 24948
rect 13354 24896 13360 24948
rect 13412 24936 13418 24948
rect 16114 24936 16120 24948
rect 13412 24908 15976 24936
rect 16075 24908 16120 24936
rect 13412 24896 13418 24908
rect 5442 24828 5448 24880
rect 5500 24868 5506 24880
rect 5500 24840 6960 24868
rect 5500 24828 5506 24840
rect 1670 24760 1676 24812
rect 1728 24800 1734 24812
rect 2133 24803 2191 24809
rect 2133 24800 2145 24803
rect 1728 24772 2145 24800
rect 1728 24760 1734 24772
rect 2133 24769 2145 24772
rect 2179 24769 2191 24803
rect 2133 24763 2191 24769
rect 2498 24760 2504 24812
rect 2556 24800 2562 24812
rect 2682 24800 2688 24812
rect 2556 24772 2688 24800
rect 2556 24760 2562 24772
rect 2682 24760 2688 24772
rect 2740 24760 2746 24812
rect 6932 24800 6960 24840
rect 12710 24828 12716 24880
rect 12768 24868 12774 24880
rect 12768 24840 13768 24868
rect 12768 24828 12774 24840
rect 7098 24800 7104 24812
rect 6932 24772 7104 24800
rect 7098 24760 7104 24772
rect 7156 24760 7162 24812
rect 7282 24800 7288 24812
rect 7243 24772 7288 24800
rect 7282 24760 7288 24772
rect 7340 24760 7346 24812
rect 7466 24800 7472 24812
rect 7427 24772 7472 24800
rect 7466 24760 7472 24772
rect 7524 24760 7530 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 13170 24800 13176 24812
rect 11931 24772 13176 24800
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 13170 24760 13176 24772
rect 13228 24760 13234 24812
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24769 13691 24803
rect 13740 24800 13768 24840
rect 13814 24828 13820 24880
rect 13872 24868 13878 24880
rect 13872 24840 15240 24868
rect 13872 24828 13878 24840
rect 14369 24803 14427 24809
rect 14369 24800 14381 24803
rect 13740 24772 14381 24800
rect 13633 24763 13691 24769
rect 14369 24769 14381 24772
rect 14415 24769 14427 24803
rect 15212 24800 15240 24840
rect 15286 24828 15292 24880
rect 15344 24868 15350 24880
rect 15948 24868 15976 24908
rect 16114 24896 16120 24908
rect 16172 24896 16178 24948
rect 17034 24896 17040 24948
rect 17092 24936 17098 24948
rect 17497 24939 17555 24945
rect 17497 24936 17509 24939
rect 17092 24908 17509 24936
rect 17092 24896 17098 24908
rect 17497 24905 17509 24908
rect 17543 24905 17555 24939
rect 18506 24936 18512 24948
rect 18467 24908 18512 24936
rect 17497 24899 17555 24905
rect 18506 24896 18512 24908
rect 18564 24896 18570 24948
rect 20622 24896 20628 24948
rect 20680 24936 20686 24948
rect 23750 24936 23756 24948
rect 20680 24908 23756 24936
rect 20680 24896 20686 24908
rect 23750 24896 23756 24908
rect 23808 24896 23814 24948
rect 24762 24936 24768 24948
rect 24723 24908 24768 24936
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 21450 24868 21456 24880
rect 15344 24840 15700 24868
rect 15948 24840 21456 24868
rect 15344 24828 15350 24840
rect 15672 24809 15700 24840
rect 21450 24828 21456 24840
rect 21508 24828 21514 24880
rect 15657 24803 15715 24809
rect 15212 24772 15608 24800
rect 14369 24763 14427 24769
rect 1949 24735 2007 24741
rect 1949 24701 1961 24735
rect 1995 24732 2007 24735
rect 2406 24732 2412 24744
rect 1995 24704 2412 24732
rect 1995 24701 2007 24704
rect 1949 24695 2007 24701
rect 2406 24692 2412 24704
rect 2464 24692 2470 24744
rect 3145 24735 3203 24741
rect 3145 24701 3157 24735
rect 3191 24732 3203 24735
rect 3234 24732 3240 24744
rect 3191 24704 3240 24732
rect 3191 24701 3203 24704
rect 3145 24695 3203 24701
rect 3234 24692 3240 24704
rect 3292 24692 3298 24744
rect 3418 24741 3424 24744
rect 3412 24732 3424 24741
rect 3379 24704 3424 24732
rect 3412 24695 3424 24704
rect 3476 24732 3482 24744
rect 4430 24732 4436 24744
rect 3476 24704 4436 24732
rect 3418 24692 3424 24695
rect 3476 24692 3482 24704
rect 4430 24692 4436 24704
rect 4488 24732 4494 24744
rect 5261 24735 5319 24741
rect 5261 24732 5273 24735
rect 4488 24704 5273 24732
rect 4488 24692 4494 24704
rect 5261 24701 5273 24704
rect 5307 24732 5319 24735
rect 5442 24732 5448 24744
rect 5307 24704 5448 24732
rect 5307 24701 5319 24704
rect 5261 24695 5319 24701
rect 5442 24692 5448 24704
rect 5500 24692 5506 24744
rect 5629 24735 5687 24741
rect 5629 24701 5641 24735
rect 5675 24732 5687 24735
rect 6273 24735 6331 24741
rect 6273 24732 6285 24735
rect 5675 24704 6285 24732
rect 5675 24701 5687 24704
rect 5629 24695 5687 24701
rect 6273 24701 6285 24704
rect 6319 24732 6331 24735
rect 6546 24732 6552 24744
rect 6319 24704 6552 24732
rect 6319 24701 6331 24704
rect 6273 24695 6331 24701
rect 6546 24692 6552 24704
rect 6604 24692 6610 24744
rect 7006 24692 7012 24744
rect 7064 24732 7070 24744
rect 8205 24735 8263 24741
rect 8205 24732 8217 24735
rect 7064 24704 8217 24732
rect 7064 24692 7070 24704
rect 8205 24701 8217 24704
rect 8251 24732 8263 24735
rect 8294 24732 8300 24744
rect 8251 24704 8300 24732
rect 8251 24701 8263 24704
rect 8205 24695 8263 24701
rect 8294 24692 8300 24704
rect 8352 24692 8358 24744
rect 8478 24732 8484 24744
rect 8439 24704 8484 24732
rect 8478 24692 8484 24704
rect 8536 24692 8542 24744
rect 11333 24735 11391 24741
rect 11333 24701 11345 24735
rect 11379 24732 11391 24735
rect 11974 24732 11980 24744
rect 11379 24704 11980 24732
rect 11379 24701 11391 24704
rect 11333 24695 11391 24701
rect 11974 24692 11980 24704
rect 12032 24692 12038 24744
rect 12253 24735 12311 24741
rect 12253 24701 12265 24735
rect 12299 24732 12311 24735
rect 13648 24732 13676 24763
rect 14921 24735 14979 24741
rect 12299 24704 12756 24732
rect 13648 24704 14044 24732
rect 12299 24701 12311 24704
rect 12253 24695 12311 24701
rect 2222 24664 2228 24676
rect 1596 24636 2228 24664
rect 1596 24605 1624 24636
rect 2222 24624 2228 24636
rect 2280 24624 2286 24676
rect 2682 24664 2688 24676
rect 2332 24636 2688 24664
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 1946 24556 1952 24608
rect 2004 24596 2010 24608
rect 2041 24599 2099 24605
rect 2041 24596 2053 24599
rect 2004 24568 2053 24596
rect 2004 24556 2010 24568
rect 2041 24565 2053 24568
rect 2087 24596 2099 24599
rect 2332 24596 2360 24636
rect 2682 24624 2688 24636
rect 2740 24624 2746 24676
rect 6641 24667 6699 24673
rect 6641 24633 6653 24667
rect 6687 24664 6699 24667
rect 6687 24636 7236 24664
rect 6687 24633 6699 24636
rect 6641 24627 6699 24633
rect 7208 24608 7236 24636
rect 8110 24624 8116 24676
rect 8168 24664 8174 24676
rect 8748 24667 8806 24673
rect 8748 24664 8760 24667
rect 8168 24636 8760 24664
rect 8168 24624 8174 24636
rect 8748 24633 8760 24636
rect 8794 24664 8806 24667
rect 9122 24664 9128 24676
rect 8794 24636 9128 24664
rect 8794 24633 8806 24636
rect 8748 24627 8806 24633
rect 9122 24624 9128 24636
rect 9180 24664 9186 24676
rect 9582 24664 9588 24676
rect 9180 24636 9588 24664
rect 9180 24624 9186 24636
rect 9582 24624 9588 24636
rect 9640 24624 9646 24676
rect 11057 24667 11115 24673
rect 11057 24633 11069 24667
rect 11103 24664 11115 24667
rect 11606 24664 11612 24676
rect 11103 24636 11612 24664
rect 11103 24633 11115 24636
rect 11057 24627 11115 24633
rect 11606 24624 11612 24636
rect 11664 24664 11670 24676
rect 12158 24664 12164 24676
rect 11664 24636 12164 24664
rect 11664 24624 11670 24636
rect 12158 24624 12164 24636
rect 12216 24624 12222 24676
rect 2087 24568 2360 24596
rect 2087 24565 2099 24568
rect 2041 24559 2099 24565
rect 2866 24556 2872 24608
rect 2924 24596 2930 24608
rect 3053 24599 3111 24605
rect 3053 24596 3065 24599
rect 2924 24568 3065 24596
rect 2924 24556 2930 24568
rect 3053 24565 3065 24568
rect 3099 24596 3111 24599
rect 3326 24596 3332 24608
rect 3099 24568 3332 24596
rect 3099 24565 3111 24568
rect 3053 24559 3111 24565
rect 3326 24556 3332 24568
rect 3384 24556 3390 24608
rect 3878 24556 3884 24608
rect 3936 24596 3942 24608
rect 4525 24599 4583 24605
rect 4525 24596 4537 24599
rect 3936 24568 4537 24596
rect 3936 24556 3942 24568
rect 4525 24565 4537 24568
rect 4571 24565 4583 24599
rect 4525 24559 4583 24565
rect 4798 24556 4804 24608
rect 4856 24596 4862 24608
rect 5813 24599 5871 24605
rect 5813 24596 5825 24599
rect 4856 24568 5825 24596
rect 4856 24556 4862 24568
rect 5813 24565 5825 24568
rect 5859 24565 5871 24599
rect 5813 24559 5871 24565
rect 6730 24556 6736 24608
rect 6788 24596 6794 24608
rect 6825 24599 6883 24605
rect 6825 24596 6837 24599
rect 6788 24568 6837 24596
rect 6788 24556 6794 24568
rect 6825 24565 6837 24568
rect 6871 24565 6883 24599
rect 7190 24596 7196 24608
rect 7151 24568 7196 24596
rect 6825 24559 6883 24565
rect 7190 24556 7196 24568
rect 7248 24556 7254 24608
rect 9858 24596 9864 24608
rect 9819 24568 9864 24596
rect 9858 24556 9864 24568
rect 9916 24556 9922 24608
rect 11514 24596 11520 24608
rect 11475 24568 11520 24596
rect 11514 24556 11520 24568
rect 11572 24556 11578 24608
rect 12728 24596 12756 24704
rect 12894 24664 12900 24676
rect 12807 24636 12900 24664
rect 12894 24624 12900 24636
rect 12952 24664 12958 24676
rect 12952 24636 13492 24664
rect 12952 24624 12958 24636
rect 13354 24596 13360 24608
rect 12728 24568 13360 24596
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 13464 24605 13492 24636
rect 14016 24608 14044 24704
rect 14921 24701 14933 24735
rect 14967 24732 14979 24735
rect 15580 24732 15608 24772
rect 15657 24769 15669 24803
rect 15703 24769 15715 24803
rect 15657 24763 15715 24769
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19981 24803 20039 24809
rect 19981 24800 19993 24803
rect 19024 24772 19993 24800
rect 19024 24760 19030 24772
rect 19981 24769 19993 24772
rect 20027 24800 20039 24803
rect 21085 24803 21143 24809
rect 21085 24800 21097 24803
rect 20027 24772 21097 24800
rect 20027 24769 20039 24772
rect 19981 24763 20039 24769
rect 21085 24769 21097 24772
rect 21131 24800 21143 24803
rect 22554 24800 22560 24812
rect 21131 24772 22560 24800
rect 21131 24769 21143 24772
rect 21085 24763 21143 24769
rect 22554 24760 22560 24772
rect 22612 24800 22618 24812
rect 22612 24772 23244 24800
rect 22612 24760 22618 24772
rect 16206 24732 16212 24744
rect 14967 24704 15516 24732
rect 15580 24704 16212 24732
rect 14967 24701 14979 24704
rect 14921 24695 14979 24701
rect 14734 24624 14740 24676
rect 14792 24664 14798 24676
rect 15381 24667 15439 24673
rect 15381 24664 15393 24667
rect 14792 24636 15393 24664
rect 14792 24624 14798 24636
rect 15381 24633 15393 24636
rect 15427 24633 15439 24667
rect 15381 24627 15439 24633
rect 15488 24608 15516 24704
rect 16206 24692 16212 24704
rect 16264 24732 16270 24744
rect 16393 24735 16451 24741
rect 16393 24732 16405 24735
rect 16264 24704 16405 24732
rect 16264 24692 16270 24704
rect 16393 24701 16405 24704
rect 16439 24701 16451 24735
rect 16574 24732 16580 24744
rect 16487 24704 16580 24732
rect 16393 24695 16451 24701
rect 16574 24692 16580 24704
rect 16632 24692 16638 24744
rect 18049 24735 18107 24741
rect 18049 24701 18061 24735
rect 18095 24732 18107 24735
rect 18138 24732 18144 24744
rect 18095 24704 18144 24732
rect 18095 24701 18107 24704
rect 18049 24695 18107 24701
rect 18138 24692 18144 24704
rect 18196 24692 18202 24744
rect 19061 24735 19119 24741
rect 19061 24732 19073 24735
rect 18892 24704 19073 24732
rect 16592 24664 16620 24692
rect 16592 24636 18276 24664
rect 13449 24599 13507 24605
rect 13449 24565 13461 24599
rect 13495 24596 13507 24599
rect 13722 24596 13728 24608
rect 13495 24568 13728 24596
rect 13495 24565 13507 24568
rect 13449 24559 13507 24565
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 13998 24596 14004 24608
rect 13959 24568 14004 24596
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 14826 24556 14832 24608
rect 14884 24596 14890 24608
rect 15013 24599 15071 24605
rect 15013 24596 15025 24599
rect 14884 24568 15025 24596
rect 14884 24556 14890 24568
rect 15013 24565 15025 24568
rect 15059 24565 15071 24599
rect 15470 24596 15476 24608
rect 15431 24568 15476 24596
rect 15013 24559 15071 24565
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 16758 24596 16764 24608
rect 16719 24568 16764 24596
rect 16758 24556 16764 24568
rect 16816 24556 16822 24608
rect 17034 24556 17040 24608
rect 17092 24596 17098 24608
rect 18248 24605 18276 24636
rect 18892 24608 18920 24704
rect 19061 24701 19073 24704
rect 19107 24701 19119 24735
rect 19061 24695 19119 24701
rect 21450 24692 21456 24744
rect 21508 24732 21514 24744
rect 22278 24732 22284 24744
rect 21508 24704 22284 24732
rect 21508 24692 21514 24704
rect 22278 24692 22284 24704
rect 22336 24732 22342 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 22336 24704 22385 24732
rect 22336 24692 22342 24704
rect 22373 24701 22385 24704
rect 22419 24732 22431 24735
rect 22646 24732 22652 24744
rect 22419 24704 22652 24732
rect 22419 24701 22431 24704
rect 22373 24695 22431 24701
rect 22646 24692 22652 24704
rect 22704 24692 22710 24744
rect 23216 24732 23244 24772
rect 23750 24760 23756 24812
rect 23808 24800 23814 24812
rect 24121 24803 24179 24809
rect 24121 24800 24133 24803
rect 23808 24772 24133 24800
rect 23808 24760 23814 24772
rect 24121 24769 24133 24772
rect 24167 24769 24179 24803
rect 24121 24763 24179 24769
rect 24213 24803 24271 24809
rect 24213 24769 24225 24803
rect 24259 24800 24271 24803
rect 24854 24800 24860 24812
rect 24259 24772 24860 24800
rect 24259 24769 24271 24772
rect 24213 24763 24271 24769
rect 24228 24732 24256 24763
rect 24854 24760 24860 24772
rect 24912 24800 24918 24812
rect 25041 24803 25099 24809
rect 25041 24800 25053 24803
rect 24912 24772 25053 24800
rect 24912 24760 24918 24772
rect 25041 24769 25053 24772
rect 25087 24769 25099 24803
rect 25041 24763 25099 24769
rect 25222 24732 25228 24744
rect 23216 24704 24256 24732
rect 25183 24704 25228 24732
rect 20901 24667 20959 24673
rect 20901 24664 20913 24667
rect 20272 24636 20913 24664
rect 17129 24599 17187 24605
rect 17129 24596 17141 24599
rect 17092 24568 17141 24596
rect 17092 24556 17098 24568
rect 17129 24565 17141 24568
rect 17175 24565 17187 24599
rect 17129 24559 17187 24565
rect 18233 24599 18291 24605
rect 18233 24565 18245 24599
rect 18279 24565 18291 24599
rect 18874 24596 18880 24608
rect 18835 24568 18880 24596
rect 18233 24559 18291 24565
rect 18874 24556 18880 24568
rect 18932 24556 18938 24608
rect 19242 24596 19248 24608
rect 19203 24568 19248 24596
rect 19242 24556 19248 24568
rect 19300 24556 19306 24608
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 20272 24605 20300 24636
rect 20901 24633 20913 24636
rect 20947 24633 20959 24667
rect 21910 24664 21916 24676
rect 21823 24636 21916 24664
rect 20901 24627 20959 24633
rect 21910 24624 21916 24636
rect 21968 24664 21974 24676
rect 22465 24667 22523 24673
rect 22465 24664 22477 24667
rect 21968 24636 22477 24664
rect 21968 24624 21974 24636
rect 22465 24633 22477 24636
rect 22511 24633 22523 24667
rect 22465 24627 22523 24633
rect 23216 24608 23244 24704
rect 25222 24692 25228 24704
rect 25280 24692 25286 24744
rect 23477 24667 23535 24673
rect 23477 24633 23489 24667
rect 23523 24664 23535 24667
rect 23934 24664 23940 24676
rect 23523 24636 23940 24664
rect 23523 24633 23535 24636
rect 23477 24627 23535 24633
rect 23934 24624 23940 24636
rect 23992 24664 23998 24676
rect 24029 24667 24087 24673
rect 24029 24664 24041 24667
rect 23992 24636 24041 24664
rect 23992 24624 23998 24636
rect 24029 24633 24041 24636
rect 24075 24633 24087 24667
rect 24029 24627 24087 24633
rect 25130 24624 25136 24676
rect 25188 24664 25194 24676
rect 25590 24664 25596 24676
rect 25188 24636 25596 24664
rect 25188 24624 25194 24636
rect 25590 24624 25596 24636
rect 25648 24664 25654 24676
rect 25777 24667 25835 24673
rect 25777 24664 25789 24667
rect 25648 24636 25789 24664
rect 25648 24624 25654 24636
rect 25777 24633 25789 24636
rect 25823 24633 25835 24667
rect 25777 24627 25835 24633
rect 20257 24599 20315 24605
rect 20257 24596 20269 24599
rect 19484 24568 20269 24596
rect 19484 24556 19490 24568
rect 20257 24565 20269 24568
rect 20303 24565 20315 24599
rect 20438 24596 20444 24608
rect 20399 24568 20444 24596
rect 20257 24559 20315 24565
rect 20438 24556 20444 24568
rect 20496 24556 20502 24608
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 20809 24599 20867 24605
rect 20809 24596 20821 24599
rect 20588 24568 20821 24596
rect 20588 24556 20594 24568
rect 20809 24565 20821 24568
rect 20855 24565 20867 24599
rect 22002 24596 22008 24608
rect 21963 24568 22008 24596
rect 20809 24559 20867 24565
rect 22002 24556 22008 24568
rect 22060 24556 22066 24608
rect 23109 24599 23167 24605
rect 23109 24565 23121 24599
rect 23155 24596 23167 24599
rect 23198 24596 23204 24608
rect 23155 24568 23204 24596
rect 23155 24565 23167 24568
rect 23109 24559 23167 24565
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23658 24596 23664 24608
rect 23619 24568 23664 24596
rect 23658 24556 23664 24568
rect 23716 24556 23722 24608
rect 25406 24596 25412 24608
rect 25367 24568 25412 24596
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1670 24352 1676 24404
rect 1728 24392 1734 24404
rect 1857 24395 1915 24401
rect 1857 24392 1869 24395
rect 1728 24364 1869 24392
rect 1728 24352 1734 24364
rect 1857 24361 1869 24364
rect 1903 24361 1915 24395
rect 1857 24355 1915 24361
rect 2317 24395 2375 24401
rect 2317 24361 2329 24395
rect 2363 24392 2375 24395
rect 3050 24392 3056 24404
rect 2363 24364 3056 24392
rect 2363 24361 2375 24364
rect 2317 24355 2375 24361
rect 3050 24352 3056 24364
rect 3108 24352 3114 24404
rect 3878 24392 3884 24404
rect 3839 24364 3884 24392
rect 3878 24352 3884 24364
rect 3936 24352 3942 24404
rect 4154 24352 4160 24404
rect 4212 24392 4218 24404
rect 4525 24395 4583 24401
rect 4525 24392 4537 24395
rect 4212 24364 4537 24392
rect 4212 24352 4218 24364
rect 4525 24361 4537 24364
rect 4571 24392 4583 24395
rect 4706 24392 4712 24404
rect 4571 24364 4712 24392
rect 4571 24361 4583 24364
rect 4525 24355 4583 24361
rect 4706 24352 4712 24364
rect 4764 24352 4770 24404
rect 6914 24352 6920 24404
rect 6972 24392 6978 24404
rect 7466 24392 7472 24404
rect 6972 24364 7472 24392
rect 6972 24352 6978 24364
rect 7466 24352 7472 24364
rect 7524 24392 7530 24404
rect 7653 24395 7711 24401
rect 7653 24392 7665 24395
rect 7524 24364 7665 24392
rect 7524 24352 7530 24364
rect 7653 24361 7665 24364
rect 7699 24361 7711 24395
rect 8110 24392 8116 24404
rect 8071 24364 8116 24392
rect 7653 24355 7711 24361
rect 8110 24352 8116 24364
rect 8168 24352 8174 24404
rect 8754 24392 8760 24404
rect 8715 24364 8760 24392
rect 8754 24352 8760 24364
rect 8812 24352 8818 24404
rect 9858 24352 9864 24404
rect 9916 24392 9922 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9916 24364 10149 24392
rect 9916 24352 9922 24364
rect 10137 24361 10149 24364
rect 10183 24361 10195 24395
rect 10686 24392 10692 24404
rect 10647 24364 10692 24392
rect 10137 24355 10195 24361
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 11146 24392 11152 24404
rect 11107 24364 11152 24392
rect 11146 24352 11152 24364
rect 11204 24352 11210 24404
rect 11790 24392 11796 24404
rect 11751 24364 11796 24392
rect 11790 24352 11796 24364
rect 11848 24352 11854 24404
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 14642 24392 14648 24404
rect 14323 24364 14648 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 14642 24352 14648 24364
rect 14700 24352 14706 24404
rect 18046 24352 18052 24404
rect 18104 24392 18110 24404
rect 18325 24395 18383 24401
rect 18325 24392 18337 24395
rect 18104 24364 18337 24392
rect 18104 24352 18110 24364
rect 18325 24361 18337 24364
rect 18371 24361 18383 24395
rect 19334 24392 19340 24404
rect 19295 24364 19340 24392
rect 18325 24355 18383 24361
rect 19334 24352 19340 24364
rect 19392 24352 19398 24404
rect 20070 24392 20076 24404
rect 20031 24364 20076 24392
rect 20070 24352 20076 24364
rect 20128 24352 20134 24404
rect 22002 24352 22008 24404
rect 22060 24392 22066 24404
rect 23109 24395 23167 24401
rect 23109 24392 23121 24395
rect 22060 24364 23121 24392
rect 22060 24352 22066 24364
rect 23109 24361 23121 24364
rect 23155 24392 23167 24395
rect 24118 24392 24124 24404
rect 23155 24364 24124 24392
rect 23155 24361 23167 24364
rect 23109 24355 23167 24361
rect 24118 24352 24124 24364
rect 24176 24352 24182 24404
rect 24210 24352 24216 24404
rect 24268 24392 24274 24404
rect 24305 24395 24363 24401
rect 24305 24392 24317 24395
rect 24268 24364 24317 24392
rect 24268 24352 24274 24364
rect 24305 24361 24317 24364
rect 24351 24361 24363 24395
rect 24305 24355 24363 24361
rect 25225 24395 25283 24401
rect 25225 24361 25237 24395
rect 25271 24392 25283 24395
rect 25314 24392 25320 24404
rect 25271 24364 25320 24392
rect 25271 24361 25283 24364
rect 25225 24355 25283 24361
rect 25314 24352 25320 24364
rect 25372 24352 25378 24404
rect 2498 24284 2504 24336
rect 2556 24324 2562 24336
rect 2777 24327 2835 24333
rect 2777 24324 2789 24327
rect 2556 24296 2789 24324
rect 2556 24284 2562 24296
rect 2777 24293 2789 24296
rect 2823 24293 2835 24327
rect 2777 24287 2835 24293
rect 2869 24327 2927 24333
rect 2869 24293 2881 24327
rect 2915 24324 2927 24327
rect 6086 24324 6092 24336
rect 2915 24296 6092 24324
rect 2915 24293 2927 24296
rect 2869 24287 2927 24293
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 1946 24216 1952 24268
rect 2004 24256 2010 24268
rect 2884 24256 2912 24287
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 10870 24284 10876 24336
rect 10928 24324 10934 24336
rect 11057 24327 11115 24333
rect 11057 24324 11069 24327
rect 10928 24296 11069 24324
rect 10928 24284 10934 24296
rect 11057 24293 11069 24296
rect 11103 24324 11115 24327
rect 11238 24324 11244 24336
rect 11103 24296 11244 24324
rect 11103 24293 11115 24296
rect 11057 24287 11115 24293
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 12066 24284 12072 24336
rect 12124 24324 12130 24336
rect 12621 24327 12679 24333
rect 12621 24324 12633 24327
rect 12124 24296 12633 24324
rect 12124 24284 12130 24296
rect 12621 24293 12633 24296
rect 12667 24293 12679 24327
rect 12621 24287 12679 24293
rect 17586 24284 17592 24336
rect 17644 24324 17650 24336
rect 17773 24327 17831 24333
rect 17773 24324 17785 24327
rect 17644 24296 17785 24324
rect 17644 24284 17650 24296
rect 17773 24293 17785 24296
rect 17819 24293 17831 24327
rect 17773 24287 17831 24293
rect 22833 24327 22891 24333
rect 22833 24293 22845 24327
rect 22879 24324 22891 24327
rect 24026 24324 24032 24336
rect 22879 24296 24032 24324
rect 22879 24293 22891 24296
rect 22833 24287 22891 24293
rect 24026 24284 24032 24296
rect 24084 24284 24090 24336
rect 5988 24259 6046 24265
rect 5988 24256 6000 24259
rect 2004 24228 2912 24256
rect 4080 24228 6000 24256
rect 2004 24216 2010 24228
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24188 3111 24191
rect 3326 24188 3332 24200
rect 3099 24160 3332 24188
rect 3099 24157 3111 24160
rect 3053 24151 3111 24157
rect 3326 24148 3332 24160
rect 3384 24188 3390 24200
rect 4080 24188 4108 24228
rect 5988 24225 6000 24228
rect 6034 24256 6046 24259
rect 6362 24256 6368 24268
rect 6034 24228 6368 24256
rect 6034 24225 6046 24228
rect 5988 24219 6046 24225
rect 6362 24216 6368 24228
rect 6420 24216 6426 24268
rect 8110 24216 8116 24268
rect 8168 24256 8174 24268
rect 8205 24259 8263 24265
rect 8205 24256 8217 24259
rect 8168 24228 8217 24256
rect 8168 24216 8174 24228
rect 8205 24225 8217 24228
rect 8251 24225 8263 24259
rect 12710 24256 12716 24268
rect 12671 24228 12716 24256
rect 8205 24219 8263 24225
rect 12710 24216 12716 24228
rect 12768 24216 12774 24268
rect 14093 24259 14151 24265
rect 14093 24225 14105 24259
rect 14139 24256 14151 24259
rect 14642 24256 14648 24268
rect 14139 24228 14648 24256
rect 14139 24225 14151 24228
rect 14093 24219 14151 24225
rect 14642 24216 14648 24228
rect 14700 24216 14706 24268
rect 16114 24256 16120 24268
rect 16075 24228 16120 24256
rect 16114 24216 16120 24228
rect 16172 24216 16178 24268
rect 17402 24216 17408 24268
rect 17460 24256 17466 24268
rect 17681 24259 17739 24265
rect 17681 24256 17693 24259
rect 17460 24228 17693 24256
rect 17460 24216 17466 24228
rect 17681 24225 17693 24228
rect 17727 24225 17739 24259
rect 17681 24219 17739 24225
rect 19058 24216 19064 24268
rect 19116 24256 19122 24268
rect 19153 24259 19211 24265
rect 19153 24256 19165 24259
rect 19116 24228 19165 24256
rect 19116 24216 19122 24228
rect 19153 24225 19165 24228
rect 19199 24225 19211 24259
rect 19153 24219 19211 24225
rect 21269 24259 21327 24265
rect 21269 24225 21281 24259
rect 21315 24256 21327 24259
rect 22097 24259 22155 24265
rect 22097 24256 22109 24259
rect 21315 24228 22109 24256
rect 21315 24225 21327 24228
rect 21269 24219 21327 24225
rect 22097 24225 22109 24228
rect 22143 24256 22155 24259
rect 22462 24256 22468 24268
rect 22143 24228 22468 24256
rect 22143 24225 22155 24228
rect 22097 24219 22155 24225
rect 22462 24216 22468 24228
rect 22520 24216 22526 24268
rect 23290 24216 23296 24268
rect 23348 24256 23354 24268
rect 23661 24259 23719 24265
rect 23661 24256 23673 24259
rect 23348 24228 23673 24256
rect 23348 24216 23354 24228
rect 23661 24225 23673 24228
rect 23707 24225 23719 24259
rect 23661 24219 23719 24225
rect 24854 24216 24860 24268
rect 24912 24256 24918 24268
rect 25317 24259 25375 24265
rect 25317 24256 25329 24259
rect 24912 24228 25329 24256
rect 24912 24216 24918 24228
rect 25317 24225 25329 24228
rect 25363 24225 25375 24259
rect 25317 24219 25375 24225
rect 4614 24188 4620 24200
rect 3384 24160 4108 24188
rect 4575 24160 4620 24188
rect 3384 24148 3390 24160
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24188 4859 24191
rect 5350 24188 5356 24200
rect 4847 24160 5356 24188
rect 4847 24157 4859 24160
rect 4801 24151 4859 24157
rect 5350 24148 5356 24160
rect 5408 24148 5414 24200
rect 5721 24191 5779 24197
rect 5721 24157 5733 24191
rect 5767 24157 5779 24191
rect 5721 24151 5779 24157
rect 5534 24120 5540 24132
rect 3160 24092 5540 24120
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 2409 24055 2467 24061
rect 2409 24021 2421 24055
rect 2455 24052 2467 24055
rect 3160 24052 3188 24092
rect 5534 24080 5540 24092
rect 5592 24080 5598 24132
rect 2455 24024 3188 24052
rect 2455 24021 2467 24024
rect 2409 24015 2467 24021
rect 3234 24012 3240 24064
rect 3292 24052 3298 24064
rect 3513 24055 3571 24061
rect 3513 24052 3525 24055
rect 3292 24024 3525 24052
rect 3292 24012 3298 24024
rect 3513 24021 3525 24024
rect 3559 24052 3571 24055
rect 3970 24052 3976 24064
rect 3559 24024 3976 24052
rect 3559 24021 3571 24024
rect 3513 24015 3571 24021
rect 3970 24012 3976 24024
rect 4028 24012 4034 24064
rect 4154 24052 4160 24064
rect 4115 24024 4160 24052
rect 4154 24012 4160 24024
rect 4212 24012 4218 24064
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5350 24052 5356 24064
rect 5307 24024 5356 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5350 24012 5356 24024
rect 5408 24012 5414 24064
rect 5736 24052 5764 24151
rect 9306 24148 9312 24200
rect 9364 24188 9370 24200
rect 9677 24191 9735 24197
rect 9677 24188 9689 24191
rect 9364 24160 9689 24188
rect 9364 24148 9370 24160
rect 9677 24157 9689 24160
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 11333 24191 11391 24197
rect 11333 24157 11345 24191
rect 11379 24188 11391 24191
rect 11790 24188 11796 24200
rect 11379 24160 11796 24188
rect 11379 24157 11391 24160
rect 11333 24151 11391 24157
rect 11790 24148 11796 24160
rect 11848 24148 11854 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 12805 24191 12863 24197
rect 12805 24188 12817 24191
rect 12207 24160 12817 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 12805 24157 12817 24160
rect 12851 24188 12863 24191
rect 13722 24188 13728 24200
rect 12851 24160 13728 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 15565 24191 15623 24197
rect 15565 24157 15577 24191
rect 15611 24188 15623 24191
rect 15746 24188 15752 24200
rect 15611 24160 15752 24188
rect 15611 24157 15623 24160
rect 15565 24151 15623 24157
rect 15746 24148 15752 24160
rect 15804 24148 15810 24200
rect 16206 24188 16212 24200
rect 16167 24160 16212 24188
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 16298 24148 16304 24200
rect 16356 24188 16362 24200
rect 17218 24188 17224 24200
rect 16356 24160 16401 24188
rect 17131 24160 17224 24188
rect 16356 24148 16362 24160
rect 17218 24148 17224 24160
rect 17276 24188 17282 24200
rect 17865 24191 17923 24197
rect 17865 24188 17877 24191
rect 17276 24160 17877 24188
rect 17276 24148 17282 24160
rect 17865 24157 17877 24160
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 21450 24148 21456 24200
rect 21508 24188 21514 24200
rect 22189 24191 22247 24197
rect 22189 24188 22201 24191
rect 21508 24160 22201 24188
rect 21508 24148 21514 24160
rect 22189 24157 22201 24160
rect 22235 24157 22247 24191
rect 22189 24151 22247 24157
rect 22281 24191 22339 24197
rect 22281 24157 22293 24191
rect 22327 24157 22339 24191
rect 22281 24151 22339 24157
rect 7098 24120 7104 24132
rect 7059 24092 7104 24120
rect 7098 24080 7104 24092
rect 7156 24080 7162 24132
rect 10778 24080 10784 24132
rect 10836 24120 10842 24132
rect 17402 24120 17408 24132
rect 10836 24092 17408 24120
rect 10836 24080 10842 24092
rect 17402 24080 17408 24092
rect 17460 24080 17466 24132
rect 21634 24120 21640 24132
rect 21595 24092 21640 24120
rect 21634 24080 21640 24092
rect 21692 24120 21698 24132
rect 22296 24120 22324 24151
rect 23566 24148 23572 24200
rect 23624 24188 23630 24200
rect 23753 24191 23811 24197
rect 23753 24188 23765 24191
rect 23624 24160 23765 24188
rect 23624 24148 23630 24160
rect 23753 24157 23765 24160
rect 23799 24157 23811 24191
rect 23753 24151 23811 24157
rect 23845 24191 23903 24197
rect 23845 24157 23857 24191
rect 23891 24188 23903 24191
rect 25409 24191 25467 24197
rect 25409 24188 25421 24191
rect 23891 24160 25421 24188
rect 23891 24157 23903 24160
rect 23845 24151 23903 24157
rect 25409 24157 25421 24160
rect 25455 24188 25467 24191
rect 25774 24188 25780 24200
rect 25455 24160 25780 24188
rect 25455 24157 25467 24160
rect 25409 24151 25467 24157
rect 21692 24092 22324 24120
rect 21692 24080 21698 24092
rect 23198 24080 23204 24132
rect 23256 24120 23262 24132
rect 23860 24120 23888 24151
rect 25774 24148 25780 24160
rect 25832 24148 25838 24200
rect 23256 24092 23888 24120
rect 23256 24080 23262 24092
rect 5994 24052 6000 24064
rect 5736 24024 6000 24052
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 8294 24012 8300 24064
rect 8352 24052 8358 24064
rect 8389 24055 8447 24061
rect 8389 24052 8401 24055
rect 8352 24024 8401 24052
rect 8352 24012 8358 24024
rect 8389 24021 8401 24024
rect 8435 24021 8447 24055
rect 9122 24052 9128 24064
rect 9083 24024 9128 24052
rect 8389 24015 8447 24021
rect 9122 24012 9128 24024
rect 9180 24012 9186 24064
rect 12250 24052 12256 24064
rect 12211 24024 12256 24052
rect 12250 24012 12256 24024
rect 12308 24012 12314 24064
rect 12986 24012 12992 24064
rect 13044 24052 13050 24064
rect 13265 24055 13323 24061
rect 13265 24052 13277 24055
rect 13044 24024 13277 24052
rect 13044 24012 13050 24024
rect 13265 24021 13277 24024
rect 13311 24021 13323 24055
rect 13265 24015 13323 24021
rect 14458 24012 14464 24064
rect 14516 24052 14522 24064
rect 14645 24055 14703 24061
rect 14645 24052 14657 24055
rect 14516 24024 14657 24052
rect 14516 24012 14522 24024
rect 14645 24021 14657 24024
rect 14691 24021 14703 24055
rect 14645 24015 14703 24021
rect 14734 24012 14740 24064
rect 14792 24052 14798 24064
rect 15013 24055 15071 24061
rect 15013 24052 15025 24055
rect 14792 24024 15025 24052
rect 14792 24012 14798 24024
rect 15013 24021 15025 24024
rect 15059 24021 15071 24055
rect 15013 24015 15071 24021
rect 15749 24055 15807 24061
rect 15749 24021 15761 24055
rect 15795 24052 15807 24055
rect 16482 24052 16488 24064
rect 15795 24024 16488 24052
rect 15795 24021 15807 24024
rect 15749 24015 15807 24021
rect 16482 24012 16488 24024
rect 16540 24012 16546 24064
rect 17310 24052 17316 24064
rect 17271 24024 17316 24052
rect 17310 24012 17316 24024
rect 17368 24012 17374 24064
rect 19058 24052 19064 24064
rect 19019 24024 19064 24052
rect 19058 24012 19064 24024
rect 19116 24012 19122 24064
rect 20530 24052 20536 24064
rect 20491 24024 20536 24052
rect 20530 24012 20536 24024
rect 20588 24012 20594 24064
rect 21726 24052 21732 24064
rect 21687 24024 21732 24052
rect 21726 24012 21732 24024
rect 21784 24012 21790 24064
rect 23293 24055 23351 24061
rect 23293 24021 23305 24055
rect 23339 24052 23351 24055
rect 23842 24052 23848 24064
rect 23339 24024 23848 24052
rect 23339 24021 23351 24024
rect 23293 24015 23351 24021
rect 23842 24012 23848 24024
rect 23900 24012 23906 24064
rect 24854 24052 24860 24064
rect 24815 24024 24860 24052
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23848 1639 23851
rect 1762 23848 1768 23860
rect 1627 23820 1768 23848
rect 1627 23817 1639 23820
rect 1581 23811 1639 23817
rect 1762 23808 1768 23820
rect 1820 23808 1826 23860
rect 1946 23848 1952 23860
rect 1907 23820 1952 23848
rect 1946 23808 1952 23820
rect 2004 23808 2010 23860
rect 8110 23848 8116 23860
rect 2884 23820 8116 23848
rect 2884 23721 2912 23820
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 9306 23848 9312 23860
rect 9267 23820 9312 23848
rect 9306 23808 9312 23820
rect 9364 23808 9370 23860
rect 11790 23848 11796 23860
rect 11751 23820 11796 23848
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 12621 23851 12679 23857
rect 12621 23848 12633 23851
rect 11900 23820 12633 23848
rect 5350 23780 5356 23792
rect 5311 23752 5356 23780
rect 5350 23740 5356 23752
rect 5408 23740 5414 23792
rect 8018 23740 8024 23792
rect 8076 23780 8082 23792
rect 8478 23780 8484 23792
rect 8076 23752 8484 23780
rect 8076 23740 8082 23752
rect 8478 23740 8484 23752
rect 8536 23780 8542 23792
rect 9122 23780 9128 23792
rect 8536 23752 9128 23780
rect 8536 23740 8542 23752
rect 9122 23740 9128 23752
rect 9180 23780 9186 23792
rect 9493 23783 9551 23789
rect 9493 23780 9505 23783
rect 9180 23752 9505 23780
rect 9180 23740 9186 23752
rect 9493 23749 9505 23752
rect 9539 23780 9551 23783
rect 9585 23783 9643 23789
rect 9585 23780 9597 23783
rect 9539 23752 9597 23780
rect 9539 23749 9551 23752
rect 9493 23743 9551 23749
rect 9585 23749 9597 23752
rect 9631 23749 9643 23783
rect 9585 23743 9643 23749
rect 11514 23740 11520 23792
rect 11572 23780 11578 23792
rect 11900 23780 11928 23820
rect 12621 23817 12633 23820
rect 12667 23848 12679 23851
rect 12710 23848 12716 23860
rect 12667 23820 12716 23848
rect 12667 23817 12679 23820
rect 12621 23811 12679 23817
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 13998 23808 14004 23860
rect 14056 23848 14062 23860
rect 14369 23851 14427 23857
rect 14369 23848 14381 23851
rect 14056 23820 14381 23848
rect 14056 23808 14062 23820
rect 14369 23817 14381 23820
rect 14415 23817 14427 23851
rect 14369 23811 14427 23817
rect 14550 23808 14556 23860
rect 14608 23848 14614 23860
rect 14921 23851 14979 23857
rect 14921 23848 14933 23851
rect 14608 23820 14933 23848
rect 14608 23808 14614 23820
rect 14921 23817 14933 23820
rect 14967 23848 14979 23851
rect 16206 23848 16212 23860
rect 14967 23820 16212 23848
rect 14967 23817 14979 23820
rect 14921 23811 14979 23817
rect 16206 23808 16212 23820
rect 16264 23808 16270 23860
rect 16390 23808 16396 23860
rect 16448 23848 16454 23860
rect 16574 23848 16580 23860
rect 16448 23820 16580 23848
rect 16448 23808 16454 23820
rect 16574 23808 16580 23820
rect 16632 23848 16638 23860
rect 16853 23851 16911 23857
rect 16853 23848 16865 23851
rect 16632 23820 16865 23848
rect 16632 23808 16638 23820
rect 16853 23817 16865 23820
rect 16899 23817 16911 23851
rect 17402 23848 17408 23860
rect 17363 23820 17408 23848
rect 16853 23811 16911 23817
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 17586 23808 17592 23860
rect 17644 23848 17650 23860
rect 17773 23851 17831 23857
rect 17773 23848 17785 23851
rect 17644 23820 17785 23848
rect 17644 23808 17650 23820
rect 17773 23817 17785 23820
rect 17819 23817 17831 23851
rect 17773 23811 17831 23817
rect 19058 23808 19064 23860
rect 19116 23848 19122 23860
rect 20073 23851 20131 23857
rect 20073 23848 20085 23851
rect 19116 23820 20085 23848
rect 19116 23808 19122 23820
rect 20073 23817 20085 23820
rect 20119 23817 20131 23851
rect 20073 23811 20131 23817
rect 22462 23808 22468 23860
rect 22520 23848 22526 23860
rect 23661 23851 23719 23857
rect 23661 23848 23673 23851
rect 22520 23820 23673 23848
rect 22520 23808 22526 23820
rect 23661 23817 23673 23820
rect 23707 23817 23719 23851
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 23661 23811 23719 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25406 23848 25412 23860
rect 25367 23820 25412 23848
rect 25406 23808 25412 23820
rect 25464 23808 25470 23860
rect 25774 23848 25780 23860
rect 25735 23820 25780 23848
rect 25774 23808 25780 23820
rect 25832 23808 25838 23860
rect 11572 23752 11928 23780
rect 11572 23740 11578 23752
rect 12066 23740 12072 23792
rect 12124 23780 12130 23792
rect 12161 23783 12219 23789
rect 12161 23780 12173 23783
rect 12124 23752 12173 23780
rect 12124 23740 12130 23752
rect 12161 23749 12173 23752
rect 12207 23749 12219 23783
rect 12161 23743 12219 23749
rect 18325 23783 18383 23789
rect 18325 23749 18337 23783
rect 18371 23780 18383 23783
rect 19334 23780 19340 23792
rect 18371 23752 19340 23780
rect 18371 23749 18383 23752
rect 18325 23743 18383 23749
rect 19334 23740 19340 23752
rect 19392 23740 19398 23792
rect 19797 23783 19855 23789
rect 19797 23749 19809 23783
rect 19843 23780 19855 23783
rect 19978 23780 19984 23792
rect 19843 23752 19984 23780
rect 19843 23749 19855 23752
rect 19797 23743 19855 23749
rect 19978 23740 19984 23752
rect 20036 23780 20042 23792
rect 20438 23780 20444 23792
rect 20036 23752 20444 23780
rect 20036 23740 20042 23752
rect 20438 23740 20444 23752
rect 20496 23740 20502 23792
rect 2317 23715 2375 23721
rect 2317 23681 2329 23715
rect 2363 23712 2375 23715
rect 2869 23715 2927 23721
rect 2869 23712 2881 23715
rect 2363 23684 2881 23712
rect 2363 23681 2375 23684
rect 2317 23675 2375 23681
rect 2869 23681 2881 23684
rect 2915 23681 2927 23715
rect 2869 23675 2927 23681
rect 3053 23715 3111 23721
rect 3053 23681 3065 23715
rect 3099 23712 3111 23715
rect 3234 23712 3240 23724
rect 3099 23684 3240 23712
rect 3099 23681 3111 23684
rect 3053 23675 3111 23681
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 3970 23712 3976 23724
rect 3931 23684 3976 23712
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 6362 23712 6368 23724
rect 6275 23684 6368 23712
rect 6362 23672 6368 23684
rect 6420 23712 6426 23724
rect 8754 23712 8760 23724
rect 6420 23684 8760 23712
rect 6420 23672 6426 23684
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 8849 23715 8907 23721
rect 8849 23681 8861 23715
rect 8895 23712 8907 23715
rect 12986 23712 12992 23724
rect 8895 23684 9904 23712
rect 8895 23681 8907 23684
rect 8849 23675 8907 23681
rect 9876 23656 9904 23684
rect 11532 23684 12992 23712
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 2130 23644 2136 23656
rect 1443 23616 2136 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2130 23604 2136 23616
rect 2188 23604 2194 23656
rect 2498 23604 2504 23656
rect 2556 23604 2562 23656
rect 2774 23604 2780 23656
rect 2832 23644 2838 23656
rect 3418 23644 3424 23656
rect 2832 23616 3424 23644
rect 2832 23604 2838 23616
rect 3418 23604 3424 23616
rect 3476 23644 3482 23656
rect 3789 23647 3847 23653
rect 3789 23644 3801 23647
rect 3476 23616 3801 23644
rect 3476 23604 3482 23616
rect 3789 23613 3801 23616
rect 3835 23613 3847 23647
rect 3789 23607 3847 23613
rect 3878 23604 3884 23656
rect 3936 23644 3942 23656
rect 4229 23647 4287 23653
rect 4229 23644 4241 23647
rect 3936 23616 4241 23644
rect 3936 23604 3942 23616
rect 4229 23613 4241 23616
rect 4275 23613 4287 23647
rect 4229 23607 4287 23613
rect 6825 23647 6883 23653
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 8573 23647 8631 23653
rect 6871 23616 7144 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 2516 23576 2544 23604
rect 3513 23579 3571 23585
rect 3513 23576 3525 23579
rect 2516 23548 3525 23576
rect 3513 23545 3525 23548
rect 3559 23576 3571 23579
rect 4522 23576 4528 23588
rect 3559 23548 4528 23576
rect 3559 23545 3571 23548
rect 3513 23539 3571 23545
rect 4522 23536 4528 23548
rect 4580 23536 4586 23588
rect 7116 23520 7144 23616
rect 8573 23613 8585 23647
rect 8619 23644 8631 23647
rect 9306 23644 9312 23656
rect 8619 23616 9312 23644
rect 8619 23613 8631 23616
rect 8573 23607 8631 23613
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 9769 23647 9827 23653
rect 9769 23613 9781 23647
rect 9815 23613 9827 23647
rect 9769 23607 9827 23613
rect 8110 23576 8116 23588
rect 8071 23548 8116 23576
rect 8110 23536 8116 23548
rect 8168 23536 8174 23588
rect 9493 23579 9551 23585
rect 9493 23545 9505 23579
rect 9539 23576 9551 23579
rect 9784 23576 9812 23607
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 10025 23647 10083 23653
rect 10025 23644 10037 23647
rect 9916 23616 10037 23644
rect 9916 23604 9922 23616
rect 10025 23613 10037 23616
rect 10071 23613 10083 23647
rect 10025 23607 10083 23613
rect 11532 23588 11560 23684
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 18230 23672 18236 23724
rect 18288 23712 18294 23724
rect 18785 23715 18843 23721
rect 18785 23712 18797 23715
rect 18288 23684 18797 23712
rect 18288 23672 18294 23684
rect 18785 23681 18797 23684
rect 18831 23681 18843 23715
rect 18966 23712 18972 23724
rect 18927 23684 18972 23712
rect 18785 23675 18843 23681
rect 18966 23672 18972 23684
rect 19024 23672 19030 23724
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23712 20407 23715
rect 24118 23712 24124 23724
rect 20395 23684 21036 23712
rect 24079 23684 24124 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 21008 23656 21036 23684
rect 24118 23672 24124 23684
rect 24176 23672 24182 23724
rect 24302 23712 24308 23724
rect 24263 23684 24308 23712
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 15378 23604 15384 23656
rect 15436 23644 15442 23656
rect 15746 23653 15752 23656
rect 15473 23647 15531 23653
rect 15473 23644 15485 23647
rect 15436 23616 15485 23644
rect 15436 23604 15442 23616
rect 15473 23613 15485 23616
rect 15519 23613 15531 23647
rect 15740 23644 15752 23653
rect 15707 23616 15752 23644
rect 15473 23607 15531 23613
rect 15740 23607 15752 23616
rect 15746 23604 15752 23607
rect 15804 23604 15810 23656
rect 18046 23604 18052 23656
rect 18104 23644 18110 23656
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18104 23616 18705 23644
rect 18104 23604 18110 23616
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 18693 23607 18751 23613
rect 19889 23647 19947 23653
rect 19889 23613 19901 23647
rect 19935 23644 19947 23647
rect 20254 23644 20260 23656
rect 19935 23616 20260 23644
rect 19935 23613 19947 23616
rect 19889 23607 19947 23613
rect 20254 23604 20260 23616
rect 20312 23604 20318 23656
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23613 20959 23647
rect 20901 23607 20959 23613
rect 11514 23576 11520 23588
rect 9539 23548 11520 23576
rect 9539 23545 9551 23548
rect 9493 23539 9551 23545
rect 11514 23536 11520 23548
rect 11572 23536 11578 23588
rect 13256 23579 13314 23585
rect 13256 23545 13268 23579
rect 13302 23576 13314 23579
rect 13538 23576 13544 23588
rect 13302 23548 13544 23576
rect 13302 23545 13314 23548
rect 13256 23539 13314 23545
rect 13538 23536 13544 23548
rect 13596 23536 13602 23588
rect 2409 23511 2467 23517
rect 2409 23477 2421 23511
rect 2455 23508 2467 23511
rect 2774 23508 2780 23520
rect 2455 23480 2780 23508
rect 2455 23477 2467 23480
rect 2409 23471 2467 23477
rect 2774 23468 2780 23480
rect 2832 23468 2838 23520
rect 3050 23468 3056 23520
rect 3108 23508 3114 23520
rect 4798 23508 4804 23520
rect 3108 23480 4804 23508
rect 3108 23468 3114 23480
rect 4798 23468 4804 23480
rect 4856 23468 4862 23520
rect 5994 23508 6000 23520
rect 5907 23480 6000 23508
rect 5994 23468 6000 23480
rect 6052 23508 6058 23520
rect 6178 23508 6184 23520
rect 6052 23480 6184 23508
rect 6052 23468 6058 23480
rect 6178 23468 6184 23480
rect 6236 23468 6242 23520
rect 7006 23508 7012 23520
rect 6967 23480 7012 23508
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 7098 23468 7104 23520
rect 7156 23508 7162 23520
rect 7377 23511 7435 23517
rect 7377 23508 7389 23511
rect 7156 23480 7389 23508
rect 7156 23468 7162 23480
rect 7377 23477 7389 23480
rect 7423 23477 7435 23511
rect 8202 23508 8208 23520
rect 8163 23480 8208 23508
rect 7377 23471 7435 23477
rect 8202 23468 8208 23480
rect 8260 23468 8266 23520
rect 8662 23508 8668 23520
rect 8623 23480 8668 23508
rect 8662 23468 8668 23480
rect 8720 23468 8726 23520
rect 11146 23508 11152 23520
rect 11059 23480 11152 23508
rect 11146 23468 11152 23480
rect 11204 23508 11210 23520
rect 11882 23508 11888 23520
rect 11204 23480 11888 23508
rect 11204 23468 11210 23480
rect 11882 23468 11888 23480
rect 11940 23468 11946 23520
rect 14918 23468 14924 23520
rect 14976 23508 14982 23520
rect 15289 23511 15347 23517
rect 15289 23508 15301 23511
rect 14976 23480 15301 23508
rect 14976 23468 14982 23480
rect 15289 23477 15301 23480
rect 15335 23508 15347 23511
rect 16114 23508 16120 23520
rect 15335 23480 16120 23508
rect 15335 23477 15347 23480
rect 15289 23471 15347 23477
rect 16114 23468 16120 23480
rect 16172 23468 16178 23520
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 20916 23508 20944 23607
rect 20990 23604 20996 23656
rect 21048 23644 21054 23656
rect 21168 23647 21226 23653
rect 21168 23644 21180 23647
rect 21048 23616 21180 23644
rect 21048 23604 21054 23616
rect 21168 23613 21180 23616
rect 21214 23644 21226 23647
rect 24026 23644 24032 23656
rect 21214 23616 23704 23644
rect 23987 23616 24032 23644
rect 21214 23613 21226 23616
rect 21168 23607 21226 23613
rect 23017 23579 23075 23585
rect 23017 23545 23029 23579
rect 23063 23576 23075 23579
rect 23566 23576 23572 23588
rect 23063 23548 23572 23576
rect 23063 23545 23075 23548
rect 23017 23539 23075 23545
rect 23566 23536 23572 23548
rect 23624 23536 23630 23588
rect 23676 23576 23704 23616
rect 24026 23604 24032 23616
rect 24084 23604 24090 23656
rect 25225 23647 25283 23653
rect 25225 23613 25237 23647
rect 25271 23644 25283 23647
rect 25590 23644 25596 23656
rect 25271 23616 25596 23644
rect 25271 23613 25283 23616
rect 25225 23607 25283 23613
rect 25590 23604 25596 23616
rect 25648 23604 25654 23656
rect 24302 23576 24308 23588
rect 23676 23548 24308 23576
rect 24302 23536 24308 23548
rect 24360 23536 24366 23588
rect 21542 23508 21548 23520
rect 20855 23480 21548 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 21634 23468 21640 23520
rect 21692 23508 21698 23520
rect 22281 23511 22339 23517
rect 22281 23508 22293 23511
rect 21692 23480 22293 23508
rect 21692 23468 21698 23480
rect 22281 23477 22293 23480
rect 22327 23477 22339 23511
rect 23290 23508 23296 23520
rect 23251 23480 23296 23508
rect 22281 23471 22339 23477
rect 23290 23468 23296 23480
rect 23348 23468 23354 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2869 23307 2927 23313
rect 2869 23273 2881 23307
rect 2915 23304 2927 23307
rect 3602 23304 3608 23316
rect 2915 23276 3608 23304
rect 2915 23273 2927 23276
rect 2869 23267 2927 23273
rect 3602 23264 3608 23276
rect 3660 23264 3666 23316
rect 4341 23307 4399 23313
rect 4341 23273 4353 23307
rect 4387 23304 4399 23307
rect 4614 23304 4620 23316
rect 4387 23276 4620 23304
rect 4387 23273 4399 23276
rect 4341 23267 4399 23273
rect 1302 23196 1308 23248
rect 1360 23236 1366 23248
rect 4356 23236 4384 23267
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 4706 23264 4712 23316
rect 4764 23304 4770 23316
rect 6273 23307 6331 23313
rect 4764 23276 4809 23304
rect 4764 23264 4770 23276
rect 6273 23273 6285 23307
rect 6319 23304 6331 23307
rect 6822 23304 6828 23316
rect 6319 23276 6828 23304
rect 6319 23273 6331 23276
rect 6273 23267 6331 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 7561 23307 7619 23313
rect 7561 23273 7573 23307
rect 7607 23304 7619 23307
rect 8202 23304 8208 23316
rect 7607 23276 8208 23304
rect 7607 23273 7619 23276
rect 7561 23267 7619 23273
rect 8202 23264 8208 23276
rect 8260 23304 8266 23316
rect 8389 23307 8447 23313
rect 8389 23304 8401 23307
rect 8260 23276 8401 23304
rect 8260 23264 8266 23276
rect 8389 23273 8401 23276
rect 8435 23273 8447 23307
rect 8389 23267 8447 23273
rect 8481 23307 8539 23313
rect 8481 23273 8493 23307
rect 8527 23304 8539 23307
rect 8570 23304 8576 23316
rect 8527 23276 8576 23304
rect 8527 23273 8539 23276
rect 8481 23267 8539 23273
rect 8570 23264 8576 23276
rect 8628 23304 8634 23316
rect 9677 23307 9735 23313
rect 9677 23304 9689 23307
rect 8628 23276 9689 23304
rect 8628 23264 8634 23276
rect 9677 23273 9689 23276
rect 9723 23273 9735 23307
rect 9677 23267 9735 23273
rect 10781 23307 10839 23313
rect 10781 23273 10793 23307
rect 10827 23304 10839 23307
rect 10870 23304 10876 23316
rect 10827 23276 10876 23304
rect 10827 23273 10839 23276
rect 10781 23267 10839 23273
rect 10870 23264 10876 23276
rect 10928 23264 10934 23316
rect 11054 23304 11060 23316
rect 11015 23276 11060 23304
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 12897 23307 12955 23313
rect 12897 23273 12909 23307
rect 12943 23304 12955 23307
rect 13170 23304 13176 23316
rect 12943 23276 13176 23304
rect 12943 23273 12955 23276
rect 12897 23267 12955 23273
rect 13170 23264 13176 23276
rect 13228 23264 13234 23316
rect 18230 23264 18236 23316
rect 18288 23304 18294 23316
rect 18325 23307 18383 23313
rect 18325 23304 18337 23307
rect 18288 23276 18337 23304
rect 18288 23264 18294 23276
rect 18325 23273 18337 23276
rect 18371 23273 18383 23307
rect 18325 23267 18383 23273
rect 18785 23307 18843 23313
rect 18785 23273 18797 23307
rect 18831 23304 18843 23307
rect 18966 23304 18972 23316
rect 18831 23276 18972 23304
rect 18831 23273 18843 23276
rect 18785 23267 18843 23273
rect 18966 23264 18972 23276
rect 19024 23264 19030 23316
rect 19334 23264 19340 23316
rect 19392 23304 19398 23316
rect 19705 23307 19763 23313
rect 19705 23304 19717 23307
rect 19392 23276 19717 23304
rect 19392 23264 19398 23276
rect 19705 23273 19717 23276
rect 19751 23273 19763 23307
rect 21450 23304 21456 23316
rect 21411 23276 21456 23304
rect 19705 23267 19763 23273
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 22922 23304 22928 23316
rect 22883 23276 22928 23304
rect 22922 23264 22928 23276
rect 22980 23264 22986 23316
rect 23658 23264 23664 23316
rect 23716 23304 23722 23316
rect 24397 23307 24455 23313
rect 24397 23304 24409 23307
rect 23716 23276 24409 23304
rect 23716 23264 23722 23276
rect 24397 23273 24409 23276
rect 24443 23273 24455 23307
rect 24397 23267 24455 23273
rect 24489 23307 24547 23313
rect 24489 23273 24501 23307
rect 24535 23304 24547 23307
rect 24854 23304 24860 23316
rect 24535 23276 24860 23304
rect 24535 23273 24547 23276
rect 24489 23267 24547 23273
rect 1360 23208 4384 23236
rect 4433 23239 4491 23245
rect 1360 23196 1366 23208
rect 4433 23205 4445 23239
rect 4479 23236 4491 23239
rect 4724 23236 4752 23264
rect 4479 23208 4752 23236
rect 4479 23205 4491 23208
rect 4433 23199 4491 23205
rect 7742 23196 7748 23248
rect 7800 23236 7806 23248
rect 7837 23239 7895 23245
rect 7837 23236 7849 23239
rect 7800 23208 7849 23236
rect 7800 23196 7806 23208
rect 7837 23205 7849 23208
rect 7883 23205 7895 23239
rect 7837 23199 7895 23205
rect 8938 23196 8944 23248
rect 8996 23236 9002 23248
rect 11790 23245 11796 23248
rect 9401 23239 9459 23245
rect 9401 23236 9413 23239
rect 8996 23208 9413 23236
rect 8996 23196 9002 23208
rect 9401 23205 9413 23208
rect 9447 23236 9459 23239
rect 10137 23239 10195 23245
rect 10137 23236 10149 23239
rect 9447 23208 10149 23236
rect 9447 23205 9459 23208
rect 9401 23199 9459 23205
rect 10137 23205 10149 23208
rect 10183 23205 10195 23239
rect 11784 23236 11796 23245
rect 11751 23208 11796 23236
rect 10137 23199 10195 23205
rect 11784 23199 11796 23208
rect 11790 23196 11796 23199
rect 11848 23196 11854 23248
rect 16206 23196 16212 23248
rect 16264 23236 16270 23248
rect 16390 23245 16396 23248
rect 16384 23236 16396 23245
rect 16264 23208 16396 23236
rect 16264 23196 16270 23208
rect 16384 23199 16396 23208
rect 16390 23196 16396 23199
rect 16448 23196 16454 23248
rect 19613 23239 19671 23245
rect 19613 23205 19625 23239
rect 19659 23236 19671 23239
rect 19978 23236 19984 23248
rect 19659 23208 19984 23236
rect 19659 23205 19671 23208
rect 19613 23199 19671 23205
rect 19978 23196 19984 23208
rect 20036 23196 20042 23248
rect 21634 23196 21640 23248
rect 21692 23236 21698 23248
rect 21790 23239 21848 23245
rect 21790 23236 21802 23239
rect 21692 23208 21802 23236
rect 21692 23196 21698 23208
rect 21790 23205 21802 23208
rect 21836 23205 21848 23239
rect 24412 23236 24440 23267
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 25133 23307 25191 23313
rect 25133 23273 25145 23307
rect 25179 23304 25191 23307
rect 25314 23304 25320 23316
rect 25179 23276 25320 23304
rect 25179 23273 25191 23276
rect 25133 23267 25191 23273
rect 25314 23264 25320 23276
rect 25372 23304 25378 23316
rect 25682 23304 25688 23316
rect 25372 23276 25688 23304
rect 25372 23264 25378 23276
rect 25682 23264 25688 23276
rect 25740 23264 25746 23316
rect 24762 23236 24768 23248
rect 24412 23208 24768 23236
rect 21790 23199 21848 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2774 23168 2780 23180
rect 1443 23140 2780 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2774 23128 2780 23140
rect 2832 23168 2838 23180
rect 2832 23140 2877 23168
rect 2832 23128 2838 23140
rect 3234 23128 3240 23180
rect 3292 23168 3298 23180
rect 3421 23171 3479 23177
rect 3421 23168 3433 23171
rect 3292 23140 3433 23168
rect 3292 23128 3298 23140
rect 3421 23137 3433 23140
rect 3467 23137 3479 23171
rect 3421 23131 3479 23137
rect 3878 23128 3884 23180
rect 3936 23128 3942 23180
rect 3970 23128 3976 23180
rect 4028 23168 4034 23180
rect 5166 23177 5172 23180
rect 4028 23140 4844 23168
rect 4028 23128 4034 23140
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23069 3111 23103
rect 3053 23063 3111 23069
rect 1946 23032 1952 23044
rect 1907 23004 1952 23032
rect 1946 22992 1952 23004
rect 2004 22992 2010 23044
rect 3068 23032 3096 23063
rect 3234 23032 3240 23044
rect 3068 23004 3240 23032
rect 3234 22992 3240 23004
rect 3292 22992 3298 23044
rect 3896 22976 3924 23128
rect 4816 23112 4844 23140
rect 5160 23131 5172 23177
rect 5224 23168 5230 23180
rect 10042 23168 10048 23180
rect 5224 23140 5260 23168
rect 10003 23140 10048 23168
rect 5166 23128 5172 23131
rect 5224 23128 5230 23140
rect 10042 23128 10048 23140
rect 10100 23128 10106 23180
rect 11330 23128 11336 23180
rect 11388 23168 11394 23180
rect 11514 23168 11520 23180
rect 11388 23140 11520 23168
rect 11388 23128 11394 23140
rect 11514 23128 11520 23140
rect 11572 23128 11578 23180
rect 13906 23128 13912 23180
rect 13964 23168 13970 23180
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 13964 23140 14105 23168
rect 13964 23128 13970 23140
rect 14093 23137 14105 23140
rect 14139 23137 14151 23171
rect 14093 23131 14151 23137
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 4433 23103 4491 23109
rect 4433 23100 4445 23103
rect 4212 23072 4445 23100
rect 4212 23060 4218 23072
rect 4433 23069 4445 23072
rect 4479 23069 4491 23103
rect 4433 23063 4491 23069
rect 4798 23060 4804 23112
rect 4856 23100 4862 23112
rect 4893 23103 4951 23109
rect 4893 23100 4905 23103
rect 4856 23072 4905 23100
rect 4856 23060 4862 23072
rect 4893 23069 4905 23072
rect 4939 23069 4951 23103
rect 8662 23100 8668 23112
rect 8623 23072 8668 23100
rect 4893 23063 4951 23069
rect 8662 23060 8668 23072
rect 8720 23060 8726 23112
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 15102 23100 15108 23112
rect 15063 23072 15108 23100
rect 10229 23063 10287 23069
rect 6638 22992 6644 23044
rect 6696 23032 6702 23044
rect 8021 23035 8079 23041
rect 8021 23032 8033 23035
rect 6696 23004 8033 23032
rect 6696 22992 6702 23004
rect 8021 23001 8033 23004
rect 8067 23001 8079 23035
rect 8021 22995 8079 23001
rect 9125 23035 9183 23041
rect 9125 23001 9137 23035
rect 9171 23032 9183 23035
rect 9490 23032 9496 23044
rect 9171 23004 9496 23032
rect 9171 23001 9183 23004
rect 9125 22995 9183 23001
rect 9490 22992 9496 23004
rect 9548 23032 9554 23044
rect 9858 23032 9864 23044
rect 9548 23004 9864 23032
rect 9548 22992 9554 23004
rect 9858 22992 9864 23004
rect 9916 23032 9922 23044
rect 10244 23032 10272 23063
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 16117 23103 16175 23109
rect 16117 23100 16129 23103
rect 15488 23072 16129 23100
rect 9916 23004 10272 23032
rect 9916 22992 9922 23004
rect 2314 22964 2320 22976
rect 2275 22936 2320 22964
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 2409 22967 2467 22973
rect 2409 22933 2421 22967
rect 2455 22964 2467 22967
rect 2498 22964 2504 22976
rect 2455 22936 2504 22964
rect 2455 22933 2467 22936
rect 2409 22927 2467 22933
rect 2498 22924 2504 22936
rect 2556 22924 2562 22976
rect 3786 22964 3792 22976
rect 3747 22936 3792 22964
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 3878 22924 3884 22976
rect 3936 22924 3942 22976
rect 6914 22964 6920 22976
rect 6875 22936 6920 22964
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 13538 22964 13544 22976
rect 13499 22936 13544 22964
rect 13538 22924 13544 22936
rect 13596 22924 13602 22976
rect 14274 22964 14280 22976
rect 14235 22936 14280 22964
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 15378 22924 15384 22976
rect 15436 22964 15442 22976
rect 15488 22973 15516 23072
rect 16117 23069 16129 23072
rect 16163 23069 16175 23103
rect 16117 23063 16175 23069
rect 19153 23103 19211 23109
rect 19153 23069 19165 23103
rect 19199 23100 19211 23103
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 19199 23072 19901 23100
rect 19199 23069 19211 23072
rect 19153 23063 19211 23069
rect 19889 23069 19901 23072
rect 19935 23100 19947 23103
rect 20990 23100 20996 23112
rect 19935 23072 20996 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20990 23060 20996 23072
rect 21048 23060 21054 23112
rect 21542 23100 21548 23112
rect 21503 23072 21548 23100
rect 21542 23060 21548 23072
rect 21600 23060 21606 23112
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 24627 23072 24661 23100
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 17494 23032 17500 23044
rect 17455 23004 17500 23032
rect 17494 22992 17500 23004
rect 17552 22992 17558 23044
rect 19245 23035 19303 23041
rect 19245 23001 19257 23035
rect 19291 23032 19303 23035
rect 21450 23032 21456 23044
rect 19291 23004 21456 23032
rect 19291 23001 19303 23004
rect 19245 22995 19303 23001
rect 21450 22992 21456 23004
rect 21508 22992 21514 23044
rect 23937 23035 23995 23041
rect 23937 23001 23949 23035
rect 23983 23032 23995 23035
rect 24302 23032 24308 23044
rect 23983 23004 24308 23032
rect 23983 23001 23995 23004
rect 23937 22995 23995 23001
rect 24302 22992 24308 23004
rect 24360 23032 24366 23044
rect 24596 23032 24624 23063
rect 24670 23032 24676 23044
rect 24360 23004 24676 23032
rect 24360 22992 24366 23004
rect 24670 22992 24676 23004
rect 24728 22992 24734 23044
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 15436 22936 15485 22964
rect 15436 22924 15442 22936
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 15473 22927 15531 22933
rect 15933 22967 15991 22973
rect 15933 22933 15945 22967
rect 15979 22964 15991 22967
rect 16298 22964 16304 22976
rect 15979 22936 16304 22964
rect 15979 22933 15991 22936
rect 15933 22927 15991 22933
rect 16298 22924 16304 22936
rect 16356 22964 16362 22976
rect 17512 22964 17540 22992
rect 20254 22964 20260 22976
rect 16356 22936 17540 22964
rect 20215 22936 20260 22964
rect 16356 22924 16362 22936
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 23198 22924 23204 22976
rect 23256 22964 23262 22976
rect 23477 22967 23535 22973
rect 23477 22964 23489 22967
rect 23256 22936 23489 22964
rect 23256 22924 23262 22936
rect 23477 22933 23489 22936
rect 23523 22933 23535 22967
rect 23477 22927 23535 22933
rect 24029 22967 24087 22973
rect 24029 22933 24041 22967
rect 24075 22964 24087 22967
rect 24118 22964 24124 22976
rect 24075 22936 24124 22964
rect 24075 22933 24087 22936
rect 24029 22927 24087 22933
rect 24118 22924 24124 22936
rect 24176 22924 24182 22976
rect 25501 22967 25559 22973
rect 25501 22933 25513 22967
rect 25547 22964 25559 22967
rect 25590 22964 25596 22976
rect 25547 22936 25596 22964
rect 25547 22933 25559 22936
rect 25501 22927 25559 22933
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2774 22720 2780 22772
rect 2832 22760 2838 22772
rect 3145 22763 3203 22769
rect 3145 22760 3157 22763
rect 2832 22732 3157 22760
rect 2832 22720 2838 22732
rect 3145 22729 3157 22732
rect 3191 22729 3203 22763
rect 3145 22723 3203 22729
rect 3329 22763 3387 22769
rect 3329 22729 3341 22763
rect 3375 22760 3387 22763
rect 3510 22760 3516 22772
rect 3375 22732 3516 22760
rect 3375 22729 3387 22732
rect 3329 22723 3387 22729
rect 3510 22720 3516 22732
rect 3568 22720 3574 22772
rect 4430 22760 4436 22772
rect 4391 22732 4436 22760
rect 4430 22720 4436 22732
rect 4488 22720 4494 22772
rect 6454 22720 6460 22772
rect 6512 22760 6518 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 6512 22732 6561 22760
rect 6512 22720 6518 22732
rect 6549 22729 6561 22732
rect 6595 22729 6607 22763
rect 6549 22723 6607 22729
rect 7929 22763 7987 22769
rect 7929 22729 7941 22763
rect 7975 22760 7987 22763
rect 8662 22760 8668 22772
rect 7975 22732 8668 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 1765 22695 1823 22701
rect 1765 22661 1777 22695
rect 1811 22692 1823 22695
rect 2869 22695 2927 22701
rect 1811 22664 2728 22692
rect 1811 22661 1823 22664
rect 1765 22655 1823 22661
rect 2314 22584 2320 22636
rect 2372 22624 2378 22636
rect 2409 22627 2467 22633
rect 2409 22624 2421 22627
rect 2372 22596 2421 22624
rect 2372 22584 2378 22596
rect 2409 22593 2421 22596
rect 2455 22624 2467 22627
rect 2498 22624 2504 22636
rect 2455 22596 2504 22624
rect 2455 22593 2467 22596
rect 2409 22587 2467 22593
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 1762 22516 1768 22568
rect 1820 22516 1826 22568
rect 1946 22516 1952 22568
rect 2004 22556 2010 22568
rect 2225 22559 2283 22565
rect 2225 22556 2237 22559
rect 2004 22528 2237 22556
rect 2004 22516 2010 22528
rect 2225 22525 2237 22528
rect 2271 22525 2283 22559
rect 2225 22519 2283 22525
rect 1673 22491 1731 22497
rect 1673 22457 1685 22491
rect 1719 22488 1731 22491
rect 1780 22488 1808 22516
rect 2133 22491 2191 22497
rect 2133 22488 2145 22491
rect 1719 22460 2145 22488
rect 1719 22457 1731 22460
rect 1673 22451 1731 22457
rect 2133 22457 2145 22460
rect 2179 22457 2191 22491
rect 2700 22488 2728 22664
rect 2869 22661 2881 22695
rect 2915 22692 2927 22695
rect 3602 22692 3608 22704
rect 2915 22664 3608 22692
rect 2915 22661 2927 22664
rect 2869 22655 2927 22661
rect 3602 22652 3608 22664
rect 3660 22652 3666 22704
rect 4893 22695 4951 22701
rect 4893 22692 4905 22695
rect 3712 22664 4905 22692
rect 2774 22584 2780 22636
rect 2832 22624 2838 22636
rect 2958 22624 2964 22636
rect 2832 22596 2964 22624
rect 2832 22584 2838 22596
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 3712 22565 3740 22664
rect 4893 22661 4905 22664
rect 4939 22692 4951 22695
rect 4982 22692 4988 22704
rect 4939 22664 4988 22692
rect 4939 22661 4951 22664
rect 4893 22655 4951 22661
rect 4982 22652 4988 22664
rect 5040 22652 5046 22704
rect 5905 22695 5963 22701
rect 5905 22692 5917 22695
rect 5368 22664 5917 22692
rect 5368 22636 5396 22664
rect 5905 22661 5917 22664
rect 5951 22661 5963 22695
rect 5905 22655 5963 22661
rect 3878 22624 3884 22636
rect 3839 22596 3884 22624
rect 3878 22584 3884 22596
rect 3936 22584 3942 22636
rect 5350 22624 5356 22636
rect 5311 22596 5356 22624
rect 5350 22584 5356 22596
rect 5408 22584 5414 22636
rect 5445 22627 5503 22633
rect 5445 22593 5457 22627
rect 5491 22593 5503 22627
rect 5445 22587 5503 22593
rect 3697 22559 3755 22565
rect 3697 22525 3709 22559
rect 3743 22525 3755 22559
rect 3697 22519 3755 22525
rect 3789 22559 3847 22565
rect 3789 22525 3801 22559
rect 3835 22556 3847 22559
rect 4062 22556 4068 22568
rect 3835 22528 4068 22556
rect 3835 22525 3847 22528
rect 3789 22519 3847 22525
rect 4062 22516 4068 22528
rect 4120 22516 4126 22568
rect 5074 22556 5080 22568
rect 4356 22528 5080 22556
rect 4356 22488 4384 22528
rect 5074 22516 5080 22528
rect 5132 22516 5138 22568
rect 5258 22556 5264 22568
rect 5219 22528 5264 22556
rect 5258 22516 5264 22528
rect 5316 22516 5322 22568
rect 2700 22460 4384 22488
rect 2133 22451 2191 22457
rect 4430 22448 4436 22500
rect 4488 22488 4494 22500
rect 5460 22488 5488 22587
rect 6564 22556 6592 22723
rect 8662 22720 8668 22732
rect 8720 22720 8726 22772
rect 8754 22720 8760 22772
rect 8812 22760 8818 22772
rect 9401 22763 9459 22769
rect 9401 22760 9413 22763
rect 8812 22732 9413 22760
rect 8812 22720 8818 22732
rect 9401 22729 9413 22732
rect 9447 22729 9459 22763
rect 9401 22723 9459 22729
rect 11330 22720 11336 22772
rect 11388 22760 11394 22772
rect 11517 22763 11575 22769
rect 11517 22760 11529 22763
rect 11388 22732 11529 22760
rect 11388 22720 11394 22732
rect 11517 22729 11529 22732
rect 11563 22729 11575 22763
rect 11517 22723 11575 22729
rect 11790 22720 11796 22772
rect 11848 22760 11854 22772
rect 11885 22763 11943 22769
rect 11885 22760 11897 22763
rect 11848 22732 11897 22760
rect 11848 22720 11854 22732
rect 11885 22729 11897 22732
rect 11931 22729 11943 22763
rect 11885 22723 11943 22729
rect 13081 22763 13139 22769
rect 13081 22729 13093 22763
rect 13127 22760 13139 22763
rect 14642 22760 14648 22772
rect 13127 22732 14648 22760
rect 13127 22729 13139 22732
rect 13081 22723 13139 22729
rect 14642 22720 14648 22732
rect 14700 22720 14706 22772
rect 16390 22760 16396 22772
rect 16351 22732 16396 22760
rect 16390 22720 16396 22732
rect 16448 22720 16454 22772
rect 18966 22720 18972 22772
rect 19024 22760 19030 22772
rect 19061 22763 19119 22769
rect 19061 22760 19073 22763
rect 19024 22732 19073 22760
rect 19024 22720 19030 22732
rect 19061 22729 19073 22732
rect 19107 22760 19119 22763
rect 19794 22760 19800 22772
rect 19107 22732 19800 22760
rect 19107 22729 19119 22732
rect 19061 22723 19119 22729
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 20990 22760 20996 22772
rect 20951 22732 20996 22760
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 22649 22763 22707 22769
rect 22649 22729 22661 22763
rect 22695 22760 22707 22763
rect 22738 22760 22744 22772
rect 22695 22732 22744 22760
rect 22695 22729 22707 22732
rect 22649 22723 22707 22729
rect 22738 22720 22744 22732
rect 22796 22720 22802 22772
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 25041 22763 25099 22769
rect 25041 22760 25053 22763
rect 24912 22732 25053 22760
rect 24912 22720 24918 22732
rect 25041 22729 25053 22732
rect 25087 22729 25099 22763
rect 25041 22723 25099 22729
rect 25409 22763 25467 22769
rect 25409 22729 25421 22763
rect 25455 22760 25467 22763
rect 26142 22760 26148 22772
rect 25455 22732 26148 22760
rect 25455 22729 25467 22732
rect 25409 22723 25467 22729
rect 26142 22720 26148 22732
rect 26200 22720 26206 22772
rect 10042 22652 10048 22704
rect 10100 22692 10106 22704
rect 10505 22695 10563 22701
rect 10505 22692 10517 22695
rect 10100 22664 10517 22692
rect 10100 22652 10106 22664
rect 10505 22661 10517 22664
rect 10551 22661 10563 22695
rect 10505 22655 10563 22661
rect 15194 22652 15200 22704
rect 15252 22692 15258 22704
rect 15289 22695 15347 22701
rect 15289 22692 15301 22695
rect 15252 22664 15301 22692
rect 15252 22652 15258 22664
rect 15289 22661 15301 22664
rect 15335 22661 15347 22695
rect 15289 22655 15347 22661
rect 16022 22652 16028 22704
rect 16080 22692 16086 22704
rect 16482 22692 16488 22704
rect 16080 22664 16488 22692
rect 16080 22652 16086 22664
rect 16482 22652 16488 22664
rect 16540 22652 16546 22704
rect 22186 22652 22192 22704
rect 22244 22692 22250 22704
rect 23661 22695 23719 22701
rect 23661 22692 23673 22695
rect 22244 22664 23673 22692
rect 22244 22652 22250 22664
rect 23661 22661 23673 22664
rect 23707 22661 23719 22695
rect 23661 22655 23719 22661
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22624 7619 22627
rect 8018 22624 8024 22636
rect 7607 22596 8024 22624
rect 7607 22593 7619 22596
rect 7561 22587 7619 22593
rect 8018 22584 8024 22596
rect 8076 22584 8082 22636
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10962 22624 10968 22636
rect 9999 22596 10968 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 11057 22627 11115 22633
rect 11057 22593 11069 22627
rect 11103 22593 11115 22627
rect 11057 22587 11115 22593
rect 6825 22559 6883 22565
rect 6825 22556 6837 22559
rect 6564 22528 6837 22556
rect 6825 22525 6837 22528
rect 6871 22525 6883 22559
rect 6825 22519 6883 22525
rect 9766 22516 9772 22568
rect 9824 22556 9830 22568
rect 11072 22556 11100 22587
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16945 22627 17003 22633
rect 16945 22624 16957 22627
rect 16632 22596 16957 22624
rect 16632 22584 16638 22596
rect 16945 22593 16957 22596
rect 16991 22593 17003 22627
rect 16945 22587 17003 22593
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22624 17739 22627
rect 18601 22627 18659 22633
rect 18601 22624 18613 22627
rect 17727 22596 18613 22624
rect 17727 22593 17739 22596
rect 17681 22587 17739 22593
rect 18601 22593 18613 22596
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 21634 22584 21640 22636
rect 21692 22624 21698 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21692 22596 22017 22624
rect 21692 22584 21698 22596
rect 22005 22593 22017 22596
rect 22051 22624 22063 22627
rect 23477 22627 23535 22633
rect 23477 22624 23489 22627
rect 22051 22596 23489 22624
rect 22051 22593 22063 22596
rect 22005 22587 22063 22593
rect 23477 22593 23489 22596
rect 23523 22624 23535 22627
rect 24213 22627 24271 22633
rect 24213 22624 24225 22627
rect 23523 22596 24225 22624
rect 23523 22593 23535 22596
rect 23477 22587 23535 22593
rect 24213 22593 24225 22596
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 9824 22528 11100 22556
rect 12897 22559 12955 22565
rect 9824 22516 9830 22528
rect 10980 22500 11008 22528
rect 12897 22525 12909 22559
rect 12943 22556 12955 22559
rect 13909 22559 13967 22565
rect 13909 22556 13921 22559
rect 12943 22528 13492 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 4488 22460 5488 22488
rect 4488 22448 4494 22460
rect 8110 22448 8116 22500
rect 8168 22488 8174 22500
rect 8266 22491 8324 22497
rect 8266 22488 8278 22491
rect 8168 22460 8278 22488
rect 8168 22448 8174 22460
rect 8266 22457 8278 22460
rect 8312 22457 8324 22491
rect 10778 22488 10784 22500
rect 8266 22451 8324 22457
rect 9784 22460 10784 22488
rect 9784 22432 9812 22460
rect 10778 22448 10784 22460
rect 10836 22448 10842 22500
rect 10962 22448 10968 22500
rect 11020 22448 11026 22500
rect 13464 22432 13492 22528
rect 13740 22528 13921 22556
rect 1302 22380 1308 22432
rect 1360 22420 1366 22432
rect 1854 22420 1860 22432
rect 1360 22392 1860 22420
rect 1360 22380 1366 22392
rect 1854 22380 1860 22392
rect 1912 22380 1918 22432
rect 3786 22380 3792 22432
rect 3844 22420 3850 22432
rect 4798 22420 4804 22432
rect 3844 22392 4804 22420
rect 3844 22380 3850 22392
rect 4798 22380 4804 22392
rect 4856 22420 4862 22432
rect 6178 22420 6184 22432
rect 4856 22392 6184 22420
rect 4856 22380 4862 22392
rect 6178 22380 6184 22392
rect 6236 22380 6242 22432
rect 7006 22420 7012 22432
rect 6967 22392 7012 22420
rect 7006 22380 7012 22392
rect 7064 22380 7070 22432
rect 9766 22380 9772 22432
rect 9824 22380 9830 22432
rect 9858 22380 9864 22432
rect 9916 22420 9922 22432
rect 10321 22423 10379 22429
rect 10321 22420 10333 22423
rect 9916 22392 10333 22420
rect 9916 22380 9922 22392
rect 10321 22389 10333 22392
rect 10367 22420 10379 22423
rect 10873 22423 10931 22429
rect 10873 22420 10885 22423
rect 10367 22392 10885 22420
rect 10367 22389 10379 22392
rect 10321 22383 10379 22389
rect 10873 22389 10885 22392
rect 10919 22389 10931 22423
rect 10873 22383 10931 22389
rect 12342 22380 12348 22432
rect 12400 22420 12406 22432
rect 12710 22420 12716 22432
rect 12400 22392 12716 22420
rect 12400 22380 12406 22392
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 13446 22420 13452 22432
rect 13407 22392 13452 22420
rect 13446 22380 13452 22392
rect 13504 22380 13510 22432
rect 13538 22380 13544 22432
rect 13596 22420 13602 22432
rect 13740 22429 13768 22528
rect 13909 22525 13921 22528
rect 13955 22556 13967 22559
rect 15378 22556 15384 22568
rect 13955 22528 15384 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 15378 22516 15384 22528
rect 15436 22556 15442 22568
rect 16117 22559 16175 22565
rect 16117 22556 16129 22559
rect 15436 22528 16129 22556
rect 15436 22516 15442 22528
rect 16117 22525 16129 22528
rect 16163 22525 16175 22559
rect 16117 22519 16175 22525
rect 16390 22516 16396 22568
rect 16448 22556 16454 22568
rect 16853 22559 16911 22565
rect 16853 22556 16865 22559
rect 16448 22528 16865 22556
rect 16448 22516 16454 22528
rect 16853 22525 16865 22528
rect 16899 22525 16911 22559
rect 16853 22519 16911 22525
rect 17770 22516 17776 22568
rect 17828 22556 17834 22568
rect 18414 22556 18420 22568
rect 17828 22528 18420 22556
rect 17828 22516 17834 22528
rect 18414 22516 18420 22528
rect 18472 22516 18478 22568
rect 19613 22559 19671 22565
rect 19613 22556 19625 22559
rect 19444 22528 19625 22556
rect 13814 22448 13820 22500
rect 13872 22488 13878 22500
rect 14154 22491 14212 22497
rect 14154 22488 14166 22491
rect 13872 22460 14166 22488
rect 13872 22448 13878 22460
rect 14154 22457 14166 22460
rect 14200 22488 14212 22491
rect 16758 22488 16764 22500
rect 14200 22460 16620 22488
rect 16719 22460 16764 22488
rect 14200 22457 14212 22460
rect 14154 22451 14212 22457
rect 13725 22423 13783 22429
rect 13725 22420 13737 22423
rect 13596 22392 13737 22420
rect 13596 22380 13602 22392
rect 13725 22389 13737 22392
rect 13771 22389 13783 22423
rect 16592 22420 16620 22460
rect 16758 22448 16764 22460
rect 16816 22448 16822 22500
rect 17497 22491 17555 22497
rect 17497 22457 17509 22491
rect 17543 22488 17555 22491
rect 17543 22460 18552 22488
rect 17543 22457 17555 22460
rect 17497 22451 17555 22457
rect 17681 22423 17739 22429
rect 17681 22420 17693 22423
rect 16592 22392 17693 22420
rect 13725 22383 13783 22389
rect 17681 22389 17693 22392
rect 17727 22420 17739 22423
rect 17773 22423 17831 22429
rect 17773 22420 17785 22423
rect 17727 22392 17785 22420
rect 17727 22389 17739 22392
rect 17681 22383 17739 22389
rect 17773 22389 17785 22392
rect 17819 22389 17831 22423
rect 18046 22420 18052 22432
rect 18007 22392 18052 22420
rect 17773 22383 17831 22389
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 18524 22429 18552 22460
rect 18509 22423 18567 22429
rect 18509 22389 18521 22423
rect 18555 22420 18567 22423
rect 18874 22420 18880 22432
rect 18555 22392 18880 22420
rect 18555 22389 18567 22392
rect 18509 22383 18567 22389
rect 18874 22380 18880 22392
rect 18932 22380 18938 22432
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19444 22429 19472 22528
rect 19613 22525 19625 22528
rect 19659 22556 19671 22559
rect 21542 22556 21548 22568
rect 19659 22528 21548 22556
rect 19659 22525 19671 22528
rect 19613 22519 19671 22525
rect 21542 22516 21548 22528
rect 21600 22516 21606 22568
rect 22465 22559 22523 22565
rect 22465 22556 22477 22559
rect 22296 22528 22477 22556
rect 19794 22448 19800 22500
rect 19852 22497 19858 22500
rect 19852 22491 19916 22497
rect 19852 22457 19870 22491
rect 19904 22457 19916 22491
rect 19852 22451 19916 22457
rect 19852 22448 19858 22451
rect 22296 22432 22324 22528
rect 22465 22525 22477 22528
rect 22511 22525 22523 22559
rect 24118 22556 24124 22568
rect 24079 22528 24124 22556
rect 22465 22519 22523 22525
rect 24118 22516 24124 22528
rect 24176 22516 24182 22568
rect 25222 22556 25228 22568
rect 25183 22528 25228 22556
rect 25222 22516 25228 22528
rect 25280 22556 25286 22568
rect 25777 22559 25835 22565
rect 25777 22556 25789 22559
rect 25280 22528 25789 22556
rect 25280 22516 25286 22528
rect 25777 22525 25789 22528
rect 25823 22525 25835 22559
rect 25777 22519 25835 22525
rect 24029 22491 24087 22497
rect 24029 22488 24041 22491
rect 23124 22460 24041 22488
rect 23124 22432 23152 22460
rect 24029 22457 24041 22460
rect 24075 22457 24087 22491
rect 24029 22451 24087 22457
rect 19429 22423 19487 22429
rect 19429 22420 19441 22423
rect 19392 22392 19441 22420
rect 19392 22380 19398 22392
rect 19429 22389 19441 22392
rect 19475 22389 19487 22423
rect 22278 22420 22284 22432
rect 22239 22392 22284 22420
rect 19429 22383 19487 22389
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 23106 22420 23112 22432
rect 23067 22392 23112 22420
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 24670 22420 24676 22432
rect 24631 22392 24676 22420
rect 24670 22380 24676 22392
rect 24728 22380 24734 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1670 22176 1676 22228
rect 1728 22216 1734 22228
rect 1949 22219 2007 22225
rect 1949 22216 1961 22219
rect 1728 22188 1961 22216
rect 1728 22176 1734 22188
rect 1949 22185 1961 22188
rect 1995 22185 2007 22219
rect 1949 22179 2007 22185
rect 2498 22176 2504 22228
rect 2556 22216 2562 22228
rect 3053 22219 3111 22225
rect 3053 22216 3065 22219
rect 2556 22188 3065 22216
rect 2556 22176 2562 22188
rect 3053 22185 3065 22188
rect 3099 22216 3111 22219
rect 3234 22216 3240 22228
rect 3099 22188 3240 22216
rect 3099 22185 3111 22188
rect 3053 22179 3111 22185
rect 3234 22176 3240 22188
rect 3292 22176 3298 22228
rect 3421 22219 3479 22225
rect 3421 22185 3433 22219
rect 3467 22216 3479 22219
rect 3878 22216 3884 22228
rect 3467 22188 3884 22216
rect 3467 22185 3479 22188
rect 3421 22179 3479 22185
rect 3878 22176 3884 22188
rect 3936 22176 3942 22228
rect 5166 22216 5172 22228
rect 5127 22188 5172 22216
rect 5166 22176 5172 22188
rect 5224 22176 5230 22228
rect 5258 22176 5264 22228
rect 5316 22216 5322 22228
rect 5445 22219 5503 22225
rect 5445 22216 5457 22219
rect 5316 22188 5457 22216
rect 5316 22176 5322 22188
rect 5445 22185 5457 22188
rect 5491 22185 5503 22219
rect 8570 22216 8576 22228
rect 8531 22188 8576 22216
rect 5445 22179 5503 22185
rect 8570 22176 8576 22188
rect 8628 22176 8634 22228
rect 9490 22216 9496 22228
rect 9451 22188 9496 22216
rect 9490 22176 9496 22188
rect 9548 22176 9554 22228
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10134 22216 10140 22228
rect 10008 22188 10140 22216
rect 10008 22176 10014 22188
rect 10134 22176 10140 22188
rect 10192 22216 10198 22228
rect 10321 22219 10379 22225
rect 10321 22216 10333 22219
rect 10192 22188 10333 22216
rect 10192 22176 10198 22188
rect 10321 22185 10333 22188
rect 10367 22185 10379 22219
rect 10962 22216 10968 22228
rect 10923 22188 10968 22216
rect 10321 22179 10379 22185
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 16206 22216 16212 22228
rect 16167 22188 16212 22216
rect 16206 22176 16212 22188
rect 16264 22176 16270 22228
rect 16758 22216 16764 22228
rect 16719 22188 16764 22216
rect 16758 22176 16764 22188
rect 16816 22176 16822 22228
rect 22186 22216 22192 22228
rect 22147 22188 22192 22216
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 23385 22219 23443 22225
rect 23385 22216 23397 22219
rect 23164 22188 23397 22216
rect 23164 22176 23170 22188
rect 23385 22185 23397 22188
rect 23431 22185 23443 22219
rect 24118 22216 24124 22228
rect 23385 22179 23443 22185
rect 23584 22188 24124 22216
rect 4430 22148 4436 22160
rect 4391 22120 4436 22148
rect 4430 22108 4436 22120
rect 4488 22108 4494 22160
rect 5994 22108 6000 22160
rect 6052 22148 6058 22160
rect 6448 22151 6506 22157
rect 6448 22148 6460 22151
rect 6052 22120 6460 22148
rect 6052 22108 6058 22120
rect 6448 22117 6460 22120
rect 6494 22148 6506 22151
rect 6822 22148 6828 22160
rect 6494 22120 6828 22148
rect 6494 22117 6506 22120
rect 6448 22111 6506 22117
rect 6822 22108 6828 22120
rect 6880 22108 6886 22160
rect 9125 22151 9183 22157
rect 9125 22117 9137 22151
rect 9171 22148 9183 22151
rect 10042 22148 10048 22160
rect 9171 22120 10048 22148
rect 9171 22117 9183 22120
rect 9125 22111 9183 22117
rect 10042 22108 10048 22120
rect 10100 22108 10106 22160
rect 10229 22151 10287 22157
rect 10229 22117 10241 22151
rect 10275 22148 10287 22151
rect 10594 22148 10600 22160
rect 10275 22120 10600 22148
rect 10275 22117 10287 22120
rect 10229 22111 10287 22117
rect 10594 22108 10600 22120
rect 10652 22108 10658 22160
rect 11692 22151 11750 22157
rect 11692 22117 11704 22151
rect 11738 22148 11750 22151
rect 12250 22148 12256 22160
rect 11738 22120 12256 22148
rect 11738 22117 11750 22120
rect 11692 22111 11750 22117
rect 12250 22108 12256 22120
rect 12308 22148 12314 22160
rect 13170 22148 13176 22160
rect 12308 22120 13176 22148
rect 12308 22108 12314 22120
rect 13170 22108 13176 22120
rect 13228 22108 13234 22160
rect 16666 22108 16672 22160
rect 16724 22148 16730 22160
rect 17129 22151 17187 22157
rect 17129 22148 17141 22151
rect 16724 22120 17141 22148
rect 16724 22108 16730 22120
rect 17129 22117 17141 22120
rect 17175 22117 17187 22151
rect 17129 22111 17187 22117
rect 1854 22040 1860 22092
rect 1912 22080 1918 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1912 22052 2053 22080
rect 1912 22040 1918 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3418 22040 3424 22092
rect 3476 22080 3482 22092
rect 3786 22080 3792 22092
rect 3476 22052 3792 22080
rect 3476 22040 3482 22052
rect 3786 22040 3792 22052
rect 3844 22040 3850 22092
rect 5905 22083 5963 22089
rect 5905 22049 5917 22083
rect 5951 22080 5963 22083
rect 6086 22080 6092 22092
rect 5951 22052 6092 22080
rect 5951 22049 5963 22052
rect 5905 22043 5963 22049
rect 6086 22040 6092 22052
rect 6144 22040 6150 22092
rect 11330 22080 11336 22092
rect 11291 22052 11336 22080
rect 11330 22040 11336 22052
rect 11388 22040 11394 22092
rect 14093 22083 14151 22089
rect 14093 22049 14105 22083
rect 14139 22080 14151 22083
rect 14550 22080 14556 22092
rect 14139 22052 14556 22080
rect 14139 22049 14151 22052
rect 14093 22043 14151 22049
rect 14550 22040 14556 22052
rect 14608 22040 14614 22092
rect 15562 22040 15568 22092
rect 15620 22080 15626 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 15620 22052 15669 22080
rect 15620 22040 15626 22052
rect 15657 22049 15669 22052
rect 15703 22049 15715 22083
rect 17770 22080 17776 22092
rect 17731 22052 17776 22080
rect 15657 22043 15715 22049
rect 17770 22040 17776 22052
rect 17828 22040 17834 22092
rect 17862 22040 17868 22092
rect 17920 22080 17926 22092
rect 18581 22083 18639 22089
rect 18581 22080 18593 22083
rect 17920 22052 18593 22080
rect 17920 22040 17926 22052
rect 18581 22049 18593 22052
rect 18627 22049 18639 22083
rect 18581 22043 18639 22049
rect 23293 22083 23351 22089
rect 23293 22049 23305 22083
rect 23339 22080 23351 22083
rect 23584 22080 23612 22188
rect 24118 22176 24124 22188
rect 24176 22176 24182 22228
rect 24762 22216 24768 22228
rect 24723 22188 24768 22216
rect 24762 22176 24768 22188
rect 24820 22176 24826 22228
rect 23842 22148 23848 22160
rect 23803 22120 23848 22148
rect 23842 22108 23848 22120
rect 23900 22108 23906 22160
rect 24670 22148 24676 22160
rect 24136 22120 24676 22148
rect 23339 22052 23612 22080
rect 23753 22083 23811 22089
rect 23339 22049 23351 22052
rect 23293 22043 23351 22049
rect 23753 22049 23765 22083
rect 23799 22049 23811 22083
rect 23753 22043 23811 22049
rect 1946 21972 1952 22024
rect 2004 22012 2010 22024
rect 2133 22015 2191 22021
rect 2133 22012 2145 22015
rect 2004 21984 2145 22012
rect 2004 21972 2010 21984
rect 2133 21981 2145 21984
rect 2179 21981 2191 22015
rect 2133 21975 2191 21981
rect 2222 21972 2228 22024
rect 2280 21972 2286 22024
rect 4522 22012 4528 22024
rect 4483 21984 4528 22012
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 22012 4767 22015
rect 5166 22012 5172 22024
rect 4755 21984 5172 22012
rect 4755 21981 4767 21984
rect 4709 21975 4767 21981
rect 5166 21972 5172 21984
rect 5224 21972 5230 22024
rect 6178 22012 6184 22024
rect 6139 21984 6184 22012
rect 6178 21972 6184 21984
rect 6236 21972 6242 22024
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 9030 22012 9036 22024
rect 8444 21984 9036 22012
rect 8444 21972 8450 21984
rect 9030 21972 9036 21984
rect 9088 21972 9094 22024
rect 10502 22012 10508 22024
rect 10463 21984 10508 22012
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 11146 21972 11152 22024
rect 11204 22012 11210 22024
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 11204 21984 11437 22012
rect 11204 21972 11210 21984
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 13906 21972 13912 22024
rect 13964 22012 13970 22024
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 13964 21984 14657 22012
rect 13964 21972 13970 21984
rect 14645 21981 14657 21984
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 15470 21972 15476 22024
rect 15528 22012 15534 22024
rect 15746 22012 15752 22024
rect 15528 21984 15752 22012
rect 15528 21972 15534 21984
rect 15746 21972 15752 21984
rect 15804 21972 15810 22024
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 17184 21984 17233 22012
rect 17184 21972 17190 21984
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 22012 17463 22015
rect 17586 22012 17592 22024
rect 17451 21984 17592 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 17586 21972 17592 21984
rect 17644 21972 17650 22024
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 18325 22015 18383 22021
rect 18325 22012 18337 22015
rect 18104 21984 18337 22012
rect 18104 21972 18110 21984
rect 18325 21981 18337 21984
rect 18371 21981 18383 22015
rect 18325 21975 18383 21981
rect 21726 21972 21732 22024
rect 21784 22012 21790 22024
rect 22002 22012 22008 22024
rect 21784 21984 22008 22012
rect 21784 21972 21790 21984
rect 22002 21972 22008 21984
rect 22060 22012 22066 22024
rect 22281 22015 22339 22021
rect 22281 22012 22293 22015
rect 22060 21984 22293 22012
rect 22060 21972 22066 21984
rect 22281 21981 22293 21984
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 22465 22015 22523 22021
rect 22465 21981 22477 22015
rect 22511 22012 22523 22015
rect 22554 22012 22560 22024
rect 22511 21984 22560 22012
rect 22511 21981 22523 21984
rect 22465 21975 22523 21981
rect 22554 21972 22560 21984
rect 22612 22012 22618 22024
rect 22922 22012 22928 22024
rect 22612 21984 22928 22012
rect 22612 21972 22618 21984
rect 22922 21972 22928 21984
rect 22980 21972 22986 22024
rect 23474 21972 23480 22024
rect 23532 22012 23538 22024
rect 23768 22012 23796 22043
rect 23532 21984 23796 22012
rect 24029 22015 24087 22021
rect 23532 21972 23538 21984
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 24136 22012 24164 22120
rect 24670 22108 24676 22120
rect 24728 22108 24734 22160
rect 24210 22040 24216 22092
rect 24268 22080 24274 22092
rect 24854 22080 24860 22092
rect 24268 22052 24860 22080
rect 24268 22040 24274 22052
rect 24854 22040 24860 22052
rect 24912 22040 24918 22092
rect 24949 22083 25007 22089
rect 24949 22049 24961 22083
rect 24995 22080 25007 22083
rect 25222 22080 25228 22092
rect 24995 22052 25228 22080
rect 24995 22049 25007 22052
rect 24949 22043 25007 22049
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 24075 21984 24164 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 1394 21904 1400 21956
rect 1452 21944 1458 21956
rect 2240 21944 2268 21972
rect 1452 21916 2268 21944
rect 1452 21904 1458 21916
rect 3418 21904 3424 21956
rect 3476 21944 3482 21956
rect 4065 21947 4123 21953
rect 4065 21944 4077 21947
rect 3476 21916 4077 21944
rect 3476 21904 3482 21916
rect 4065 21913 4077 21916
rect 4111 21913 4123 21947
rect 4065 21907 4123 21913
rect 12434 21904 12440 21956
rect 12492 21944 12498 21956
rect 13357 21947 13415 21953
rect 13357 21944 13369 21947
rect 12492 21916 13369 21944
rect 12492 21904 12498 21916
rect 13357 21913 13369 21916
rect 13403 21913 13415 21947
rect 13357 21907 13415 21913
rect 14277 21947 14335 21953
rect 14277 21913 14289 21947
rect 14323 21944 14335 21947
rect 14366 21944 14372 21956
rect 14323 21916 14372 21944
rect 14323 21913 14335 21916
rect 14277 21907 14335 21913
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 15105 21947 15163 21953
rect 15105 21913 15117 21947
rect 15151 21944 15163 21947
rect 15378 21944 15384 21956
rect 15151 21916 15384 21944
rect 15151 21913 15163 21916
rect 15105 21907 15163 21913
rect 15378 21904 15384 21916
rect 15436 21904 15442 21956
rect 15838 21944 15844 21956
rect 15799 21916 15844 21944
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 19702 21944 19708 21956
rect 19663 21916 19708 21944
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 21542 21944 21548 21956
rect 21503 21916 21548 21944
rect 21542 21904 21548 21916
rect 21600 21904 21606 21956
rect 25133 21947 25191 21953
rect 25133 21913 25145 21947
rect 25179 21944 25191 21947
rect 25866 21944 25872 21956
rect 25179 21916 25872 21944
rect 25179 21913 25191 21916
rect 25133 21907 25191 21913
rect 25866 21904 25872 21916
rect 25924 21904 25930 21956
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 2222 21876 2228 21888
rect 1627 21848 2228 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 2222 21836 2228 21848
rect 2280 21836 2286 21888
rect 2498 21836 2504 21888
rect 2556 21876 2562 21888
rect 2593 21879 2651 21885
rect 2593 21876 2605 21879
rect 2556 21848 2605 21876
rect 2556 21836 2562 21848
rect 2593 21845 2605 21848
rect 2639 21845 2651 21879
rect 2593 21839 2651 21845
rect 3602 21836 3608 21888
rect 3660 21876 3666 21888
rect 3697 21879 3755 21885
rect 3697 21876 3709 21879
rect 3660 21848 3709 21876
rect 3660 21836 3666 21848
rect 3697 21845 3709 21848
rect 3743 21845 3755 21879
rect 7558 21876 7564 21888
rect 7519 21848 7564 21876
rect 3697 21839 3755 21845
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 8110 21876 8116 21888
rect 8071 21848 8116 21876
rect 8110 21836 8116 21848
rect 8168 21836 8174 21888
rect 9861 21879 9919 21885
rect 9861 21845 9873 21879
rect 9907 21876 9919 21879
rect 10870 21876 10876 21888
rect 9907 21848 10876 21876
rect 9907 21845 9919 21848
rect 9861 21839 9919 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 12526 21876 12532 21888
rect 12216 21848 12532 21876
rect 12216 21836 12222 21848
rect 12526 21836 12532 21848
rect 12584 21876 12590 21888
rect 12805 21879 12863 21885
rect 12805 21876 12817 21879
rect 12584 21848 12817 21876
rect 12584 21836 12590 21848
rect 12805 21845 12817 21848
rect 12851 21845 12863 21879
rect 12805 21839 12863 21845
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 13909 21879 13967 21885
rect 13909 21876 13921 21879
rect 13872 21848 13921 21876
rect 13872 21836 13878 21848
rect 13909 21845 13921 21848
rect 13955 21845 13967 21879
rect 15470 21876 15476 21888
rect 15431 21848 15476 21876
rect 13909 21839 13967 21845
rect 15470 21836 15476 21848
rect 15528 21836 15534 21888
rect 16574 21836 16580 21888
rect 16632 21876 16638 21888
rect 16669 21879 16727 21885
rect 16669 21876 16681 21879
rect 16632 21848 16681 21876
rect 16632 21836 16638 21848
rect 16669 21845 16681 21848
rect 16715 21876 16727 21879
rect 17770 21876 17776 21888
rect 16715 21848 17776 21876
rect 16715 21845 16727 21848
rect 16669 21839 16727 21845
rect 17770 21836 17776 21848
rect 17828 21836 17834 21888
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21876 18291 21879
rect 18690 21876 18696 21888
rect 18279 21848 18696 21876
rect 18279 21845 18291 21848
rect 18233 21839 18291 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 19518 21836 19524 21888
rect 19576 21876 19582 21888
rect 20257 21879 20315 21885
rect 20257 21876 20269 21879
rect 19576 21848 20269 21876
rect 19576 21836 19582 21848
rect 20257 21845 20269 21848
rect 20303 21845 20315 21879
rect 20257 21839 20315 21845
rect 21174 21836 21180 21888
rect 21232 21876 21238 21888
rect 21821 21879 21879 21885
rect 21821 21876 21833 21879
rect 21232 21848 21833 21876
rect 21232 21836 21238 21848
rect 21821 21845 21833 21848
rect 21867 21845 21879 21879
rect 21821 21839 21879 21845
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 23934 21876 23940 21888
rect 23716 21848 23940 21876
rect 23716 21836 23722 21848
rect 23934 21836 23940 21848
rect 23992 21836 23998 21888
rect 24489 21879 24547 21885
rect 24489 21845 24501 21879
rect 24535 21876 24547 21879
rect 24762 21876 24768 21888
rect 24535 21848 24768 21876
rect 24535 21845 24547 21848
rect 24489 21839 24547 21845
rect 24762 21836 24768 21848
rect 24820 21836 24826 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1670 21632 1676 21684
rect 1728 21672 1734 21684
rect 2593 21675 2651 21681
rect 2593 21672 2605 21675
rect 1728 21644 2605 21672
rect 1728 21632 1734 21644
rect 2593 21641 2605 21644
rect 2639 21672 2651 21675
rect 2682 21672 2688 21684
rect 2639 21644 2688 21672
rect 2639 21641 2651 21644
rect 2593 21635 2651 21641
rect 2682 21632 2688 21644
rect 2740 21632 2746 21684
rect 4709 21675 4767 21681
rect 4709 21641 4721 21675
rect 4755 21672 4767 21675
rect 5166 21672 5172 21684
rect 4755 21644 5172 21672
rect 4755 21641 4767 21644
rect 4709 21635 4767 21641
rect 5166 21632 5172 21644
rect 5224 21672 5230 21684
rect 5261 21675 5319 21681
rect 5261 21672 5273 21675
rect 5224 21644 5273 21672
rect 5224 21632 5230 21644
rect 5261 21641 5273 21644
rect 5307 21641 5319 21675
rect 5261 21635 5319 21641
rect 5905 21675 5963 21681
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 5994 21672 6000 21684
rect 5951 21644 6000 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 5994 21632 6000 21644
rect 6052 21632 6058 21684
rect 8294 21672 8300 21684
rect 8255 21644 8300 21672
rect 8294 21632 8300 21644
rect 8352 21632 8358 21684
rect 10226 21672 10232 21684
rect 10187 21644 10232 21672
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 10594 21672 10600 21684
rect 10555 21644 10600 21672
rect 10594 21632 10600 21644
rect 10652 21632 10658 21684
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11793 21675 11851 21681
rect 11793 21672 11805 21675
rect 11204 21644 11805 21672
rect 11204 21632 11210 21644
rect 11793 21641 11805 21644
rect 11839 21641 11851 21675
rect 12250 21672 12256 21684
rect 12211 21644 12256 21672
rect 11793 21635 11851 21641
rect 1946 21564 1952 21616
rect 2004 21604 2010 21616
rect 11808 21604 11836 21635
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 13081 21675 13139 21681
rect 13081 21672 13093 21675
rect 12360 21644 13093 21672
rect 12158 21604 12164 21616
rect 2004 21576 2176 21604
rect 11808 21576 12164 21604
rect 2004 21564 2010 21576
rect 2038 21536 2044 21548
rect 1999 21508 2044 21536
rect 2038 21496 2044 21508
rect 2096 21496 2102 21548
rect 2148 21545 2176 21576
rect 12158 21564 12164 21576
rect 12216 21604 12222 21616
rect 12360 21604 12388 21644
rect 13081 21641 13093 21644
rect 13127 21672 13139 21675
rect 13538 21672 13544 21684
rect 13127 21644 13544 21672
rect 13127 21641 13139 21644
rect 13081 21635 13139 21641
rect 12216 21576 12388 21604
rect 12216 21564 12222 21576
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21505 2191 21539
rect 2133 21499 2191 21505
rect 6178 21496 6184 21548
rect 6236 21496 6242 21548
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21536 7527 21539
rect 7558 21536 7564 21548
rect 7515 21508 7564 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 7558 21496 7564 21508
rect 7616 21536 7622 21548
rect 7742 21536 7748 21548
rect 7616 21508 7748 21536
rect 7616 21496 7622 21508
rect 7742 21496 7748 21508
rect 7800 21536 7806 21548
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 7800 21508 7849 21536
rect 7800 21496 7806 21508
rect 7837 21505 7849 21508
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 9398 21496 9404 21548
rect 9456 21536 9462 21548
rect 9677 21539 9735 21545
rect 9677 21536 9689 21539
rect 9456 21508 9689 21536
rect 9456 21496 9462 21508
rect 9677 21505 9689 21508
rect 9723 21505 9735 21539
rect 9677 21499 9735 21505
rect 9861 21539 9919 21545
rect 9861 21505 9873 21539
rect 9907 21536 9919 21539
rect 9950 21536 9956 21548
rect 9907 21508 9956 21536
rect 9907 21505 9919 21508
rect 9861 21499 9919 21505
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 1949 21471 2007 21477
rect 1949 21468 1961 21471
rect 1452 21440 1961 21468
rect 1452 21428 1458 21440
rect 1949 21437 1961 21440
rect 1995 21468 2007 21471
rect 2498 21468 2504 21480
rect 1995 21440 2504 21468
rect 1995 21437 2007 21440
rect 1949 21431 2007 21437
rect 2498 21428 2504 21440
rect 2556 21428 2562 21480
rect 3329 21471 3387 21477
rect 3329 21437 3341 21471
rect 3375 21437 3387 21471
rect 3329 21431 3387 21437
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 1762 21332 1768 21344
rect 1627 21304 1768 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 1762 21292 1768 21304
rect 1820 21292 1826 21344
rect 3237 21335 3295 21341
rect 3237 21301 3249 21335
rect 3283 21332 3295 21335
rect 3344 21332 3372 21431
rect 3602 21409 3608 21412
rect 3596 21400 3608 21409
rect 3563 21372 3608 21400
rect 3596 21363 3608 21372
rect 3602 21360 3608 21363
rect 3660 21360 3666 21412
rect 3694 21332 3700 21344
rect 3283 21304 3700 21332
rect 3283 21301 3295 21304
rect 3237 21295 3295 21301
rect 3694 21292 3700 21304
rect 3752 21292 3758 21344
rect 6196 21332 6224 21496
rect 6641 21471 6699 21477
rect 6641 21437 6653 21471
rect 6687 21468 6699 21471
rect 7190 21468 7196 21480
rect 6687 21440 7196 21468
rect 6687 21437 6699 21440
rect 6641 21431 6699 21437
rect 7190 21428 7196 21440
rect 7248 21428 7254 21480
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 8757 21471 8815 21477
rect 7340 21440 7385 21468
rect 7340 21428 7346 21440
rect 8757 21437 8769 21471
rect 8803 21468 8815 21471
rect 9876 21468 9904 21499
rect 9950 21496 9956 21508
rect 10008 21536 10014 21548
rect 10502 21536 10508 21548
rect 10008 21508 10508 21536
rect 10008 21496 10014 21508
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 11330 21536 11336 21548
rect 11291 21508 11336 21536
rect 11330 21496 11336 21508
rect 11388 21496 11394 21548
rect 13280 21545 13308 21644
rect 13538 21632 13544 21644
rect 13596 21632 13602 21684
rect 15378 21632 15384 21684
rect 15436 21672 15442 21684
rect 16390 21672 16396 21684
rect 15436 21644 16396 21672
rect 15436 21632 15442 21644
rect 16390 21632 16396 21644
rect 16448 21632 16454 21684
rect 17862 21672 17868 21684
rect 17823 21644 17868 21672
rect 17862 21632 17868 21644
rect 17920 21632 17926 21684
rect 21450 21672 21456 21684
rect 21411 21644 21456 21672
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 22554 21672 22560 21684
rect 22515 21644 22560 21672
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 23474 21632 23480 21684
rect 23532 21672 23538 21684
rect 23934 21672 23940 21684
rect 23532 21644 23940 21672
rect 23532 21632 23538 21644
rect 23934 21632 23940 21644
rect 23992 21632 23998 21684
rect 24670 21632 24676 21684
rect 24728 21672 24734 21684
rect 24765 21675 24823 21681
rect 24765 21672 24777 21675
rect 24728 21644 24777 21672
rect 24728 21632 24734 21644
rect 24765 21641 24777 21644
rect 24811 21641 24823 21675
rect 25498 21672 25504 21684
rect 25459 21644 25504 21672
rect 24765 21635 24823 21641
rect 25498 21632 25504 21644
rect 25556 21632 25562 21684
rect 23753 21607 23811 21613
rect 23753 21573 23765 21607
rect 23799 21573 23811 21607
rect 23753 21567 23811 21573
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 15470 21496 15476 21548
rect 15528 21536 15534 21548
rect 15565 21539 15623 21545
rect 15565 21536 15577 21539
rect 15528 21508 15577 21536
rect 15528 21496 15534 21508
rect 15565 21505 15577 21508
rect 15611 21536 15623 21539
rect 17034 21536 17040 21548
rect 15611 21508 17040 21536
rect 15611 21505 15623 21508
rect 15565 21499 15623 21505
rect 17034 21496 17040 21508
rect 17092 21536 17098 21548
rect 17586 21536 17592 21548
rect 17092 21508 17592 21536
rect 17092 21496 17098 21508
rect 17586 21496 17592 21508
rect 17644 21496 17650 21548
rect 20898 21536 20904 21548
rect 20859 21508 20904 21536
rect 20898 21496 20904 21508
rect 20956 21536 20962 21548
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 20956 21508 22017 21536
rect 20956 21496 20962 21508
rect 22005 21505 22017 21508
rect 22051 21536 22063 21539
rect 22094 21536 22100 21548
rect 22051 21508 22100 21536
rect 22051 21505 22063 21508
rect 22005 21499 22063 21505
rect 22094 21496 22100 21508
rect 22152 21496 22158 21548
rect 23768 21536 23796 21567
rect 23400 21508 23796 21536
rect 23400 21480 23428 21508
rect 24302 21496 24308 21548
rect 24360 21536 24366 21548
rect 24762 21536 24768 21548
rect 24360 21508 24768 21536
rect 24360 21496 24366 21508
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 11238 21468 11244 21480
rect 8803 21440 9904 21468
rect 11151 21440 11244 21468
rect 8803 21437 8815 21440
rect 8757 21431 8815 21437
rect 11238 21428 11244 21440
rect 11296 21468 11302 21480
rect 12434 21468 12440 21480
rect 11296 21440 12440 21468
rect 11296 21428 11302 21440
rect 12434 21428 12440 21440
rect 12492 21428 12498 21480
rect 12618 21468 12624 21480
rect 12579 21440 12624 21468
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 13354 21428 13360 21480
rect 13412 21468 13418 21480
rect 13521 21471 13579 21477
rect 13521 21468 13533 21471
rect 13412 21440 13533 21468
rect 13412 21428 13418 21440
rect 13521 21437 13533 21440
rect 13567 21437 13579 21471
rect 13521 21431 13579 21437
rect 15933 21471 15991 21477
rect 15933 21437 15945 21471
rect 15979 21468 15991 21471
rect 16666 21468 16672 21480
rect 15979 21440 16672 21468
rect 15979 21437 15991 21440
rect 15933 21431 15991 21437
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 18969 21471 19027 21477
rect 18969 21468 18981 21471
rect 18616 21440 18981 21468
rect 9125 21403 9183 21409
rect 9125 21369 9137 21403
rect 9171 21400 9183 21403
rect 9582 21400 9588 21412
rect 9171 21372 9588 21400
rect 9171 21369 9183 21372
rect 9125 21363 9183 21369
rect 9582 21360 9588 21372
rect 9640 21360 9646 21412
rect 11149 21403 11207 21409
rect 11149 21369 11161 21403
rect 11195 21400 11207 21403
rect 12342 21400 12348 21412
rect 11195 21372 12348 21400
rect 11195 21369 11207 21372
rect 11149 21363 11207 21369
rect 12342 21360 12348 21372
rect 12400 21360 12406 21412
rect 16390 21360 16396 21412
rect 16448 21400 16454 21412
rect 16853 21403 16911 21409
rect 16853 21400 16865 21403
rect 16448 21372 16865 21400
rect 16448 21360 16454 21372
rect 16853 21369 16865 21372
rect 16899 21369 16911 21403
rect 16853 21363 16911 21369
rect 6273 21335 6331 21341
rect 6273 21332 6285 21335
rect 6196 21304 6285 21332
rect 6273 21301 6285 21304
rect 6319 21332 6331 21335
rect 6362 21332 6368 21344
rect 6319 21304 6368 21332
rect 6319 21301 6331 21304
rect 6273 21295 6331 21301
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 6454 21292 6460 21344
rect 6512 21332 6518 21344
rect 6825 21335 6883 21341
rect 6825 21332 6837 21335
rect 6512 21304 6837 21332
rect 6512 21292 6518 21304
rect 6825 21301 6837 21304
rect 6871 21301 6883 21335
rect 9214 21332 9220 21344
rect 9175 21304 9220 21332
rect 6825 21295 6883 21301
rect 9214 21292 9220 21304
rect 9272 21292 9278 21344
rect 9766 21292 9772 21344
rect 9824 21332 9830 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 9824 21304 10793 21332
rect 9824 21292 9830 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 10781 21295 10839 21301
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 14645 21335 14703 21341
rect 14645 21332 14657 21335
rect 13872 21304 14657 21332
rect 13872 21292 13878 21304
rect 14645 21301 14657 21304
rect 14691 21301 14703 21335
rect 14645 21295 14703 21301
rect 16301 21335 16359 21341
rect 16301 21301 16313 21335
rect 16347 21332 16359 21335
rect 16761 21335 16819 21341
rect 16761 21332 16773 21335
rect 16347 21304 16773 21332
rect 16347 21301 16359 21304
rect 16301 21295 16359 21301
rect 16761 21301 16773 21304
rect 16807 21332 16819 21335
rect 16942 21332 16948 21344
rect 16807 21304 16948 21332
rect 16807 21301 16819 21304
rect 16761 21295 16819 21301
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 17126 21292 17132 21344
rect 17184 21332 17190 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 17184 21304 17417 21332
rect 17184 21292 17190 21304
rect 17405 21301 17417 21304
rect 17451 21301 17463 21335
rect 17405 21295 17463 21301
rect 18046 21292 18052 21344
rect 18104 21332 18110 21344
rect 18325 21335 18383 21341
rect 18325 21332 18337 21335
rect 18104 21304 18337 21332
rect 18104 21292 18110 21304
rect 18325 21301 18337 21304
rect 18371 21332 18383 21335
rect 18616 21332 18644 21440
rect 18969 21437 18981 21440
rect 19015 21468 19027 21471
rect 19058 21468 19064 21480
rect 19015 21440 19064 21468
rect 19015 21437 19027 21440
rect 18969 21431 19027 21437
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 20530 21428 20536 21480
rect 20588 21468 20594 21480
rect 21910 21468 21916 21480
rect 20588 21440 21916 21468
rect 20588 21428 20594 21440
rect 21910 21428 21916 21440
rect 21968 21468 21974 21480
rect 21968 21440 22048 21468
rect 21968 21428 21974 21440
rect 18690 21360 18696 21412
rect 18748 21400 18754 21412
rect 19214 21403 19272 21409
rect 19214 21400 19226 21403
rect 18748 21372 19226 21400
rect 18748 21360 18754 21372
rect 19214 21369 19226 21372
rect 19260 21400 19272 21403
rect 19426 21400 19432 21412
rect 19260 21372 19432 21400
rect 19260 21369 19272 21372
rect 19214 21363 19272 21369
rect 19426 21360 19432 21372
rect 19484 21360 19490 21412
rect 21542 21360 21548 21412
rect 21600 21400 21606 21412
rect 21600 21372 21956 21400
rect 21600 21360 21606 21372
rect 18785 21335 18843 21341
rect 18785 21332 18797 21335
rect 18371 21304 18797 21332
rect 18371 21301 18383 21304
rect 18325 21295 18383 21301
rect 18785 21301 18797 21304
rect 18831 21301 18843 21335
rect 20346 21332 20352 21344
rect 20307 21304 20352 21332
rect 18785 21295 18843 21301
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 21361 21335 21419 21341
rect 21361 21301 21373 21335
rect 21407 21332 21419 21335
rect 21634 21332 21640 21344
rect 21407 21304 21640 21332
rect 21407 21301 21419 21304
rect 21361 21295 21419 21301
rect 21634 21292 21640 21304
rect 21692 21332 21698 21344
rect 21928 21341 21956 21372
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 21692 21304 21833 21332
rect 21692 21292 21698 21304
rect 21821 21301 21833 21304
rect 21867 21301 21879 21335
rect 21821 21295 21879 21301
rect 21913 21335 21971 21341
rect 21913 21301 21925 21335
rect 21959 21301 21971 21335
rect 22020 21332 22048 21440
rect 23382 21428 23388 21480
rect 23440 21428 23446 21480
rect 24121 21471 24179 21477
rect 24121 21468 24133 21471
rect 23676 21440 24133 21468
rect 23109 21403 23167 21409
rect 23109 21369 23121 21403
rect 23155 21400 23167 21403
rect 23474 21400 23480 21412
rect 23155 21372 23480 21400
rect 23155 21369 23167 21372
rect 23109 21363 23167 21369
rect 23474 21360 23480 21372
rect 23532 21400 23538 21412
rect 23676 21400 23704 21440
rect 24121 21437 24133 21440
rect 24167 21468 24179 21471
rect 24854 21468 24860 21480
rect 24167 21440 24860 21468
rect 24167 21437 24179 21440
rect 24121 21431 24179 21437
rect 24854 21428 24860 21440
rect 24912 21428 24918 21480
rect 25314 21468 25320 21480
rect 25275 21440 25320 21468
rect 25314 21428 25320 21440
rect 25372 21468 25378 21480
rect 25869 21471 25927 21477
rect 25869 21468 25881 21471
rect 25372 21440 25881 21468
rect 25372 21428 25378 21440
rect 25869 21437 25881 21440
rect 25915 21437 25927 21471
rect 25869 21431 25927 21437
rect 23532 21372 23704 21400
rect 23532 21360 23538 21372
rect 23842 21360 23848 21412
rect 23900 21400 23906 21412
rect 25133 21403 25191 21409
rect 25133 21400 25145 21403
rect 23900 21372 25145 21400
rect 23900 21360 23906 21372
rect 25133 21369 25145 21372
rect 25179 21369 25191 21403
rect 25133 21363 25191 21369
rect 23385 21335 23443 21341
rect 23385 21332 23397 21335
rect 22020 21304 23397 21332
rect 21913 21295 21971 21301
rect 23385 21301 23397 21304
rect 23431 21332 23443 21335
rect 24213 21335 24271 21341
rect 24213 21332 24225 21335
rect 23431 21304 24225 21332
rect 23431 21301 23443 21304
rect 23385 21295 23443 21301
rect 24213 21301 24225 21304
rect 24259 21332 24271 21335
rect 25774 21332 25780 21344
rect 24259 21304 25780 21332
rect 24259 21301 24271 21304
rect 24213 21295 24271 21301
rect 25774 21292 25780 21304
rect 25832 21292 25838 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1394 21128 1400 21140
rect 1355 21100 1400 21128
rect 1394 21088 1400 21100
rect 1452 21088 1458 21140
rect 1854 21128 1860 21140
rect 1815 21100 1860 21128
rect 1854 21088 1860 21100
rect 1912 21088 1918 21140
rect 2038 21088 2044 21140
rect 2096 21128 2102 21140
rect 2225 21131 2283 21137
rect 2225 21128 2237 21131
rect 2096 21100 2237 21128
rect 2096 21088 2102 21100
rect 2225 21097 2237 21100
rect 2271 21097 2283 21131
rect 2406 21128 2412 21140
rect 2367 21100 2412 21128
rect 2225 21091 2283 21097
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 3326 21088 3332 21140
rect 3384 21128 3390 21140
rect 6178 21128 6184 21140
rect 3384 21100 6184 21128
rect 3384 21088 3390 21100
rect 6178 21088 6184 21100
rect 6236 21088 6242 21140
rect 6270 21088 6276 21140
rect 6328 21128 6334 21140
rect 7374 21128 7380 21140
rect 6328 21100 7380 21128
rect 6328 21088 6334 21100
rect 7374 21088 7380 21100
rect 7432 21128 7438 21140
rect 7926 21128 7932 21140
rect 7432 21100 7604 21128
rect 7887 21100 7932 21128
rect 7432 21088 7438 21100
rect 2777 21063 2835 21069
rect 2777 21029 2789 21063
rect 2823 21060 2835 21063
rect 4062 21060 4068 21072
rect 2823 21032 4068 21060
rect 2823 21029 2835 21032
rect 2777 21023 2835 21029
rect 4062 21020 4068 21032
rect 4120 21020 4126 21072
rect 5994 21060 6000 21072
rect 5955 21032 6000 21060
rect 5994 21020 6000 21032
rect 6052 21020 6058 21072
rect 7466 21020 7472 21072
rect 7524 21020 7530 21072
rect 7576 21060 7604 21100
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 9309 21131 9367 21137
rect 9309 21097 9321 21131
rect 9355 21128 9367 21131
rect 9398 21128 9404 21140
rect 9355 21100 9404 21128
rect 9355 21097 9367 21100
rect 9309 21091 9367 21097
rect 9398 21088 9404 21100
rect 9456 21088 9462 21140
rect 9950 21128 9956 21140
rect 9911 21100 9956 21128
rect 9950 21088 9956 21100
rect 10008 21088 10014 21140
rect 10042 21088 10048 21140
rect 10100 21128 10106 21140
rect 10229 21131 10287 21137
rect 10229 21128 10241 21131
rect 10100 21100 10241 21128
rect 10100 21088 10106 21100
rect 10229 21097 10241 21100
rect 10275 21097 10287 21131
rect 10229 21091 10287 21097
rect 10505 21131 10563 21137
rect 10505 21097 10517 21131
rect 10551 21128 10563 21131
rect 11238 21128 11244 21140
rect 10551 21100 11244 21128
rect 10551 21097 10563 21100
rect 10505 21091 10563 21097
rect 11238 21088 11244 21100
rect 11296 21088 11302 21140
rect 11790 21088 11796 21140
rect 11848 21128 11854 21140
rect 11885 21131 11943 21137
rect 11885 21128 11897 21131
rect 11848 21100 11897 21128
rect 11848 21088 11854 21100
rect 11885 21097 11897 21100
rect 11931 21097 11943 21131
rect 12066 21128 12072 21140
rect 12027 21100 12072 21128
rect 11885 21091 11943 21097
rect 7834 21060 7840 21072
rect 7576 21032 7840 21060
rect 7834 21020 7840 21032
rect 7892 21020 7898 21072
rect 10962 21020 10968 21072
rect 11020 21020 11026 21072
rect 11900 21060 11928 21091
rect 12066 21088 12072 21100
rect 12124 21088 12130 21140
rect 13354 21128 13360 21140
rect 13315 21100 13360 21128
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 13630 21128 13636 21140
rect 13591 21100 13636 21128
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 15841 21131 15899 21137
rect 15841 21097 15853 21131
rect 15887 21128 15899 21131
rect 15930 21128 15936 21140
rect 15887 21100 15936 21128
rect 15887 21097 15899 21100
rect 15841 21091 15899 21097
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 16390 21128 16396 21140
rect 16351 21100 16396 21128
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 19061 21131 19119 21137
rect 19061 21128 19073 21131
rect 17920 21100 19073 21128
rect 17920 21088 17926 21100
rect 19061 21097 19073 21100
rect 19107 21097 19119 21131
rect 19242 21128 19248 21140
rect 19203 21100 19248 21128
rect 19061 21091 19119 21097
rect 14001 21063 14059 21069
rect 11900 21032 12756 21060
rect 3602 20992 3608 21004
rect 3344 20964 3608 20992
rect 2866 20924 2872 20936
rect 2827 20896 2872 20924
rect 2866 20884 2872 20896
rect 2924 20884 2930 20936
rect 3344 20933 3372 20964
rect 3602 20952 3608 20964
rect 3660 20952 3666 21004
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4321 20995 4379 21001
rect 4321 20992 4333 20995
rect 4212 20964 4333 20992
rect 4212 20952 4218 20964
rect 4321 20961 4333 20964
rect 4367 20961 4379 20995
rect 4321 20955 4379 20961
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 7285 20995 7343 21001
rect 7285 20992 7297 20995
rect 6972 20964 7297 20992
rect 6972 20952 6978 20964
rect 7285 20961 7297 20964
rect 7331 20992 7343 20995
rect 7484 20992 7512 21020
rect 7331 20964 7512 20992
rect 8481 20995 8539 21001
rect 7331 20961 7343 20964
rect 7285 20955 7343 20961
rect 8481 20961 8493 20995
rect 8527 20992 8539 20995
rect 8570 20992 8576 21004
rect 8527 20964 8576 20992
rect 8527 20961 8539 20964
rect 8481 20955 8539 20961
rect 8570 20952 8576 20964
rect 8628 20952 8634 21004
rect 10870 20992 10876 21004
rect 10831 20964 10876 20992
rect 10870 20952 10876 20964
rect 10928 20952 10934 21004
rect 10980 20992 11008 21020
rect 10980 20964 11100 20992
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 3329 20927 3387 20933
rect 3329 20924 3341 20927
rect 3007 20896 3341 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 3329 20893 3341 20896
rect 3375 20893 3387 20927
rect 3329 20887 3387 20893
rect 3694 20884 3700 20936
rect 3752 20924 3758 20936
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 3752 20896 4077 20924
rect 3752 20884 3758 20896
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 4065 20887 4123 20893
rect 7561 20927 7619 20933
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 7834 20924 7840 20936
rect 7607 20896 7840 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 9214 20884 9220 20936
rect 9272 20924 9278 20936
rect 11072 20933 11100 20964
rect 11698 20952 11704 21004
rect 11756 20992 11762 21004
rect 12437 20995 12495 21001
rect 12437 20992 12449 20995
rect 11756 20964 12449 20992
rect 11756 20952 11762 20964
rect 12437 20961 12449 20964
rect 12483 20961 12495 20995
rect 12437 20955 12495 20961
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 9272 20896 10977 20924
rect 9272 20884 9278 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11057 20927 11115 20933
rect 11057 20893 11069 20927
rect 11103 20893 11115 20927
rect 11057 20887 11115 20893
rect 1854 20816 1860 20868
rect 1912 20856 1918 20868
rect 3050 20856 3056 20868
rect 1912 20828 3056 20856
rect 1912 20816 1918 20828
rect 3050 20816 3056 20828
rect 3108 20816 3114 20868
rect 3789 20859 3847 20865
rect 3789 20856 3801 20859
rect 3252 20828 3801 20856
rect 2590 20748 2596 20800
rect 2648 20788 2654 20800
rect 3252 20788 3280 20828
rect 3789 20825 3801 20828
rect 3835 20825 3847 20859
rect 3789 20819 3847 20825
rect 6457 20859 6515 20865
rect 6457 20825 6469 20859
rect 6503 20856 6515 20859
rect 6917 20859 6975 20865
rect 6917 20856 6929 20859
rect 6503 20828 6929 20856
rect 6503 20825 6515 20828
rect 6457 20819 6515 20825
rect 6917 20825 6929 20828
rect 6963 20856 6975 20859
rect 7282 20856 7288 20868
rect 6963 20828 7288 20856
rect 6963 20825 6975 20828
rect 6917 20819 6975 20825
rect 7282 20816 7288 20828
rect 7340 20816 7346 20868
rect 8662 20856 8668 20868
rect 8623 20828 8668 20856
rect 8662 20816 8668 20828
rect 8720 20816 8726 20868
rect 10980 20856 11008 20887
rect 12066 20884 12072 20936
rect 12124 20924 12130 20936
rect 12728 20933 12756 21032
rect 14001 21029 14013 21063
rect 14047 21060 14059 21063
rect 14366 21060 14372 21072
rect 14047 21032 14372 21060
rect 14047 21029 14059 21032
rect 14001 21023 14059 21029
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 15565 21063 15623 21069
rect 15565 21029 15577 21063
rect 15611 21060 15623 21063
rect 15746 21060 15752 21072
rect 15611 21032 15752 21060
rect 15611 21029 15623 21032
rect 15565 21023 15623 21029
rect 15746 21020 15752 21032
rect 15804 21060 15810 21072
rect 16574 21060 16580 21072
rect 15804 21032 16580 21060
rect 15804 21020 15810 21032
rect 16574 21020 16580 21032
rect 16632 21020 16638 21072
rect 17034 21069 17040 21072
rect 17028 21060 17040 21069
rect 16995 21032 17040 21060
rect 17028 21023 17040 21032
rect 17034 21020 17040 21023
rect 17092 21020 17098 21072
rect 18690 21060 18696 21072
rect 18651 21032 18696 21060
rect 18690 21020 18696 21032
rect 18748 21020 18754 21072
rect 19076 21060 19104 21091
rect 19242 21088 19248 21100
rect 19300 21088 19306 21140
rect 21269 21131 21327 21137
rect 21269 21097 21281 21131
rect 21315 21128 21327 21131
rect 21542 21128 21548 21140
rect 21315 21100 21548 21128
rect 21315 21097 21327 21100
rect 21269 21091 21327 21097
rect 21542 21088 21548 21100
rect 21600 21088 21606 21140
rect 22002 21128 22008 21140
rect 21963 21100 22008 21128
rect 22002 21088 22008 21100
rect 22060 21088 22066 21140
rect 22186 21088 22192 21140
rect 22244 21128 22250 21140
rect 22281 21131 22339 21137
rect 22281 21128 22293 21131
rect 22244 21100 22293 21128
rect 22244 21088 22250 21100
rect 22281 21097 22293 21100
rect 22327 21097 22339 21131
rect 22281 21091 22339 21097
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 24305 21131 24363 21137
rect 24305 21128 24317 21131
rect 23716 21100 24317 21128
rect 23716 21088 23722 21100
rect 24305 21097 24317 21100
rect 24351 21097 24363 21131
rect 24305 21091 24363 21097
rect 19794 21060 19800 21072
rect 19076 21032 19800 21060
rect 19794 21020 19800 21032
rect 19852 21060 19858 21072
rect 20346 21060 20352 21072
rect 19852 21032 20352 21060
rect 19852 21020 19858 21032
rect 20346 21020 20352 21032
rect 20404 21020 20410 21072
rect 21358 21060 21364 21072
rect 21319 21032 21364 21060
rect 21358 21020 21364 21032
rect 21416 21020 21422 21072
rect 14093 20995 14151 21001
rect 14093 20961 14105 20995
rect 14139 20992 14151 20995
rect 14826 20992 14832 21004
rect 14139 20964 14832 20992
rect 14139 20961 14151 20964
rect 14093 20955 14151 20961
rect 14826 20952 14832 20964
rect 14884 20952 14890 21004
rect 15657 20995 15715 21001
rect 15657 20961 15669 20995
rect 15703 20992 15715 20995
rect 16390 20992 16396 21004
rect 15703 20964 16396 20992
rect 15703 20961 15715 20964
rect 15657 20955 15715 20961
rect 16390 20952 16396 20964
rect 16448 20952 16454 21004
rect 19242 20952 19248 21004
rect 19300 20992 19306 21004
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 19300 20964 19625 20992
rect 19300 20952 19306 20964
rect 19613 20961 19625 20964
rect 19659 20992 19671 20995
rect 20625 20995 20683 21001
rect 20625 20992 20637 20995
rect 19659 20964 20637 20992
rect 19659 20961 19671 20964
rect 19613 20955 19671 20961
rect 20625 20961 20637 20964
rect 20671 20961 20683 20995
rect 20625 20955 20683 20961
rect 22741 20995 22799 21001
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 23290 20992 23296 21004
rect 22787 20964 23296 20992
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 23290 20952 23296 20964
rect 23348 20952 23354 21004
rect 24213 20995 24271 21001
rect 24213 20961 24225 20995
rect 24259 20992 24271 20995
rect 24670 20992 24676 21004
rect 24259 20964 24676 20992
rect 24259 20961 24271 20964
rect 24213 20955 24271 20961
rect 24670 20952 24676 20964
rect 24728 20952 24734 21004
rect 12529 20927 12587 20933
rect 12529 20924 12541 20927
rect 12124 20896 12541 20924
rect 12124 20884 12130 20896
rect 12529 20893 12541 20896
rect 12575 20893 12587 20927
rect 12529 20887 12587 20893
rect 12713 20927 12771 20933
rect 12713 20893 12725 20927
rect 12759 20893 12771 20927
rect 12713 20887 12771 20893
rect 14185 20927 14243 20933
rect 14185 20893 14197 20927
rect 14231 20893 14243 20927
rect 16758 20924 16764 20936
rect 16719 20896 16764 20924
rect 14185 20887 14243 20893
rect 11146 20856 11152 20868
rect 10980 20828 11152 20856
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 12728 20856 12756 20887
rect 13538 20856 13544 20868
rect 12728 20828 13544 20856
rect 13538 20816 13544 20828
rect 13596 20856 13602 20868
rect 14200 20856 14228 20887
rect 16758 20884 16764 20896
rect 16816 20884 16822 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19705 20927 19763 20933
rect 19705 20924 19717 20927
rect 19392 20896 19717 20924
rect 19392 20884 19398 20896
rect 19705 20893 19717 20896
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 13596 20828 14228 20856
rect 15105 20859 15163 20865
rect 13596 20816 13602 20828
rect 15105 20825 15117 20859
rect 15151 20856 15163 20859
rect 15562 20856 15568 20868
rect 15151 20828 15568 20856
rect 15151 20825 15163 20828
rect 15105 20819 15163 20825
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 17770 20816 17776 20868
rect 17828 20856 17834 20868
rect 18141 20859 18199 20865
rect 18141 20856 18153 20859
rect 17828 20828 18153 20856
rect 17828 20816 17834 20828
rect 18141 20825 18153 20828
rect 18187 20825 18199 20859
rect 19720 20856 19748 20887
rect 19794 20884 19800 20936
rect 19852 20924 19858 20936
rect 19852 20896 19897 20924
rect 19852 20884 19858 20896
rect 21450 20884 21456 20936
rect 21508 20924 21514 20936
rect 24397 20927 24455 20933
rect 21508 20896 21553 20924
rect 21508 20884 21514 20896
rect 24397 20893 24409 20927
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 20257 20859 20315 20865
rect 20257 20856 20269 20859
rect 19720 20828 20269 20856
rect 18141 20819 18199 20825
rect 20257 20825 20269 20828
rect 20303 20825 20315 20859
rect 22922 20856 22928 20868
rect 22883 20828 22928 20856
rect 20257 20819 20315 20825
rect 22922 20816 22928 20828
rect 22980 20816 22986 20868
rect 23477 20859 23535 20865
rect 23477 20825 23489 20859
rect 23523 20856 23535 20859
rect 23934 20856 23940 20868
rect 23523 20828 23940 20856
rect 23523 20825 23535 20828
rect 23477 20819 23535 20825
rect 23934 20816 23940 20828
rect 23992 20816 23998 20868
rect 24210 20816 24216 20868
rect 24268 20856 24274 20868
rect 24412 20856 24440 20887
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 25409 20927 25467 20933
rect 25409 20924 25421 20927
rect 24912 20896 25421 20924
rect 24912 20884 24918 20896
rect 25409 20893 25421 20896
rect 25455 20893 25467 20927
rect 25409 20887 25467 20893
rect 24268 20828 24440 20856
rect 24268 20816 24274 20828
rect 2648 20760 3280 20788
rect 3329 20791 3387 20797
rect 2648 20748 2654 20760
rect 3329 20757 3341 20791
rect 3375 20788 3387 20791
rect 3513 20791 3571 20797
rect 3513 20788 3525 20791
rect 3375 20760 3525 20788
rect 3375 20757 3387 20760
rect 3329 20751 3387 20757
rect 3513 20757 3525 20760
rect 3559 20788 3571 20791
rect 5442 20788 5448 20800
rect 3559 20760 5448 20788
rect 3559 20757 3571 20760
rect 3513 20751 3571 20757
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 6730 20788 6736 20800
rect 5592 20760 6736 20788
rect 5592 20748 5598 20760
rect 6730 20748 6736 20760
rect 6788 20748 6794 20800
rect 8294 20788 8300 20800
rect 8255 20760 8300 20788
rect 8294 20748 8300 20760
rect 8352 20748 8358 20800
rect 11514 20788 11520 20800
rect 11475 20760 11520 20788
rect 11514 20748 11520 20760
rect 11572 20748 11578 20800
rect 14550 20748 14556 20800
rect 14608 20788 14614 20800
rect 14645 20791 14703 20797
rect 14645 20788 14657 20791
rect 14608 20760 14657 20788
rect 14608 20748 14614 20760
rect 14645 20757 14657 20760
rect 14691 20757 14703 20791
rect 14645 20751 14703 20757
rect 20901 20791 20959 20797
rect 20901 20757 20913 20791
rect 20947 20788 20959 20791
rect 21266 20788 21272 20800
rect 20947 20760 21272 20788
rect 20947 20757 20959 20760
rect 20901 20751 20959 20757
rect 21266 20748 21272 20760
rect 21324 20748 21330 20800
rect 23842 20788 23848 20800
rect 23803 20760 23848 20788
rect 23842 20748 23848 20760
rect 23900 20748 23906 20800
rect 24946 20788 24952 20800
rect 24907 20760 24952 20788
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 25314 20788 25320 20800
rect 25275 20760 25320 20788
rect 25314 20748 25320 20760
rect 25372 20748 25378 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2041 20587 2099 20593
rect 2041 20553 2053 20587
rect 2087 20584 2099 20587
rect 2314 20584 2320 20596
rect 2087 20556 2320 20584
rect 2087 20553 2099 20556
rect 2041 20547 2099 20553
rect 1394 20380 1400 20392
rect 1452 20389 1458 20392
rect 1452 20383 1480 20389
rect 1332 20352 1400 20380
rect 1394 20340 1400 20352
rect 1468 20380 1480 20383
rect 2056 20380 2084 20547
rect 2314 20544 2320 20556
rect 2372 20544 2378 20596
rect 3142 20544 3148 20596
rect 3200 20584 3206 20596
rect 3510 20584 3516 20596
rect 3200 20556 3516 20584
rect 3200 20544 3206 20556
rect 3510 20544 3516 20556
rect 3568 20544 3574 20596
rect 4433 20587 4491 20593
rect 4433 20553 4445 20587
rect 4479 20584 4491 20587
rect 4522 20584 4528 20596
rect 4479 20556 4528 20584
rect 4479 20553 4491 20556
rect 4433 20547 4491 20553
rect 4522 20544 4528 20556
rect 4580 20544 4586 20596
rect 5442 20544 5448 20596
rect 5500 20584 5506 20596
rect 5813 20587 5871 20593
rect 5813 20584 5825 20587
rect 5500 20556 5825 20584
rect 5500 20544 5506 20556
rect 5813 20553 5825 20556
rect 5859 20553 5871 20587
rect 6270 20584 6276 20596
rect 6231 20556 6276 20584
rect 5813 20547 5871 20553
rect 6270 20544 6276 20556
rect 6328 20544 6334 20596
rect 6822 20584 6828 20596
rect 6783 20556 6828 20584
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 8110 20544 8116 20596
rect 8168 20584 8174 20596
rect 9953 20587 10011 20593
rect 9953 20584 9965 20587
rect 8168 20556 9965 20584
rect 8168 20544 8174 20556
rect 9953 20553 9965 20556
rect 9999 20553 10011 20587
rect 9953 20547 10011 20553
rect 10597 20587 10655 20593
rect 10597 20553 10609 20587
rect 10643 20584 10655 20587
rect 10962 20584 10968 20596
rect 10643 20556 10968 20584
rect 10643 20553 10655 20556
rect 10597 20547 10655 20553
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 11698 20584 11704 20596
rect 11659 20556 11704 20584
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 14366 20584 14372 20596
rect 14327 20556 14372 20584
rect 14366 20544 14372 20556
rect 14424 20544 14430 20596
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 18322 20584 18328 20596
rect 18279 20556 18328 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 18322 20544 18328 20556
rect 18380 20544 18386 20596
rect 19153 20587 19211 20593
rect 19153 20553 19165 20587
rect 19199 20584 19211 20587
rect 19242 20584 19248 20596
rect 19199 20556 19248 20584
rect 19199 20553 19211 20556
rect 19153 20547 19211 20553
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19518 20544 19524 20596
rect 19576 20544 19582 20596
rect 20530 20584 20536 20596
rect 20443 20556 20536 20584
rect 20530 20544 20536 20556
rect 20588 20584 20594 20596
rect 21358 20584 21364 20596
rect 20588 20556 21364 20584
rect 20588 20544 20594 20556
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 22094 20544 22100 20596
rect 22152 20584 22158 20596
rect 22373 20587 22431 20593
rect 22373 20584 22385 20587
rect 22152 20556 22385 20584
rect 22152 20544 22158 20556
rect 22373 20553 22385 20556
rect 22419 20553 22431 20587
rect 22373 20547 22431 20553
rect 23017 20587 23075 20593
rect 23017 20553 23029 20587
rect 23063 20584 23075 20587
rect 23290 20584 23296 20596
rect 23063 20556 23296 20584
rect 23063 20553 23075 20556
rect 23017 20547 23075 20553
rect 3970 20516 3976 20528
rect 1468 20352 2084 20380
rect 2700 20488 3976 20516
rect 2700 20380 2728 20488
rect 3970 20476 3976 20488
rect 4028 20476 4034 20528
rect 3421 20451 3479 20457
rect 3421 20448 3433 20451
rect 3160 20420 3433 20448
rect 2774 20380 2780 20392
rect 2700 20352 2780 20380
rect 1468 20349 1480 20352
rect 1452 20343 1480 20349
rect 1452 20340 1458 20343
rect 2774 20340 2780 20352
rect 2832 20340 2838 20392
rect 3160 20312 3188 20420
rect 3421 20417 3433 20420
rect 3467 20448 3479 20451
rect 4154 20448 4160 20460
rect 3467 20420 4160 20448
rect 3467 20417 3479 20420
rect 3421 20411 3479 20417
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 5077 20451 5135 20457
rect 5077 20417 5089 20451
rect 5123 20448 5135 20451
rect 5460 20448 5488 20544
rect 6730 20476 6736 20528
rect 6788 20516 6794 20528
rect 19536 20516 19564 20544
rect 6788 20488 7420 20516
rect 6788 20476 6794 20488
rect 7282 20448 7288 20460
rect 5123 20420 5488 20448
rect 7243 20420 7288 20448
rect 5123 20417 5135 20420
rect 5077 20411 5135 20417
rect 7282 20408 7288 20420
rect 7340 20408 7346 20460
rect 7392 20457 7420 20488
rect 18064 20488 19564 20516
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12437 20451 12495 20457
rect 12437 20448 12449 20451
rect 12216 20420 12449 20448
rect 12216 20408 12222 20420
rect 12437 20417 12449 20420
rect 12483 20417 12495 20451
rect 12437 20411 12495 20417
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 3292 20352 3337 20380
rect 3292 20340 3298 20352
rect 3510 20340 3516 20392
rect 3568 20380 3574 20392
rect 3970 20380 3976 20392
rect 3568 20352 3976 20380
rect 3568 20340 3574 20352
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 4893 20383 4951 20389
rect 4893 20349 4905 20383
rect 4939 20380 4951 20383
rect 6822 20380 6828 20392
rect 4939 20352 6828 20380
rect 4939 20349 4951 20352
rect 4893 20343 4951 20349
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 8573 20383 8631 20389
rect 8573 20380 8585 20383
rect 8159 20352 8585 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 8573 20349 8585 20352
rect 8619 20380 8631 20383
rect 8662 20380 8668 20392
rect 8619 20352 8668 20380
rect 8619 20349 8631 20352
rect 8573 20343 8631 20349
rect 8662 20340 8668 20352
rect 8720 20340 8726 20392
rect 10870 20380 10876 20392
rect 10831 20352 10876 20380
rect 10870 20340 10876 20352
rect 10928 20340 10934 20392
rect 15381 20383 15439 20389
rect 15381 20380 15393 20383
rect 15212 20352 15393 20380
rect 3326 20312 3332 20324
rect 2792 20284 3188 20312
rect 3287 20284 3332 20312
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 1854 20204 1860 20256
rect 1912 20244 1918 20256
rect 2792 20253 2820 20284
rect 3326 20272 3332 20284
rect 3384 20272 3390 20324
rect 3694 20272 3700 20324
rect 3752 20312 3758 20324
rect 4157 20315 4215 20321
rect 4157 20312 4169 20315
rect 3752 20284 4169 20312
rect 3752 20272 3758 20284
rect 4157 20281 4169 20284
rect 4203 20312 4215 20315
rect 4246 20312 4252 20324
rect 4203 20284 4252 20312
rect 4203 20281 4215 20284
rect 4157 20275 4215 20281
rect 4246 20272 4252 20284
rect 4304 20312 4310 20324
rect 6362 20312 6368 20324
rect 4304 20284 6368 20312
rect 4304 20272 4310 20284
rect 6362 20272 6368 20284
rect 6420 20272 6426 20324
rect 8754 20272 8760 20324
rect 8812 20321 8818 20324
rect 8812 20315 8876 20321
rect 8812 20281 8830 20315
rect 8864 20281 8876 20315
rect 8812 20275 8876 20281
rect 8812 20272 8818 20275
rect 12618 20272 12624 20324
rect 12676 20321 12682 20324
rect 12676 20315 12740 20321
rect 12676 20281 12694 20315
rect 12728 20281 12740 20315
rect 12676 20275 12740 20281
rect 12676 20272 12682 20275
rect 2317 20247 2375 20253
rect 2317 20244 2329 20247
rect 1912 20216 2329 20244
rect 1912 20204 1918 20216
rect 2317 20213 2329 20216
rect 2363 20213 2375 20247
rect 2317 20207 2375 20213
rect 2777 20247 2835 20253
rect 2777 20213 2789 20247
rect 2823 20213 2835 20247
rect 2777 20207 2835 20213
rect 2866 20204 2872 20256
rect 2924 20244 2930 20256
rect 3510 20244 3516 20256
rect 2924 20216 3516 20244
rect 2924 20204 2930 20216
rect 3510 20204 3516 20216
rect 3568 20204 3574 20256
rect 4801 20247 4859 20253
rect 4801 20213 4813 20247
rect 4847 20244 4859 20247
rect 5166 20244 5172 20256
rect 4847 20216 5172 20244
rect 4847 20213 4859 20216
rect 4801 20207 4859 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 5442 20244 5448 20256
rect 5403 20216 5448 20244
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 6641 20247 6699 20253
rect 6641 20213 6653 20247
rect 6687 20244 6699 20247
rect 6822 20244 6828 20256
rect 6687 20216 6828 20244
rect 6687 20213 6699 20216
rect 6641 20207 6699 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7190 20244 7196 20256
rect 7151 20216 7196 20244
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 8481 20247 8539 20253
rect 8481 20213 8493 20247
rect 8527 20244 8539 20247
rect 8570 20244 8576 20256
rect 8527 20216 8576 20244
rect 8527 20213 8539 20216
rect 8481 20207 8539 20213
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 11054 20244 11060 20256
rect 11015 20216 11060 20244
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 12066 20244 12072 20256
rect 12027 20216 12072 20244
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 13817 20247 13875 20253
rect 13817 20213 13829 20247
rect 13863 20244 13875 20247
rect 13906 20244 13912 20256
rect 13863 20216 13912 20244
rect 13863 20213 13875 20216
rect 13817 20207 13875 20213
rect 13906 20204 13912 20216
rect 13964 20204 13970 20256
rect 14826 20244 14832 20256
rect 14787 20216 14832 20244
rect 14826 20204 14832 20216
rect 14884 20204 14890 20256
rect 14918 20204 14924 20256
rect 14976 20244 14982 20256
rect 15212 20253 15240 20352
rect 15381 20349 15393 20352
rect 15427 20380 15439 20383
rect 16758 20380 16764 20392
rect 15427 20352 16764 20380
rect 15427 20349 15439 20352
rect 15381 20343 15439 20349
rect 16758 20340 16764 20352
rect 16816 20380 16822 20392
rect 17310 20380 17316 20392
rect 16816 20352 17316 20380
rect 16816 20340 16822 20352
rect 17310 20340 17316 20352
rect 17368 20340 17374 20392
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18064 20389 18092 20488
rect 19426 20408 19432 20460
rect 19484 20448 19490 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19484 20420 19717 20448
rect 19484 20408 19490 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 18049 20383 18107 20389
rect 18049 20380 18061 20383
rect 18012 20352 18061 20380
rect 18012 20340 18018 20352
rect 18049 20349 18061 20352
rect 18095 20349 18107 20383
rect 18049 20343 18107 20349
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 19518 20380 19524 20392
rect 18739 20352 19524 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 19518 20340 19524 20352
rect 19576 20340 19582 20392
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20956 20352 21005 20380
rect 20956 20340 20962 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 23032 20380 23060 20547
rect 23290 20544 23296 20556
rect 23348 20544 23354 20596
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 23658 20584 23664 20596
rect 23523 20556 23664 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 23658 20544 23664 20556
rect 23716 20584 23722 20596
rect 24026 20584 24032 20596
rect 23716 20556 24032 20584
rect 23716 20544 23722 20556
rect 24026 20544 24032 20556
rect 24084 20544 24090 20596
rect 25406 20584 25412 20596
rect 25367 20556 25412 20584
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 23900 20420 24133 20448
rect 23900 20408 23906 20420
rect 24121 20417 24133 20420
rect 24167 20417 24179 20451
rect 24302 20448 24308 20460
rect 24263 20420 24308 20448
rect 24121 20411 24179 20417
rect 20993 20343 21051 20349
rect 21192 20352 23060 20380
rect 24136 20380 24164 20411
rect 24302 20408 24308 20420
rect 24360 20408 24366 20460
rect 25041 20383 25099 20389
rect 25041 20380 25053 20383
rect 24136 20352 25053 20380
rect 15648 20315 15706 20321
rect 15648 20281 15660 20315
rect 15694 20312 15706 20315
rect 15746 20312 15752 20324
rect 15694 20284 15752 20312
rect 15694 20281 15706 20284
rect 15648 20275 15706 20281
rect 15746 20272 15752 20284
rect 15804 20272 15810 20324
rect 21192 20312 21220 20352
rect 25041 20349 25053 20352
rect 25087 20349 25099 20383
rect 25222 20380 25228 20392
rect 25183 20352 25228 20380
rect 25041 20343 25099 20349
rect 25222 20340 25228 20352
rect 25280 20380 25286 20392
rect 25777 20383 25835 20389
rect 25777 20380 25789 20383
rect 25280 20352 25789 20380
rect 25280 20340 25286 20352
rect 25777 20349 25789 20352
rect 25823 20349 25835 20383
rect 25777 20343 25835 20349
rect 19628 20284 21220 20312
rect 21260 20315 21318 20321
rect 15197 20247 15255 20253
rect 15197 20244 15209 20247
rect 14976 20216 15209 20244
rect 14976 20204 14982 20216
rect 15197 20213 15209 20216
rect 15243 20213 15255 20247
rect 16758 20244 16764 20256
rect 16719 20216 16764 20244
rect 15197 20207 15255 20213
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 17770 20244 17776 20256
rect 17731 20216 17776 20244
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 18966 20244 18972 20256
rect 18927 20216 18972 20244
rect 18966 20204 18972 20216
rect 19024 20244 19030 20256
rect 19628 20253 19656 20284
rect 21260 20281 21272 20315
rect 21306 20312 21318 20315
rect 21910 20312 21916 20324
rect 21306 20284 21916 20312
rect 21306 20281 21318 20284
rect 21260 20275 21318 20281
rect 21910 20272 21916 20284
rect 21968 20272 21974 20324
rect 24029 20315 24087 20321
rect 24029 20281 24041 20315
rect 24075 20312 24087 20315
rect 24762 20312 24768 20324
rect 24075 20284 24768 20312
rect 24075 20281 24087 20284
rect 24029 20275 24087 20281
rect 24762 20272 24768 20284
rect 24820 20272 24826 20324
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19024 20216 19625 20244
rect 19024 20204 19030 20216
rect 19613 20213 19625 20216
rect 19659 20213 19671 20247
rect 20898 20244 20904 20256
rect 20859 20216 20904 20244
rect 19613 20207 19671 20213
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 23661 20247 23719 20253
rect 23661 20213 23673 20247
rect 23707 20244 23719 20247
rect 23750 20244 23756 20256
rect 23707 20216 23756 20244
rect 23707 20213 23719 20216
rect 23661 20207 23719 20213
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 24670 20244 24676 20256
rect 24583 20216 24676 20244
rect 24670 20204 24676 20216
rect 24728 20244 24734 20256
rect 25866 20244 25872 20256
rect 24728 20216 25872 20244
rect 24728 20204 24734 20216
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2406 20040 2412 20052
rect 2367 20012 2412 20040
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 2869 20043 2927 20049
rect 2869 20009 2881 20043
rect 2915 20040 2927 20043
rect 3050 20040 3056 20052
rect 2915 20012 3056 20040
rect 2915 20009 2927 20012
rect 2869 20003 2927 20009
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 4062 20040 4068 20052
rect 4023 20012 4068 20040
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7248 20012 8125 20040
rect 7248 20000 7254 20012
rect 8113 20009 8125 20012
rect 8159 20009 8171 20043
rect 8113 20003 8171 20009
rect 8754 20000 8760 20052
rect 8812 20040 8818 20052
rect 11057 20043 11115 20049
rect 11057 20040 11069 20043
rect 8812 20012 11069 20040
rect 8812 20000 8818 20012
rect 11057 20009 11069 20012
rect 11103 20009 11115 20043
rect 11057 20003 11115 20009
rect 12161 20043 12219 20049
rect 12161 20009 12173 20043
rect 12207 20040 12219 20043
rect 12618 20040 12624 20052
rect 12207 20012 12624 20040
rect 12207 20009 12219 20012
rect 12161 20003 12219 20009
rect 12618 20000 12624 20012
rect 12676 20000 12682 20052
rect 13538 20040 13544 20052
rect 13499 20012 13544 20040
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 13630 20000 13636 20052
rect 13688 20040 13694 20052
rect 14642 20040 14648 20052
rect 13688 20012 13733 20040
rect 14603 20012 14648 20040
rect 13688 20000 13694 20012
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 16853 20043 16911 20049
rect 16853 20009 16865 20043
rect 16899 20040 16911 20043
rect 17034 20040 17040 20052
rect 16899 20012 17040 20040
rect 16899 20009 16911 20012
rect 16853 20003 16911 20009
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 17402 20040 17408 20052
rect 17363 20012 17408 20040
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19484 20012 19717 20040
rect 19484 20000 19490 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 21082 20040 21088 20052
rect 21043 20012 21088 20040
rect 19705 20003 19763 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21542 20040 21548 20052
rect 21503 20012 21548 20040
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 24857 20043 24915 20049
rect 24857 20040 24869 20043
rect 23440 20012 24869 20040
rect 23440 20000 23446 20012
rect 24857 20009 24869 20012
rect 24903 20009 24915 20043
rect 24857 20003 24915 20009
rect 24949 20043 25007 20049
rect 24949 20009 24961 20043
rect 24995 20040 25007 20043
rect 25038 20040 25044 20052
rect 24995 20012 25044 20040
rect 24995 20009 25007 20012
rect 24949 20003 25007 20009
rect 2130 19932 2136 19984
rect 2188 19972 2194 19984
rect 3326 19972 3332 19984
rect 2188 19944 3332 19972
rect 2188 19932 2194 19944
rect 3326 19932 3332 19944
rect 3384 19932 3390 19984
rect 4433 19975 4491 19981
rect 4433 19941 4445 19975
rect 4479 19972 4491 19975
rect 4614 19972 4620 19984
rect 4479 19944 4620 19972
rect 4479 19941 4491 19944
rect 4433 19935 4491 19941
rect 4614 19932 4620 19944
rect 4672 19932 4678 19984
rect 6080 19975 6138 19981
rect 6080 19941 6092 19975
rect 6126 19972 6138 19975
rect 7834 19972 7840 19984
rect 6126 19944 7840 19972
rect 6126 19941 6138 19944
rect 6080 19935 6138 19941
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 9674 19932 9680 19984
rect 9732 19972 9738 19984
rect 9922 19975 9980 19981
rect 9922 19972 9934 19975
rect 9732 19944 9934 19972
rect 9732 19932 9738 19944
rect 9922 19941 9934 19944
rect 9968 19941 9980 19975
rect 9922 19935 9980 19941
rect 12066 19932 12072 19984
rect 12124 19972 12130 19984
rect 20717 19975 20775 19981
rect 12124 19944 17264 19972
rect 12124 19932 12130 19944
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2590 19904 2596 19916
rect 1443 19876 2596 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2590 19864 2596 19876
rect 2648 19864 2654 19916
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 2832 19876 2877 19904
rect 2832 19864 2838 19876
rect 4154 19864 4160 19916
rect 4212 19904 4218 19916
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 4212 19876 5181 19904
rect 4212 19864 4218 19876
rect 2866 19796 2872 19848
rect 2924 19836 2930 19848
rect 3053 19839 3111 19845
rect 3053 19836 3065 19839
rect 2924 19808 3065 19836
rect 2924 19796 2930 19808
rect 3053 19805 3065 19808
rect 3099 19836 3111 19839
rect 4522 19836 4528 19848
rect 3099 19808 3740 19836
rect 4483 19808 4528 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 1581 19771 1639 19777
rect 1581 19737 1593 19771
rect 1627 19768 1639 19771
rect 2406 19768 2412 19780
rect 1627 19740 2412 19768
rect 1627 19737 1639 19740
rect 1581 19731 1639 19737
rect 2406 19728 2412 19740
rect 2464 19728 2470 19780
rect 3712 19712 3740 19808
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4632 19845 4660 19876
rect 5169 19873 5181 19876
rect 5215 19904 5227 19907
rect 5442 19904 5448 19916
rect 5215 19876 5448 19904
rect 5215 19873 5227 19876
rect 5169 19867 5227 19873
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 5813 19907 5871 19913
rect 5813 19873 5825 19907
rect 5859 19904 5871 19907
rect 6362 19904 6368 19916
rect 5859 19876 6368 19904
rect 5859 19873 5871 19876
rect 5813 19867 5871 19873
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 8297 19907 8355 19913
rect 8297 19873 8309 19907
rect 8343 19904 8355 19907
rect 8846 19904 8852 19916
rect 8343 19876 8852 19904
rect 8343 19873 8355 19876
rect 8297 19867 8355 19873
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 9692 19904 9720 19932
rect 17236 19916 17264 19944
rect 20717 19941 20729 19975
rect 20763 19972 20775 19975
rect 21450 19972 21456 19984
rect 20763 19944 21456 19972
rect 20763 19941 20775 19944
rect 20717 19935 20775 19941
rect 21450 19932 21456 19944
rect 21508 19932 21514 19984
rect 24872 19972 24900 20003
rect 25038 20000 25044 20012
rect 25096 20000 25102 20052
rect 25501 19975 25559 19981
rect 25501 19972 25513 19975
rect 24872 19944 25513 19972
rect 25501 19941 25513 19944
rect 25547 19941 25559 19975
rect 25501 19935 25559 19941
rect 9272 19876 9720 19904
rect 9272 19864 9278 19876
rect 12158 19864 12164 19916
rect 12216 19904 12222 19916
rect 12437 19907 12495 19913
rect 12437 19904 12449 19907
rect 12216 19876 12449 19904
rect 12216 19864 12222 19876
rect 12437 19873 12449 19876
rect 12483 19904 12495 19907
rect 13630 19904 13636 19916
rect 12483 19876 13636 19904
rect 12483 19873 12495 19876
rect 12437 19867 12495 19873
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 13998 19904 14004 19916
rect 13959 19876 14004 19904
rect 13998 19864 14004 19876
rect 14056 19864 14062 19916
rect 14093 19907 14151 19913
rect 14093 19873 14105 19907
rect 14139 19904 14151 19907
rect 15013 19907 15071 19913
rect 15013 19904 15025 19907
rect 14139 19876 15025 19904
rect 14139 19873 14151 19876
rect 14093 19867 14151 19873
rect 15013 19873 15025 19876
rect 15059 19873 15071 19907
rect 15013 19867 15071 19873
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 8662 19796 8668 19848
rect 8720 19836 8726 19848
rect 9674 19836 9680 19848
rect 8720 19808 9680 19836
rect 8720 19796 8726 19808
rect 9674 19796 9680 19808
rect 9732 19836 9738 19848
rect 11606 19836 11612 19848
rect 9732 19808 9777 19836
rect 11567 19808 11612 19836
rect 9732 19796 9738 19808
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 12618 19836 12624 19848
rect 12579 19808 12624 19836
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 13814 19796 13820 19848
rect 13872 19836 13878 19848
rect 14108 19836 14136 19867
rect 15286 19864 15292 19916
rect 15344 19904 15350 19916
rect 15657 19907 15715 19913
rect 15657 19904 15669 19907
rect 15344 19876 15669 19904
rect 15344 19864 15350 19876
rect 15657 19873 15669 19876
rect 15703 19873 15715 19907
rect 15838 19904 15844 19916
rect 15657 19867 15715 19873
rect 15764 19876 15844 19904
rect 14274 19836 14280 19848
rect 13872 19808 14136 19836
rect 14235 19808 14280 19836
rect 13872 19796 13878 19808
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 15470 19796 15476 19848
rect 15528 19836 15534 19848
rect 15764 19845 15792 19876
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 17218 19904 17224 19916
rect 17131 19876 17224 19904
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 18598 19913 18604 19916
rect 18592 19904 18604 19913
rect 18559 19876 18604 19904
rect 18592 19867 18604 19876
rect 18598 19864 18604 19867
rect 18656 19864 18662 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 22272 19907 22330 19913
rect 22272 19873 22284 19907
rect 22318 19904 22330 19907
rect 23014 19904 23020 19916
rect 22318 19876 23020 19904
rect 22318 19873 22330 19876
rect 22272 19867 22330 19873
rect 23014 19864 23020 19876
rect 23072 19904 23078 19916
rect 23290 19904 23296 19916
rect 23072 19876 23296 19904
rect 23072 19864 23078 19876
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 15749 19839 15807 19845
rect 15749 19836 15761 19839
rect 15528 19808 15761 19836
rect 15528 19796 15534 19808
rect 15749 19805 15761 19808
rect 15795 19805 15807 19839
rect 15930 19836 15936 19848
rect 15843 19808 15936 19836
rect 15749 19799 15807 19805
rect 15930 19796 15936 19808
rect 15988 19836 15994 19848
rect 16758 19836 16764 19848
rect 15988 19808 16764 19836
rect 15988 19796 15994 19808
rect 16758 19796 16764 19808
rect 16816 19796 16822 19848
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 18064 19808 18337 19836
rect 6822 19728 6828 19780
rect 6880 19768 6886 19780
rect 8754 19768 8760 19780
rect 6880 19740 8760 19768
rect 6880 19728 6886 19740
rect 8754 19728 8760 19740
rect 8812 19768 8818 19780
rect 8849 19771 8907 19777
rect 8849 19768 8861 19771
rect 8812 19740 8861 19768
rect 8812 19728 8818 19740
rect 8849 19737 8861 19740
rect 8895 19737 8907 19771
rect 8849 19731 8907 19737
rect 18064 19712 18092 19808
rect 18325 19805 18337 19808
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19978 19836 19984 19848
rect 19392 19808 19984 19836
rect 19392 19796 19398 19808
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19805 22063 19839
rect 24302 19836 24308 19848
rect 22005 19799 22063 19805
rect 23400 19808 24308 19836
rect 20898 19728 20904 19780
rect 20956 19768 20962 19780
rect 22020 19768 22048 19799
rect 23400 19777 23428 19808
rect 24302 19796 24308 19808
rect 24360 19836 24366 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 24360 19808 24409 19836
rect 24360 19796 24366 19808
rect 24397 19805 24409 19808
rect 24443 19836 24455 19839
rect 25130 19836 25136 19848
rect 24443 19808 25136 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 25130 19796 25136 19808
rect 25188 19796 25194 19848
rect 20956 19740 22048 19768
rect 23385 19771 23443 19777
rect 20956 19728 20962 19740
rect 23385 19737 23397 19771
rect 23431 19737 23443 19771
rect 23385 19731 23443 19737
rect 23658 19728 23664 19780
rect 23716 19768 23722 19780
rect 24489 19771 24547 19777
rect 24489 19768 24501 19771
rect 23716 19740 24501 19768
rect 23716 19728 23722 19740
rect 24489 19737 24501 19740
rect 24535 19737 24547 19771
rect 24489 19731 24547 19737
rect 1486 19660 1492 19712
rect 1544 19700 1550 19712
rect 1854 19700 1860 19712
rect 1544 19672 1860 19700
rect 1544 19660 1550 19672
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 2038 19660 2044 19712
rect 2096 19700 2102 19712
rect 2225 19703 2283 19709
rect 2225 19700 2237 19703
rect 2096 19672 2237 19700
rect 2096 19660 2102 19672
rect 2225 19669 2237 19672
rect 2271 19669 2283 19703
rect 3694 19700 3700 19712
rect 3655 19672 3700 19700
rect 2225 19663 2283 19669
rect 3694 19660 3700 19672
rect 3752 19660 3758 19712
rect 5534 19700 5540 19712
rect 5495 19672 5540 19700
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 7193 19703 7251 19709
rect 7193 19700 7205 19703
rect 6788 19672 7205 19700
rect 6788 19660 6794 19672
rect 7193 19669 7205 19672
rect 7239 19669 7251 19703
rect 7193 19663 7251 19669
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 8481 19703 8539 19709
rect 8481 19700 8493 19703
rect 7340 19672 8493 19700
rect 7340 19660 7346 19672
rect 8481 19669 8493 19672
rect 8527 19669 8539 19703
rect 9306 19700 9312 19712
rect 9267 19672 9312 19700
rect 8481 19663 8539 19669
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 13170 19700 13176 19712
rect 13083 19672 13176 19700
rect 13170 19660 13176 19672
rect 13228 19700 13234 19712
rect 13446 19700 13452 19712
rect 13228 19672 13452 19700
rect 13228 19660 13234 19672
rect 13446 19660 13452 19672
rect 13504 19660 13510 19712
rect 13998 19660 14004 19712
rect 14056 19700 14062 19712
rect 15289 19703 15347 19709
rect 15289 19700 15301 19703
rect 14056 19672 15301 19700
rect 14056 19660 14062 19672
rect 15289 19669 15301 19672
rect 15335 19669 15347 19703
rect 16390 19700 16396 19712
rect 16351 19672 16396 19700
rect 15289 19663 15347 19669
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 18046 19700 18052 19712
rect 18007 19672 18052 19700
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 19978 19660 19984 19712
rect 20036 19700 20042 19712
rect 20257 19703 20315 19709
rect 20257 19700 20269 19703
rect 20036 19672 20269 19700
rect 20036 19660 20042 19672
rect 20257 19669 20269 19672
rect 20303 19669 20315 19703
rect 21910 19700 21916 19712
rect 21871 19672 21916 19700
rect 20257 19663 20315 19669
rect 21910 19660 21916 19672
rect 21968 19660 21974 19712
rect 23290 19660 23296 19712
rect 23348 19700 23354 19712
rect 23937 19703 23995 19709
rect 23937 19700 23949 19703
rect 23348 19672 23949 19700
rect 23348 19660 23354 19672
rect 23937 19669 23949 19672
rect 23983 19700 23995 19703
rect 24210 19700 24216 19712
rect 23983 19672 24216 19700
rect 23983 19669 23995 19672
rect 23937 19663 23995 19669
rect 24210 19660 24216 19672
rect 24268 19660 24274 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2961 19499 3019 19505
rect 2961 19465 2973 19499
rect 3007 19496 3019 19499
rect 3050 19496 3056 19508
rect 3007 19468 3056 19496
rect 3007 19465 3019 19468
rect 2961 19459 3019 19465
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 5166 19496 5172 19508
rect 3712 19468 5028 19496
rect 5127 19468 5172 19496
rect 1118 19388 1124 19440
rect 1176 19428 1182 19440
rect 3712 19428 3740 19468
rect 1176 19400 3740 19428
rect 1176 19388 1182 19400
rect 3786 19388 3792 19440
rect 3844 19428 3850 19440
rect 4062 19428 4068 19440
rect 3844 19400 4068 19428
rect 3844 19388 3850 19400
rect 4062 19388 4068 19400
rect 4120 19388 4126 19440
rect 5000 19428 5028 19468
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 6273 19499 6331 19505
rect 6273 19465 6285 19499
rect 6319 19496 6331 19499
rect 6362 19496 6368 19508
rect 6319 19468 6368 19496
rect 6319 19465 6331 19468
rect 6273 19459 6331 19465
rect 6362 19456 6368 19468
rect 6420 19496 6426 19508
rect 8662 19496 8668 19508
rect 6420 19468 8668 19496
rect 6420 19456 6426 19468
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 9732 19468 10241 19496
rect 9732 19456 9738 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 10229 19459 10287 19465
rect 13630 19456 13636 19508
rect 13688 19496 13694 19508
rect 14369 19499 14427 19505
rect 14369 19496 14381 19499
rect 13688 19468 14381 19496
rect 13688 19456 13694 19468
rect 14369 19465 14381 19468
rect 14415 19496 14427 19499
rect 14826 19496 14832 19508
rect 14415 19468 14832 19496
rect 14415 19465 14427 19468
rect 14369 19459 14427 19465
rect 7282 19428 7288 19440
rect 5000 19400 7288 19428
rect 7282 19388 7288 19400
rect 7340 19388 7346 19440
rect 7834 19428 7840 19440
rect 7484 19400 7840 19428
rect 7484 19372 7512 19400
rect 7834 19388 7840 19400
rect 7892 19388 7898 19440
rect 9306 19388 9312 19440
rect 9364 19428 9370 19440
rect 9364 19400 9812 19428
rect 9364 19388 9370 19400
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 2038 19360 2044 19372
rect 1719 19332 2044 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 2038 19320 2044 19332
rect 2096 19360 2102 19372
rect 2409 19363 2467 19369
rect 2409 19360 2421 19363
rect 2096 19332 2421 19360
rect 2096 19320 2102 19332
rect 2409 19329 2421 19332
rect 2455 19329 2467 19363
rect 2409 19323 2467 19329
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 4249 19363 4307 19369
rect 4249 19360 4261 19363
rect 3752 19332 4261 19360
rect 3752 19320 3758 19332
rect 4249 19329 4261 19332
rect 4295 19329 4307 19363
rect 4249 19323 4307 19329
rect 1854 19252 1860 19304
rect 1912 19292 1918 19304
rect 2314 19292 2320 19304
rect 1912 19264 2320 19292
rect 1912 19252 1918 19264
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 3936 19264 4077 19292
rect 3936 19252 3942 19264
rect 4065 19261 4077 19264
rect 4111 19261 4123 19295
rect 4264 19292 4292 19323
rect 5350 19320 5356 19372
rect 5408 19360 5414 19372
rect 5721 19363 5779 19369
rect 5721 19360 5733 19363
rect 5408 19332 5733 19360
rect 5408 19320 5414 19332
rect 5721 19329 5733 19332
rect 5767 19329 5779 19363
rect 7466 19360 7472 19372
rect 7379 19332 7472 19360
rect 5721 19323 5779 19329
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 9784 19369 9812 19400
rect 9677 19363 9735 19369
rect 9677 19360 9689 19363
rect 9640 19332 9689 19360
rect 9640 19320 9646 19332
rect 9677 19329 9689 19332
rect 9723 19329 9735 19363
rect 9677 19323 9735 19329
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 9858 19360 9864 19372
rect 9815 19332 9864 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 11425 19363 11483 19369
rect 11425 19360 11437 19363
rect 11072 19332 11437 19360
rect 5534 19292 5540 19304
rect 4264 19264 5120 19292
rect 5495 19264 5540 19292
rect 4065 19255 4123 19261
rect 1670 19184 1676 19236
rect 1728 19224 1734 19236
rect 2222 19224 2228 19236
rect 1728 19196 2228 19224
rect 1728 19184 1734 19196
rect 2222 19184 2228 19196
rect 2280 19184 2286 19236
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19224 3571 19227
rect 3786 19224 3792 19236
rect 3559 19196 3792 19224
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 3786 19184 3792 19196
rect 3844 19224 3850 19236
rect 3973 19227 4031 19233
rect 3973 19224 3985 19227
rect 3844 19196 3985 19224
rect 3844 19184 3850 19196
rect 3973 19193 3985 19196
rect 4019 19193 4031 19227
rect 3973 19187 4031 19193
rect 5092 19168 5120 19264
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 7282 19292 7288 19304
rect 6687 19264 7288 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 7834 19292 7840 19304
rect 7795 19264 7840 19292
rect 7834 19252 7840 19264
rect 7892 19252 7898 19304
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9214 19292 9220 19304
rect 9171 19264 9220 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 9490 19252 9496 19304
rect 9548 19292 9554 19304
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 9548 19264 10701 19292
rect 9548 19252 9554 19264
rect 10689 19261 10701 19264
rect 10735 19292 10747 19295
rect 11072 19292 11100 19332
rect 11425 19329 11437 19332
rect 11471 19360 11483 19363
rect 12342 19360 12348 19372
rect 11471 19332 12348 19360
rect 11471 19329 11483 19332
rect 11425 19323 11483 19329
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 13633 19363 13691 19369
rect 13633 19360 13645 19363
rect 12452 19332 13645 19360
rect 10735 19264 11100 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 11146 19252 11152 19304
rect 11204 19292 11210 19304
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11204 19264 11805 19292
rect 11204 19252 11210 19264
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 11793 19255 11851 19261
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12452 19292 12480 19332
rect 13633 19329 13645 19332
rect 13679 19360 13691 19363
rect 14384 19360 14412 19459
rect 14826 19456 14832 19468
rect 14884 19456 14890 19508
rect 15286 19456 15292 19508
rect 15344 19496 15350 19508
rect 16485 19499 16543 19505
rect 16485 19496 16497 19499
rect 15344 19468 16497 19496
rect 15344 19456 15350 19468
rect 16485 19465 16497 19468
rect 16531 19465 16543 19499
rect 16485 19459 16543 19465
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 16853 19499 16911 19505
rect 16853 19496 16865 19499
rect 16816 19468 16865 19496
rect 16816 19456 16822 19468
rect 16853 19465 16865 19468
rect 16899 19465 16911 19499
rect 17218 19496 17224 19508
rect 17179 19468 17224 19496
rect 16853 19459 16911 19465
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 17310 19456 17316 19508
rect 17368 19496 17374 19508
rect 17773 19499 17831 19505
rect 17773 19496 17785 19499
rect 17368 19468 17785 19496
rect 17368 19456 17374 19468
rect 17773 19465 17785 19468
rect 17819 19465 17831 19499
rect 17773 19459 17831 19465
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 13679 19332 13860 19360
rect 14384 19332 14565 19360
rect 13679 19329 13691 19332
rect 13633 19323 13691 19329
rect 12299 19264 12480 19292
rect 12897 19295 12955 19301
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 13078 19292 13084 19304
rect 12943 19264 13084 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 13446 19292 13452 19304
rect 13407 19264 13452 19292
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 13832 19292 13860 19332
rect 14553 19329 14565 19332
rect 14599 19329 14611 19363
rect 15930 19360 15936 19372
rect 14553 19323 14611 19329
rect 15571 19332 15936 19360
rect 14826 19301 14832 19304
rect 14820 19292 14832 19301
rect 13832 19264 14832 19292
rect 14820 19255 14832 19264
rect 14884 19292 14890 19304
rect 15571 19292 15599 19332
rect 15930 19320 15936 19332
rect 15988 19320 15994 19372
rect 17788 19360 17816 19459
rect 25038 19456 25044 19508
rect 25096 19496 25102 19508
rect 25961 19499 26019 19505
rect 25961 19496 25973 19499
rect 25096 19468 25973 19496
rect 25096 19456 25102 19468
rect 25961 19465 25973 19468
rect 26007 19465 26019 19499
rect 25961 19459 26019 19465
rect 25130 19388 25136 19440
rect 25188 19428 25194 19440
rect 25593 19431 25651 19437
rect 25593 19428 25605 19431
rect 25188 19400 25605 19428
rect 25188 19388 25194 19400
rect 25593 19397 25605 19400
rect 25639 19397 25651 19431
rect 25593 19391 25651 19397
rect 18046 19360 18052 19372
rect 17788 19332 18052 19360
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 14884 19264 15599 19292
rect 18064 19292 18092 19320
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 18064 19264 20361 19292
rect 14826 19252 14832 19255
rect 14884 19252 14890 19264
rect 20349 19261 20361 19264
rect 20395 19292 20407 19295
rect 20898 19292 20904 19304
rect 20395 19264 20904 19292
rect 20395 19261 20407 19264
rect 20349 19255 20407 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 23661 19295 23719 19301
rect 23661 19292 23673 19295
rect 23400 19264 23673 19292
rect 5629 19227 5687 19233
rect 5629 19193 5641 19227
rect 5675 19224 5687 19227
rect 8665 19227 8723 19233
rect 8665 19224 8677 19227
rect 5675 19196 8677 19224
rect 5675 19193 5687 19196
rect 5629 19187 5687 19193
rect 1857 19159 1915 19165
rect 1857 19125 1869 19159
rect 1903 19156 1915 19159
rect 1946 19156 1952 19168
rect 1903 19128 1952 19156
rect 1903 19125 1915 19128
rect 1857 19119 1915 19125
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 3602 19156 3608 19168
rect 3563 19128 3608 19156
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 4614 19156 4620 19168
rect 4575 19128 4620 19156
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 5074 19156 5080 19168
rect 5035 19128 5080 19156
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 6840 19165 6868 19196
rect 8665 19193 8677 19196
rect 8711 19193 8723 19227
rect 11241 19227 11299 19233
rect 11241 19224 11253 19227
rect 8665 19187 8723 19193
rect 9232 19196 11253 19224
rect 6825 19159 6883 19165
rect 6825 19125 6837 19159
rect 6871 19125 6883 19159
rect 6825 19119 6883 19125
rect 7006 19116 7012 19168
rect 7064 19156 7070 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 7064 19128 7205 19156
rect 7064 19116 7070 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7193 19119 7251 19125
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 8202 19156 8208 19168
rect 7340 19128 8208 19156
rect 7340 19116 7346 19128
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8389 19159 8447 19165
rect 8389 19125 8401 19159
rect 8435 19156 8447 19159
rect 8846 19156 8852 19168
rect 8435 19128 8852 19156
rect 8435 19125 8447 19128
rect 8389 19119 8447 19125
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 9232 19165 9260 19196
rect 11241 19193 11253 19196
rect 11287 19224 11299 19227
rect 12158 19224 12164 19236
rect 11287 19196 12164 19224
rect 11287 19193 11299 19196
rect 11241 19187 11299 19193
rect 12158 19184 12164 19196
rect 12216 19184 12222 19236
rect 13722 19224 13728 19236
rect 13004 19196 13728 19224
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19125 9275 19159
rect 9217 19119 9275 19125
rect 9398 19116 9404 19168
rect 9456 19156 9462 19168
rect 9585 19159 9643 19165
rect 9585 19156 9597 19159
rect 9456 19128 9597 19156
rect 9456 19116 9462 19128
rect 9585 19125 9597 19128
rect 9631 19125 9643 19159
rect 9585 19119 9643 19125
rect 10686 19116 10692 19168
rect 10744 19156 10750 19168
rect 10781 19159 10839 19165
rect 10781 19156 10793 19159
rect 10744 19128 10793 19156
rect 10744 19116 10750 19128
rect 10781 19125 10793 19128
rect 10827 19125 10839 19159
rect 11146 19156 11152 19168
rect 11107 19128 11152 19156
rect 10781 19119 10839 19125
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 13004 19165 13032 19196
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 14093 19227 14151 19233
rect 14093 19193 14105 19227
rect 14139 19224 14151 19227
rect 14274 19224 14280 19236
rect 14139 19196 14280 19224
rect 14139 19193 14151 19196
rect 14093 19187 14151 19193
rect 14274 19184 14280 19196
rect 14332 19224 14338 19236
rect 18316 19227 18374 19233
rect 14332 19196 14688 19224
rect 14332 19184 14338 19196
rect 12989 19159 13047 19165
rect 12989 19125 13001 19159
rect 13035 19125 13047 19159
rect 12989 19119 13047 19125
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 13357 19159 13415 19165
rect 13357 19156 13369 19159
rect 13136 19128 13369 19156
rect 13136 19116 13142 19128
rect 13357 19125 13369 19128
rect 13403 19125 13415 19159
rect 13357 19119 13415 19125
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 14660 19156 14688 19196
rect 18316 19193 18328 19227
rect 18362 19224 18374 19227
rect 18506 19224 18512 19236
rect 18362 19196 18512 19224
rect 18362 19193 18374 19196
rect 18316 19187 18374 19193
rect 18506 19184 18512 19196
rect 18564 19184 18570 19236
rect 20073 19227 20131 19233
rect 20073 19193 20085 19227
rect 20119 19224 20131 19227
rect 20438 19224 20444 19236
rect 20119 19196 20444 19224
rect 20119 19193 20131 19196
rect 20073 19187 20131 19193
rect 20438 19184 20444 19196
rect 20496 19184 20502 19236
rect 21174 19233 21180 19236
rect 21168 19224 21180 19233
rect 21135 19196 21180 19224
rect 21168 19187 21180 19196
rect 21174 19184 21180 19187
rect 21232 19184 21238 19236
rect 23198 19224 23204 19236
rect 22296 19196 23204 19224
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 14608 19128 15945 19156
rect 14608 19116 14614 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 18598 19116 18604 19168
rect 18656 19156 18662 19168
rect 19429 19159 19487 19165
rect 19429 19156 19441 19159
rect 18656 19128 19441 19156
rect 18656 19116 18662 19128
rect 19429 19125 19441 19128
rect 19475 19125 19487 19159
rect 20806 19156 20812 19168
rect 20767 19128 20812 19156
rect 19429 19119 19487 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 22296 19165 22324 19196
rect 23198 19184 23204 19196
rect 23256 19184 23262 19236
rect 22281 19159 22339 19165
rect 22281 19125 22293 19159
rect 22327 19125 22339 19159
rect 22281 19119 22339 19125
rect 22925 19159 22983 19165
rect 22925 19125 22937 19159
rect 22971 19156 22983 19159
rect 23014 19156 23020 19168
rect 22971 19128 23020 19156
rect 22971 19125 22983 19128
rect 22925 19119 22983 19125
rect 23014 19116 23020 19128
rect 23072 19156 23078 19168
rect 23400 19165 23428 19264
rect 23661 19261 23673 19264
rect 23707 19261 23719 19295
rect 23661 19255 23719 19261
rect 23928 19295 23986 19301
rect 23928 19261 23940 19295
rect 23974 19292 23986 19295
rect 25130 19292 25136 19304
rect 23974 19264 25136 19292
rect 23974 19261 23986 19264
rect 23928 19255 23986 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 23385 19159 23443 19165
rect 23385 19156 23397 19159
rect 23072 19128 23397 19156
rect 23072 19116 23078 19128
rect 23385 19125 23397 19128
rect 23431 19125 23443 19159
rect 23385 19119 23443 19125
rect 23842 19116 23848 19168
rect 23900 19156 23906 19168
rect 25041 19159 25099 19165
rect 25041 19156 25053 19159
rect 23900 19128 25053 19156
rect 23900 19116 23906 19128
rect 25041 19125 25053 19128
rect 25087 19125 25099 19159
rect 25041 19119 25099 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1857 18955 1915 18961
rect 1857 18921 1869 18955
rect 1903 18952 1915 18955
rect 2130 18952 2136 18964
rect 1903 18924 2136 18952
rect 1903 18921 1915 18924
rect 1857 18915 1915 18921
rect 2130 18912 2136 18924
rect 2188 18912 2194 18964
rect 2866 18952 2872 18964
rect 2827 18924 2872 18952
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 2961 18955 3019 18961
rect 2961 18921 2973 18955
rect 3007 18952 3019 18955
rect 4614 18952 4620 18964
rect 3007 18924 4620 18952
rect 3007 18921 3019 18924
rect 2961 18915 3019 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 5169 18955 5227 18961
rect 5169 18921 5181 18955
rect 5215 18952 5227 18955
rect 5350 18952 5356 18964
rect 5215 18924 5356 18952
rect 5215 18921 5227 18924
rect 5169 18915 5227 18921
rect 5350 18912 5356 18924
rect 5408 18912 5414 18964
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 5813 18955 5871 18961
rect 5813 18952 5825 18955
rect 5592 18924 5825 18952
rect 5592 18912 5598 18924
rect 5813 18921 5825 18924
rect 5859 18921 5871 18955
rect 5813 18915 5871 18921
rect 6178 18912 6184 18964
rect 6236 18952 6242 18964
rect 7006 18952 7012 18964
rect 6236 18924 7012 18952
rect 6236 18912 6242 18924
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 7190 18912 7196 18964
rect 7248 18952 7254 18964
rect 7377 18955 7435 18961
rect 7377 18952 7389 18955
rect 7248 18924 7389 18952
rect 7248 18912 7254 18924
rect 7377 18921 7389 18924
rect 7423 18921 7435 18955
rect 7834 18952 7840 18964
rect 7795 18924 7840 18952
rect 7377 18915 7435 18921
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 9861 18955 9919 18961
rect 9861 18921 9873 18955
rect 9907 18952 9919 18955
rect 11146 18952 11152 18964
rect 9907 18924 11152 18952
rect 9907 18921 9919 18924
rect 9861 18915 9919 18921
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 13354 18952 13360 18964
rect 13315 18924 13360 18952
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 14737 18955 14795 18961
rect 14737 18921 14749 18955
rect 14783 18952 14795 18955
rect 14826 18952 14832 18964
rect 14783 18924 14832 18952
rect 14783 18921 14795 18924
rect 14737 18915 14795 18921
rect 14826 18912 14832 18924
rect 14884 18912 14890 18964
rect 15010 18952 15016 18964
rect 14971 18924 15016 18952
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 17494 18952 17500 18964
rect 17455 18924 17500 18952
rect 17494 18912 17500 18924
rect 17552 18912 17558 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 17865 18955 17923 18961
rect 17865 18952 17877 18955
rect 17828 18924 17877 18952
rect 17828 18912 17834 18924
rect 17865 18921 17877 18924
rect 17911 18921 17923 18955
rect 18598 18952 18604 18964
rect 18559 18924 18604 18952
rect 17865 18915 17923 18921
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 19061 18955 19119 18961
rect 19061 18921 19073 18955
rect 19107 18952 19119 18955
rect 19242 18952 19248 18964
rect 19107 18924 19248 18952
rect 19107 18921 19119 18924
rect 19061 18915 19119 18921
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 21726 18912 21732 18964
rect 21784 18952 21790 18964
rect 22002 18952 22008 18964
rect 21784 18924 22008 18952
rect 21784 18912 21790 18924
rect 22002 18912 22008 18924
rect 22060 18952 22066 18964
rect 22097 18955 22155 18961
rect 22097 18952 22109 18955
rect 22060 18924 22109 18952
rect 22060 18912 22066 18924
rect 22097 18921 22109 18924
rect 22143 18921 22155 18955
rect 24762 18952 24768 18964
rect 24723 18924 24768 18952
rect 22097 18915 22155 18921
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 25222 18952 25228 18964
rect 25183 18924 25228 18952
rect 25222 18912 25228 18924
rect 25280 18912 25286 18964
rect 3697 18887 3755 18893
rect 3697 18853 3709 18887
rect 3743 18884 3755 18887
rect 3878 18884 3884 18896
rect 3743 18856 3884 18884
rect 3743 18853 3755 18856
rect 3697 18847 3755 18853
rect 3878 18844 3884 18856
rect 3936 18844 3942 18896
rect 4338 18844 4344 18896
rect 4396 18884 4402 18896
rect 4433 18887 4491 18893
rect 4433 18884 4445 18887
rect 4396 18856 4445 18884
rect 4396 18844 4402 18856
rect 4433 18853 4445 18856
rect 4479 18853 4491 18887
rect 4433 18847 4491 18853
rect 7285 18887 7343 18893
rect 7285 18853 7297 18887
rect 7331 18884 7343 18887
rect 7466 18884 7472 18896
rect 7331 18856 7472 18884
rect 7331 18853 7343 18856
rect 7285 18847 7343 18853
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2501 18819 2559 18825
rect 2501 18785 2513 18819
rect 2547 18816 2559 18819
rect 2682 18816 2688 18828
rect 2547 18788 2688 18816
rect 2547 18785 2559 18788
rect 2501 18779 2559 18785
rect 2682 18776 2688 18788
rect 2740 18816 2746 18828
rect 2958 18816 2964 18828
rect 2740 18788 2964 18816
rect 2740 18776 2746 18788
rect 2958 18776 2964 18788
rect 3016 18776 3022 18828
rect 6178 18816 6184 18828
rect 6139 18788 6184 18816
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 6273 18819 6331 18825
rect 6273 18785 6285 18819
rect 6319 18816 6331 18819
rect 6546 18816 6552 18828
rect 6319 18788 6552 18816
rect 6319 18785 6331 18788
rect 6273 18779 6331 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 2038 18748 2044 18760
rect 1999 18720 2044 18748
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 4430 18708 4436 18760
rect 4488 18748 4494 18760
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4488 18720 4537 18748
rect 4488 18708 4494 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18748 6515 18751
rect 7098 18748 7104 18760
rect 6503 18720 7104 18748
rect 6503 18717 6515 18720
rect 6457 18711 6515 18717
rect 3234 18640 3240 18692
rect 3292 18680 3298 18692
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 3292 18652 4077 18680
rect 3292 18640 3298 18652
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4724 18680 4752 18711
rect 5074 18680 5080 18692
rect 4724 18652 5080 18680
rect 4065 18643 4123 18649
rect 5074 18640 5080 18652
rect 5132 18680 5138 18692
rect 5721 18683 5779 18689
rect 5721 18680 5733 18683
rect 5132 18652 5733 18680
rect 5132 18640 5138 18652
rect 5721 18649 5733 18652
rect 5767 18680 5779 18683
rect 6472 18680 6500 18711
rect 7098 18708 7104 18720
rect 7156 18748 7162 18760
rect 7300 18748 7328 18847
rect 7466 18844 7472 18856
rect 7524 18884 7530 18896
rect 8754 18884 8760 18896
rect 7524 18856 7972 18884
rect 8715 18856 8760 18884
rect 7524 18844 7530 18856
rect 7745 18819 7803 18825
rect 7745 18785 7757 18819
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 7156 18720 7328 18748
rect 7156 18708 7162 18720
rect 5767 18652 6500 18680
rect 7760 18680 7788 18779
rect 7944 18757 7972 18856
rect 8754 18844 8760 18856
rect 8812 18844 8818 18896
rect 9674 18844 9680 18896
rect 9732 18884 9738 18896
rect 10873 18887 10931 18893
rect 10873 18884 10885 18887
rect 9732 18856 10885 18884
rect 9732 18844 9738 18856
rect 10873 18853 10885 18856
rect 10919 18853 10931 18887
rect 10873 18847 10931 18853
rect 14185 18887 14243 18893
rect 14185 18853 14197 18887
rect 14231 18884 14243 18887
rect 15286 18884 15292 18896
rect 14231 18856 15292 18884
rect 14231 18853 14243 18856
rect 14185 18847 14243 18853
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 23569 18887 23627 18893
rect 21468 18856 22140 18884
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 9692 18788 10241 18816
rect 9692 18760 9720 18788
rect 10229 18785 10241 18788
rect 10275 18785 10287 18819
rect 10229 18779 10287 18785
rect 10321 18819 10379 18825
rect 10321 18785 10333 18819
rect 10367 18816 10379 18819
rect 10962 18816 10968 18828
rect 10367 18788 10968 18816
rect 10367 18785 10379 18788
rect 10321 18779 10379 18785
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 11681 18819 11739 18825
rect 11681 18816 11693 18819
rect 11204 18788 11693 18816
rect 11204 18776 11210 18788
rect 11681 18785 11693 18788
rect 11727 18816 11739 18819
rect 13906 18816 13912 18828
rect 11727 18788 13912 18816
rect 11727 18785 11739 18788
rect 11681 18779 11739 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 16298 18816 16304 18828
rect 16259 18788 16304 18816
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18816 17463 18819
rect 17451 18788 18184 18816
rect 17451 18785 17463 18788
rect 17405 18779 17463 18785
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18717 7987 18751
rect 7929 18711 7987 18717
rect 9674 18708 9680 18760
rect 9732 18708 9738 18760
rect 9858 18708 9864 18760
rect 9916 18748 9922 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 9916 18720 10425 18748
rect 9916 18708 9922 18720
rect 10413 18717 10425 18720
rect 10459 18748 10471 18751
rect 11054 18748 11060 18760
rect 10459 18720 11060 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 11238 18748 11244 18760
rect 11199 18720 11244 18748
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 11422 18748 11428 18760
rect 11383 18720 11428 18748
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 16264 18720 16405 18748
rect 16264 18708 16270 18720
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 16485 18751 16543 18757
rect 16485 18717 16497 18751
rect 16531 18748 16543 18751
rect 16574 18748 16580 18760
rect 16531 18720 16580 18748
rect 16531 18717 16543 18720
rect 16485 18711 16543 18717
rect 16574 18708 16580 18720
rect 16632 18708 16638 18760
rect 18156 18757 18184 18788
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19116 18788 19441 18816
rect 19116 18776 19122 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 19429 18779 19487 18785
rect 21358 18776 21364 18828
rect 21416 18816 21422 18828
rect 21468 18825 21496 18856
rect 21453 18819 21511 18825
rect 21453 18816 21465 18819
rect 21416 18788 21465 18816
rect 21416 18776 21422 18788
rect 21453 18785 21465 18788
rect 21499 18785 21511 18819
rect 21453 18779 21511 18785
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 22005 18819 22063 18825
rect 22005 18816 22017 18819
rect 21876 18788 22017 18816
rect 21876 18776 21882 18788
rect 22005 18785 22017 18788
rect 22051 18785 22063 18819
rect 22112 18816 22140 18856
rect 23569 18853 23581 18887
rect 23615 18884 23627 18887
rect 23750 18884 23756 18896
rect 23615 18856 23756 18884
rect 23615 18853 23627 18856
rect 23569 18847 23627 18853
rect 23750 18844 23756 18856
rect 23808 18884 23814 18896
rect 25777 18887 25835 18893
rect 25777 18884 25789 18887
rect 23808 18856 25789 18884
rect 23808 18844 23814 18856
rect 25777 18853 25789 18856
rect 25823 18853 25835 18887
rect 25777 18847 25835 18853
rect 23109 18819 23167 18825
rect 22112 18788 22324 18816
rect 22005 18779 22063 18785
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 17083 18720 17969 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17957 18717 17969 18720
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18748 18199 18751
rect 18598 18748 18604 18760
rect 18187 18720 18604 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 8018 18680 8024 18692
rect 7760 18652 8024 18680
rect 5767 18649 5779 18652
rect 5721 18643 5779 18649
rect 8018 18640 8024 18652
rect 8076 18640 8082 18692
rect 9490 18680 9496 18692
rect 9451 18652 9496 18680
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 15933 18683 15991 18689
rect 15933 18649 15945 18683
rect 15979 18680 15991 18683
rect 17052 18680 17080 18711
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 19518 18748 19524 18760
rect 19479 18720 19524 18748
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 21174 18748 21180 18760
rect 21087 18720 21180 18748
rect 19613 18711 19671 18717
rect 15979 18652 17080 18680
rect 15979 18649 15991 18652
rect 15933 18643 15991 18649
rect 19426 18640 19432 18692
rect 19484 18680 19490 18692
rect 19628 18680 19656 18711
rect 21174 18708 21180 18720
rect 21232 18748 21238 18760
rect 21910 18748 21916 18760
rect 21232 18720 21916 18748
rect 21232 18708 21238 18720
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22296 18757 22324 18788
rect 23109 18785 23121 18819
rect 23155 18816 23167 18819
rect 23290 18816 23296 18828
rect 23155 18788 23296 18816
rect 23155 18785 23167 18788
rect 23109 18779 23167 18785
rect 23290 18776 23296 18788
rect 23348 18816 23354 18828
rect 23348 18788 24900 18816
rect 23348 18776 23354 18788
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18717 22339 18751
rect 23658 18748 23664 18760
rect 23619 18720 23664 18748
rect 22281 18711 22339 18717
rect 23658 18708 23664 18720
rect 23716 18708 23722 18760
rect 23842 18748 23848 18760
rect 23803 18720 23848 18748
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 24872 18748 24900 18788
rect 24946 18776 24952 18828
rect 25004 18816 25010 18828
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 25004 18788 25145 18816
rect 25004 18776 25010 18788
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 25409 18751 25467 18757
rect 25409 18748 25421 18751
rect 24872 18720 25421 18748
rect 25409 18717 25421 18720
rect 25455 18748 25467 18751
rect 25774 18748 25780 18760
rect 25455 18720 25780 18748
rect 25455 18717 25467 18720
rect 25409 18711 25467 18717
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 19484 18652 19656 18680
rect 20717 18683 20775 18689
rect 19484 18640 19490 18652
rect 20717 18649 20729 18683
rect 20763 18680 20775 18683
rect 21634 18680 21640 18692
rect 20763 18652 21640 18680
rect 20763 18649 20775 18652
rect 20717 18643 20775 18649
rect 21634 18640 21640 18652
rect 21692 18640 21698 18692
rect 22738 18640 22744 18692
rect 22796 18680 22802 18692
rect 23201 18683 23259 18689
rect 23201 18680 23213 18683
rect 22796 18652 23213 18680
rect 22796 18640 22802 18652
rect 23201 18649 23213 18652
rect 23247 18649 23259 18683
rect 23201 18643 23259 18649
rect 23382 18640 23388 18692
rect 23440 18680 23446 18692
rect 23860 18680 23888 18708
rect 24302 18680 24308 18692
rect 23440 18652 23888 18680
rect 24044 18652 24308 18680
rect 23440 18640 23446 18652
rect 1397 18615 1455 18621
rect 1397 18581 1409 18615
rect 1443 18612 1455 18615
rect 2130 18612 2136 18624
rect 1443 18584 2136 18612
rect 1443 18581 1455 18584
rect 1397 18575 1455 18581
rect 2130 18572 2136 18584
rect 2188 18572 2194 18624
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7006 18612 7012 18624
rect 6963 18584 7012 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7006 18572 7012 18584
rect 7064 18612 7070 18624
rect 7282 18612 7288 18624
rect 7064 18584 7288 18612
rect 7064 18572 7070 18584
rect 7282 18572 7288 18584
rect 7340 18572 7346 18624
rect 8481 18615 8539 18621
rect 8481 18581 8493 18615
rect 8527 18612 8539 18615
rect 8662 18612 8668 18624
rect 8527 18584 8668 18612
rect 8527 18581 8539 18584
rect 8481 18575 8539 18581
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 12805 18615 12863 18621
rect 12805 18612 12817 18615
rect 12124 18584 12817 18612
rect 12124 18572 12130 18584
rect 12805 18581 12817 18584
rect 12851 18581 12863 18615
rect 13814 18612 13820 18624
rect 13775 18584 13820 18612
rect 12805 18575 12863 18581
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 15470 18612 15476 18624
rect 15431 18584 15476 18612
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 18877 18615 18935 18621
rect 18877 18612 18889 18615
rect 18656 18584 18889 18612
rect 18656 18572 18662 18584
rect 18877 18581 18889 18584
rect 18923 18581 18935 18615
rect 20162 18612 20168 18624
rect 20123 18584 20168 18612
rect 18877 18575 18935 18581
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 22554 18572 22560 18624
rect 22612 18612 22618 18624
rect 22649 18615 22707 18621
rect 22649 18612 22661 18615
rect 22612 18584 22661 18612
rect 22612 18572 22618 18584
rect 22649 18581 22661 18584
rect 22695 18581 22707 18615
rect 22649 18575 22707 18581
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24044 18612 24072 18652
rect 24302 18640 24308 18652
rect 24360 18640 24366 18692
rect 24673 18683 24731 18689
rect 24673 18649 24685 18683
rect 24719 18680 24731 18683
rect 25130 18680 25136 18692
rect 24719 18652 25136 18680
rect 24719 18649 24731 18652
rect 24673 18643 24731 18649
rect 25130 18640 25136 18652
rect 25188 18640 25194 18692
rect 24210 18612 24216 18624
rect 23900 18584 24072 18612
rect 24171 18584 24216 18612
rect 23900 18572 23906 18584
rect 24210 18572 24216 18584
rect 24268 18572 24274 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 4525 18411 4583 18417
rect 4525 18408 4537 18411
rect 4120 18380 4537 18408
rect 4120 18368 4126 18380
rect 4525 18377 4537 18380
rect 4571 18408 4583 18411
rect 5074 18408 5080 18420
rect 4571 18380 5080 18408
rect 4571 18377 4583 18380
rect 4525 18371 4583 18377
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 7837 18411 7895 18417
rect 7837 18377 7849 18411
rect 7883 18408 7895 18411
rect 9582 18408 9588 18420
rect 7883 18380 9588 18408
rect 7883 18377 7895 18380
rect 7837 18371 7895 18377
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 12526 18408 12532 18420
rect 12483 18380 12532 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 12526 18368 12532 18380
rect 12584 18368 12590 18420
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 13688 18380 14105 18408
rect 13688 18368 13694 18380
rect 14093 18377 14105 18380
rect 14139 18377 14151 18411
rect 17402 18408 17408 18420
rect 17363 18380 17408 18408
rect 14093 18371 14151 18377
rect 5537 18343 5595 18349
rect 5537 18309 5549 18343
rect 5583 18340 5595 18343
rect 6546 18340 6552 18352
rect 5583 18312 6552 18340
rect 5583 18309 5595 18312
rect 5537 18303 5595 18309
rect 6546 18300 6552 18312
rect 6604 18300 6610 18352
rect 12253 18343 12311 18349
rect 12253 18309 12265 18343
rect 12299 18340 12311 18343
rect 12710 18340 12716 18352
rect 12299 18312 12716 18340
rect 12299 18309 12311 18312
rect 12253 18303 12311 18309
rect 12710 18300 12716 18312
rect 12768 18300 12774 18352
rect 1946 18272 1952 18284
rect 1907 18244 1952 18272
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2593 18275 2651 18281
rect 2593 18272 2605 18275
rect 2179 18244 2605 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2593 18241 2605 18244
rect 2639 18272 2651 18275
rect 2639 18244 3280 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 3145 18207 3203 18213
rect 3145 18204 3157 18207
rect 2976 18176 3157 18204
rect 1946 18136 1952 18148
rect 1504 18108 1952 18136
rect 1504 18077 1532 18108
rect 1946 18096 1952 18108
rect 2004 18096 2010 18148
rect 1489 18071 1547 18077
rect 1489 18037 1501 18071
rect 1535 18037 1547 18071
rect 1489 18031 1547 18037
rect 1857 18071 1915 18077
rect 1857 18037 1869 18071
rect 1903 18068 1915 18071
rect 2130 18068 2136 18080
rect 1903 18040 2136 18068
rect 1903 18037 1915 18040
rect 1857 18031 1915 18037
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 2774 18028 2780 18080
rect 2832 18068 2838 18080
rect 2976 18077 3004 18176
rect 3145 18173 3157 18176
rect 3191 18173 3203 18207
rect 3252 18204 3280 18244
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 5077 18275 5135 18281
rect 5077 18272 5089 18275
rect 4212 18244 5089 18272
rect 4212 18232 4218 18244
rect 5077 18241 5089 18244
rect 5123 18272 5135 18275
rect 6178 18272 6184 18284
rect 5123 18244 6184 18272
rect 5123 18241 5135 18244
rect 5077 18235 5135 18241
rect 6178 18232 6184 18244
rect 6236 18232 6242 18284
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 7834 18272 7840 18284
rect 6687 18244 7840 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8481 18275 8539 18281
rect 8481 18241 8493 18275
rect 8527 18272 8539 18275
rect 8662 18272 8668 18284
rect 8527 18244 8668 18272
rect 8527 18241 8539 18244
rect 8481 18235 8539 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 13081 18275 13139 18281
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 13449 18275 13507 18281
rect 13449 18272 13461 18275
rect 13127 18244 13461 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13449 18241 13461 18244
rect 13495 18272 13507 18275
rect 13722 18272 13728 18284
rect 13495 18244 13728 18272
rect 13495 18241 13507 18244
rect 13449 18235 13507 18241
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14108 18272 14136 18371
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 17770 18368 17776 18420
rect 17828 18408 17834 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17828 18380 18061 18408
rect 17828 18368 17834 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 21726 18408 21732 18420
rect 21687 18380 21732 18408
rect 18049 18371 18107 18377
rect 21726 18368 21732 18380
rect 21784 18368 21790 18420
rect 23474 18408 23480 18420
rect 23435 18380 23480 18408
rect 23474 18368 23480 18380
rect 23532 18408 23538 18420
rect 24857 18411 24915 18417
rect 23532 18380 24164 18408
rect 23532 18368 23538 18380
rect 19981 18343 20039 18349
rect 19981 18309 19993 18343
rect 20027 18340 20039 18343
rect 21361 18343 21419 18349
rect 20027 18312 20668 18340
rect 20027 18309 20039 18312
rect 19981 18303 20039 18309
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 14108 18244 14289 18272
rect 14277 18241 14289 18244
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 16666 18232 16672 18284
rect 16724 18272 16730 18284
rect 16945 18275 17003 18281
rect 16945 18272 16957 18275
rect 16724 18244 16957 18272
rect 16724 18232 16730 18244
rect 16945 18241 16957 18244
rect 16991 18241 17003 18275
rect 18598 18272 18604 18284
rect 18559 18244 18604 18272
rect 16945 18235 17003 18241
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 20162 18232 20168 18284
rect 20220 18272 20226 18284
rect 20640 18281 20668 18312
rect 21361 18309 21373 18343
rect 21407 18340 21419 18343
rect 21818 18340 21824 18352
rect 21407 18312 21824 18340
rect 21407 18309 21419 18312
rect 21361 18303 21419 18309
rect 21818 18300 21824 18312
rect 21876 18300 21882 18352
rect 20533 18275 20591 18281
rect 20533 18272 20545 18275
rect 20220 18244 20545 18272
rect 20220 18232 20226 18244
rect 20533 18241 20545 18244
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18272 20683 18275
rect 21174 18272 21180 18284
rect 20671 18244 21180 18272
rect 20671 18241 20683 18244
rect 20625 18235 20683 18241
rect 3418 18213 3424 18216
rect 3401 18207 3424 18213
rect 3401 18204 3413 18207
rect 3252 18176 3413 18204
rect 3145 18167 3203 18173
rect 3401 18173 3413 18176
rect 3476 18204 3482 18216
rect 5629 18207 5687 18213
rect 3476 18176 3549 18204
rect 3401 18167 3424 18173
rect 3418 18164 3424 18167
rect 3476 18164 3482 18176
rect 5629 18173 5641 18207
rect 5675 18204 5687 18207
rect 5994 18204 6000 18216
rect 5675 18176 6000 18204
rect 5675 18173 5687 18176
rect 5629 18167 5687 18173
rect 5994 18164 6000 18176
rect 6052 18204 6058 18216
rect 6052 18176 6316 18204
rect 6052 18164 6058 18176
rect 2961 18071 3019 18077
rect 2961 18068 2973 18071
rect 2832 18040 2973 18068
rect 2832 18028 2838 18040
rect 2961 18037 2973 18040
rect 3007 18037 3019 18071
rect 5810 18068 5816 18080
rect 5771 18040 5816 18068
rect 2961 18031 3019 18037
rect 5810 18028 5816 18040
rect 5868 18028 5874 18080
rect 6288 18077 6316 18176
rect 7374 18164 7380 18216
rect 7432 18204 7438 18216
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 7432 18176 8309 18204
rect 7432 18164 7438 18176
rect 8297 18173 8309 18176
rect 8343 18204 8355 18207
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 8343 18176 8861 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 8849 18173 8861 18176
rect 8895 18173 8907 18207
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 8849 18167 8907 18173
rect 8956 18176 9413 18204
rect 6914 18096 6920 18148
rect 6972 18136 6978 18148
rect 6972 18108 8248 18136
rect 6972 18096 6978 18108
rect 8220 18080 8248 18108
rect 6273 18071 6331 18077
rect 6273 18037 6285 18071
rect 6319 18068 6331 18071
rect 6362 18068 6368 18080
rect 6319 18040 6368 18068
rect 6319 18037 6331 18040
rect 6273 18031 6331 18037
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 6638 18028 6644 18080
rect 6696 18068 6702 18080
rect 6825 18071 6883 18077
rect 6825 18068 6837 18071
rect 6696 18040 6837 18068
rect 6696 18028 6702 18040
rect 6825 18037 6837 18040
rect 6871 18037 6883 18071
rect 6825 18031 6883 18037
rect 7469 18071 7527 18077
rect 7469 18037 7481 18071
rect 7515 18068 7527 18071
rect 8018 18068 8024 18080
rect 7515 18040 8024 18068
rect 7515 18037 7527 18040
rect 7469 18031 7527 18037
rect 8018 18028 8024 18040
rect 8076 18028 8082 18080
rect 8202 18068 8208 18080
rect 8163 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 8956 18068 8984 18176
rect 9401 18173 9413 18176
rect 9447 18173 9459 18207
rect 9401 18167 9459 18173
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 9657 18207 9715 18213
rect 9657 18204 9669 18207
rect 9548 18176 9669 18204
rect 9548 18164 9554 18176
rect 9657 18173 9669 18176
rect 9703 18173 9715 18207
rect 9657 18167 9715 18173
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10192 18176 11928 18204
rect 10192 18164 10198 18176
rect 9030 18096 9036 18148
rect 9088 18136 9094 18148
rect 11793 18139 11851 18145
rect 11793 18136 11805 18139
rect 9088 18108 11805 18136
rect 9088 18096 9094 18108
rect 11793 18105 11805 18108
rect 11839 18105 11851 18139
rect 11900 18136 11928 18176
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 14550 18213 14556 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12768 18176 12817 18204
rect 12768 18164 12774 18176
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 14544 18204 14556 18213
rect 14511 18176 14556 18204
rect 12805 18167 12863 18173
rect 14544 18167 14556 18176
rect 14550 18164 14556 18167
rect 14608 18164 14614 18216
rect 15654 18204 15660 18216
rect 14660 18176 15660 18204
rect 14660 18136 14688 18176
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 17460 18176 18429 18204
rect 17460 18164 17466 18176
rect 18417 18173 18429 18176
rect 18463 18173 18475 18207
rect 20548 18204 20576 18235
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 22370 18272 22376 18284
rect 22331 18244 22376 18272
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 22554 18272 22560 18284
rect 22515 18244 22560 18272
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 24136 18281 24164 18380
rect 24857 18377 24869 18411
rect 24903 18408 24915 18411
rect 25222 18408 25228 18420
rect 24903 18380 25228 18408
rect 24903 18377 24915 18380
rect 24857 18371 24915 18377
rect 25222 18368 25228 18380
rect 25280 18368 25286 18420
rect 25409 18411 25467 18417
rect 25409 18377 25421 18411
rect 25455 18408 25467 18411
rect 25498 18408 25504 18420
rect 25455 18380 25504 18408
rect 25455 18377 25467 18380
rect 25409 18371 25467 18377
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 25774 18408 25780 18420
rect 25735 18380 25780 18408
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 26234 18408 26240 18420
rect 26195 18380 26240 18408
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24210 18232 24216 18284
rect 24268 18272 24274 18284
rect 24268 18244 24361 18272
rect 24268 18232 24274 18244
rect 20714 18204 20720 18216
rect 20548 18176 20720 18204
rect 18417 18167 18475 18173
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 21634 18164 21640 18216
rect 21692 18204 21698 18216
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 21692 18176 22293 18204
rect 21692 18164 21698 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22572 18204 22600 18232
rect 23106 18204 23112 18216
rect 22572 18176 23112 18204
rect 22281 18167 22339 18173
rect 23106 18164 23112 18176
rect 23164 18204 23170 18216
rect 24228 18204 24256 18232
rect 25222 18204 25228 18216
rect 23164 18176 24256 18204
rect 25183 18176 25228 18204
rect 23164 18164 23170 18176
rect 25222 18164 25228 18176
rect 25280 18164 25286 18216
rect 11900 18108 14688 18136
rect 11793 18099 11851 18105
rect 9217 18071 9275 18077
rect 9217 18068 9229 18071
rect 8628 18040 9229 18068
rect 8628 18028 8634 18040
rect 9217 18037 9229 18040
rect 9263 18037 9275 18071
rect 9217 18031 9275 18037
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 10100 18040 10793 18068
rect 10100 18028 10106 18040
rect 10781 18037 10793 18040
rect 10827 18037 10839 18071
rect 11514 18068 11520 18080
rect 11475 18040 11520 18068
rect 10781 18031 10839 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 11808 18068 11836 18099
rect 15286 18096 15292 18148
rect 15344 18136 15350 18148
rect 16206 18136 16212 18148
rect 15344 18108 16212 18136
rect 15344 18096 15350 18108
rect 16206 18096 16212 18108
rect 16264 18136 16270 18148
rect 16577 18139 16635 18145
rect 16577 18136 16589 18139
rect 16264 18108 16589 18136
rect 16264 18096 16270 18108
rect 16577 18105 16589 18108
rect 16623 18105 16635 18139
rect 16577 18099 16635 18105
rect 18322 18096 18328 18148
rect 18380 18136 18386 18148
rect 19058 18136 19064 18148
rect 18380 18108 19064 18136
rect 18380 18096 18386 18108
rect 19058 18096 19064 18108
rect 19116 18136 19122 18148
rect 20162 18136 20168 18148
rect 19116 18108 20168 18136
rect 19116 18096 19122 18108
rect 20162 18096 20168 18108
rect 20220 18096 20226 18148
rect 22922 18096 22928 18148
rect 22980 18136 22986 18148
rect 23017 18139 23075 18145
rect 23017 18136 23029 18139
rect 22980 18108 23029 18136
rect 22980 18096 22986 18108
rect 23017 18105 23029 18108
rect 23063 18136 23075 18139
rect 23842 18136 23848 18148
rect 23063 18108 23848 18136
rect 23063 18105 23075 18108
rect 23017 18099 23075 18105
rect 23842 18096 23848 18108
rect 23900 18136 23906 18148
rect 24029 18139 24087 18145
rect 24029 18136 24041 18139
rect 23900 18108 24041 18136
rect 23900 18096 23906 18108
rect 24029 18105 24041 18108
rect 24075 18105 24087 18139
rect 24029 18099 24087 18105
rect 12897 18071 12955 18077
rect 12897 18068 12909 18071
rect 11808 18040 12909 18068
rect 12897 18037 12909 18040
rect 12943 18037 12955 18071
rect 12897 18031 12955 18037
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 13964 18040 15669 18068
rect 13964 18028 13970 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 16298 18068 16304 18080
rect 16259 18040 16304 18068
rect 15657 18031 15715 18037
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 17310 18028 17316 18080
rect 17368 18068 17374 18080
rect 17773 18071 17831 18077
rect 17773 18068 17785 18071
rect 17368 18040 17785 18068
rect 17368 18028 17374 18040
rect 17773 18037 17785 18040
rect 17819 18068 17831 18071
rect 18506 18068 18512 18080
rect 17819 18040 18512 18068
rect 17819 18037 17831 18040
rect 17773 18031 17831 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 19518 18068 19524 18080
rect 19479 18040 19524 18068
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 20073 18071 20131 18077
rect 20073 18037 20085 18071
rect 20119 18068 20131 18071
rect 20254 18068 20260 18080
rect 20119 18040 20260 18068
rect 20119 18037 20131 18040
rect 20073 18031 20131 18037
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 20438 18068 20444 18080
rect 20399 18040 20444 18068
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 21358 18028 21364 18080
rect 21416 18068 21422 18080
rect 21634 18068 21640 18080
rect 21416 18040 21640 18068
rect 21416 18028 21422 18040
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 21913 18071 21971 18077
rect 21913 18037 21925 18071
rect 21959 18068 21971 18071
rect 22002 18068 22008 18080
rect 21959 18040 22008 18068
rect 21959 18037 21971 18040
rect 21913 18031 21971 18037
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 23658 18068 23664 18080
rect 23619 18040 23664 18068
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2866 17864 2872 17876
rect 2096 17836 2872 17864
rect 2096 17824 2102 17836
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 4062 17864 4068 17876
rect 3927 17836 4068 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4617 17867 4675 17873
rect 4617 17864 4629 17867
rect 4396 17836 4629 17864
rect 4396 17824 4402 17836
rect 4617 17833 4629 17836
rect 4663 17833 4675 17867
rect 6730 17864 6736 17876
rect 6691 17836 6736 17864
rect 4617 17827 4675 17833
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 7098 17864 7104 17876
rect 7059 17836 7104 17864
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 8202 17824 8208 17876
rect 8260 17864 8266 17876
rect 8297 17867 8355 17873
rect 8297 17864 8309 17867
rect 8260 17836 8309 17864
rect 8260 17824 8266 17836
rect 8297 17833 8309 17836
rect 8343 17833 8355 17867
rect 8297 17827 8355 17833
rect 9125 17867 9183 17873
rect 9125 17833 9137 17867
rect 9171 17864 9183 17867
rect 9306 17864 9312 17876
rect 9171 17836 9312 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 10778 17864 10784 17876
rect 10739 17836 10784 17864
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 12805 17867 12863 17873
rect 12805 17864 12817 17867
rect 12492 17836 12817 17864
rect 12492 17824 12498 17836
rect 12805 17833 12817 17836
rect 12851 17833 12863 17867
rect 12805 17827 12863 17833
rect 13817 17867 13875 17873
rect 13817 17833 13829 17867
rect 13863 17864 13875 17867
rect 13998 17864 14004 17876
rect 13863 17836 14004 17864
rect 13863 17833 13875 17836
rect 13817 17827 13875 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 14550 17824 14556 17876
rect 14608 17864 14614 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14608 17836 14657 17864
rect 14608 17824 14614 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 16574 17824 16580 17876
rect 16632 17864 16638 17876
rect 16761 17867 16819 17873
rect 16761 17864 16773 17867
rect 16632 17836 16773 17864
rect 16632 17824 16638 17836
rect 16761 17833 16773 17836
rect 16807 17864 16819 17867
rect 18325 17867 18383 17873
rect 18325 17864 18337 17867
rect 16807 17836 18337 17864
rect 16807 17833 16819 17836
rect 16761 17827 16819 17833
rect 18325 17833 18337 17836
rect 18371 17864 18383 17867
rect 18598 17864 18604 17876
rect 18371 17836 18604 17864
rect 18371 17833 18383 17836
rect 18325 17827 18383 17833
rect 18598 17824 18604 17836
rect 18656 17864 18662 17876
rect 18877 17867 18935 17873
rect 18877 17864 18889 17867
rect 18656 17836 18889 17864
rect 18656 17824 18662 17836
rect 18877 17833 18889 17836
rect 18923 17833 18935 17867
rect 18877 17827 18935 17833
rect 19337 17867 19395 17873
rect 19337 17833 19349 17867
rect 19383 17864 19395 17867
rect 19426 17864 19432 17876
rect 19383 17836 19432 17864
rect 19383 17833 19395 17836
rect 19337 17827 19395 17833
rect 19426 17824 19432 17836
rect 19484 17824 19490 17876
rect 19889 17867 19947 17873
rect 19889 17833 19901 17867
rect 19935 17864 19947 17867
rect 20070 17864 20076 17876
rect 19935 17836 20076 17864
rect 19935 17833 19947 17836
rect 19889 17827 19947 17833
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22281 17867 22339 17873
rect 22281 17864 22293 17867
rect 22244 17836 22293 17864
rect 22244 17824 22250 17836
rect 22281 17833 22293 17836
rect 22327 17833 22339 17867
rect 22281 17827 22339 17833
rect 22370 17824 22376 17876
rect 22428 17864 22434 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 22428 17836 22845 17864
rect 22428 17824 22434 17836
rect 22833 17833 22845 17836
rect 22879 17833 22891 17867
rect 22833 17827 22891 17833
rect 23293 17867 23351 17873
rect 23293 17833 23305 17867
rect 23339 17864 23351 17867
rect 23382 17864 23388 17876
rect 23339 17836 23388 17864
rect 23339 17833 23351 17836
rect 23293 17827 23351 17833
rect 23382 17824 23388 17836
rect 23440 17824 23446 17876
rect 1486 17756 1492 17808
rect 1544 17756 1550 17808
rect 7282 17756 7288 17808
rect 7340 17796 7346 17808
rect 7745 17799 7803 17805
rect 7745 17796 7757 17799
rect 7340 17768 7757 17796
rect 7340 17756 7346 17768
rect 7745 17765 7757 17768
rect 7791 17765 7803 17799
rect 7745 17759 7803 17765
rect 11054 17756 11060 17808
rect 11112 17796 11118 17808
rect 11670 17799 11728 17805
rect 11670 17796 11682 17799
rect 11112 17768 11682 17796
rect 11112 17756 11118 17768
rect 11670 17765 11682 17768
rect 11716 17796 11728 17799
rect 12066 17796 12072 17808
rect 11716 17768 12072 17796
rect 11716 17765 11728 17768
rect 11670 17759 11728 17765
rect 12066 17756 12072 17768
rect 12124 17756 12130 17808
rect 12158 17756 12164 17808
rect 12216 17796 12222 17808
rect 13357 17799 13415 17805
rect 13357 17796 13369 17799
rect 12216 17768 13369 17796
rect 12216 17756 12222 17768
rect 13357 17765 13369 17768
rect 13403 17765 13415 17799
rect 13357 17759 13415 17765
rect 14182 17756 14188 17808
rect 14240 17796 14246 17808
rect 16485 17799 16543 17805
rect 14240 17768 16335 17796
rect 14240 17756 14246 17768
rect 1504 17728 1532 17756
rect 1756 17731 1814 17737
rect 1756 17728 1768 17731
rect 1504 17700 1768 17728
rect 1756 17697 1768 17700
rect 1802 17728 1814 17731
rect 2222 17728 2228 17740
rect 1802 17700 2228 17728
rect 1802 17697 1814 17700
rect 1756 17691 1814 17697
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 5074 17737 5080 17740
rect 5068 17728 5080 17737
rect 5035 17700 5080 17728
rect 5068 17691 5080 17700
rect 5074 17688 5080 17691
rect 5132 17688 5138 17740
rect 7650 17728 7656 17740
rect 7611 17700 7656 17728
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9180 17700 10057 17728
rect 9180 17688 9186 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 11425 17731 11483 17737
rect 11425 17697 11437 17731
rect 11471 17728 11483 17731
rect 11514 17728 11520 17740
rect 11471 17700 11520 17728
rect 11471 17697 11483 17700
rect 11425 17691 11483 17697
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 15654 17688 15660 17740
rect 15712 17728 15718 17740
rect 15749 17731 15807 17737
rect 15749 17728 15761 17731
rect 15712 17700 15761 17728
rect 15712 17688 15718 17700
rect 15749 17697 15761 17700
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 15841 17731 15899 17737
rect 15841 17697 15853 17731
rect 15887 17728 15899 17731
rect 16114 17728 16120 17740
rect 15887 17700 16120 17728
rect 15887 17697 15899 17700
rect 15841 17691 15899 17697
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 16307 17728 16335 17768
rect 16485 17765 16497 17799
rect 16531 17796 16543 17799
rect 17034 17796 17040 17808
rect 16531 17768 17040 17796
rect 16531 17765 16543 17768
rect 16485 17759 16543 17765
rect 17034 17756 17040 17768
rect 17092 17796 17098 17808
rect 17190 17799 17248 17805
rect 17190 17796 17202 17799
rect 17092 17768 17202 17796
rect 17092 17756 17098 17768
rect 17190 17765 17202 17768
rect 17236 17765 17248 17799
rect 17190 17759 17248 17765
rect 20717 17799 20775 17805
rect 20717 17765 20729 17799
rect 20763 17796 20775 17799
rect 21168 17799 21226 17805
rect 21168 17796 21180 17799
rect 20763 17768 21180 17796
rect 20763 17765 20775 17768
rect 20717 17759 20775 17765
rect 21168 17765 21180 17768
rect 21214 17796 21226 17799
rect 21450 17796 21456 17808
rect 21214 17768 21456 17796
rect 21214 17765 21226 17768
rect 21168 17759 21226 17765
rect 21450 17756 21456 17768
rect 21508 17796 21514 17808
rect 22462 17796 22468 17808
rect 21508 17768 22468 17796
rect 21508 17756 21514 17768
rect 22462 17756 22468 17768
rect 22520 17756 22526 17808
rect 18138 17728 18144 17740
rect 16307 17700 18144 17728
rect 18138 17688 18144 17700
rect 18196 17688 18202 17740
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19484 17700 19717 17728
rect 19484 17688 19490 17700
rect 19705 17697 19717 17700
rect 19751 17728 19763 17731
rect 19978 17728 19984 17740
rect 19751 17700 19984 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 22554 17688 22560 17740
rect 22612 17728 22618 17740
rect 23658 17728 23664 17740
rect 22612 17700 23664 17728
rect 22612 17688 22618 17700
rect 23658 17688 23664 17700
rect 23716 17728 23722 17740
rect 23753 17731 23811 17737
rect 23753 17728 23765 17731
rect 23716 17700 23765 17728
rect 23716 17688 23722 17700
rect 23753 17697 23765 17700
rect 23799 17697 23811 17731
rect 23753 17691 23811 17697
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17728 25007 17731
rect 25314 17728 25320 17740
rect 24995 17700 25320 17728
rect 24995 17697 25007 17700
rect 24949 17691 25007 17697
rect 25314 17688 25320 17700
rect 25372 17688 25378 17740
rect 1486 17660 1492 17672
rect 1447 17632 1492 17660
rect 1486 17620 1492 17632
rect 1544 17620 1550 17672
rect 4798 17660 4804 17672
rect 4759 17632 4804 17660
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 6822 17620 6828 17672
rect 6880 17660 6886 17672
rect 7742 17660 7748 17672
rect 6880 17632 7748 17660
rect 6880 17620 6886 17632
rect 7742 17620 7748 17632
rect 7800 17660 7806 17672
rect 7837 17663 7895 17669
rect 7837 17660 7849 17663
rect 7800 17632 7849 17660
rect 7800 17620 7806 17632
rect 7837 17629 7849 17632
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 10137 17663 10195 17669
rect 10137 17629 10149 17663
rect 10183 17660 10195 17663
rect 10226 17660 10232 17672
rect 10183 17632 10232 17660
rect 10183 17629 10195 17632
rect 10137 17623 10195 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 11330 17660 11336 17672
rect 10367 17632 11336 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 14182 17660 14188 17672
rect 14143 17632 14188 17660
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 15102 17660 15108 17672
rect 15063 17632 15108 17660
rect 15102 17620 15108 17632
rect 15160 17620 15166 17672
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17660 16083 17663
rect 16574 17660 16580 17672
rect 16071 17632 16580 17660
rect 16071 17629 16083 17632
rect 16025 17623 16083 17629
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17629 17003 17663
rect 20898 17660 20904 17672
rect 20859 17632 20904 17660
rect 16945 17623 17003 17629
rect 15746 17552 15752 17604
rect 15804 17592 15810 17604
rect 16850 17592 16856 17604
rect 15804 17564 16856 17592
rect 15804 17552 15810 17564
rect 16850 17552 16856 17564
rect 16908 17592 16914 17604
rect 16960 17592 16988 17623
rect 20898 17620 20904 17632
rect 20956 17620 20962 17672
rect 22094 17620 22100 17672
rect 22152 17660 22158 17672
rect 22922 17660 22928 17672
rect 22152 17632 22928 17660
rect 22152 17620 22158 17632
rect 22922 17620 22928 17632
rect 22980 17660 22986 17672
rect 23845 17663 23903 17669
rect 23845 17660 23857 17663
rect 22980 17632 23857 17660
rect 22980 17620 22986 17632
rect 23845 17629 23857 17632
rect 23891 17629 23903 17663
rect 23845 17623 23903 17629
rect 24029 17663 24087 17669
rect 24029 17629 24041 17663
rect 24075 17660 24087 17663
rect 24075 17632 24256 17660
rect 24075 17629 24087 17632
rect 24029 17623 24087 17629
rect 16908 17564 16988 17592
rect 16908 17552 16914 17564
rect 24228 17536 24256 17632
rect 2866 17524 2872 17536
rect 2827 17496 2872 17524
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4430 17524 4436 17536
rect 4387 17496 4436 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 6178 17524 6184 17536
rect 6139 17496 6184 17524
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 7285 17527 7343 17533
rect 7285 17524 7297 17527
rect 6972 17496 7297 17524
rect 6972 17484 6978 17496
rect 7285 17493 7297 17496
rect 7331 17493 7343 17527
rect 7285 17487 7343 17493
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 8665 17527 8723 17533
rect 8665 17524 8677 17527
rect 8628 17496 8677 17524
rect 8628 17484 8634 17496
rect 8665 17493 8677 17496
rect 8711 17493 8723 17527
rect 9398 17524 9404 17536
rect 9359 17496 9404 17524
rect 8665 17487 8723 17493
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9674 17524 9680 17536
rect 9635 17496 9680 17524
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 11204 17496 11253 17524
rect 11204 17484 11210 17496
rect 11241 17493 11253 17496
rect 11287 17493 11299 17527
rect 15378 17524 15384 17536
rect 15339 17496 15384 17524
rect 11241 17487 11299 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 20346 17524 20352 17536
rect 20307 17496 20352 17524
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 23198 17484 23204 17536
rect 23256 17524 23262 17536
rect 23385 17527 23443 17533
rect 23385 17524 23397 17527
rect 23256 17496 23397 17524
rect 23256 17484 23262 17496
rect 23385 17493 23397 17496
rect 23431 17493 23443 17527
rect 23385 17487 23443 17493
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 24268 17496 24409 17524
rect 24268 17484 24274 17496
rect 24397 17493 24409 17496
rect 24443 17493 24455 17527
rect 24397 17487 24455 17493
rect 24857 17527 24915 17533
rect 24857 17493 24869 17527
rect 24903 17524 24915 17527
rect 24946 17524 24952 17536
rect 24903 17496 24952 17524
rect 24903 17493 24915 17496
rect 24857 17487 24915 17493
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 25130 17524 25136 17536
rect 25091 17496 25136 17524
rect 25130 17484 25136 17496
rect 25188 17484 25194 17536
rect 25222 17484 25228 17536
rect 25280 17524 25286 17536
rect 25593 17527 25651 17533
rect 25593 17524 25605 17527
rect 25280 17496 25605 17524
rect 25280 17484 25286 17496
rect 25593 17493 25605 17496
rect 25639 17524 25651 17527
rect 25958 17524 25964 17536
rect 25639 17496 25964 17524
rect 25639 17493 25651 17496
rect 25593 17487 25651 17493
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1486 17280 1492 17332
rect 1544 17320 1550 17332
rect 1857 17323 1915 17329
rect 1857 17320 1869 17323
rect 1544 17292 1869 17320
rect 1544 17280 1550 17292
rect 1857 17289 1869 17292
rect 1903 17320 1915 17323
rect 2774 17320 2780 17332
rect 1903 17292 2780 17320
rect 1903 17289 1915 17292
rect 1857 17283 1915 17289
rect 1872 17184 1900 17283
rect 2774 17280 2780 17292
rect 2832 17320 2838 17332
rect 3418 17320 3424 17332
rect 2832 17292 3280 17320
rect 3379 17292 3424 17320
rect 2832 17280 2838 17292
rect 3252 17252 3280 17292
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 4706 17320 4712 17332
rect 4667 17292 4712 17320
rect 4706 17280 4712 17292
rect 4764 17320 4770 17332
rect 5350 17320 5356 17332
rect 4764 17292 5356 17320
rect 4764 17280 4770 17292
rect 5350 17280 5356 17292
rect 5408 17280 5414 17332
rect 6270 17280 6276 17332
rect 6328 17320 6334 17332
rect 6641 17323 6699 17329
rect 6641 17320 6653 17323
rect 6328 17292 6653 17320
rect 6328 17280 6334 17292
rect 6641 17289 6653 17292
rect 6687 17320 6699 17323
rect 6822 17320 6828 17332
rect 6687 17292 6828 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7006 17320 7012 17332
rect 6967 17292 7012 17320
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 11793 17323 11851 17329
rect 11793 17320 11805 17323
rect 11572 17292 11805 17320
rect 11572 17280 11578 17292
rect 11793 17289 11805 17292
rect 11839 17289 11851 17323
rect 11793 17283 11851 17289
rect 12066 17280 12072 17332
rect 12124 17320 12130 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 12124 17292 12173 17320
rect 12124 17280 12130 17292
rect 12161 17289 12173 17292
rect 12207 17289 12219 17323
rect 12161 17283 12219 17289
rect 12621 17323 12679 17329
rect 12621 17289 12633 17323
rect 12667 17320 12679 17323
rect 13262 17320 13268 17332
rect 12667 17292 13268 17320
rect 12667 17289 12679 17292
rect 12621 17283 12679 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13538 17320 13544 17332
rect 13499 17292 13544 17320
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 16393 17323 16451 17329
rect 16393 17289 16405 17323
rect 16439 17320 16451 17323
rect 16482 17320 16488 17332
rect 16439 17292 16488 17320
rect 16439 17289 16451 17292
rect 16393 17283 16451 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 16908 17292 17417 17320
rect 16908 17280 16914 17292
rect 17405 17289 17417 17292
rect 17451 17320 17463 17323
rect 18417 17323 18475 17329
rect 18417 17320 18429 17323
rect 17451 17292 18429 17320
rect 17451 17289 17463 17292
rect 17405 17283 17463 17289
rect 18417 17289 18429 17292
rect 18463 17320 18475 17323
rect 19981 17323 20039 17329
rect 18463 17292 19564 17320
rect 18463 17289 18475 17292
rect 18417 17283 18475 17289
rect 4246 17252 4252 17264
rect 3252 17224 4252 17252
rect 4246 17212 4252 17224
rect 4304 17252 4310 17264
rect 4341 17255 4399 17261
rect 4341 17252 4353 17255
rect 4304 17224 4353 17252
rect 4304 17212 4310 17224
rect 4341 17221 4353 17224
rect 4387 17252 4399 17255
rect 4798 17252 4804 17264
rect 4387 17224 4804 17252
rect 4387 17221 4399 17224
rect 4341 17215 4399 17221
rect 4798 17212 4804 17224
rect 4856 17212 4862 17264
rect 2038 17184 2044 17196
rect 1872 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 5368 17193 5396 17280
rect 5353 17187 5411 17193
rect 5353 17153 5365 17187
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 11422 17184 11428 17196
rect 5500 17156 5545 17184
rect 11383 17156 11428 17184
rect 5500 17144 5506 17156
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 13556 17184 13584 17280
rect 13725 17187 13783 17193
rect 13725 17184 13737 17187
rect 13556 17156 13737 17184
rect 13725 17153 13737 17156
rect 13771 17153 13783 17187
rect 13725 17147 13783 17153
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 15436 17156 16865 17184
rect 15436 17144 15442 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 17034 17184 17040 17196
rect 16995 17156 17040 17184
rect 16853 17147 16911 17153
rect 17034 17144 17040 17156
rect 17092 17184 17098 17196
rect 17678 17184 17684 17196
rect 17092 17156 17684 17184
rect 17092 17144 17098 17156
rect 17678 17144 17684 17156
rect 17736 17184 17742 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17736 17156 17785 17184
rect 17736 17144 17742 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 18432 17184 18460 17283
rect 19536 17252 19564 17292
rect 19981 17289 19993 17323
rect 20027 17320 20039 17323
rect 21358 17320 21364 17332
rect 20027 17292 21364 17320
rect 20027 17289 20039 17292
rect 19981 17283 20039 17289
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 22462 17320 22468 17332
rect 22423 17292 22468 17320
rect 22462 17280 22468 17292
rect 22520 17280 22526 17332
rect 20533 17255 20591 17261
rect 20533 17252 20545 17255
rect 19536 17224 20545 17252
rect 20533 17221 20545 17224
rect 20579 17252 20591 17255
rect 20898 17252 20904 17264
rect 20579 17224 20904 17252
rect 20579 17221 20591 17224
rect 20533 17215 20591 17221
rect 20898 17212 20904 17224
rect 20956 17252 20962 17264
rect 20956 17224 21128 17252
rect 20956 17212 20962 17224
rect 21100 17193 21128 17224
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 18432 17156 18613 17184
rect 17773 17147 17831 17153
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 2308 17119 2366 17125
rect 2308 17085 2320 17119
rect 2354 17116 2366 17119
rect 2866 17116 2872 17128
rect 2354 17088 2872 17116
rect 2354 17085 2366 17088
rect 2308 17079 2366 17085
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 4338 17076 4344 17128
rect 4396 17116 4402 17128
rect 5261 17119 5319 17125
rect 5261 17116 5273 17119
rect 4396 17088 5273 17116
rect 4396 17076 4402 17088
rect 5261 17085 5273 17088
rect 5307 17085 5319 17119
rect 5261 17079 5319 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 7374 17116 7380 17128
rect 6871 17088 7380 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7558 17076 7564 17128
rect 7616 17116 7622 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7616 17088 8033 17116
rect 7616 17076 7622 17088
rect 8021 17085 8033 17088
rect 8067 17116 8079 17119
rect 8570 17116 8576 17128
rect 8067 17088 8576 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 9398 17076 9404 17128
rect 9456 17076 9462 17128
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10008 17088 10609 17116
rect 10008 17076 10014 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 4065 17051 4123 17057
rect 4065 17048 4077 17051
rect 3200 17020 4077 17048
rect 3200 17008 3206 17020
rect 4065 17017 4077 17020
rect 4111 17048 4123 17051
rect 5074 17048 5080 17060
rect 4111 17020 5080 17048
rect 4111 17017 4123 17020
rect 4065 17011 4123 17017
rect 5074 17008 5080 17020
rect 5132 17008 5138 17060
rect 5166 17008 5172 17060
rect 5224 17048 5230 17060
rect 7282 17048 7288 17060
rect 5224 17020 7288 17048
rect 5224 17008 5230 17020
rect 7282 17008 7288 17020
rect 7340 17048 7346 17060
rect 7745 17051 7803 17057
rect 7745 17048 7757 17051
rect 7340 17020 7757 17048
rect 7340 17008 7346 17020
rect 7745 17017 7757 17020
rect 7791 17017 7803 17051
rect 7745 17011 7803 17017
rect 7834 17008 7840 17060
rect 7892 17048 7898 17060
rect 8288 17051 8346 17057
rect 8288 17048 8300 17051
rect 7892 17020 8300 17048
rect 7892 17008 7898 17020
rect 8288 17017 8300 17020
rect 8334 17048 8346 17051
rect 9416 17048 9444 17076
rect 10042 17048 10048 17060
rect 8334 17020 10048 17048
rect 8334 17017 8346 17020
rect 8288 17011 8346 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10226 17008 10232 17060
rect 10284 17008 10290 17060
rect 10612 17048 10640 17079
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 10836 17088 11161 17116
rect 10836 17076 10842 17088
rect 11149 17085 11161 17088
rect 11195 17085 11207 17119
rect 11149 17079 11207 17085
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 13998 17125 14004 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12492 17088 12909 17116
rect 12492 17076 12498 17088
rect 12897 17085 12909 17088
rect 12943 17085 12955 17119
rect 13992 17116 14004 17125
rect 13959 17088 14004 17116
rect 12897 17079 12955 17085
rect 13992 17079 14004 17088
rect 13998 17076 14004 17079
rect 14056 17076 14062 17128
rect 16482 17076 16488 17128
rect 16540 17116 16546 17128
rect 16758 17116 16764 17128
rect 16540 17088 16764 17116
rect 16540 17076 16546 17088
rect 16758 17076 16764 17088
rect 16816 17076 16822 17128
rect 18690 17076 18696 17128
rect 18748 17116 18754 17128
rect 18857 17119 18915 17125
rect 18857 17116 18869 17119
rect 18748 17088 18869 17116
rect 18748 17076 18754 17088
rect 18857 17085 18869 17088
rect 18903 17085 18915 17119
rect 18857 17079 18915 17085
rect 11241 17051 11299 17057
rect 11241 17048 11253 17051
rect 10612 17020 11253 17048
rect 11241 17017 11253 17020
rect 11287 17048 11299 17051
rect 12802 17048 12808 17060
rect 11287 17020 12808 17048
rect 11287 17017 11299 17020
rect 11241 17011 11299 17017
rect 12802 17008 12808 17020
rect 12860 17008 12866 17060
rect 15654 17048 15660 17060
rect 12912 17020 15660 17048
rect 4890 16980 4896 16992
rect 4851 16952 4896 16980
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 5592 16952 5917 16980
rect 5592 16940 5598 16952
rect 5905 16949 5917 16952
rect 5951 16949 5963 16983
rect 5905 16943 5963 16949
rect 8570 16940 8576 16992
rect 8628 16980 8634 16992
rect 9401 16983 9459 16989
rect 9401 16980 9413 16983
rect 8628 16952 9413 16980
rect 8628 16940 8634 16952
rect 9401 16949 9413 16952
rect 9447 16949 9459 16983
rect 9401 16943 9459 16949
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9732 16952 9965 16980
rect 9732 16940 9738 16952
rect 9953 16949 9965 16952
rect 9999 16980 10011 16983
rect 10244 16980 10272 17008
rect 12912 16992 12940 17020
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 10778 16980 10784 16992
rect 9999 16952 10272 16980
rect 10739 16952 10784 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 12894 16940 12900 16992
rect 12952 16940 12958 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 14608 16952 15117 16980
rect 14608 16940 14614 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 15672 16980 15700 17008
rect 15930 16980 15936 16992
rect 15672 16952 15936 16980
rect 15105 16943 15163 16949
rect 15930 16940 15936 16952
rect 15988 16940 15994 16992
rect 16114 16980 16120 16992
rect 16075 16952 16120 16980
rect 16114 16940 16120 16952
rect 16172 16940 16178 16992
rect 21100 16980 21128 17147
rect 21358 17125 21364 17128
rect 21352 17116 21364 17125
rect 21319 17088 21364 17116
rect 21352 17079 21364 17088
rect 21358 17076 21364 17079
rect 21416 17076 21422 17128
rect 23293 17119 23351 17125
rect 23293 17085 23305 17119
rect 23339 17116 23351 17119
rect 23661 17119 23719 17125
rect 23661 17116 23673 17119
rect 23339 17088 23673 17116
rect 23339 17085 23351 17088
rect 23293 17079 23351 17085
rect 23661 17085 23673 17088
rect 23707 17085 23719 17119
rect 23661 17079 23719 17085
rect 23109 17051 23167 17057
rect 23109 17017 23121 17051
rect 23155 17048 23167 17051
rect 23928 17051 23986 17057
rect 23928 17048 23940 17051
rect 23155 17020 23940 17048
rect 23155 17017 23167 17020
rect 23109 17011 23167 17017
rect 23928 17017 23940 17020
rect 23974 17048 23986 17051
rect 24210 17048 24216 17060
rect 23974 17020 24216 17048
rect 23974 17017 23986 17020
rect 23928 17011 23986 17017
rect 24210 17008 24216 17020
rect 24268 17008 24274 17060
rect 22094 16980 22100 16992
rect 21100 16952 22100 16980
rect 22094 16940 22100 16952
rect 22152 16940 22158 16992
rect 23014 16940 23020 16992
rect 23072 16980 23078 16992
rect 23293 16983 23351 16989
rect 23293 16980 23305 16983
rect 23072 16952 23305 16980
rect 23072 16940 23078 16952
rect 23293 16949 23305 16952
rect 23339 16980 23351 16983
rect 23385 16983 23443 16989
rect 23385 16980 23397 16983
rect 23339 16952 23397 16980
rect 23339 16949 23351 16952
rect 23293 16943 23351 16949
rect 23385 16949 23397 16952
rect 23431 16949 23443 16983
rect 25038 16980 25044 16992
rect 24999 16952 25044 16980
rect 23385 16943 23443 16949
rect 25038 16940 25044 16952
rect 25096 16940 25102 16992
rect 25314 16940 25320 16992
rect 25372 16980 25378 16992
rect 25593 16983 25651 16989
rect 25593 16980 25605 16983
rect 25372 16952 25605 16980
rect 25372 16940 25378 16952
rect 25593 16949 25605 16952
rect 25639 16949 25651 16983
rect 25593 16943 25651 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1397 16779 1455 16785
rect 1397 16745 1409 16779
rect 1443 16776 1455 16779
rect 1578 16776 1584 16788
rect 1443 16748 1584 16776
rect 1443 16745 1455 16748
rect 1397 16739 1455 16745
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 2038 16776 2044 16788
rect 1995 16748 2044 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3421 16779 3479 16785
rect 3421 16776 3433 16779
rect 2924 16748 3433 16776
rect 2924 16736 2930 16748
rect 3421 16745 3433 16748
rect 3467 16745 3479 16779
rect 4246 16776 4252 16788
rect 4207 16748 4252 16776
rect 3421 16739 3479 16745
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 4893 16779 4951 16785
rect 4893 16776 4905 16779
rect 4396 16748 4905 16776
rect 4396 16736 4402 16748
rect 4893 16745 4905 16748
rect 4939 16745 4951 16779
rect 4893 16739 4951 16745
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5258 16776 5264 16788
rect 5132 16748 5264 16776
rect 5132 16736 5138 16748
rect 5258 16736 5264 16748
rect 5316 16776 5322 16788
rect 6825 16779 6883 16785
rect 6825 16776 6837 16779
rect 5316 16748 6837 16776
rect 5316 16736 5322 16748
rect 6825 16745 6837 16748
rect 6871 16745 6883 16779
rect 6825 16739 6883 16745
rect 7469 16779 7527 16785
rect 7469 16745 7481 16779
rect 7515 16776 7527 16779
rect 7650 16776 7656 16788
rect 7515 16748 7656 16776
rect 7515 16745 7527 16748
rect 7469 16739 7527 16745
rect 7650 16736 7656 16748
rect 7708 16736 7714 16788
rect 7926 16776 7932 16788
rect 7887 16748 7932 16776
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8294 16776 8300 16788
rect 8255 16748 8300 16776
rect 8294 16736 8300 16748
rect 8352 16736 8358 16788
rect 9125 16779 9183 16785
rect 9125 16745 9137 16779
rect 9171 16776 9183 16779
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 9171 16748 10977 16776
rect 9171 16745 9183 16748
rect 9125 16739 9183 16745
rect 10965 16745 10977 16748
rect 11011 16776 11023 16779
rect 11422 16776 11428 16788
rect 11011 16748 11428 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 11422 16736 11428 16748
rect 11480 16736 11486 16788
rect 15105 16779 15163 16785
rect 15105 16745 15117 16779
rect 15151 16776 15163 16779
rect 15378 16776 15384 16788
rect 15151 16748 15384 16776
rect 15151 16745 15163 16748
rect 15105 16739 15163 16745
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 17678 16776 17684 16788
rect 17639 16748 17684 16776
rect 17678 16736 17684 16748
rect 17736 16736 17742 16788
rect 18690 16776 18696 16788
rect 18651 16748 18696 16776
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 18785 16779 18843 16785
rect 18785 16745 18797 16779
rect 18831 16745 18843 16779
rect 19150 16776 19156 16788
rect 19111 16748 19156 16776
rect 18785 16739 18843 16745
rect 1210 16668 1216 16720
rect 1268 16708 1274 16720
rect 4522 16708 4528 16720
rect 1268 16680 4528 16708
rect 1268 16668 1274 16680
rect 4522 16668 4528 16680
rect 4580 16668 4586 16720
rect 5353 16711 5411 16717
rect 5353 16677 5365 16711
rect 5399 16708 5411 16711
rect 5442 16708 5448 16720
rect 5399 16680 5448 16708
rect 5399 16677 5411 16680
rect 5353 16671 5411 16677
rect 5442 16668 5448 16680
rect 5500 16708 5506 16720
rect 5690 16711 5748 16717
rect 5690 16708 5702 16711
rect 5500 16680 5702 16708
rect 5500 16668 5506 16680
rect 5690 16677 5702 16680
rect 5736 16677 5748 16711
rect 7834 16708 7840 16720
rect 7795 16680 7840 16708
rect 5690 16671 5748 16677
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 10229 16711 10287 16717
rect 10229 16708 10241 16711
rect 9692 16680 10241 16708
rect 2590 16600 2596 16652
rect 2648 16600 2654 16652
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3878 16640 3884 16652
rect 2823 16612 3884 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 3878 16600 3884 16612
rect 3936 16600 3942 16652
rect 4062 16640 4068 16652
rect 4023 16612 4068 16640
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 6236 16612 6868 16640
rect 6236 16600 6242 16612
rect 2608 16572 2636 16600
rect 2682 16572 2688 16584
rect 2608 16544 2688 16572
rect 2682 16532 2688 16544
rect 2740 16532 2746 16584
rect 2866 16572 2872 16584
rect 2827 16544 2872 16572
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3142 16572 3148 16584
rect 3099 16544 3148 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 5350 16572 5356 16584
rect 4856 16544 5356 16572
rect 4856 16532 4862 16544
rect 5350 16532 5356 16544
rect 5408 16572 5414 16584
rect 5445 16575 5503 16581
rect 5445 16572 5457 16575
rect 5408 16544 5457 16572
rect 5408 16532 5414 16544
rect 5445 16541 5457 16544
rect 5491 16541 5503 16575
rect 6840 16572 6868 16612
rect 7650 16600 7656 16652
rect 7708 16640 7714 16652
rect 9030 16640 9036 16652
rect 7708 16612 9036 16640
rect 7708 16600 7714 16612
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9122 16600 9128 16652
rect 9180 16640 9186 16652
rect 9401 16643 9459 16649
rect 9401 16640 9413 16643
rect 9180 16612 9413 16640
rect 9180 16600 9186 16612
rect 9401 16609 9413 16612
rect 9447 16609 9459 16643
rect 9692 16640 9720 16680
rect 10229 16677 10241 16680
rect 10275 16708 10287 16711
rect 10870 16708 10876 16720
rect 10275 16680 10876 16708
rect 10275 16677 10287 16680
rect 10229 16671 10287 16677
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 18800 16708 18828 16739
rect 19150 16736 19156 16748
rect 19208 16776 19214 16788
rect 19797 16779 19855 16785
rect 19797 16776 19809 16779
rect 19208 16748 19809 16776
rect 19208 16736 19214 16748
rect 19797 16745 19809 16748
rect 19843 16745 19855 16779
rect 19797 16739 19855 16745
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 20901 16779 20959 16785
rect 20901 16776 20913 16779
rect 20772 16748 20913 16776
rect 20772 16736 20778 16748
rect 20901 16745 20913 16748
rect 20947 16745 20959 16779
rect 21266 16776 21272 16788
rect 21227 16748 21272 16776
rect 20901 16739 20959 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 22554 16776 22560 16788
rect 22515 16748 22560 16776
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 22922 16776 22928 16788
rect 22883 16748 22928 16776
rect 22922 16736 22928 16748
rect 22980 16736 22986 16788
rect 24394 16776 24400 16788
rect 24355 16748 24400 16776
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 20806 16708 20812 16720
rect 18800 16680 20812 16708
rect 20806 16668 20812 16680
rect 20864 16708 20870 16720
rect 23290 16717 23296 16720
rect 21361 16711 21419 16717
rect 21361 16708 21373 16711
rect 20864 16680 21373 16708
rect 20864 16668 20870 16680
rect 21361 16677 21373 16680
rect 21407 16677 21419 16711
rect 23284 16708 23296 16717
rect 23251 16680 23296 16708
rect 21361 16671 21419 16677
rect 23284 16671 23296 16680
rect 23290 16668 23296 16671
rect 23348 16668 23354 16720
rect 9401 16603 9459 16609
rect 9600 16612 9720 16640
rect 7098 16572 7104 16584
rect 6840 16544 7104 16572
rect 5445 16535 5503 16541
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16541 8447 16575
rect 8570 16572 8576 16584
rect 8531 16544 8576 16572
rect 8389 16535 8447 16541
rect 290 16464 296 16516
rect 348 16504 354 16516
rect 348 16476 2544 16504
rect 348 16464 354 16476
rect 1394 16396 1400 16448
rect 1452 16436 1458 16448
rect 2222 16436 2228 16448
rect 1452 16408 2228 16436
rect 1452 16396 1458 16408
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 2406 16436 2412 16448
rect 2367 16408 2412 16436
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 2516 16436 2544 16476
rect 8294 16464 8300 16516
rect 8352 16504 8358 16516
rect 8404 16504 8432 16535
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 9490 16532 9496 16584
rect 9548 16572 9554 16584
rect 9600 16572 9628 16612
rect 9858 16600 9864 16652
rect 9916 16600 9922 16652
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11241 16643 11299 16649
rect 11241 16640 11253 16643
rect 11112 16612 11253 16640
rect 11112 16600 11118 16612
rect 11241 16609 11253 16612
rect 11287 16640 11299 16643
rect 11330 16640 11336 16652
rect 11287 16612 11336 16640
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11698 16649 11704 16652
rect 11692 16640 11704 16649
rect 11659 16612 11704 16640
rect 11692 16603 11704 16612
rect 11698 16600 11704 16603
rect 11756 16600 11762 16652
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13872 16612 13921 16640
rect 13872 16600 13878 16612
rect 13909 16609 13921 16612
rect 13955 16609 13967 16643
rect 13909 16603 13967 16609
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15654 16640 15660 16652
rect 15335 16612 15660 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 15746 16600 15752 16652
rect 15804 16640 15810 16652
rect 16574 16649 16580 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 15804 16612 16313 16640
rect 15804 16600 15810 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16568 16640 16580 16649
rect 16535 16612 16580 16640
rect 16301 16603 16359 16609
rect 16568 16603 16580 16612
rect 16574 16600 16580 16603
rect 16632 16600 16638 16652
rect 19242 16640 19248 16652
rect 19203 16612 19248 16640
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 20349 16643 20407 16649
rect 20349 16609 20361 16643
rect 20395 16640 20407 16643
rect 21266 16640 21272 16652
rect 20395 16612 21272 16640
rect 20395 16609 20407 16612
rect 20349 16603 20407 16609
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 9548 16544 9628 16572
rect 9548 16532 9554 16544
rect 9876 16513 9904 16600
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 10321 16575 10379 16581
rect 10321 16572 10333 16575
rect 10284 16544 10333 16572
rect 10284 16532 10290 16544
rect 10321 16541 10333 16544
rect 10367 16541 10379 16575
rect 10321 16535 10379 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16572 10563 16575
rect 10962 16572 10968 16584
rect 10551 16544 10968 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11422 16572 11428 16584
rect 11383 16544 11428 16572
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 21450 16572 21456 16584
rect 21411 16544 21456 16572
rect 19429 16535 19487 16541
rect 8352 16476 8432 16504
rect 9861 16507 9919 16513
rect 8352 16464 8358 16476
rect 9861 16473 9873 16507
rect 9907 16473 9919 16507
rect 9861 16467 9919 16473
rect 19150 16464 19156 16516
rect 19208 16504 19214 16516
rect 19444 16504 19472 16535
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 23014 16572 23020 16584
rect 22975 16544 23020 16572
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 20717 16507 20775 16513
rect 20717 16504 20729 16507
rect 19208 16476 20729 16504
rect 19208 16464 19214 16476
rect 20717 16473 20729 16476
rect 20763 16504 20775 16507
rect 21358 16504 21364 16516
rect 20763 16476 21364 16504
rect 20763 16473 20775 16476
rect 20717 16467 20775 16473
rect 21358 16464 21364 16476
rect 21416 16504 21422 16516
rect 21913 16507 21971 16513
rect 21913 16504 21925 16507
rect 21416 16476 21925 16504
rect 21416 16464 21422 16476
rect 21913 16473 21925 16476
rect 21959 16504 21971 16507
rect 22002 16504 22008 16516
rect 21959 16476 22008 16504
rect 21959 16473 21971 16476
rect 21913 16467 21971 16473
rect 22002 16464 22008 16476
rect 22060 16464 22066 16516
rect 7282 16436 7288 16448
rect 2516 16408 7288 16436
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 12805 16439 12863 16445
rect 12805 16436 12817 16439
rect 12124 16408 12817 16436
rect 12124 16396 12130 16408
rect 12805 16405 12817 16408
rect 12851 16405 12863 16439
rect 12805 16399 12863 16405
rect 13817 16439 13875 16445
rect 13817 16405 13829 16439
rect 13863 16436 13875 16439
rect 13998 16436 14004 16448
rect 13863 16408 14004 16436
rect 13863 16405 13875 16408
rect 13817 16399 13875 16405
rect 13998 16396 14004 16408
rect 14056 16396 14062 16448
rect 14366 16436 14372 16448
rect 14327 16408 14372 16436
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 15841 16439 15899 16445
rect 15841 16405 15853 16439
rect 15887 16436 15899 16439
rect 16209 16439 16267 16445
rect 16209 16436 16221 16439
rect 15887 16408 16221 16436
rect 15887 16405 15899 16408
rect 15841 16399 15899 16405
rect 16209 16405 16221 16408
rect 16255 16436 16267 16439
rect 16574 16436 16580 16448
rect 16255 16408 16580 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 16574 16396 16580 16408
rect 16632 16436 16638 16448
rect 17034 16436 17040 16448
rect 16632 16408 17040 16436
rect 16632 16396 16638 16408
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 18325 16439 18383 16445
rect 18325 16405 18337 16439
rect 18371 16436 18383 16439
rect 18598 16436 18604 16448
rect 18371 16408 18604 16436
rect 18371 16405 18383 16408
rect 18325 16399 18383 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2409 16235 2467 16241
rect 2409 16232 2421 16235
rect 2096 16204 2421 16232
rect 2096 16192 2102 16204
rect 2409 16201 2421 16204
rect 2455 16201 2467 16235
rect 2409 16195 2467 16201
rect 2424 16096 2452 16195
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 5994 16232 6000 16244
rect 5408 16204 6000 16232
rect 5408 16192 5414 16204
rect 5994 16192 6000 16204
rect 6052 16232 6058 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 6052 16204 6193 16232
rect 6052 16192 6058 16204
rect 6181 16201 6193 16204
rect 6227 16232 6239 16235
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6227 16204 6561 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6549 16201 6561 16204
rect 6595 16232 6607 16235
rect 7558 16232 7564 16244
rect 6595 16204 7564 16232
rect 6595 16201 6607 16204
rect 6549 16195 6607 16201
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 2424 16068 2605 16096
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2593 16059 2651 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5442 16096 5448 16108
rect 5123 16068 5448 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 5442 16056 5448 16068
rect 5500 16096 5506 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5500 16068 5733 16096
rect 5500 16056 5506 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 6564 16096 6592 16195
rect 7558 16192 7564 16204
rect 7616 16232 7622 16244
rect 7616 16204 7788 16232
rect 7616 16192 7622 16204
rect 7760 16164 7788 16204
rect 8386 16192 8392 16244
rect 8444 16232 8450 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8444 16204 8769 16232
rect 8444 16192 8450 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 10226 16232 10232 16244
rect 9815 16204 10232 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 13906 16232 13912 16244
rect 12492 16204 12537 16232
rect 13867 16204 13912 16232
rect 12492 16192 12498 16204
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 14090 16232 14096 16244
rect 14047 16204 14096 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 15746 16192 15752 16244
rect 15804 16232 15810 16244
rect 15841 16235 15899 16241
rect 15841 16232 15853 16235
rect 15804 16204 15853 16232
rect 15804 16192 15810 16204
rect 15841 16201 15853 16204
rect 15887 16201 15899 16235
rect 15841 16195 15899 16201
rect 16393 16235 16451 16241
rect 16393 16201 16405 16235
rect 16439 16232 16451 16235
rect 16482 16232 16488 16244
rect 16439 16204 16488 16232
rect 16439 16201 16451 16204
rect 16393 16195 16451 16201
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 19150 16232 19156 16244
rect 19111 16204 19156 16232
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 19889 16235 19947 16241
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 20438 16232 20444 16244
rect 19935 16204 20444 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 21174 16192 21180 16244
rect 21232 16232 21238 16244
rect 21269 16235 21327 16241
rect 21269 16232 21281 16235
rect 21232 16204 21281 16232
rect 21232 16192 21238 16204
rect 21269 16201 21281 16204
rect 21315 16232 21327 16235
rect 21910 16232 21916 16244
rect 21315 16204 21916 16232
rect 21315 16201 21327 16204
rect 21269 16195 21327 16201
rect 21910 16192 21916 16204
rect 21968 16192 21974 16244
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 23014 16232 23020 16244
rect 22152 16204 23020 16232
rect 22152 16192 22158 16204
rect 23014 16192 23020 16204
rect 23072 16232 23078 16244
rect 23385 16235 23443 16241
rect 23385 16232 23397 16235
rect 23072 16204 23397 16232
rect 23072 16192 23078 16204
rect 23385 16201 23397 16204
rect 23431 16201 23443 16235
rect 23385 16195 23443 16201
rect 9309 16167 9367 16173
rect 9309 16164 9321 16167
rect 7760 16136 9321 16164
rect 9309 16133 9321 16136
rect 9355 16133 9367 16167
rect 9309 16127 9367 16133
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6564 16068 6837 16096
rect 5721 16059 5779 16065
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 1412 15960 1440 15991
rect 3234 15988 3240 16040
rect 3292 16028 3298 16040
rect 7374 16028 7380 16040
rect 3292 16000 7380 16028
rect 3292 15988 3298 16000
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 9324 16028 9352 16127
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12860 16068 13001 16096
rect 12860 16056 12866 16068
rect 12989 16065 13001 16068
rect 13035 16096 13047 16099
rect 13449 16099 13507 16105
rect 13449 16096 13461 16099
rect 13035 16068 13461 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 13449 16065 13461 16068
rect 13495 16065 13507 16099
rect 13924 16096 13952 16192
rect 19797 16167 19855 16173
rect 19797 16133 19809 16167
rect 19843 16164 19855 16167
rect 22741 16167 22799 16173
rect 19843 16136 20576 16164
rect 19843 16133 19855 16136
rect 19797 16127 19855 16133
rect 14550 16096 14556 16108
rect 13924 16068 14556 16096
rect 13449 16059 13507 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 17034 16096 17040 16108
rect 16995 16068 17040 16096
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 18598 16096 18604 16108
rect 18559 16068 18604 16096
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 20346 16096 20352 16108
rect 20307 16068 20352 16096
rect 20346 16056 20352 16068
rect 20404 16056 20410 16108
rect 20548 16105 20576 16136
rect 22741 16133 22753 16167
rect 22787 16164 22799 16167
rect 23290 16164 23296 16176
rect 22787 16136 23296 16164
rect 22787 16133 22799 16136
rect 22741 16127 22799 16133
rect 23290 16124 23296 16136
rect 23348 16124 23354 16176
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16096 20591 16099
rect 21450 16096 21456 16108
rect 20579 16068 21456 16096
rect 20579 16065 20591 16068
rect 20533 16059 20591 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 9861 16031 9919 16037
rect 9861 16028 9873 16031
rect 9324 16000 9873 16028
rect 9861 15997 9873 16000
rect 9907 16028 9919 16031
rect 11422 16028 11428 16040
rect 9907 16000 11428 16028
rect 9907 15997 9919 16000
rect 9861 15991 9919 15997
rect 11422 15988 11428 16000
rect 11480 16028 11486 16040
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11480 16000 11805 16028
rect 11480 15988 11486 16000
rect 11793 15997 11805 16000
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 14182 15988 14188 16040
rect 14240 16028 14246 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 14240 16000 17785 16028
rect 14240 15988 14246 16000
rect 17773 15997 17785 16000
rect 17819 16028 17831 16031
rect 18506 16028 18512 16040
rect 17819 16000 18512 16028
rect 17819 15997 17831 16000
rect 17773 15991 17831 15997
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 20990 15988 20996 16040
rect 21048 16028 21054 16040
rect 21910 16028 21916 16040
rect 21048 16000 21588 16028
rect 21871 16000 21916 16028
rect 21048 15988 21054 16000
rect 2038 15960 2044 15972
rect 1412 15932 2044 15960
rect 2038 15920 2044 15932
rect 2096 15920 2102 15972
rect 2860 15963 2918 15969
rect 2860 15929 2872 15963
rect 2906 15960 2918 15963
rect 3510 15960 3516 15972
rect 2906 15932 3516 15960
rect 2906 15929 2918 15932
rect 2860 15923 2918 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 7098 15969 7104 15972
rect 4709 15963 4767 15969
rect 4709 15929 4721 15963
rect 4755 15960 4767 15963
rect 5629 15963 5687 15969
rect 5629 15960 5641 15963
rect 4755 15932 5641 15960
rect 4755 15929 4767 15932
rect 4709 15923 4767 15929
rect 5629 15929 5641 15932
rect 5675 15960 5687 15963
rect 7092 15960 7104 15969
rect 5675 15932 6684 15960
rect 7059 15932 7104 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 3970 15892 3976 15904
rect 3931 15864 3976 15892
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6656 15892 6684 15932
rect 7092 15923 7104 15932
rect 7098 15920 7104 15923
rect 7156 15920 7162 15972
rect 10128 15963 10186 15969
rect 10128 15929 10140 15963
rect 10174 15960 10186 15963
rect 10962 15960 10968 15972
rect 10174 15932 10968 15960
rect 10174 15929 10186 15932
rect 10128 15923 10186 15929
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 12253 15963 12311 15969
rect 12253 15929 12265 15963
rect 12299 15960 12311 15963
rect 12805 15963 12863 15969
rect 12805 15960 12817 15963
rect 12299 15932 12817 15960
rect 12299 15929 12311 15932
rect 12253 15923 12311 15929
rect 12805 15929 12817 15932
rect 12851 15960 12863 15963
rect 13722 15960 13728 15972
rect 12851 15932 13728 15960
rect 12851 15929 12863 15932
rect 12805 15923 12863 15929
rect 13722 15920 13728 15932
rect 13780 15920 13786 15972
rect 16761 15963 16819 15969
rect 16761 15960 16773 15963
rect 15488 15932 16773 15960
rect 15488 15904 15516 15932
rect 16761 15929 16773 15932
rect 16807 15929 16819 15963
rect 18417 15963 18475 15969
rect 18417 15960 18429 15963
rect 16761 15923 16819 15929
rect 17420 15932 18429 15960
rect 17420 15904 17448 15932
rect 18417 15929 18429 15932
rect 18463 15929 18475 15963
rect 18417 15923 18475 15929
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15960 20315 15963
rect 20530 15960 20536 15972
rect 20303 15932 20536 15960
rect 20303 15929 20315 15932
rect 20257 15923 20315 15929
rect 20530 15920 20536 15932
rect 20588 15960 20594 15972
rect 21560 15960 21588 16000
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 23308 16028 23336 16124
rect 23400 16096 23428 16195
rect 23661 16099 23719 16105
rect 23661 16096 23673 16099
rect 23400 16068 23673 16096
rect 23661 16065 23673 16068
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 23566 16028 23572 16040
rect 23308 16000 23572 16028
rect 23566 15988 23572 16000
rect 23624 15988 23630 16040
rect 21821 15963 21879 15969
rect 21821 15960 21833 15963
rect 20588 15932 21496 15960
rect 21560 15932 21833 15960
rect 20588 15920 20594 15932
rect 7190 15892 7196 15904
rect 6656 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7524 15864 8217 15892
rect 7524 15852 7530 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 11238 15892 11244 15904
rect 11199 15864 11244 15892
rect 8205 15855 8263 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13354 15892 13360 15904
rect 12943 15864 13360 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14366 15892 14372 15904
rect 14327 15864 14372 15892
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 15470 15892 15476 15904
rect 14516 15864 14561 15892
rect 15431 15864 15476 15892
rect 14516 15852 14522 15864
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16850 15892 16856 15904
rect 16347 15864 16856 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 17402 15892 17408 15904
rect 17363 15864 17408 15892
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 18046 15892 18052 15904
rect 18007 15864 18052 15892
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 20990 15892 20996 15904
rect 20951 15864 20996 15892
rect 20990 15852 20996 15864
rect 21048 15852 21054 15904
rect 21468 15901 21496 15932
rect 21821 15929 21833 15932
rect 21867 15929 21879 15963
rect 21821 15923 21879 15929
rect 23106 15920 23112 15972
rect 23164 15960 23170 15972
rect 23906 15963 23964 15969
rect 23906 15960 23918 15963
rect 23164 15932 23918 15960
rect 23164 15920 23170 15932
rect 23906 15929 23918 15932
rect 23952 15929 23964 15963
rect 23906 15923 23964 15929
rect 21453 15895 21511 15901
rect 21453 15861 21465 15895
rect 21499 15861 21511 15895
rect 21453 15855 21511 15861
rect 24210 15852 24216 15904
rect 24268 15892 24274 15904
rect 25041 15895 25099 15901
rect 25041 15892 25053 15895
rect 24268 15864 25053 15892
rect 24268 15852 24274 15864
rect 25041 15861 25053 15864
rect 25087 15892 25099 15895
rect 25222 15892 25228 15904
rect 25087 15864 25228 15892
rect 25087 15861 25099 15864
rect 25041 15855 25099 15861
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 2041 15691 2099 15697
rect 2041 15688 2053 15691
rect 1728 15660 2053 15688
rect 1728 15648 1734 15660
rect 2041 15657 2053 15660
rect 2087 15657 2099 15691
rect 2041 15651 2099 15657
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 2774 15688 2780 15700
rect 2556 15660 2780 15688
rect 2556 15648 2562 15660
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 2924 15660 3801 15688
rect 2924 15648 2930 15660
rect 3789 15657 3801 15660
rect 3835 15688 3847 15691
rect 5166 15688 5172 15700
rect 3835 15660 5172 15688
rect 3835 15657 3847 15660
rect 3789 15651 3847 15657
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 5537 15691 5595 15697
rect 5537 15688 5549 15691
rect 5500 15660 5549 15688
rect 5500 15648 5506 15660
rect 5537 15657 5549 15660
rect 5583 15688 5595 15691
rect 6086 15688 6092 15700
rect 5583 15660 6092 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 6086 15648 6092 15660
rect 6144 15688 6150 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 6144 15660 8033 15688
rect 6144 15648 6150 15660
rect 8021 15657 8033 15660
rect 8067 15688 8079 15691
rect 8570 15688 8576 15700
rect 8067 15660 8576 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 8754 15688 8760 15700
rect 8715 15660 8760 15688
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 9490 15688 9496 15700
rect 9451 15660 9496 15688
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9861 15691 9919 15697
rect 9861 15657 9873 15691
rect 9907 15688 9919 15691
rect 10778 15688 10784 15700
rect 9907 15660 10784 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 10962 15688 10968 15700
rect 10923 15660 10968 15688
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 11333 15691 11391 15697
rect 11333 15657 11345 15691
rect 11379 15688 11391 15691
rect 11698 15688 11704 15700
rect 11379 15660 11704 15688
rect 11379 15657 11391 15660
rect 11333 15651 11391 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 12802 15688 12808 15700
rect 12763 15660 12808 15688
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 14093 15691 14151 15697
rect 14093 15657 14105 15691
rect 14139 15688 14151 15691
rect 14826 15688 14832 15700
rect 14139 15660 14832 15688
rect 14139 15657 14151 15660
rect 14093 15651 14151 15657
rect 14826 15648 14832 15660
rect 14884 15648 14890 15700
rect 15657 15691 15715 15697
rect 15657 15657 15669 15691
rect 15703 15688 15715 15691
rect 16022 15688 16028 15700
rect 15703 15660 16028 15688
rect 15703 15657 15715 15660
rect 15657 15651 15715 15657
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 16393 15691 16451 15697
rect 16393 15657 16405 15691
rect 16439 15688 16451 15691
rect 17034 15688 17040 15700
rect 16439 15660 17040 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 17034 15648 17040 15660
rect 17092 15688 17098 15700
rect 17865 15691 17923 15697
rect 17865 15688 17877 15691
rect 17092 15660 17877 15688
rect 17092 15648 17098 15660
rect 17865 15657 17877 15660
rect 17911 15657 17923 15691
rect 19150 15688 19156 15700
rect 19111 15660 19156 15688
rect 17865 15651 17923 15657
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 19245 15691 19303 15697
rect 19245 15657 19257 15691
rect 19291 15688 19303 15691
rect 20346 15688 20352 15700
rect 19291 15660 20352 15688
rect 19291 15657 19303 15660
rect 19245 15651 19303 15657
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 20806 15688 20812 15700
rect 20763 15660 20812 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 21177 15691 21235 15697
rect 21177 15657 21189 15691
rect 21223 15688 21235 15691
rect 21450 15688 21456 15700
rect 21223 15660 21456 15688
rect 21223 15657 21235 15660
rect 21177 15651 21235 15657
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 22925 15691 22983 15697
rect 22925 15657 22937 15691
rect 22971 15688 22983 15691
rect 23106 15688 23112 15700
rect 22971 15660 23112 15688
rect 22971 15657 22983 15660
rect 22925 15651 22983 15657
rect 23106 15648 23112 15660
rect 23164 15688 23170 15700
rect 23477 15691 23535 15697
rect 23477 15688 23489 15691
rect 23164 15660 23489 15688
rect 23164 15648 23170 15660
rect 23477 15657 23489 15660
rect 23523 15657 23535 15691
rect 23477 15651 23535 15657
rect 2409 15623 2467 15629
rect 2409 15589 2421 15623
rect 2455 15620 2467 15623
rect 2590 15620 2596 15632
rect 2455 15592 2596 15620
rect 2455 15589 2467 15592
rect 2409 15583 2467 15589
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 3142 15620 3148 15632
rect 3103 15592 3148 15620
rect 3142 15580 3148 15592
rect 3200 15580 3206 15632
rect 4798 15620 4804 15632
rect 4711 15592 4804 15620
rect 4798 15580 4804 15592
rect 4856 15620 4862 15632
rect 6172 15623 6230 15629
rect 4856 15592 5212 15620
rect 4856 15580 4862 15592
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 3510 15552 3516 15564
rect 1452 15524 2728 15552
rect 3471 15524 3516 15552
rect 1452 15512 1458 15524
rect 2498 15484 2504 15496
rect 2459 15456 2504 15484
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2700 15493 2728 15524
rect 3510 15512 3516 15524
rect 3568 15512 3574 15564
rect 4706 15552 4712 15564
rect 4667 15524 4712 15552
rect 4706 15512 4712 15524
rect 4764 15552 4770 15564
rect 5074 15552 5080 15564
rect 4764 15524 5080 15552
rect 4764 15512 4770 15524
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 4982 15484 4988 15496
rect 4943 15456 4988 15484
rect 2685 15447 2743 15453
rect 2700 15416 2728 15447
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 3970 15416 3976 15428
rect 2700 15388 3976 15416
rect 3970 15376 3976 15388
rect 4028 15376 4034 15428
rect 4338 15416 4344 15428
rect 4299 15388 4344 15416
rect 4338 15376 4344 15388
rect 4396 15376 4402 15428
rect 1394 15308 1400 15360
rect 1452 15348 1458 15360
rect 1581 15351 1639 15357
rect 1581 15348 1593 15351
rect 1452 15320 1593 15348
rect 1452 15308 1458 15320
rect 1581 15317 1593 15320
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 5000 15348 5028 15444
rect 4212 15320 5028 15348
rect 5184 15348 5212 15592
rect 6172 15589 6184 15623
rect 6218 15620 6230 15623
rect 6270 15620 6276 15632
rect 6218 15592 6276 15620
rect 6218 15589 6230 15592
rect 6172 15583 6230 15589
rect 6270 15580 6276 15592
rect 6328 15580 6334 15632
rect 6362 15580 6368 15632
rect 6420 15580 6426 15632
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 9640 15592 10241 15620
rect 9640 15580 9646 15592
rect 10229 15589 10241 15592
rect 10275 15620 10287 15623
rect 10870 15620 10876 15632
rect 10275 15592 10876 15620
rect 10275 15589 10287 15592
rect 10229 15583 10287 15589
rect 10870 15580 10876 15592
rect 10928 15580 10934 15632
rect 19168 15620 19196 15648
rect 23492 15620 23520 15651
rect 24118 15620 24124 15632
rect 19168 15592 19748 15620
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 5994 15552 6000 15564
rect 5951 15524 6000 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 5994 15512 6000 15524
rect 6052 15552 6058 15564
rect 6380 15552 6408 15580
rect 8570 15552 8576 15564
rect 6052 15524 6408 15552
rect 8531 15524 8576 15552
rect 6052 15512 6058 15524
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 8662 15512 8668 15564
rect 8720 15552 8726 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 8720 15524 9137 15552
rect 8720 15512 8726 15524
rect 9125 15521 9137 15524
rect 9171 15552 9183 15555
rect 10962 15552 10968 15564
rect 9171 15524 10968 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11422 15552 11428 15564
rect 11383 15524 11428 15552
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 11692 15555 11750 15561
rect 11692 15552 11704 15555
rect 11572 15524 11704 15552
rect 11572 15512 11578 15524
rect 11692 15521 11704 15524
rect 11738 15552 11750 15555
rect 12066 15552 12072 15564
rect 11738 15524 12072 15552
rect 11738 15521 11750 15524
rect 11692 15515 11750 15521
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 13906 15552 13912 15564
rect 13867 15524 13912 15552
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 15470 15552 15476 15564
rect 15431 15524 15476 15552
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 16758 15561 16764 15564
rect 16485 15555 16543 15561
rect 16485 15552 16497 15555
rect 15804 15524 16497 15552
rect 15804 15512 15810 15524
rect 16485 15521 16497 15524
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 16752 15515 16764 15561
rect 16816 15552 16822 15564
rect 18785 15555 18843 15561
rect 16816 15524 16852 15552
rect 16758 15512 16764 15515
rect 16816 15512 16822 15524
rect 18785 15521 18797 15555
rect 18831 15552 18843 15555
rect 19242 15552 19248 15564
rect 18831 15524 19248 15552
rect 18831 15521 18843 15524
rect 18785 15515 18843 15521
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 19392 15524 19625 15552
rect 19392 15512 19398 15524
rect 19613 15521 19625 15524
rect 19659 15521 19671 15555
rect 19720 15552 19748 15592
rect 21560 15592 21956 15620
rect 23492 15592 24124 15620
rect 19720 15524 19840 15552
rect 19613 15515 19671 15521
rect 8294 15484 8300 15496
rect 8255 15456 8300 15484
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 10192 15456 10333 15484
rect 10192 15444 10198 15456
rect 10321 15453 10333 15456
rect 10367 15453 10379 15487
rect 10321 15447 10379 15453
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15453 10471 15487
rect 10413 15447 10471 15453
rect 9030 15416 9036 15428
rect 6840 15388 9036 15416
rect 6840 15348 6868 15388
rect 9030 15376 9036 15388
rect 9088 15376 9094 15428
rect 9950 15376 9956 15428
rect 10008 15416 10014 15428
rect 10428 15416 10456 15447
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15764 15484 15792 15512
rect 19812 15493 19840 15524
rect 21560 15496 21588 15592
rect 21634 15512 21640 15564
rect 21692 15552 21698 15564
rect 21801 15555 21859 15561
rect 21801 15552 21813 15555
rect 21692 15524 21813 15552
rect 21692 15512 21698 15524
rect 21801 15521 21813 15524
rect 21847 15521 21859 15555
rect 21928 15552 21956 15592
rect 24118 15580 24124 15592
rect 24176 15580 24182 15632
rect 22094 15552 22100 15564
rect 21928 15524 22100 15552
rect 21801 15515 21859 15521
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 23842 15512 23848 15564
rect 23900 15552 23906 15564
rect 24397 15555 24455 15561
rect 24397 15552 24409 15555
rect 23900 15524 24409 15552
rect 23900 15512 23906 15524
rect 24397 15521 24409 15524
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 24489 15555 24547 15561
rect 24489 15521 24501 15555
rect 24535 15552 24547 15555
rect 24762 15552 24768 15564
rect 24535 15524 24768 15552
rect 24535 15521 24547 15524
rect 24489 15515 24547 15521
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 15436 15456 15792 15484
rect 19705 15487 19763 15493
rect 15436 15444 15442 15456
rect 19705 15453 19717 15487
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15453 19855 15487
rect 21542 15484 21548 15496
rect 21503 15456 21548 15484
rect 19797 15447 19855 15453
rect 10008 15388 10456 15416
rect 10008 15376 10014 15388
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 13872 15388 14381 15416
rect 13872 15376 13878 15388
rect 14369 15385 14381 15388
rect 14415 15416 14427 15419
rect 14458 15416 14464 15428
rect 14415 15388 14464 15416
rect 14415 15385 14427 15388
rect 14369 15379 14427 15385
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 19720 15416 19748 15447
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 23658 15444 23664 15496
rect 23716 15484 23722 15496
rect 24026 15484 24032 15496
rect 23716 15456 24032 15484
rect 23716 15444 23722 15456
rect 24026 15444 24032 15456
rect 24084 15444 24090 15496
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 25222 15484 25228 15496
rect 24719 15456 25228 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 20622 15416 20628 15428
rect 19720 15388 20628 15416
rect 20622 15376 20628 15388
rect 20680 15376 20686 15428
rect 23014 15376 23020 15428
rect 23072 15416 23078 15428
rect 23474 15416 23480 15428
rect 23072 15388 23480 15416
rect 23072 15376 23078 15388
rect 23474 15376 23480 15388
rect 23532 15376 23538 15428
rect 23937 15419 23995 15425
rect 23937 15385 23949 15419
rect 23983 15416 23995 15419
rect 24210 15416 24216 15428
rect 23983 15388 24216 15416
rect 23983 15385 23995 15388
rect 23937 15379 23995 15385
rect 24210 15376 24216 15388
rect 24268 15376 24274 15428
rect 5184 15320 6868 15348
rect 4212 15308 4218 15320
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7285 15351 7343 15357
rect 7285 15348 7297 15351
rect 7064 15320 7297 15348
rect 7064 15308 7070 15320
rect 7285 15317 7297 15320
rect 7331 15317 7343 15351
rect 13354 15348 13360 15360
rect 13315 15320 13360 15348
rect 7285 15311 7343 15317
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 20128 15320 20269 15348
rect 20128 15308 20134 15320
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 24026 15348 24032 15360
rect 23987 15320 24032 15348
rect 20257 15311 20315 15317
rect 24026 15308 24032 15320
rect 24084 15308 24090 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1578 15144 1584 15156
rect 1539 15116 1584 15144
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 2133 15147 2191 15153
rect 2133 15113 2145 15147
rect 2179 15144 2191 15147
rect 2498 15144 2504 15156
rect 2179 15116 2504 15144
rect 2179 15113 2191 15116
rect 2133 15107 2191 15113
rect 2498 15104 2504 15116
rect 2556 15104 2562 15156
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15144 4123 15147
rect 4154 15144 4160 15156
rect 4111 15116 4160 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 4433 15147 4491 15153
rect 4433 15144 4445 15147
rect 4396 15116 4445 15144
rect 4396 15104 4402 15116
rect 4433 15113 4445 15116
rect 4479 15144 4491 15147
rect 4798 15144 4804 15156
rect 4479 15116 4804 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 6270 15104 6276 15156
rect 6328 15144 6334 15156
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 6328 15116 6561 15144
rect 6328 15104 6334 15116
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 6549 15107 6607 15113
rect 9953 15147 10011 15153
rect 9953 15113 9965 15147
rect 9999 15144 10011 15147
rect 10134 15144 10140 15156
rect 9999 15116 10140 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 10778 15144 10784 15156
rect 10739 15116 10784 15144
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 11790 15144 11796 15156
rect 11480 15116 11796 15144
rect 11480 15104 11486 15116
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 14553 15147 14611 15153
rect 14553 15113 14565 15147
rect 14599 15144 14611 15147
rect 15378 15144 15384 15156
rect 14599 15116 15384 15144
rect 14599 15113 14611 15116
rect 14553 15107 14611 15113
rect 1854 15036 1860 15088
rect 1912 15076 1918 15088
rect 2685 15079 2743 15085
rect 2685 15076 2697 15079
rect 1912 15048 2697 15076
rect 1912 15036 1918 15048
rect 2685 15045 2697 15048
rect 2731 15045 2743 15079
rect 4706 15076 4712 15088
rect 4667 15048 4712 15076
rect 2685 15039 2743 15045
rect 4706 15036 4712 15048
rect 4764 15036 4770 15088
rect 11330 15036 11336 15088
rect 11388 15076 11394 15088
rect 12713 15079 12771 15085
rect 12713 15076 12725 15079
rect 11388 15048 12725 15076
rect 11388 15036 11394 15048
rect 12713 15045 12725 15048
rect 12759 15045 12771 15079
rect 12713 15039 12771 15045
rect 3329 15011 3387 15017
rect 3329 14977 3341 15011
rect 3375 15008 3387 15011
rect 3970 15008 3976 15020
rect 3375 14980 3976 15008
rect 3375 14977 3387 14980
rect 3329 14971 3387 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 5810 15008 5816 15020
rect 5771 14980 5816 15008
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 6273 15011 6331 15017
rect 6273 14977 6285 15011
rect 6319 15008 6331 15011
rect 6362 15008 6368 15020
rect 6319 14980 6368 15008
rect 6319 14977 6331 14980
rect 6273 14971 6331 14977
rect 6362 14968 6368 14980
rect 6420 15008 6426 15020
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 6420 14980 7573 15008
rect 6420 14968 6426 14980
rect 7561 14977 7573 14980
rect 7607 15008 7619 15011
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7607 14980 7757 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 11425 15011 11483 15017
rect 11425 14977 11437 15011
rect 11471 15008 11483 15011
rect 11514 15008 11520 15020
rect 11471 14980 11520 15008
rect 11471 14977 11483 14980
rect 11425 14971 11483 14977
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 13262 15008 13268 15020
rect 13223 14980 13268 15008
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13538 14968 13544 15020
rect 13596 15008 13602 15020
rect 14660 15017 14688 15116
rect 15378 15104 15384 15116
rect 15436 15144 15442 15156
rect 16206 15144 16212 15156
rect 15436 15116 16212 15144
rect 15436 15104 15442 15116
rect 16206 15104 16212 15116
rect 16264 15144 16270 15156
rect 16577 15147 16635 15153
rect 16577 15144 16589 15147
rect 16264 15116 16589 15144
rect 16264 15104 16270 15116
rect 16577 15113 16589 15116
rect 16623 15113 16635 15147
rect 16577 15107 16635 15113
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 16945 15147 17003 15153
rect 16945 15144 16957 15147
rect 16816 15116 16957 15144
rect 16816 15104 16822 15116
rect 16945 15113 16957 15116
rect 16991 15113 17003 15147
rect 16945 15107 17003 15113
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 18046 15144 18052 15156
rect 17543 15116 18052 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 16960 15076 16988 15107
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21634 15144 21640 15156
rect 21039 15116 21640 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21634 15104 21640 15116
rect 21692 15144 21698 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21692 15116 21925 15144
rect 21692 15104 21698 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 21913 15107 21971 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 23842 15144 23848 15156
rect 23803 15116 23848 15144
rect 23842 15104 23848 15116
rect 23900 15104 23906 15156
rect 24670 15104 24676 15156
rect 24728 15144 24734 15156
rect 25593 15147 25651 15153
rect 25593 15144 25605 15147
rect 24728 15116 25605 15144
rect 24728 15104 24734 15116
rect 25593 15113 25605 15116
rect 25639 15113 25651 15147
rect 25593 15107 25651 15113
rect 17586 15076 17592 15088
rect 16960 15048 17592 15076
rect 17586 15036 17592 15048
rect 17644 15076 17650 15088
rect 17773 15079 17831 15085
rect 17773 15076 17785 15079
rect 17644 15048 17785 15076
rect 17644 15036 17650 15048
rect 17773 15045 17785 15048
rect 17819 15076 17831 15079
rect 22649 15079 22707 15085
rect 17819 15048 18644 15076
rect 17819 15045 17831 15048
rect 17773 15039 17831 15045
rect 18616 15017 18644 15048
rect 22649 15045 22661 15079
rect 22695 15076 22707 15079
rect 23382 15076 23388 15088
rect 22695 15048 23388 15076
rect 22695 15045 22707 15048
rect 22649 15039 22707 15045
rect 23382 15036 23388 15048
rect 23440 15036 23446 15088
rect 14645 15011 14703 15017
rect 14645 15008 14657 15011
rect 13596 14980 14657 15008
rect 13596 14968 13602 14980
rect 14645 14977 14657 14980
rect 14691 14977 14703 15011
rect 14645 14971 14703 14977
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 14977 18659 15011
rect 23492 15008 23520 15104
rect 24118 15036 24124 15088
rect 24176 15076 24182 15088
rect 24857 15079 24915 15085
rect 24857 15076 24869 15079
rect 24176 15048 24869 15076
rect 24176 15036 24182 15048
rect 24412 15017 24440 15048
rect 24857 15045 24869 15048
rect 24903 15045 24915 15079
rect 25222 15076 25228 15088
rect 25183 15048 25228 15076
rect 24857 15039 24915 15045
rect 25222 15036 25228 15048
rect 25280 15036 25286 15088
rect 24305 15011 24363 15017
rect 24305 15008 24317 15011
rect 23492 14980 24317 15008
rect 18601 14971 18659 14977
rect 24305 14977 24317 14980
rect 24351 14977 24363 15011
rect 24305 14971 24363 14977
rect 24397 15011 24455 15017
rect 24397 14977 24409 15011
rect 24443 14977 24455 15011
rect 24397 14971 24455 14977
rect 1394 14940 1400 14952
rect 1307 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14940 1458 14952
rect 3145 14943 3203 14949
rect 1452 14912 2636 14940
rect 1452 14900 1458 14912
rect 2608 14813 2636 14912
rect 3145 14909 3157 14943
rect 3191 14940 3203 14943
rect 4706 14940 4712 14952
rect 3191 14912 4712 14940
rect 3191 14909 3203 14912
rect 3145 14903 3203 14909
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 5537 14943 5595 14949
rect 5537 14940 5549 14943
rect 5224 14912 5549 14940
rect 5224 14900 5230 14912
rect 5537 14909 5549 14912
rect 5583 14909 5595 14943
rect 5537 14903 5595 14909
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 13170 14940 13176 14952
rect 12299 14912 13176 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 13170 14900 13176 14912
rect 13228 14900 13234 14952
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 16666 14940 16672 14952
rect 13504 14912 16672 14940
rect 13504 14900 13510 14912
rect 16666 14900 16672 14912
rect 16724 14900 16730 14952
rect 18046 14900 18052 14952
rect 18104 14940 18110 14952
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 18104 14912 18429 14940
rect 18104 14900 18110 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18417 14903 18475 14909
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 22462 14940 22468 14952
rect 19659 14912 20944 14940
rect 22423 14912 22468 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 3878 14832 3884 14884
rect 3936 14872 3942 14884
rect 7009 14875 7067 14881
rect 7009 14872 7021 14875
rect 3936 14844 7021 14872
rect 3936 14832 3942 14844
rect 7009 14841 7021 14844
rect 7055 14872 7067 14875
rect 7098 14872 7104 14884
rect 7055 14844 7104 14872
rect 7055 14841 7067 14844
rect 7009 14835 7067 14841
rect 7098 14832 7104 14844
rect 7156 14832 7162 14884
rect 7990 14875 8048 14881
rect 7990 14872 8002 14875
rect 7760 14844 8002 14872
rect 7760 14816 7788 14844
rect 7990 14841 8002 14844
rect 8036 14841 8048 14875
rect 10594 14872 10600 14884
rect 10555 14844 10600 14872
rect 7990 14835 8048 14841
rect 10594 14832 10600 14844
rect 10652 14872 10658 14884
rect 11149 14875 11207 14881
rect 11149 14872 11161 14875
rect 10652 14844 11161 14872
rect 10652 14832 10658 14844
rect 11149 14841 11161 14844
rect 11195 14841 11207 14875
rect 14182 14872 14188 14884
rect 11149 14835 11207 14841
rect 13096 14844 14188 14872
rect 2593 14807 2651 14813
rect 2593 14773 2605 14807
rect 2639 14804 2651 14807
rect 3053 14807 3111 14813
rect 3053 14804 3065 14807
rect 2639 14776 3065 14804
rect 2639 14773 2651 14776
rect 2593 14767 2651 14773
rect 3053 14773 3065 14776
rect 3099 14804 3111 14807
rect 3694 14804 3700 14816
rect 3099 14776 3700 14804
rect 3099 14773 3111 14776
rect 3053 14767 3111 14773
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 5169 14807 5227 14813
rect 5169 14804 5181 14807
rect 5132 14776 5181 14804
rect 5132 14764 5138 14776
rect 5169 14773 5181 14776
rect 5215 14773 5227 14807
rect 5626 14804 5632 14816
rect 5587 14776 5632 14804
rect 5169 14767 5227 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 7742 14764 7748 14816
rect 7800 14764 7806 14816
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9214 14804 9220 14816
rect 9171 14776 9220 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10229 14807 10287 14813
rect 10229 14804 10241 14807
rect 10192 14776 10241 14804
rect 10192 14764 10198 14776
rect 10229 14773 10241 14776
rect 10275 14804 10287 14807
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 10275 14776 11253 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 11241 14773 11253 14776
rect 11287 14804 11299 14807
rect 11422 14804 11428 14816
rect 11287 14776 11428 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13096 14813 13124 14844
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 14826 14832 14832 14884
rect 14884 14881 14890 14884
rect 14884 14875 14948 14881
rect 14884 14841 14902 14875
rect 14936 14841 14948 14875
rect 14884 14835 14948 14841
rect 19880 14875 19938 14881
rect 19880 14841 19892 14875
rect 19926 14872 19938 14875
rect 20070 14872 20076 14884
rect 19926 14844 20076 14872
rect 19926 14841 19938 14844
rect 19880 14835 19938 14841
rect 14884 14832 14890 14835
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 20916 14816 20944 14912
rect 22462 14900 22468 14912
rect 22520 14940 22526 14952
rect 23017 14943 23075 14949
rect 23017 14940 23029 14943
rect 22520 14912 23029 14940
rect 22520 14900 22526 14912
rect 23017 14909 23029 14912
rect 23063 14909 23075 14943
rect 24320 14940 24348 14971
rect 25409 14943 25467 14949
rect 25409 14940 25421 14943
rect 24320 14912 25421 14940
rect 23017 14903 23075 14909
rect 25409 14909 25421 14912
rect 25455 14940 25467 14943
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25455 14912 25973 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 25961 14909 25973 14912
rect 26007 14909 26019 14943
rect 25961 14903 26019 14909
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 12676 14776 13093 14804
rect 12676 14764 12682 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 13081 14767 13139 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 16025 14807 16083 14813
rect 16025 14773 16037 14807
rect 16071 14804 16083 14807
rect 16390 14804 16396 14816
rect 16071 14776 16396 14804
rect 16071 14773 16083 14776
rect 16025 14767 16083 14773
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18414 14804 18420 14816
rect 18095 14776 18420 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 18509 14807 18567 14813
rect 18509 14773 18521 14807
rect 18555 14804 18567 14807
rect 18690 14804 18696 14816
rect 18555 14776 18696 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 19334 14804 19340 14816
rect 19295 14776 19340 14804
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 21542 14804 21548 14816
rect 20956 14776 21548 14804
rect 20956 14764 20962 14776
rect 21542 14764 21548 14776
rect 21600 14764 21606 14816
rect 24210 14804 24216 14816
rect 24171 14776 24216 14804
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2133 14603 2191 14609
rect 2133 14569 2145 14603
rect 2179 14600 2191 14603
rect 2590 14600 2596 14612
rect 2179 14572 2596 14600
rect 2179 14569 2191 14572
rect 2133 14563 2191 14569
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 3513 14603 3571 14609
rect 3513 14569 3525 14603
rect 3559 14600 3571 14603
rect 3881 14603 3939 14609
rect 3881 14600 3893 14603
rect 3559 14572 3893 14600
rect 3559 14569 3571 14572
rect 3513 14563 3571 14569
rect 3881 14569 3893 14572
rect 3927 14600 3939 14603
rect 3970 14600 3976 14612
rect 3927 14572 3976 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 4120 14572 4261 14600
rect 4120 14560 4126 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 5626 14560 5632 14612
rect 5684 14600 5690 14612
rect 6273 14603 6331 14609
rect 6273 14600 6285 14603
rect 5684 14572 6285 14600
rect 5684 14560 5690 14572
rect 6273 14569 6285 14572
rect 6319 14600 6331 14603
rect 6914 14600 6920 14612
rect 6319 14572 6920 14600
rect 6319 14569 6331 14572
rect 6273 14563 6331 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9582 14600 9588 14612
rect 9539 14572 9588 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 11514 14560 11520 14612
rect 11572 14600 11578 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 11572 14572 11621 14600
rect 11572 14560 11578 14572
rect 11609 14569 11621 14572
rect 11655 14600 11667 14603
rect 11977 14603 12035 14609
rect 11977 14600 11989 14603
rect 11655 14572 11989 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 11977 14569 11989 14572
rect 12023 14569 12035 14603
rect 11977 14563 12035 14569
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13262 14600 13268 14612
rect 13219 14572 13268 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13633 14603 13691 14609
rect 13633 14569 13645 14603
rect 13679 14600 13691 14603
rect 13814 14600 13820 14612
rect 13679 14572 13820 14600
rect 13679 14569 13691 14572
rect 13633 14563 13691 14569
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 17586 14600 17592 14612
rect 17547 14572 17592 14600
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 18233 14603 18291 14609
rect 18233 14569 18245 14603
rect 18279 14600 18291 14603
rect 18690 14600 18696 14612
rect 18279 14572 18696 14600
rect 18279 14569 18291 14572
rect 18233 14563 18291 14569
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 20530 14600 20536 14612
rect 19300 14572 20208 14600
rect 20491 14572 20536 14600
rect 19300 14560 19306 14572
rect 1486 14492 1492 14544
rect 1544 14532 1550 14544
rect 1854 14532 1860 14544
rect 1544 14504 1860 14532
rect 1544 14492 1550 14504
rect 1854 14492 1860 14504
rect 1912 14532 1918 14544
rect 2869 14535 2927 14541
rect 2869 14532 2881 14535
rect 1912 14504 2881 14532
rect 1912 14492 1918 14504
rect 2869 14501 2881 14504
rect 2915 14501 2927 14535
rect 2869 14495 2927 14501
rect 5810 14492 5816 14544
rect 5868 14532 5874 14544
rect 5905 14535 5963 14541
rect 5905 14532 5917 14535
rect 5868 14504 5917 14532
rect 5868 14492 5874 14504
rect 5905 14501 5917 14504
rect 5951 14532 5963 14535
rect 6632 14535 6690 14541
rect 6632 14532 6644 14535
rect 5951 14504 6644 14532
rect 5951 14501 5963 14504
rect 5905 14495 5963 14501
rect 6632 14501 6644 14504
rect 6678 14532 6690 14535
rect 7006 14532 7012 14544
rect 6678 14504 7012 14532
rect 6678 14501 6690 14504
rect 6632 14495 6690 14501
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 13556 14532 13584 14560
rect 11848 14504 13584 14532
rect 11848 14492 11854 14504
rect 18322 14492 18328 14544
rect 18380 14532 18386 14544
rect 20180 14541 20208 14572
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 22278 14600 22284 14612
rect 22239 14572 22284 14600
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 23845 14603 23903 14609
rect 23845 14569 23857 14603
rect 23891 14600 23903 14603
rect 24762 14600 24768 14612
rect 23891 14572 24768 14600
rect 23891 14569 23903 14572
rect 23845 14563 23903 14569
rect 24762 14560 24768 14572
rect 24820 14600 24826 14612
rect 24857 14603 24915 14609
rect 24857 14600 24869 14603
rect 24820 14572 24869 14600
rect 24820 14560 24826 14572
rect 24857 14569 24869 14572
rect 24903 14569 24915 14603
rect 25590 14600 25596 14612
rect 25551 14572 25596 14600
rect 24857 14563 24915 14569
rect 25590 14560 25596 14572
rect 25648 14560 25654 14612
rect 19061 14535 19119 14541
rect 19061 14532 19073 14535
rect 18380 14504 19073 14532
rect 18380 14492 18386 14504
rect 19061 14501 19073 14504
rect 19107 14501 19119 14535
rect 19061 14495 19119 14501
rect 20165 14535 20223 14541
rect 20165 14501 20177 14535
rect 20211 14532 20223 14535
rect 20622 14532 20628 14544
rect 20211 14504 20628 14532
rect 20211 14501 20223 14504
rect 20165 14495 20223 14501
rect 20622 14492 20628 14504
rect 20680 14492 20686 14544
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 24305 14535 24363 14541
rect 24305 14532 24317 14535
rect 23716 14504 24317 14532
rect 23716 14492 23722 14504
rect 24305 14501 24317 14504
rect 24351 14501 24363 14535
rect 24305 14495 24363 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14433 1455 14467
rect 1397 14427 1455 14433
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 3142 14464 3148 14476
rect 2823 14436 3148 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 1412 14328 1440 14427
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 5074 14464 5080 14476
rect 4672 14436 5080 14464
rect 4672 14424 4678 14436
rect 5074 14424 5080 14436
rect 5132 14464 5138 14476
rect 5169 14467 5227 14473
rect 5169 14464 5181 14467
rect 5132 14436 5181 14464
rect 5132 14424 5138 14436
rect 5169 14433 5181 14436
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5442 14464 5448 14476
rect 5307 14436 5448 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 6362 14464 6368 14476
rect 6323 14436 6368 14464
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 8662 14424 8668 14476
rect 8720 14464 8726 14476
rect 9944 14467 10002 14473
rect 9944 14464 9956 14467
rect 8720 14436 9956 14464
rect 8720 14424 8726 14436
rect 9944 14433 9956 14436
rect 9990 14464 10002 14467
rect 11238 14464 11244 14476
rect 9990 14436 11244 14464
rect 9990 14433 10002 14436
rect 9944 14427 10002 14433
rect 11238 14424 11244 14436
rect 11296 14424 11302 14476
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 12124 14436 12173 14464
rect 12124 14424 12130 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12161 14427 12219 14433
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13446 14464 13452 14476
rect 13044 14436 13452 14464
rect 13044 14424 13050 14436
rect 13446 14424 13452 14436
rect 13504 14464 13510 14476
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13504 14436 14013 14464
rect 13504 14424 13510 14436
rect 14001 14433 14013 14436
rect 14047 14464 14059 14467
rect 15378 14464 15384 14476
rect 14047 14436 15384 14464
rect 14047 14433 14059 14436
rect 14001 14427 14059 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16206 14464 16212 14476
rect 16167 14436 16212 14464
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 21174 14473 21180 14476
rect 16465 14467 16523 14473
rect 16465 14464 16477 14467
rect 16356 14436 16477 14464
rect 16356 14424 16362 14436
rect 16465 14433 16477 14436
rect 16511 14433 16523 14467
rect 16465 14427 16523 14433
rect 21168 14427 21180 14473
rect 21232 14464 21238 14476
rect 23385 14467 23443 14473
rect 21232 14436 21268 14464
rect 21174 14424 21180 14427
rect 21232 14424 21238 14436
rect 23385 14433 23397 14467
rect 23431 14464 23443 14467
rect 23842 14464 23848 14476
rect 23431 14436 23848 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 24213 14467 24271 14473
rect 24213 14433 24225 14467
rect 24259 14464 24271 14467
rect 24670 14464 24676 14476
rect 24259 14436 24676 14464
rect 24259 14433 24271 14436
rect 24213 14427 24271 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 25130 14424 25136 14476
rect 25188 14464 25194 14476
rect 25409 14467 25467 14473
rect 25409 14464 25421 14467
rect 25188 14436 25421 14464
rect 25188 14424 25194 14436
rect 25409 14433 25421 14436
rect 25455 14433 25467 14467
rect 25409 14427 25467 14433
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2924 14368 2973 14396
rect 2924 14356 2930 14368
rect 2961 14365 2973 14368
rect 3007 14365 3019 14399
rect 5350 14396 5356 14408
rect 5311 14368 5356 14396
rect 2961 14359 3019 14365
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 9490 14356 9496 14408
rect 9548 14396 9554 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9548 14368 9689 14396
rect 9548 14356 9554 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 14090 14396 14096 14408
rect 14051 14368 14096 14396
rect 9677 14359 9735 14365
rect 14090 14356 14096 14368
rect 14148 14356 14154 14408
rect 14182 14356 14188 14408
rect 14240 14396 14246 14408
rect 19150 14396 19156 14408
rect 14240 14368 14285 14396
rect 19111 14368 19156 14396
rect 14240 14356 14246 14368
rect 19150 14356 19156 14368
rect 19208 14356 19214 14408
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 19797 14399 19855 14405
rect 19300 14368 19345 14396
rect 19300 14356 19306 14368
rect 19797 14365 19809 14399
rect 19843 14396 19855 14399
rect 20898 14396 20904 14408
rect 19843 14368 20904 14396
rect 19843 14365 19855 14368
rect 19797 14359 19855 14365
rect 20898 14356 20904 14368
rect 20956 14356 20962 14408
rect 24118 14356 24124 14408
rect 24176 14396 24182 14408
rect 24397 14399 24455 14405
rect 24397 14396 24409 14399
rect 24176 14368 24409 14396
rect 24176 14356 24182 14368
rect 24397 14365 24409 14368
rect 24443 14365 24455 14399
rect 24397 14359 24455 14365
rect 3234 14328 3240 14340
rect 1412 14300 3240 14328
rect 3234 14288 3240 14300
rect 3292 14328 3298 14340
rect 4801 14331 4859 14337
rect 4801 14328 4813 14331
rect 3292 14300 4813 14328
rect 3292 14288 3298 14300
rect 4801 14297 4813 14300
rect 4847 14297 4859 14331
rect 7742 14328 7748 14340
rect 7703 14300 7748 14328
rect 4801 14291 4859 14297
rect 7742 14288 7748 14300
rect 7800 14328 7806 14340
rect 8297 14331 8355 14337
rect 8297 14328 8309 14331
rect 7800 14300 8309 14328
rect 7800 14288 7806 14300
rect 8297 14297 8309 14300
rect 8343 14297 8355 14331
rect 12342 14328 12348 14340
rect 12303 14300 12348 14328
rect 8297 14291 8355 14297
rect 12342 14288 12348 14300
rect 12400 14288 12406 14340
rect 1394 14220 1400 14272
rect 1452 14260 1458 14272
rect 1581 14263 1639 14269
rect 1581 14260 1593 14263
rect 1452 14232 1593 14260
rect 1452 14220 1458 14232
rect 1581 14229 1593 14232
rect 1627 14229 1639 14263
rect 1581 14223 1639 14229
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 2682 14260 2688 14272
rect 2455 14232 2688 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 4706 14260 4712 14272
rect 4667 14232 4712 14260
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 8754 14260 8760 14272
rect 8715 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9582 14260 9588 14272
rect 9171 14232 9588 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 11054 14260 11060 14272
rect 11015 14232 11060 14260
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 12713 14263 12771 14269
rect 12713 14260 12725 14263
rect 12676 14232 12725 14260
rect 12676 14220 12682 14232
rect 12713 14229 12725 14232
rect 12759 14229 12771 14263
rect 12713 14223 12771 14229
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 14516 14232 14657 14260
rect 14516 14220 14522 14232
rect 14645 14229 14657 14232
rect 14691 14260 14703 14263
rect 14826 14260 14832 14272
rect 14691 14232 14832 14260
rect 14691 14229 14703 14232
rect 14645 14223 14703 14229
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 16022 14260 16028 14272
rect 15983 14232 16028 14260
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 18601 14263 18659 14269
rect 18601 14229 18613 14263
rect 18647 14260 18659 14263
rect 18782 14260 18788 14272
rect 18647 14232 18788 14260
rect 18647 14229 18659 14232
rect 18601 14223 18659 14229
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 23017 14263 23075 14269
rect 23017 14229 23029 14263
rect 23063 14260 23075 14263
rect 23290 14260 23296 14272
rect 23063 14232 23296 14260
rect 23063 14229 23075 14232
rect 23017 14223 23075 14229
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 23750 14260 23756 14272
rect 23711 14232 23756 14260
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1578 14056 1584 14068
rect 1539 14028 1584 14056
rect 1578 14016 1584 14028
rect 1636 14016 1642 14068
rect 1854 14016 1860 14068
rect 1912 14056 1918 14068
rect 1949 14059 2007 14065
rect 1949 14056 1961 14059
rect 1912 14028 1961 14056
rect 1912 14016 1918 14028
rect 1949 14025 1961 14028
rect 1995 14025 2007 14059
rect 1949 14019 2007 14025
rect 2222 14016 2228 14068
rect 2280 14056 2286 14068
rect 2685 14059 2743 14065
rect 2685 14056 2697 14059
rect 2280 14028 2697 14056
rect 2280 14016 2286 14028
rect 2685 14025 2697 14028
rect 2731 14025 2743 14059
rect 2685 14019 2743 14025
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 3786 14056 3792 14068
rect 3476 14028 3792 14056
rect 3476 14016 3482 14028
rect 3786 14016 3792 14028
rect 3844 14056 3850 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 3844 14028 4997 14056
rect 3844 14016 3850 14028
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 6362 14056 6368 14068
rect 6323 14028 6368 14056
rect 4985 14019 5043 14025
rect 2409 13991 2467 13997
rect 2409 13957 2421 13991
rect 2455 13988 2467 13991
rect 2866 13988 2872 14000
rect 2455 13960 2872 13988
rect 2455 13957 2467 13960
rect 2409 13951 2467 13957
rect 2866 13948 2872 13960
rect 2924 13948 2930 14000
rect 5000 13932 5028 14019
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 7469 14059 7527 14065
rect 7469 14056 7481 14059
rect 7432 14028 7481 14056
rect 7432 14016 7438 14028
rect 7469 14025 7481 14028
rect 7515 14025 7527 14059
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 7469 14019 7527 14025
rect 7576 14028 9045 14056
rect 5166 13988 5172 14000
rect 5127 13960 5172 13988
rect 5166 13948 5172 13960
rect 5224 13948 5230 14000
rect 6380 13988 6408 14016
rect 7576 13988 7604 14028
rect 9033 14025 9045 14028
rect 9079 14056 9091 14059
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 9079 14028 9413 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9401 14025 9413 14028
rect 9447 14056 9459 14059
rect 9490 14056 9496 14068
rect 9447 14028 9496 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 11238 14016 11244 14068
rect 11296 14056 11302 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 11296 14028 11529 14056
rect 11296 14016 11302 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12216 14028 12909 14056
rect 12216 14016 12222 14028
rect 12897 14025 12909 14028
rect 12943 14056 12955 14059
rect 14090 14056 14096 14068
rect 12943 14028 14096 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 15841 14059 15899 14065
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 16298 14056 16304 14068
rect 15887 14028 16304 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 16298 14016 16304 14028
rect 16356 14056 16362 14068
rect 17865 14059 17923 14065
rect 17865 14056 17877 14059
rect 16356 14028 17877 14056
rect 16356 14016 16362 14028
rect 17865 14025 17877 14028
rect 17911 14056 17923 14059
rect 18598 14056 18604 14068
rect 17911 14028 18604 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 18598 14016 18604 14028
rect 18656 14056 18662 14068
rect 19242 14056 19248 14068
rect 18656 14028 19248 14056
rect 18656 14016 18662 14028
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 21453 14059 21511 14065
rect 21453 14025 21465 14059
rect 21499 14056 21511 14059
rect 23290 14056 23296 14068
rect 21499 14028 23296 14056
rect 21499 14025 21511 14028
rect 21453 14019 21511 14025
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25409 14059 25467 14065
rect 25409 14056 25421 14059
rect 24912 14028 25421 14056
rect 24912 14016 24918 14028
rect 25409 14025 25421 14028
rect 25455 14025 25467 14059
rect 25409 14019 25467 14025
rect 6380 13960 7604 13988
rect 8021 13991 8079 13997
rect 8021 13957 8033 13991
rect 8067 13988 8079 13991
rect 8202 13988 8208 14000
rect 8067 13960 8208 13988
rect 8067 13957 8079 13960
rect 8021 13951 8079 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 13446 13988 13452 14000
rect 13403 13960 13452 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 13446 13948 13452 13960
rect 13504 13948 13510 14000
rect 14458 13948 14464 14000
rect 14516 13988 14522 14000
rect 14829 13991 14887 13997
rect 14829 13988 14841 13991
rect 14516 13960 14841 13988
rect 14516 13948 14522 13960
rect 14829 13957 14841 13960
rect 14875 13957 14887 13991
rect 14829 13951 14887 13957
rect 16206 13948 16212 14000
rect 16264 13988 16270 14000
rect 16758 13988 16764 14000
rect 16264 13960 16764 13988
rect 16264 13948 16270 13960
rect 16758 13948 16764 13960
rect 16816 13988 16822 14000
rect 16945 13991 17003 13997
rect 16945 13988 16957 13991
rect 16816 13960 16957 13988
rect 16816 13948 16822 13960
rect 16945 13957 16957 13960
rect 16991 13957 17003 13991
rect 16945 13951 17003 13957
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 2222 13920 2228 13932
rect 1728 13892 2228 13920
rect 1728 13880 1734 13892
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 3878 13920 3884 13932
rect 3559 13892 3884 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 3878 13880 3884 13892
rect 3936 13920 3942 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 3936 13892 4169 13920
rect 3936 13880 3942 13892
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 4982 13920 4988 13932
rect 4895 13892 4988 13920
rect 4157 13883 4215 13889
rect 4982 13880 4988 13892
rect 5040 13920 5046 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5040 13892 5641 13920
rect 5040 13880 5046 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5810 13920 5816 13932
rect 5723 13892 5816 13920
rect 5629 13883 5687 13889
rect 5810 13880 5816 13892
rect 5868 13920 5874 13932
rect 6270 13920 6276 13932
rect 5868 13892 6276 13920
rect 5868 13880 5874 13892
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8662 13920 8668 13932
rect 8168 13892 8668 13920
rect 8168 13880 8174 13892
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 8812 13892 9720 13920
rect 8812 13880 8818 13892
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 3050 13852 3056 13864
rect 2547 13824 3056 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3602 13812 3608 13864
rect 3660 13852 3666 13864
rect 4709 13855 4767 13861
rect 3660 13824 4200 13852
rect 3660 13812 3666 13824
rect 3510 13744 3516 13796
rect 3568 13784 3574 13796
rect 4065 13787 4123 13793
rect 4065 13784 4077 13787
rect 3568 13756 4077 13784
rect 3568 13744 3574 13756
rect 4065 13753 4077 13756
rect 4111 13753 4123 13787
rect 4065 13747 4123 13753
rect 3602 13716 3608 13728
rect 3563 13688 3608 13716
rect 3602 13676 3608 13688
rect 3660 13676 3666 13728
rect 3970 13716 3976 13728
rect 3931 13688 3976 13716
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4172 13716 4200 13824
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 7834 13852 7840 13864
rect 4755 13824 5488 13852
rect 7795 13824 7840 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 5460 13784 5488 13824
rect 7834 13812 7840 13824
rect 7892 13852 7898 13864
rect 7892 13824 8248 13852
rect 7892 13812 7898 13824
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5460 13756 5549 13784
rect 5537 13753 5549 13756
rect 5583 13784 5595 13787
rect 6825 13787 6883 13793
rect 6825 13784 6837 13787
rect 5583 13756 6837 13784
rect 5583 13753 5595 13756
rect 5537 13747 5595 13753
rect 6825 13753 6837 13756
rect 6871 13753 6883 13787
rect 8220 13784 8248 13824
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9548 13824 9597 13852
rect 9548 13812 9554 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9692 13852 9720 13892
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 16485 13923 16543 13929
rect 16485 13920 16497 13923
rect 16080 13892 16497 13920
rect 16080 13880 16086 13892
rect 16485 13889 16497 13892
rect 16531 13889 16543 13923
rect 16485 13883 16543 13889
rect 9841 13855 9899 13861
rect 9841 13852 9853 13855
rect 9692 13824 9853 13852
rect 9585 13815 9643 13821
rect 9841 13821 9853 13824
rect 9887 13852 9899 13855
rect 10134 13852 10140 13864
rect 9887 13824 10140 13852
rect 9887 13821 9899 13824
rect 9841 13815 9899 13821
rect 10134 13812 10140 13824
rect 10192 13852 10198 13864
rect 11054 13852 11060 13864
rect 10192 13824 11060 13852
rect 10192 13812 10198 13824
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 13446 13852 13452 13864
rect 13407 13824 13452 13852
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 15378 13852 15384 13864
rect 15339 13824 15384 13852
rect 15378 13812 15384 13824
rect 15436 13852 15442 13864
rect 16393 13855 16451 13861
rect 16393 13852 16405 13855
rect 15436 13824 16405 13852
rect 15436 13812 15442 13824
rect 16393 13821 16405 13824
rect 16439 13821 16451 13855
rect 16960 13852 16988 13951
rect 18322 13948 18328 14000
rect 18380 13988 18386 14000
rect 18417 13991 18475 13997
rect 18417 13988 18429 13991
rect 18380 13960 18429 13988
rect 18380 13948 18386 13960
rect 18417 13957 18429 13960
rect 18463 13957 18475 13991
rect 18417 13951 18475 13957
rect 19981 13991 20039 13997
rect 19981 13957 19993 13991
rect 20027 13988 20039 13991
rect 20070 13988 20076 14000
rect 20027 13960 20076 13988
rect 20027 13957 20039 13960
rect 19981 13951 20039 13957
rect 18432 13920 18460 13951
rect 20070 13948 20076 13960
rect 20128 13948 20134 14000
rect 23109 13991 23167 13997
rect 23109 13957 23121 13991
rect 23155 13988 23167 13991
rect 24118 13988 24124 14000
rect 23155 13960 24124 13988
rect 23155 13957 23167 13960
rect 23109 13951 23167 13957
rect 24118 13948 24124 13960
rect 24176 13948 24182 14000
rect 22002 13920 22008 13932
rect 18432 13892 18736 13920
rect 21963 13892 22008 13920
rect 18708 13864 18736 13892
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 23382 13880 23388 13932
rect 23440 13920 23446 13932
rect 23750 13920 23756 13932
rect 23440 13892 23756 13920
rect 23440 13880 23446 13892
rect 23750 13880 23756 13892
rect 23808 13920 23814 13932
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 23808 13892 24225 13920
rect 23808 13880 23814 13892
rect 24213 13889 24225 13892
rect 24259 13889 24271 13923
rect 24213 13883 24271 13889
rect 25130 13880 25136 13932
rect 25188 13920 25194 13932
rect 26145 13923 26203 13929
rect 26145 13920 26157 13923
rect 25188 13892 26157 13920
rect 25188 13880 25194 13892
rect 26145 13889 26157 13892
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 18598 13852 18604 13864
rect 16960 13824 18604 13852
rect 16393 13815 16451 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 18690 13812 18696 13864
rect 18748 13812 18754 13864
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 8389 13787 8447 13793
rect 8389 13784 8401 13787
rect 8220 13756 8401 13784
rect 6825 13747 6883 13753
rect 8389 13753 8401 13756
rect 8435 13753 8447 13787
rect 8389 13747 8447 13753
rect 8481 13787 8539 13793
rect 8481 13753 8493 13787
rect 8527 13784 8539 13787
rect 11146 13784 11152 13796
rect 8527 13756 11152 13784
rect 8527 13753 8539 13756
rect 8481 13747 8539 13753
rect 6914 13716 6920 13728
rect 4172 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 7374 13676 7380 13728
rect 7432 13716 7438 13728
rect 8496 13716 8524 13747
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 13694 13787 13752 13793
rect 13694 13784 13706 13787
rect 12268 13756 13706 13784
rect 12268 13728 12296 13756
rect 13694 13753 13706 13756
rect 13740 13784 13752 13787
rect 13814 13784 13820 13796
rect 13740 13756 13820 13784
rect 13740 13753 13752 13756
rect 13694 13747 13752 13753
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 18782 13744 18788 13796
rect 18840 13793 18846 13796
rect 18840 13787 18904 13793
rect 18840 13753 18858 13787
rect 18892 13753 18904 13787
rect 18840 13747 18904 13753
rect 18840 13744 18846 13747
rect 19242 13744 19248 13796
rect 19300 13784 19306 13796
rect 19518 13784 19524 13796
rect 19300 13756 19524 13784
rect 19300 13744 19306 13756
rect 19518 13744 19524 13756
rect 19576 13744 19582 13796
rect 20640 13784 20668 13815
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 21913 13855 21971 13861
rect 21913 13852 21925 13855
rect 21324 13824 21925 13852
rect 21324 13812 21330 13824
rect 21913 13821 21925 13824
rect 21959 13852 21971 13855
rect 22462 13852 22468 13864
rect 21959 13824 22468 13852
rect 21959 13821 21971 13824
rect 21913 13815 21971 13821
rect 22462 13812 22468 13824
rect 22520 13812 22526 13864
rect 23477 13855 23535 13861
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 23658 13852 23664 13864
rect 23523 13824 23664 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 24118 13852 24124 13864
rect 24079 13824 24124 13852
rect 24118 13812 24124 13824
rect 24176 13852 24182 13864
rect 25041 13855 25099 13861
rect 25041 13852 25053 13855
rect 24176 13824 25053 13852
rect 24176 13812 24182 13824
rect 25041 13821 25053 13824
rect 25087 13821 25099 13855
rect 25222 13852 25228 13864
rect 25183 13824 25228 13852
rect 25041 13815 25099 13821
rect 25222 13812 25228 13824
rect 25280 13852 25286 13864
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25280 13824 25789 13852
rect 25280 13812 25286 13824
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 25777 13815 25835 13821
rect 21542 13784 21548 13796
rect 20640 13756 21548 13784
rect 21542 13744 21548 13756
rect 21600 13784 21606 13796
rect 21821 13787 21879 13793
rect 21821 13784 21833 13787
rect 21600 13756 21833 13784
rect 21600 13744 21606 13756
rect 21821 13753 21833 13756
rect 21867 13753 21879 13787
rect 21821 13747 21879 13753
rect 22094 13744 22100 13796
rect 22152 13784 22158 13796
rect 22152 13756 22600 13784
rect 22152 13744 22158 13756
rect 10962 13716 10968 13728
rect 7432 13688 8524 13716
rect 10923 13688 10968 13716
rect 7432 13676 7438 13688
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 12250 13716 12256 13728
rect 12211 13688 12256 13716
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 12437 13719 12495 13725
rect 12437 13685 12449 13719
rect 12483 13716 12495 13719
rect 12526 13716 12532 13728
rect 12483 13688 12532 13716
rect 12483 13685 12495 13688
rect 12437 13679 12495 13685
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 15930 13716 15936 13728
rect 15891 13688 15936 13716
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16298 13716 16304 13728
rect 16259 13688 16304 13716
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 20898 13676 20904 13728
rect 20956 13716 20962 13728
rect 20993 13719 21051 13725
rect 20993 13716 21005 13719
rect 20956 13688 21005 13716
rect 20956 13676 20962 13688
rect 20993 13685 21005 13688
rect 21039 13716 21051 13719
rect 21266 13716 21272 13728
rect 21039 13688 21272 13716
rect 21039 13685 21051 13688
rect 20993 13679 21051 13685
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 22002 13676 22008 13728
rect 22060 13716 22066 13728
rect 22465 13719 22523 13725
rect 22465 13716 22477 13719
rect 22060 13688 22477 13716
rect 22060 13676 22066 13688
rect 22465 13685 22477 13688
rect 22511 13685 22523 13719
rect 22572 13716 22600 13756
rect 23290 13744 23296 13796
rect 23348 13784 23354 13796
rect 24029 13787 24087 13793
rect 24029 13784 24041 13787
rect 23348 13756 24041 13784
rect 23348 13744 23354 13756
rect 24029 13753 24041 13756
rect 24075 13753 24087 13787
rect 24029 13747 24087 13753
rect 23661 13719 23719 13725
rect 23661 13716 23673 13719
rect 22572 13688 23673 13716
rect 22465 13679 22523 13685
rect 23661 13685 23673 13688
rect 23707 13685 23719 13719
rect 24670 13716 24676 13728
rect 24631 13688 24676 13716
rect 23661 13679 23719 13685
rect 24670 13676 24676 13688
rect 24728 13676 24734 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1762 13472 1768 13524
rect 1820 13512 1826 13524
rect 1949 13515 2007 13521
rect 1949 13512 1961 13515
rect 1820 13484 1961 13512
rect 1820 13472 1826 13484
rect 1949 13481 1961 13484
rect 1995 13481 2007 13515
rect 1949 13475 2007 13481
rect 2130 13472 2136 13524
rect 2188 13512 2194 13524
rect 2317 13515 2375 13521
rect 2317 13512 2329 13515
rect 2188 13484 2329 13512
rect 2188 13472 2194 13484
rect 2317 13481 2329 13484
rect 2363 13481 2375 13515
rect 2317 13475 2375 13481
rect 2685 13515 2743 13521
rect 2685 13481 2697 13515
rect 2731 13512 2743 13515
rect 2774 13512 2780 13524
rect 2731 13484 2780 13512
rect 2731 13481 2743 13484
rect 2685 13475 2743 13481
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 3510 13472 3516 13524
rect 3568 13512 3574 13524
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 3568 13484 3617 13512
rect 3568 13472 3574 13484
rect 3605 13481 3617 13484
rect 3651 13481 3663 13515
rect 3605 13475 3663 13481
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 4028 13484 4261 13512
rect 4028 13472 4034 13484
rect 4249 13481 4261 13484
rect 4295 13512 4307 13515
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4295 13484 4445 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 4433 13481 4445 13484
rect 4479 13481 4491 13515
rect 4890 13512 4896 13524
rect 4851 13484 4896 13512
rect 4433 13475 4491 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 5408 13484 5457 13512
rect 5408 13472 5414 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5445 13475 5503 13481
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5592 13484 6009 13512
rect 5592 13472 5598 13484
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 6454 13512 6460 13524
rect 6415 13484 6460 13512
rect 5997 13475 6055 13481
rect 6454 13472 6460 13484
rect 6512 13472 6518 13524
rect 7006 13512 7012 13524
rect 6967 13484 7012 13512
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 8110 13512 8116 13524
rect 7975 13484 8116 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 8478 13512 8484 13524
rect 8435 13484 8484 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 8478 13472 8484 13484
rect 8536 13512 8542 13524
rect 9030 13512 9036 13524
rect 8536 13484 9036 13512
rect 8536 13472 8542 13484
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9398 13512 9404 13524
rect 9359 13484 9404 13512
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 11054 13512 11060 13524
rect 10744 13484 11060 13512
rect 10744 13472 10750 13484
rect 11054 13472 11060 13484
rect 11112 13472 11118 13524
rect 13814 13512 13820 13524
rect 13775 13484 13820 13512
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14369 13515 14427 13521
rect 14369 13512 14381 13515
rect 14240 13484 14381 13512
rect 14240 13472 14246 13484
rect 14369 13481 14381 13484
rect 14415 13481 14427 13515
rect 14369 13475 14427 13481
rect 18598 13472 18604 13524
rect 18656 13512 18662 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 18656 13484 18705 13512
rect 18656 13472 18662 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 19150 13512 19156 13524
rect 19111 13484 19156 13512
rect 18693 13475 18751 13481
rect 19150 13472 19156 13484
rect 19208 13472 19214 13524
rect 21174 13512 21180 13524
rect 21135 13484 21180 13512
rect 21174 13472 21180 13484
rect 21232 13512 21238 13524
rect 22649 13515 22707 13521
rect 22649 13512 22661 13515
rect 21232 13484 22661 13512
rect 21232 13472 21238 13484
rect 22649 13481 22661 13484
rect 22695 13512 22707 13515
rect 23382 13512 23388 13524
rect 22695 13484 23388 13512
rect 22695 13481 22707 13484
rect 22649 13475 22707 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 23661 13515 23719 13521
rect 23661 13481 23673 13515
rect 23707 13512 23719 13515
rect 24026 13512 24032 13524
rect 23707 13484 24032 13512
rect 23707 13481 23719 13484
rect 23661 13475 23719 13481
rect 24026 13472 24032 13484
rect 24084 13512 24090 13524
rect 24121 13515 24179 13521
rect 24121 13512 24133 13515
rect 24084 13484 24133 13512
rect 24084 13472 24090 13484
rect 24121 13481 24133 13484
rect 24167 13481 24179 13515
rect 24121 13475 24179 13481
rect 5810 13444 5816 13456
rect 5771 13416 5816 13444
rect 5810 13404 5816 13416
rect 5868 13404 5874 13456
rect 6472 13444 6500 13472
rect 7377 13447 7435 13453
rect 7377 13444 7389 13447
rect 6472 13416 7389 13444
rect 7377 13413 7389 13416
rect 7423 13413 7435 13447
rect 7377 13407 7435 13413
rect 16390 13404 16396 13456
rect 16448 13444 16454 13456
rect 17006 13447 17064 13453
rect 17006 13444 17018 13447
rect 16448 13416 17018 13444
rect 16448 13404 16454 13416
rect 17006 13413 17018 13416
rect 17052 13413 17064 13447
rect 19702 13444 19708 13456
rect 19615 13416 19708 13444
rect 17006 13407 17064 13413
rect 19702 13404 19708 13416
rect 19760 13444 19766 13456
rect 19760 13416 22692 13444
rect 19760 13404 19766 13416
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2130 13376 2136 13388
rect 1443 13348 2136 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2130 13336 2136 13348
rect 2188 13336 2194 13388
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2774 13376 2780 13388
rect 2547 13348 2780 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 4798 13376 4804 13388
rect 4759 13348 4804 13376
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 6362 13376 6368 13388
rect 6323 13348 6368 13376
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 8110 13376 8116 13388
rect 6972 13348 8116 13376
rect 6972 13336 6978 13348
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8352 13348 8493 13376
rect 8352 13336 8358 13348
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 10220 13379 10278 13385
rect 10220 13345 10232 13379
rect 10266 13376 10278 13379
rect 10962 13376 10968 13388
rect 10266 13348 10968 13376
rect 10266 13345 10278 13348
rect 10220 13339 10278 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 12710 13385 12716 13388
rect 12704 13339 12716 13385
rect 12768 13376 12774 13388
rect 15746 13376 15752 13388
rect 12768 13348 12804 13376
rect 15707 13348 15752 13376
rect 12710 13336 12716 13339
rect 12768 13336 12774 13348
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 16758 13376 16764 13388
rect 16719 13348 16764 13376
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13376 19671 13379
rect 20622 13376 20628 13388
rect 19659 13348 20628 13376
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 21536 13379 21594 13385
rect 21536 13345 21548 13379
rect 21582 13376 21594 13379
rect 22002 13376 22008 13388
rect 21582 13348 22008 13376
rect 21582 13345 21594 13348
rect 21536 13339 21594 13345
rect 22002 13336 22008 13348
rect 22060 13336 22066 13388
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 5258 13308 5264 13320
rect 5123 13280 5264 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 6604 13280 6653 13308
rect 6604 13268 6610 13280
rect 6641 13277 6653 13280
rect 6687 13308 6699 13311
rect 7006 13308 7012 13320
rect 6687 13280 7012 13308
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 8754 13308 8760 13320
rect 8711 13280 8760 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 8754 13268 8760 13280
rect 8812 13308 8818 13320
rect 9398 13308 9404 13320
rect 8812 13280 9404 13308
rect 8812 13268 8818 13280
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 9950 13308 9956 13320
rect 9911 13280 9956 13308
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 19889 13311 19947 13317
rect 12492 13280 12537 13308
rect 12492 13268 12498 13280
rect 19889 13277 19901 13311
rect 19935 13308 19947 13311
rect 20438 13308 20444 13320
rect 19935 13280 20444 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 21266 13308 21272 13320
rect 21227 13280 21272 13308
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 7190 13200 7196 13252
rect 7248 13240 7254 13252
rect 8021 13243 8079 13249
rect 8021 13240 8033 13243
rect 7248 13212 8033 13240
rect 7248 13200 7254 13212
rect 8021 13209 8033 13212
rect 8067 13209 8079 13243
rect 8021 13203 8079 13209
rect 18141 13243 18199 13249
rect 18141 13209 18153 13243
rect 18187 13240 18199 13243
rect 18782 13240 18788 13252
rect 18187 13212 18788 13240
rect 18187 13209 18199 13212
rect 18141 13203 18199 13209
rect 18782 13200 18788 13212
rect 18840 13200 18846 13252
rect 22664 13240 22692 13416
rect 23198 13404 23204 13456
rect 23256 13444 23262 13456
rect 24213 13447 24271 13453
rect 24213 13444 24225 13447
rect 23256 13416 24225 13444
rect 23256 13404 23262 13416
rect 24213 13413 24225 13416
rect 24259 13444 24271 13447
rect 25038 13444 25044 13456
rect 24259 13416 25044 13444
rect 24259 13413 24271 13416
rect 24213 13407 24271 13413
rect 25038 13404 25044 13416
rect 25096 13404 25102 13456
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 24026 13376 24032 13388
rect 23624 13348 24032 13376
rect 23624 13336 23630 13348
rect 24026 13336 24032 13348
rect 24084 13376 24090 13388
rect 24084 13348 24348 13376
rect 24084 13336 24090 13348
rect 24320 13317 24348 13348
rect 25222 13336 25228 13388
rect 25280 13376 25286 13388
rect 25317 13379 25375 13385
rect 25317 13376 25329 13379
rect 25280 13348 25329 13376
rect 25280 13336 25286 13348
rect 25317 13345 25329 13348
rect 25363 13345 25375 13379
rect 25317 13339 25375 13345
rect 24305 13311 24363 13317
rect 24305 13277 24317 13311
rect 24351 13277 24363 13311
rect 24305 13271 24363 13277
rect 25866 13240 25872 13252
rect 22664 13212 25872 13240
rect 25866 13200 25872 13212
rect 25924 13200 25930 13252
rect 3142 13172 3148 13184
rect 3103 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 11330 13172 11336 13184
rect 11291 13144 11336 13172
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12161 13175 12219 13181
rect 12161 13172 12173 13175
rect 12124 13144 12173 13172
rect 12124 13132 12130 13144
rect 12161 13141 12173 13144
rect 12207 13141 12219 13175
rect 15470 13172 15476 13184
rect 15431 13144 15476 13172
rect 12161 13135 12219 13141
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 16298 13172 16304 13184
rect 16259 13144 16304 13172
rect 16298 13132 16304 13144
rect 16356 13132 16362 13184
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 19208 13144 19257 13172
rect 19208 13132 19214 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 20254 13172 20260 13184
rect 20215 13144 20260 13172
rect 19245 13135 19303 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 23290 13172 23296 13184
rect 23251 13144 23296 13172
rect 23290 13132 23296 13144
rect 23348 13132 23354 13184
rect 23750 13172 23756 13184
rect 23711 13144 23756 13172
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 25498 13172 25504 13184
rect 25459 13144 25504 13172
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 1544 12940 1593 12968
rect 1544 12928 1550 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 3513 12971 3571 12977
rect 3513 12937 3525 12971
rect 3559 12968 3571 12971
rect 3602 12968 3608 12980
rect 3559 12940 3608 12968
rect 3559 12937 3571 12940
rect 3513 12931 3571 12937
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 4798 12928 4804 12980
rect 4856 12968 4862 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4856 12940 5181 12968
rect 4856 12928 4862 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 6270 12968 6276 12980
rect 6231 12940 6276 12968
rect 5169 12931 5227 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6822 12968 6828 12980
rect 6420 12940 6828 12968
rect 6420 12928 6426 12940
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8294 12968 8300 12980
rect 8159 12940 8300 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 8478 12968 8484 12980
rect 8439 12940 8484 12968
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 8846 12928 8852 12980
rect 8904 12968 8910 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 8904 12940 9321 12968
rect 8904 12928 8910 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 10008 12940 10333 12968
rect 10008 12928 10014 12940
rect 10321 12937 10333 12940
rect 10367 12968 10379 12971
rect 10686 12968 10692 12980
rect 10367 12940 10692 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 10962 12968 10968 12980
rect 10827 12940 10968 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12986 12968 12992 12980
rect 12492 12940 12992 12968
rect 12492 12928 12498 12940
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15059 12940 15608 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 2682 12900 2688 12912
rect 2643 12872 2688 12900
rect 2682 12860 2688 12872
rect 2740 12860 2746 12912
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3145 12903 3203 12909
rect 3145 12900 3157 12903
rect 2832 12872 3157 12900
rect 2832 12860 2838 12872
rect 3145 12869 3157 12872
rect 3191 12900 3203 12903
rect 4338 12900 4344 12912
rect 3191 12872 4344 12900
rect 3191 12869 3203 12872
rect 3145 12863 3203 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 4982 12900 4988 12912
rect 4943 12872 4988 12900
rect 4982 12860 4988 12872
rect 5040 12900 5046 12912
rect 6288 12900 6316 12928
rect 5040 12872 5672 12900
rect 6288 12872 7420 12900
rect 5040 12860 5046 12872
rect 5644 12841 5672 12872
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 6086 12832 6092 12844
rect 5859 12804 6092 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6086 12792 6092 12804
rect 6144 12792 6150 12844
rect 6178 12792 6184 12844
rect 6236 12832 6242 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6236 12804 6561 12832
rect 6236 12792 6242 12804
rect 6549 12801 6561 12804
rect 6595 12832 6607 12835
rect 6595 12804 6868 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12733 1455 12767
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 1397 12727 1455 12733
rect 2332 12736 2513 12764
rect 1412 12696 1440 12727
rect 2038 12696 2044 12708
rect 1412 12668 2044 12696
rect 2038 12656 2044 12668
rect 2096 12656 2102 12708
rect 2332 12640 2360 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 3602 12764 3608 12776
rect 3563 12736 3608 12764
rect 2501 12727 2559 12733
rect 3602 12724 3608 12736
rect 3660 12724 3666 12776
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 5258 12764 5264 12776
rect 4387 12736 5264 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 5534 12764 5540 12776
rect 5447 12736 5540 12764
rect 5534 12724 5540 12736
rect 5592 12764 5598 12776
rect 6638 12764 6644 12776
rect 5592 12736 6644 12764
rect 5592 12724 5598 12736
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 6840 12764 6868 12804
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 7282 12832 7288 12844
rect 6972 12804 7288 12832
rect 6972 12792 6978 12804
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7392 12841 7420 12872
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 15105 12903 15163 12909
rect 15105 12900 15117 12903
rect 14884 12872 15117 12900
rect 14884 12860 14890 12872
rect 15105 12869 15117 12872
rect 15151 12869 15163 12903
rect 15580 12900 15608 12940
rect 16206 12928 16212 12980
rect 16264 12968 16270 12980
rect 16390 12968 16396 12980
rect 16264 12940 16396 12968
rect 16264 12928 16270 12940
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16758 12968 16764 12980
rect 16719 12940 16764 12968
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17129 12971 17187 12977
rect 17129 12937 17141 12971
rect 17175 12968 17187 12971
rect 17862 12968 17868 12980
rect 17175 12940 17868 12968
rect 17175 12937 17187 12940
rect 17129 12931 17187 12937
rect 17862 12928 17868 12940
rect 17920 12928 17926 12980
rect 18046 12968 18052 12980
rect 18007 12940 18052 12968
rect 18046 12928 18052 12940
rect 18104 12928 18110 12980
rect 19337 12971 19395 12977
rect 19337 12937 19349 12971
rect 19383 12968 19395 12971
rect 19702 12968 19708 12980
rect 19383 12940 19708 12968
rect 19383 12937 19395 12940
rect 19337 12931 19395 12937
rect 19702 12928 19708 12940
rect 19760 12968 19766 12980
rect 20162 12968 20168 12980
rect 19760 12940 20168 12968
rect 19760 12928 19766 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20622 12968 20628 12980
rect 20583 12940 20628 12968
rect 20622 12928 20628 12940
rect 20680 12968 20686 12980
rect 20898 12968 20904 12980
rect 20680 12940 20904 12968
rect 20680 12928 20686 12940
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21910 12968 21916 12980
rect 21871 12940 21916 12968
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 23290 12968 23296 12980
rect 22388 12940 23296 12968
rect 15580 12872 15700 12900
rect 15105 12863 15163 12869
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9456 12804 9873 12832
rect 9456 12792 9462 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 13722 12832 13728 12844
rect 12575 12804 13728 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 15672 12841 15700 12872
rect 20346 12860 20352 12912
rect 20404 12900 20410 12912
rect 22094 12900 22100 12912
rect 20404 12872 22100 12900
rect 20404 12860 20410 12872
rect 22094 12860 22100 12872
rect 22152 12860 22158 12912
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12832 14703 12835
rect 15657 12835 15715 12841
rect 14691 12804 15608 12832
rect 14691 12801 14703 12804
rect 14645 12795 14703 12801
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6840 12736 7205 12764
rect 7193 12733 7205 12736
rect 7239 12764 7251 12767
rect 8110 12764 8116 12776
rect 7239 12736 8116 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 9140 12736 9689 12764
rect 9140 12708 9168 12736
rect 9677 12733 9689 12736
rect 9723 12764 9735 12767
rect 9950 12764 9956 12776
rect 9723 12736 9956 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 9950 12724 9956 12736
rect 10008 12724 10014 12776
rect 13446 12764 13452 12776
rect 13359 12736 13452 12764
rect 13446 12724 13452 12736
rect 13504 12764 13510 12776
rect 13998 12764 14004 12776
rect 13504 12736 14004 12764
rect 13504 12724 13510 12736
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 15470 12764 15476 12776
rect 15431 12736 15476 12764
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 15580 12773 15608 12804
rect 15657 12801 15669 12835
rect 15703 12832 15715 12835
rect 16298 12832 16304 12844
rect 15703 12804 16304 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 18230 12832 18236 12844
rect 17543 12804 18236 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 18230 12792 18236 12804
rect 18288 12832 18294 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18288 12804 18613 12832
rect 18288 12792 18294 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 18601 12795 18659 12801
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12832 21879 12835
rect 22278 12832 22284 12844
rect 21867 12804 22284 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 22388 12841 22416 12940
rect 23290 12928 23296 12940
rect 23348 12968 23354 12980
rect 23661 12971 23719 12977
rect 23661 12968 23673 12971
rect 23348 12940 23673 12968
rect 23348 12928 23354 12940
rect 23661 12937 23673 12940
rect 23707 12937 23719 12971
rect 23661 12931 23719 12937
rect 24026 12928 24032 12980
rect 24084 12968 24090 12980
rect 24673 12971 24731 12977
rect 24673 12968 24685 12971
rect 24084 12940 24685 12968
rect 24084 12928 24090 12940
rect 24673 12937 24685 12940
rect 24719 12937 24731 12971
rect 25038 12968 25044 12980
rect 24999 12940 25044 12968
rect 24673 12931 24731 12937
rect 25038 12928 25044 12940
rect 25096 12928 25102 12980
rect 25222 12928 25228 12980
rect 25280 12968 25286 12980
rect 26145 12971 26203 12977
rect 26145 12968 26157 12971
rect 25280 12940 26157 12968
rect 25280 12928 25286 12940
rect 26145 12937 26157 12940
rect 26191 12937 26203 12971
rect 26145 12931 26203 12937
rect 22738 12860 22744 12912
rect 22796 12900 22802 12912
rect 22922 12900 22928 12912
rect 22796 12872 22928 12900
rect 22796 12860 22802 12872
rect 22922 12860 22928 12872
rect 22980 12900 22986 12912
rect 23017 12903 23075 12909
rect 23017 12900 23029 12903
rect 22980 12872 23029 12900
rect 22980 12860 22986 12872
rect 23017 12869 23029 12872
rect 23063 12900 23075 12903
rect 24486 12900 24492 12912
rect 23063 12872 24492 12900
rect 23063 12869 23075 12872
rect 23017 12863 23075 12869
rect 22373 12835 22431 12841
rect 22373 12801 22385 12835
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12832 22615 12835
rect 23382 12832 23388 12844
rect 22603 12804 23388 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 15565 12767 15623 12773
rect 15565 12733 15577 12767
rect 15611 12764 15623 12767
rect 15930 12764 15936 12776
rect 15611 12736 15936 12764
rect 15611 12733 15623 12736
rect 15565 12727 15623 12733
rect 15930 12724 15936 12736
rect 15988 12724 15994 12776
rect 16942 12764 16948 12776
rect 16903 12736 16948 12764
rect 16942 12724 16948 12736
rect 17000 12724 17006 12776
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 20622 12764 20628 12776
rect 20119 12736 20628 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 20622 12724 20628 12736
rect 20680 12724 20686 12776
rect 22002 12724 22008 12776
rect 22060 12764 22066 12776
rect 22572 12764 22600 12795
rect 23382 12792 23388 12804
rect 23440 12792 23446 12844
rect 24136 12841 24164 12872
rect 24486 12860 24492 12872
rect 24544 12860 24550 12912
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24302 12832 24308 12844
rect 24263 12804 24308 12832
rect 24121 12795 24179 12801
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 22060 12736 22600 12764
rect 22060 12724 22066 12736
rect 25038 12724 25044 12776
rect 25096 12764 25102 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 25096 12736 25237 12764
rect 25096 12724 25102 12736
rect 25225 12733 25237 12736
rect 25271 12764 25283 12767
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 25271 12736 25789 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25777 12733 25789 12736
rect 25823 12733 25835 12767
rect 25777 12727 25835 12733
rect 2590 12656 2596 12708
rect 2648 12696 2654 12708
rect 4709 12699 4767 12705
rect 2648 12668 3832 12696
rect 2648 12656 2654 12668
rect 2314 12628 2320 12640
rect 2275 12600 2320 12628
rect 2314 12588 2320 12600
rect 2372 12588 2378 12640
rect 3804 12637 3832 12668
rect 4709 12665 4721 12699
rect 4755 12696 4767 12699
rect 6086 12696 6092 12708
rect 4755 12668 6092 12696
rect 4755 12665 4767 12668
rect 4709 12659 4767 12665
rect 6086 12656 6092 12668
rect 6144 12656 6150 12708
rect 9122 12696 9128 12708
rect 9083 12668 9128 12696
rect 9122 12656 9128 12668
rect 9180 12656 9186 12708
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 9640 12668 10977 12696
rect 9640 12656 9646 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 10965 12659 11023 12665
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 11204 12668 12848 12696
rect 11204 12656 11210 12668
rect 3789 12631 3847 12637
rect 3789 12597 3801 12631
rect 3835 12597 3847 12631
rect 3789 12591 3847 12597
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12628 9827 12631
rect 9858 12628 9864 12640
rect 9815 12600 9864 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 11664 12600 12173 12628
rect 11664 12588 11670 12600
rect 12161 12597 12173 12600
rect 12207 12628 12219 12631
rect 12434 12628 12440 12640
rect 12207 12600 12440 12628
rect 12207 12597 12219 12600
rect 12161 12591 12219 12597
rect 12434 12588 12440 12600
rect 12492 12628 12498 12640
rect 12710 12628 12716 12640
rect 12492 12600 12716 12628
rect 12492 12588 12498 12600
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 12820 12628 12848 12668
rect 18322 12656 18328 12708
rect 18380 12696 18386 12708
rect 18417 12699 18475 12705
rect 18417 12696 18429 12699
rect 18380 12668 18429 12696
rect 18380 12656 18386 12668
rect 18417 12665 18429 12668
rect 18463 12665 18475 12699
rect 18417 12659 18475 12665
rect 19981 12699 20039 12705
rect 19981 12665 19993 12699
rect 20027 12696 20039 12699
rect 20714 12696 20720 12708
rect 20027 12668 20720 12696
rect 20027 12665 20039 12668
rect 19981 12659 20039 12665
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 22278 12696 22284 12708
rect 22239 12668 22284 12696
rect 22278 12656 22284 12668
rect 22336 12656 22342 12708
rect 22370 12656 22376 12708
rect 22428 12696 22434 12708
rect 23385 12699 23443 12705
rect 23385 12696 23397 12699
rect 22428 12668 23397 12696
rect 22428 12656 22434 12668
rect 23385 12665 23397 12668
rect 23431 12696 23443 12699
rect 24029 12699 24087 12705
rect 24029 12696 24041 12699
rect 23431 12668 24041 12696
rect 23431 12665 23443 12668
rect 23385 12659 23443 12665
rect 24029 12665 24041 12668
rect 24075 12665 24087 12699
rect 24029 12659 24087 12665
rect 13814 12628 13820 12640
rect 12820 12600 13820 12628
rect 13814 12588 13820 12600
rect 13872 12628 13878 12640
rect 13909 12631 13967 12637
rect 13909 12628 13921 12631
rect 13872 12600 13921 12628
rect 13872 12588 13878 12600
rect 13909 12597 13921 12600
rect 13955 12628 13967 12631
rect 16114 12628 16120 12640
rect 13955 12600 16120 12628
rect 13955 12597 13967 12600
rect 13909 12591 13967 12597
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 17460 12600 17785 12628
rect 17460 12588 17466 12600
rect 17773 12597 17785 12600
rect 17819 12628 17831 12631
rect 18506 12628 18512 12640
rect 17819 12600 18512 12628
rect 17819 12597 17831 12600
rect 17773 12591 17831 12597
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 19518 12588 19524 12640
rect 19576 12628 19582 12640
rect 19613 12631 19671 12637
rect 19613 12628 19625 12631
rect 19576 12600 19625 12628
rect 19576 12588 19582 12600
rect 19613 12597 19625 12600
rect 19659 12597 19671 12631
rect 19613 12591 19671 12597
rect 21266 12588 21272 12640
rect 21324 12628 21330 12640
rect 21361 12631 21419 12637
rect 21361 12628 21373 12631
rect 21324 12600 21373 12628
rect 21324 12588 21330 12600
rect 21361 12597 21373 12600
rect 21407 12628 21419 12631
rect 21910 12628 21916 12640
rect 21407 12600 21916 12628
rect 21407 12597 21419 12600
rect 21361 12591 21419 12597
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 25406 12628 25412 12640
rect 25367 12600 25412 12628
rect 25406 12588 25412 12600
rect 25464 12588 25470 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1762 12424 1768 12436
rect 1723 12396 1768 12424
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 2130 12424 2136 12436
rect 2091 12396 2136 12424
rect 2130 12384 2136 12396
rect 2188 12424 2194 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2188 12396 2881 12424
rect 2188 12384 2194 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 3234 12424 3240 12436
rect 3195 12396 3240 12424
rect 2869 12387 2927 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4614 12424 4620 12436
rect 3927 12396 4620 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 4798 12424 4804 12436
rect 4759 12396 4804 12424
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5626 12424 5632 12436
rect 5587 12396 5632 12424
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 7156 12396 7205 12424
rect 7156 12384 7162 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7193 12387 7251 12393
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8352 12396 8953 12424
rect 8352 12384 8358 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 8941 12387 8999 12393
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9858 12424 9864 12436
rect 9447 12396 9864 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 1394 12316 1400 12368
rect 1452 12356 1458 12368
rect 2501 12359 2559 12365
rect 2501 12356 2513 12359
rect 1452 12328 2513 12356
rect 1452 12316 1458 12328
rect 2501 12325 2513 12328
rect 2547 12325 2559 12359
rect 2501 12319 2559 12325
rect 4525 12359 4583 12365
rect 4525 12325 4537 12359
rect 4571 12356 4583 12359
rect 4890 12356 4896 12368
rect 4571 12328 4896 12356
rect 4571 12325 4583 12328
rect 4525 12319 4583 12325
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 8956 12356 8984 12387
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12492 12396 12909 12424
rect 12492 12384 12498 12396
rect 12897 12393 12909 12396
rect 12943 12393 12955 12427
rect 12897 12387 12955 12393
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 18049 12427 18107 12433
rect 18049 12424 18061 12427
rect 16724 12396 18061 12424
rect 16724 12384 16730 12396
rect 18049 12393 18061 12396
rect 18095 12424 18107 12427
rect 18322 12424 18328 12436
rect 18095 12396 18328 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 18656 12396 19717 12424
rect 18656 12384 18662 12396
rect 19705 12393 19717 12396
rect 19751 12424 19763 12427
rect 20254 12424 20260 12436
rect 19751 12396 20260 12424
rect 19751 12393 19763 12396
rect 19705 12387 19763 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 21450 12424 21456 12436
rect 21411 12396 21456 12424
rect 21450 12384 21456 12396
rect 21508 12384 21514 12436
rect 22002 12424 22008 12436
rect 21928 12396 22008 12424
rect 10137 12359 10195 12365
rect 10137 12356 10149 12359
rect 8956 12328 10149 12356
rect 10137 12325 10149 12328
rect 10183 12325 10195 12359
rect 10137 12319 10195 12325
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11388 12328 11652 12356
rect 11388 12316 11394 12328
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12288 1639 12291
rect 1854 12288 1860 12300
rect 1627 12260 1860 12288
rect 1627 12257 1639 12260
rect 1581 12251 1639 12257
rect 1854 12248 1860 12260
rect 1912 12288 1918 12300
rect 2590 12288 2596 12300
rect 1912 12260 2596 12288
rect 1912 12248 1918 12260
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 2685 12291 2743 12297
rect 2685 12257 2697 12291
rect 2731 12288 2743 12291
rect 2774 12288 2780 12300
rect 2731 12260 2780 12288
rect 2731 12257 2743 12260
rect 2685 12251 2743 12257
rect 2774 12248 2780 12260
rect 2832 12288 2838 12300
rect 3326 12288 3332 12300
rect 2832 12260 3332 12288
rect 2832 12248 2838 12260
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5442 12288 5448 12300
rect 5307 12260 5448 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5994 12288 6000 12300
rect 5955 12260 6000 12288
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 6362 12288 6368 12300
rect 6135 12260 6368 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 7558 12288 7564 12300
rect 7519 12260 7564 12288
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10686 12248 10692 12300
rect 10744 12288 10750 12300
rect 11514 12288 11520 12300
rect 10744 12260 11520 12288
rect 10744 12248 10750 12260
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 11624 12288 11652 12328
rect 14642 12316 14648 12368
rect 14700 12356 14706 12368
rect 18340 12356 18368 12384
rect 18874 12356 18880 12368
rect 14700 12328 15599 12356
rect 18340 12328 18880 12356
rect 14700 12316 14706 12328
rect 11790 12297 11796 12300
rect 11784 12288 11796 12297
rect 11624 12260 11796 12288
rect 11784 12251 11796 12260
rect 11790 12248 11796 12251
rect 11848 12248 11854 12300
rect 14001 12291 14059 12297
rect 14001 12257 14013 12291
rect 14047 12288 14059 12291
rect 14090 12288 14096 12300
rect 14047 12260 14096 12288
rect 14047 12257 14059 12260
rect 14001 12251 14059 12257
rect 14090 12248 14096 12260
rect 14148 12288 14154 12300
rect 14660 12288 14688 12316
rect 14148 12260 14688 12288
rect 15289 12291 15347 12297
rect 14148 12248 14154 12260
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15378 12288 15384 12300
rect 15335 12260 15384 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15571 12297 15599 12328
rect 18874 12316 18880 12328
rect 18932 12316 18938 12368
rect 15556 12291 15614 12297
rect 15556 12257 15568 12291
rect 15602 12288 15614 12291
rect 16850 12288 16856 12300
rect 15602 12260 16856 12288
rect 15602 12257 15614 12260
rect 15556 12251 15614 12257
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 17770 12248 17776 12300
rect 17828 12288 17834 12300
rect 18592 12291 18650 12297
rect 18592 12288 18604 12291
rect 17828 12260 18604 12288
rect 17828 12248 17834 12260
rect 18592 12257 18604 12260
rect 18638 12288 18650 12291
rect 20438 12288 20444 12300
rect 18638 12260 20444 12288
rect 18638 12257 18650 12260
rect 18592 12251 18650 12257
rect 20438 12248 20444 12260
rect 20496 12248 20502 12300
rect 20714 12288 20720 12300
rect 20675 12260 20720 12288
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 21266 12288 21272 12300
rect 21227 12260 21272 12288
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 6270 12220 6276 12232
rect 6183 12192 6276 12220
rect 6270 12180 6276 12192
rect 6328 12220 6334 12232
rect 6730 12220 6736 12232
rect 6328 12192 6736 12220
rect 6328 12180 6334 12192
rect 6730 12180 6736 12192
rect 6788 12180 6794 12232
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 7650 12220 7656 12232
rect 7340 12192 7656 12220
rect 7340 12180 7346 12192
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 6638 12112 6644 12164
rect 6696 12152 6702 12164
rect 7466 12152 7472 12164
rect 6696 12124 7472 12152
rect 6696 12112 6702 12124
rect 7466 12112 7472 12124
rect 7524 12152 7530 12164
rect 7760 12152 7788 12183
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10192 12192 10241 12220
rect 10192 12180 10198 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 14182 12220 14188 12232
rect 14143 12192 14188 12220
rect 10229 12183 10287 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 18322 12220 18328 12232
rect 18283 12192 18328 12220
rect 18322 12180 18328 12192
rect 18380 12180 18386 12232
rect 21928 12229 21956 12396
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 23382 12384 23388 12436
rect 23440 12424 23446 12436
rect 23753 12427 23811 12433
rect 23753 12424 23765 12427
rect 23440 12396 23765 12424
rect 23440 12384 23446 12396
rect 23753 12393 23765 12396
rect 23799 12393 23811 12427
rect 24302 12424 24308 12436
rect 24263 12396 24308 12424
rect 23753 12387 23811 12393
rect 24302 12384 24308 12396
rect 24360 12384 24366 12436
rect 24670 12384 24676 12436
rect 24728 12424 24734 12436
rect 25317 12427 25375 12433
rect 25317 12424 25329 12427
rect 24728 12396 25329 12424
rect 24728 12384 24734 12396
rect 22640 12359 22698 12365
rect 22640 12325 22652 12359
rect 22686 12356 22698 12359
rect 23198 12356 23204 12368
rect 22686 12328 23204 12356
rect 22686 12325 22698 12328
rect 22640 12319 22698 12325
rect 23198 12316 23204 12328
rect 23256 12356 23262 12368
rect 24320 12356 24348 12384
rect 23256 12328 24348 12356
rect 23256 12316 23262 12328
rect 25056 12232 25084 12396
rect 25317 12393 25329 12396
rect 25363 12393 25375 12427
rect 25317 12387 25375 12393
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 25590 12288 25596 12300
rect 25271 12260 25596 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 25590 12248 25596 12260
rect 25648 12248 25654 12300
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12220 21235 12223
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21223 12192 21925 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 22094 12180 22100 12232
rect 22152 12220 22158 12232
rect 22373 12223 22431 12229
rect 22373 12220 22385 12223
rect 22152 12192 22385 12220
rect 22152 12180 22158 12192
rect 22373 12189 22385 12192
rect 22419 12189 22431 12223
rect 22373 12183 22431 12189
rect 25038 12180 25044 12232
rect 25096 12180 25102 12232
rect 25406 12220 25412 12232
rect 25367 12192 25412 12220
rect 25406 12180 25412 12192
rect 25464 12180 25470 12232
rect 7524 12124 7788 12152
rect 7524 12112 7530 12124
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 8665 12155 8723 12161
rect 8665 12152 8677 12155
rect 8628 12124 8677 12152
rect 8628 12112 8634 12124
rect 8665 12121 8677 12124
rect 8711 12152 8723 12155
rect 9677 12155 9735 12161
rect 9677 12152 9689 12155
rect 8711 12124 9689 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 9677 12121 9689 12124
rect 9723 12121 9735 12155
rect 9677 12115 9735 12121
rect 10873 12155 10931 12161
rect 10873 12121 10885 12155
rect 10919 12152 10931 12155
rect 11422 12152 11428 12164
rect 10919 12124 11428 12152
rect 10919 12121 10931 12124
rect 10873 12115 10931 12121
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 24394 12112 24400 12164
rect 24452 12152 24458 12164
rect 24857 12155 24915 12161
rect 24857 12152 24869 12155
rect 24452 12124 24869 12152
rect 24452 12112 24458 12124
rect 24857 12121 24869 12124
rect 24903 12121 24915 12155
rect 24857 12115 24915 12121
rect 6914 12084 6920 12096
rect 6875 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 8294 12084 8300 12096
rect 8255 12056 8300 12084
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 11238 12084 11244 12096
rect 11199 12056 11244 12084
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 13633 12087 13691 12093
rect 13633 12053 13645 12087
rect 13679 12084 13691 12087
rect 13814 12084 13820 12096
rect 13679 12056 13820 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 16206 12084 16212 12096
rect 15151 12056 16212 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16666 12084 16672 12096
rect 16627 12056 16672 12084
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17313 12087 17371 12093
rect 17313 12084 17325 12087
rect 17000 12056 17325 12084
rect 17000 12044 17006 12056
rect 17313 12053 17325 12056
rect 17359 12084 17371 12087
rect 17862 12084 17868 12096
rect 17359 12056 17868 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 20349 12087 20407 12093
rect 20349 12053 20361 12087
rect 20395 12084 20407 12087
rect 20438 12084 20444 12096
rect 20395 12056 20444 12084
rect 20395 12053 20407 12056
rect 20349 12047 20407 12053
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 22738 12084 22744 12096
rect 21416 12056 22744 12084
rect 21416 12044 21422 12056
rect 22738 12044 22744 12056
rect 22796 12044 22802 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2314 11880 2320 11892
rect 1627 11852 2320 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 4985 11883 5043 11889
rect 2832 11852 2877 11880
rect 2832 11840 2838 11852
rect 4985 11849 4997 11883
rect 5031 11880 5043 11883
rect 5166 11880 5172 11892
rect 5031 11852 5172 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 6089 11883 6147 11889
rect 6089 11849 6101 11883
rect 6135 11880 6147 11883
rect 6454 11880 6460 11892
rect 6135 11852 6460 11880
rect 6135 11849 6147 11852
rect 6089 11843 6147 11849
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 6638 11880 6644 11892
rect 6599 11852 6644 11880
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 7193 11883 7251 11889
rect 7193 11849 7205 11883
rect 7239 11880 7251 11883
rect 7558 11880 7564 11892
rect 7239 11852 7564 11880
rect 7239 11849 7251 11852
rect 7193 11843 7251 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9217 11883 9275 11889
rect 9217 11880 9229 11883
rect 9088 11852 9229 11880
rect 9088 11840 9094 11852
rect 9217 11849 9229 11852
rect 9263 11849 9275 11883
rect 9217 11843 9275 11849
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10100 11852 10241 11880
rect 10100 11840 10106 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 10778 11880 10784 11892
rect 10739 11852 10784 11880
rect 10229 11843 10287 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11572 11852 11805 11880
rect 11572 11840 11578 11852
rect 11793 11849 11805 11852
rect 11839 11880 11851 11883
rect 12158 11880 12164 11892
rect 11839 11852 12164 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 12158 11840 12164 11852
rect 12216 11880 12222 11892
rect 12986 11880 12992 11892
rect 12216 11852 12992 11880
rect 12216 11840 12222 11852
rect 12986 11840 12992 11852
rect 13044 11880 13050 11892
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 13044 11852 13093 11880
rect 13044 11840 13050 11852
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 13081 11843 13139 11849
rect 1854 11812 1860 11824
rect 1815 11784 1860 11812
rect 1854 11772 1860 11784
rect 1912 11772 1918 11824
rect 1946 11772 1952 11824
rect 2004 11812 2010 11824
rect 2225 11815 2283 11821
rect 2225 11812 2237 11815
rect 2004 11784 2237 11812
rect 2004 11772 2010 11784
rect 2225 11781 2237 11784
rect 2271 11781 2283 11815
rect 2225 11775 2283 11781
rect 4617 11815 4675 11821
rect 4617 11781 4629 11815
rect 4663 11812 4675 11815
rect 5350 11812 5356 11824
rect 4663 11784 5356 11812
rect 4663 11781 4675 11784
rect 4617 11775 4675 11781
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 5721 11815 5779 11821
rect 5721 11781 5733 11815
rect 5767 11812 5779 11815
rect 6270 11812 6276 11824
rect 5767 11784 6276 11812
rect 5767 11781 5779 11784
rect 5721 11775 5779 11781
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 7653 11815 7711 11821
rect 7653 11812 7665 11815
rect 6420 11784 7665 11812
rect 6420 11772 6426 11784
rect 7653 11781 7665 11784
rect 7699 11781 7711 11815
rect 12250 11812 12256 11824
rect 7653 11775 7711 11781
rect 9784 11784 12256 11812
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1964 11676 1992 11772
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 6380 11744 6408 11772
rect 5307 11716 6408 11744
rect 7561 11747 7619 11753
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 7561 11713 7573 11747
rect 7607 11744 7619 11747
rect 7742 11744 7748 11756
rect 7607 11716 7748 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 7742 11704 7748 11716
rect 7800 11744 7806 11756
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7800 11716 8125 11744
rect 7800 11704 7806 11716
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 8570 11744 8576 11756
rect 8343 11716 8576 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8570 11704 8576 11716
rect 8628 11744 8634 11756
rect 8757 11747 8815 11753
rect 8757 11744 8769 11747
rect 8628 11716 8769 11744
rect 8628 11704 8634 11716
rect 8757 11713 8769 11716
rect 8803 11744 8815 11747
rect 9214 11744 9220 11756
rect 8803 11716 9220 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 9784 11753 9812 11784
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9364 11716 9781 11744
rect 9364 11704 9370 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11054 11744 11060 11756
rect 10836 11716 11060 11744
rect 10836 11704 10842 11716
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 11238 11744 11244 11756
rect 11199 11716 11244 11744
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11422 11744 11428 11756
rect 11383 11716 11428 11744
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 13096 11744 13124 11843
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 15528 11852 15761 11880
rect 15528 11840 15534 11852
rect 15749 11849 15761 11852
rect 15795 11849 15807 11883
rect 22646 11880 22652 11892
rect 22607 11852 22652 11880
rect 15749 11843 15807 11849
rect 22646 11840 22652 11852
rect 22704 11840 22710 11892
rect 23474 11880 23480 11892
rect 23435 11852 23480 11880
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 23658 11880 23664 11892
rect 23619 11852 23664 11880
rect 23658 11840 23664 11852
rect 23716 11840 23722 11892
rect 24949 11883 25007 11889
rect 24949 11849 24961 11883
rect 24995 11880 25007 11883
rect 25038 11880 25044 11892
rect 24995 11852 25044 11880
rect 24995 11849 25007 11852
rect 24949 11843 25007 11849
rect 25038 11840 25044 11852
rect 25096 11840 25102 11892
rect 25409 11883 25467 11889
rect 25409 11849 25421 11883
rect 25455 11880 25467 11883
rect 25682 11880 25688 11892
rect 25455 11852 25688 11880
rect 25455 11849 25467 11852
rect 25409 11843 25467 11849
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 16080 11784 16436 11812
rect 16080 11772 16086 11784
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 13096 11716 13277 11744
rect 13265 11713 13277 11716
rect 13311 11713 13323 11747
rect 16206 11744 16212 11756
rect 16167 11716 16212 11744
rect 13265 11707 13323 11713
rect 1443 11648 1992 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 8021 11679 8079 11685
rect 8021 11676 8033 11679
rect 7984 11648 8033 11676
rect 7984 11636 7990 11648
rect 8021 11645 8033 11648
rect 8067 11645 8079 11679
rect 8021 11639 8079 11645
rect 9125 11679 9183 11685
rect 9125 11645 9137 11679
rect 9171 11676 9183 11679
rect 9490 11676 9496 11688
rect 9171 11648 9496 11676
rect 9171 11645 9183 11648
rect 9125 11639 9183 11645
rect 9490 11636 9496 11648
rect 9548 11676 9554 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9548 11648 9597 11676
rect 9548 11636 9554 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 11146 11676 11152 11688
rect 10735 11648 11152 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 13280 11676 13308 11707
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 16408 11753 16436 11784
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 18049 11815 18107 11821
rect 18049 11812 18061 11815
rect 18012 11784 18061 11812
rect 18012 11772 18018 11784
rect 18049 11781 18061 11784
rect 18095 11781 18107 11815
rect 18049 11775 18107 11781
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11744 16451 11747
rect 16666 11744 16672 11756
rect 16439 11716 16672 11744
rect 16439 11713 16451 11716
rect 16393 11707 16451 11713
rect 16666 11704 16672 11716
rect 16724 11704 16730 11756
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17497 11747 17555 11753
rect 17497 11744 17509 11747
rect 16908 11716 17509 11744
rect 16908 11704 16914 11716
rect 17497 11713 17509 11716
rect 17543 11744 17555 11747
rect 18230 11744 18236 11756
rect 17543 11716 18236 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 18230 11704 18236 11716
rect 18288 11744 18294 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18288 11716 18613 11744
rect 18288 11704 18294 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11744 22063 11747
rect 23198 11744 23204 11756
rect 22051 11716 23204 11744
rect 22051 11713 22063 11716
rect 22005 11707 22063 11713
rect 23198 11704 23204 11716
rect 23256 11704 23262 11756
rect 23492 11744 23520 11840
rect 24121 11747 24179 11753
rect 24121 11744 24133 11747
rect 23492 11716 24133 11744
rect 24121 11713 24133 11716
rect 24167 11713 24179 11747
rect 24302 11744 24308 11756
rect 24263 11716 24308 11744
rect 24121 11707 24179 11713
rect 24302 11704 24308 11716
rect 24360 11744 24366 11756
rect 25406 11744 25412 11756
rect 24360 11716 25412 11744
rect 24360 11704 24366 11716
rect 25406 11704 25412 11716
rect 25464 11744 25470 11756
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25464 11716 26157 11744
rect 25464 11704 25470 11716
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 15289 11679 15347 11685
rect 15289 11676 15301 11679
rect 13280 11648 15301 11676
rect 15289 11645 15301 11648
rect 15335 11676 15347 11679
rect 15378 11676 15384 11688
rect 15335 11648 15384 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 15378 11636 15384 11648
rect 15436 11636 15442 11688
rect 16114 11676 16120 11688
rect 16075 11648 16120 11676
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 17954 11636 17960 11688
rect 18012 11676 18018 11688
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 18012 11648 18429 11676
rect 18012 11636 18018 11648
rect 18417 11645 18429 11648
rect 18463 11645 18475 11679
rect 18417 11639 18475 11645
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11645 19947 11679
rect 22462 11676 22468 11688
rect 22423 11648 22468 11676
rect 19889 11639 19947 11645
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 9674 11608 9680 11620
rect 8352 11580 9680 11608
rect 8352 11568 8358 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 11790 11568 11796 11620
rect 11848 11608 11854 11620
rect 12161 11611 12219 11617
rect 12161 11608 12173 11611
rect 11848 11580 12173 11608
rect 11848 11568 11854 11580
rect 12161 11577 12173 11580
rect 12207 11577 12219 11611
rect 12161 11571 12219 11577
rect 12805 11611 12863 11617
rect 12805 11577 12817 11611
rect 12851 11608 12863 11611
rect 13532 11611 13590 11617
rect 13532 11608 13544 11611
rect 12851 11580 13544 11608
rect 12851 11577 12863 11580
rect 12805 11571 12863 11577
rect 13532 11577 13544 11580
rect 13578 11608 13590 11611
rect 13722 11608 13728 11620
rect 13578 11580 13728 11608
rect 13578 11577 13590 11580
rect 13532 11571 13590 11577
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 19061 11611 19119 11617
rect 19061 11608 19073 11611
rect 18380 11580 19073 11608
rect 18380 11568 18386 11580
rect 19061 11577 19073 11580
rect 19107 11608 19119 11611
rect 19705 11611 19763 11617
rect 19705 11608 19717 11611
rect 19107 11580 19717 11608
rect 19107 11577 19119 11580
rect 19061 11571 19119 11577
rect 19705 11577 19717 11580
rect 19751 11608 19763 11611
rect 19904 11608 19932 11639
rect 22462 11636 22468 11648
rect 22520 11676 22526 11688
rect 23017 11679 23075 11685
rect 23017 11676 23029 11679
rect 22520 11648 23029 11676
rect 22520 11636 22526 11648
rect 23017 11645 23029 11648
rect 23063 11645 23075 11679
rect 24026 11676 24032 11688
rect 23987 11648 24032 11676
rect 23017 11639 23075 11645
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 25225 11679 25283 11685
rect 25225 11645 25237 11679
rect 25271 11676 25283 11679
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25271 11648 25789 11676
rect 25271 11645 25283 11648
rect 25225 11639 25283 11645
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 20162 11617 20168 11620
rect 20156 11608 20168 11617
rect 19751 11580 19932 11608
rect 20123 11580 20168 11608
rect 19751 11577 19763 11580
rect 19705 11571 19763 11577
rect 20156 11571 20168 11580
rect 20162 11568 20168 11571
rect 20220 11568 20226 11620
rect 22738 11568 22744 11620
rect 22796 11608 22802 11620
rect 25240 11608 25268 11639
rect 22796 11580 25268 11608
rect 22796 11568 22802 11580
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 17402 11540 17408 11552
rect 11388 11512 17408 11540
rect 11388 11500 11394 11512
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17552 11512 17785 11540
rect 17552 11500 17558 11512
rect 17773 11509 17785 11512
rect 17819 11540 17831 11543
rect 18509 11543 18567 11549
rect 18509 11540 18521 11543
rect 17819 11512 18521 11540
rect 17819 11509 17831 11512
rect 17773 11503 17831 11509
rect 18509 11509 18521 11512
rect 18555 11540 18567 11543
rect 19334 11540 19340 11552
rect 18555 11512 19340 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21450 11540 21456 11552
rect 21315 11512 21456 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22281 11543 22339 11549
rect 22281 11540 22293 11543
rect 22152 11512 22293 11540
rect 22152 11500 22158 11512
rect 22281 11509 22293 11512
rect 22327 11509 22339 11543
rect 22281 11503 22339 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 6089 11339 6147 11345
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 6822 11336 6828 11348
rect 6135 11308 6828 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7282 11336 7288 11348
rect 7243 11308 7288 11336
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7745 11339 7803 11345
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 7926 11336 7932 11348
rect 7791 11308 7932 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 8389 11339 8447 11345
rect 8389 11305 8401 11339
rect 8435 11336 8447 11339
rect 8478 11336 8484 11348
rect 8435 11308 8484 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 8478 11296 8484 11308
rect 8536 11336 8542 11348
rect 8938 11336 8944 11348
rect 8536 11308 8944 11336
rect 8536 11296 8542 11308
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9306 11336 9312 11348
rect 9267 11308 9312 11336
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 10965 11339 11023 11345
rect 10965 11305 10977 11339
rect 11011 11336 11023 11339
rect 11238 11336 11244 11348
rect 11011 11308 11244 11336
rect 11011 11305 11023 11308
rect 10965 11299 11023 11305
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 14366 11336 14372 11348
rect 14231 11308 14372 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16356 11308 16681 11336
rect 16356 11296 16362 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 17770 11336 17776 11348
rect 17731 11308 17776 11336
rect 16669 11299 16727 11305
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18049 11339 18107 11345
rect 18049 11336 18061 11339
rect 18012 11308 18061 11336
rect 18012 11296 18018 11308
rect 18049 11305 18061 11308
rect 18095 11305 18107 11339
rect 18049 11299 18107 11305
rect 18506 11296 18512 11348
rect 18564 11336 18570 11348
rect 18782 11336 18788 11348
rect 18564 11308 18788 11336
rect 18564 11296 18570 11308
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 21266 11296 21272 11348
rect 21324 11336 21330 11348
rect 21545 11339 21603 11345
rect 21545 11336 21557 11339
rect 21324 11308 21557 11336
rect 21324 11296 21330 11308
rect 21545 11305 21557 11308
rect 21591 11305 21603 11339
rect 21545 11299 21603 11305
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 23477 11339 23535 11345
rect 23477 11336 23489 11339
rect 23256 11308 23489 11336
rect 23256 11296 23262 11308
rect 23477 11305 23489 11308
rect 23523 11305 23535 11339
rect 24026 11336 24032 11348
rect 23987 11308 24032 11336
rect 23477 11299 23535 11305
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24302 11296 24308 11348
rect 24360 11336 24366 11348
rect 24397 11339 24455 11345
rect 24397 11336 24409 11339
rect 24360 11308 24409 11336
rect 24360 11296 24366 11308
rect 24397 11305 24409 11308
rect 24443 11305 24455 11339
rect 24397 11299 24455 11305
rect 24949 11339 25007 11345
rect 24949 11305 24961 11339
rect 24995 11336 25007 11339
rect 25222 11336 25228 11348
rect 24995 11308 25228 11336
rect 24995 11305 25007 11308
rect 24949 11299 25007 11305
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 9677 11271 9735 11277
rect 9677 11237 9689 11271
rect 9723 11268 9735 11271
rect 10042 11268 10048 11280
rect 9723 11240 10048 11268
rect 9723 11237 9735 11240
rect 9677 11231 9735 11237
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 11422 11228 11428 11280
rect 11480 11268 11486 11280
rect 11882 11268 11888 11280
rect 11480 11240 11888 11268
rect 11480 11228 11486 11240
rect 11882 11228 11888 11240
rect 11940 11228 11946 11280
rect 15562 11277 15568 11280
rect 15105 11271 15163 11277
rect 15105 11237 15117 11271
rect 15151 11268 15163 11271
rect 15556 11268 15568 11277
rect 15151 11240 15568 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 15556 11231 15568 11240
rect 15620 11268 15626 11280
rect 16022 11268 16028 11280
rect 15620 11240 16028 11268
rect 15562 11228 15568 11231
rect 15620 11228 15626 11240
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 18598 11277 18604 11280
rect 18592 11268 18604 11277
rect 18559 11240 18604 11268
rect 18592 11231 18604 11240
rect 18598 11228 18604 11231
rect 18656 11228 18662 11280
rect 25130 11228 25136 11280
rect 25188 11228 25194 11280
rect 25590 11268 25596 11280
rect 25551 11240 25596 11268
rect 25590 11228 25596 11240
rect 25648 11228 25654 11280
rect 8386 11160 8392 11212
rect 8444 11200 8450 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 8444 11172 8493 11200
rect 8444 11160 8450 11172
rect 8481 11169 8493 11172
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 10781 11203 10839 11209
rect 10781 11200 10793 11203
rect 8720 11172 10793 11200
rect 8720 11160 8726 11172
rect 10781 11169 10793 11172
rect 10827 11200 10839 11203
rect 11238 11200 11244 11212
rect 10827 11172 11244 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11790 11200 11796 11212
rect 11379 11172 11796 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 12894 11200 12900 11212
rect 12855 11172 12900 11200
rect 12894 11160 12900 11172
rect 12952 11200 12958 11212
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 12952 11172 13553 11200
rect 12952 11160 12958 11172
rect 13541 11169 13553 11172
rect 13587 11169 13599 11203
rect 13541 11163 13599 11169
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15378 11200 15384 11212
rect 15335 11172 15384 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15378 11160 15384 11172
rect 15436 11160 15442 11212
rect 22353 11203 22411 11209
rect 22353 11200 22365 11203
rect 22020 11172 22365 11200
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 11422 11132 11428 11144
rect 8628 11104 8673 11132
rect 11383 11104 11428 11132
rect 8628 11092 8634 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11132 11667 11135
rect 11698 11132 11704 11144
rect 11655 11104 11704 11132
rect 11655 11101 11667 11104
rect 11609 11095 11667 11101
rect 5721 11067 5779 11073
rect 5721 11033 5733 11067
rect 5767 11064 5779 11067
rect 5994 11064 6000 11076
rect 5767 11036 6000 11064
rect 5767 11033 5779 11036
rect 5721 11027 5779 11033
rect 5994 11024 6000 11036
rect 6052 11064 6058 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 6052 11036 8033 11064
rect 6052 11024 6058 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 8588 11064 8616 11092
rect 11624 11064 11652 11095
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11132 12127 11135
rect 12986 11132 12992 11144
rect 12115 11104 12992 11132
rect 12115 11101 12127 11104
rect 12069 11095 12127 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11132 13231 11135
rect 13722 11132 13728 11144
rect 13219 11104 13728 11132
rect 13219 11101 13231 11104
rect 13173 11095 13231 11101
rect 8168 11036 8616 11064
rect 11072 11036 11652 11064
rect 12437 11067 12495 11073
rect 8168 11024 8174 11036
rect 10870 10956 10876 11008
rect 10928 10996 10934 11008
rect 11072 10996 11100 11036
rect 12437 11033 12449 11067
rect 12483 11064 12495 11067
rect 13188 11064 13216 11095
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 18322 11132 18328 11144
rect 18283 11104 18328 11132
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 21085 11135 21143 11141
rect 21085 11101 21097 11135
rect 21131 11132 21143 11135
rect 21910 11132 21916 11144
rect 21131 11104 21916 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 12483 11036 13216 11064
rect 17405 11067 17463 11073
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 17405 11033 17417 11067
rect 17451 11064 17463 11067
rect 17954 11064 17960 11076
rect 17451 11036 17960 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 19705 11067 19763 11073
rect 19705 11064 19717 11067
rect 19392 11036 19717 11064
rect 19392 11024 19398 11036
rect 19705 11033 19717 11036
rect 19751 11064 19763 11067
rect 20162 11064 20168 11076
rect 19751 11036 20168 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20162 11024 20168 11036
rect 20220 11064 20226 11076
rect 20257 11067 20315 11073
rect 20257 11064 20269 11067
rect 20220 11036 20269 11064
rect 20220 11024 20226 11036
rect 20257 11033 20269 11036
rect 20303 11033 20315 11067
rect 20257 11027 20315 11033
rect 21818 11024 21824 11076
rect 21876 11064 21882 11076
rect 22020 11073 22048 11172
rect 22353 11169 22365 11172
rect 22399 11169 22411 11203
rect 25148 11200 25176 11228
rect 22353 11163 22411 11169
rect 24872 11172 25176 11200
rect 22094 11092 22100 11144
rect 22152 11132 22158 11144
rect 22152 11104 22197 11132
rect 22152 11092 22158 11104
rect 22005 11067 22063 11073
rect 22005 11064 22017 11067
rect 21876 11036 22017 11064
rect 21876 11024 21882 11036
rect 22005 11033 22017 11036
rect 22051 11033 22063 11067
rect 22005 11027 22063 11033
rect 24210 11024 24216 11076
rect 24268 11064 24274 11076
rect 24581 11067 24639 11073
rect 24581 11064 24593 11067
rect 24268 11036 24593 11064
rect 24268 11024 24274 11036
rect 24581 11033 24593 11036
rect 24627 11033 24639 11067
rect 24581 11027 24639 11033
rect 12526 10996 12532 11008
rect 10928 10968 11100 10996
rect 12487 10968 12532 10996
rect 10928 10956 10934 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 24026 10956 24032 11008
rect 24084 10996 24090 11008
rect 24872 10996 24900 11172
rect 25041 11135 25099 11141
rect 25041 11132 25053 11135
rect 24964 11104 25053 11132
rect 24964 11008 24992 11104
rect 25041 11101 25053 11104
rect 25087 11101 25099 11135
rect 25041 11095 25099 11101
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11101 25191 11135
rect 25133 11095 25191 11101
rect 25148 11008 25176 11095
rect 24084 10968 24900 10996
rect 24084 10956 24090 10968
rect 24946 10956 24952 11008
rect 25004 10956 25010 11008
rect 25130 10956 25136 11008
rect 25188 10956 25194 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 7745 10795 7803 10801
rect 7745 10761 7757 10795
rect 7791 10792 7803 10795
rect 8110 10792 8116 10804
rect 7791 10764 8116 10792
rect 7791 10761 7803 10764
rect 7745 10755 7803 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8478 10792 8484 10804
rect 8439 10764 8484 10792
rect 8478 10752 8484 10764
rect 8536 10752 8542 10804
rect 9214 10792 9220 10804
rect 9175 10764 9220 10792
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 9732 10764 10793 10792
rect 9732 10752 9738 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 13814 10792 13820 10804
rect 13775 10764 13820 10792
rect 10781 10755 10839 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15436 10764 15945 10792
rect 15436 10752 15442 10764
rect 15933 10761 15945 10764
rect 15979 10792 15991 10795
rect 16022 10792 16028 10804
rect 15979 10764 16028 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16022 10752 16028 10764
rect 16080 10752 16086 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 16172 10764 16313 10792
rect 16172 10752 16178 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 17037 10795 17095 10801
rect 17037 10792 17049 10795
rect 16632 10764 17049 10792
rect 16632 10752 16638 10764
rect 17037 10761 17049 10764
rect 17083 10761 17095 10795
rect 17037 10755 17095 10761
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18104 10764 18245 10792
rect 18104 10752 18110 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 19518 10792 19524 10804
rect 18233 10755 18291 10761
rect 18708 10764 19524 10792
rect 12158 10724 12164 10736
rect 12119 10696 12164 10724
rect 12158 10684 12164 10696
rect 12216 10684 12222 10736
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 13964 10696 14933 10724
rect 13964 10684 13970 10696
rect 14921 10693 14933 10696
rect 14967 10693 14979 10727
rect 14921 10687 14979 10693
rect 17497 10727 17555 10733
rect 17497 10693 17509 10727
rect 17543 10724 17555 10727
rect 18598 10724 18604 10736
rect 17543 10696 18604 10724
rect 17543 10693 17555 10696
rect 17497 10687 17555 10693
rect 18598 10684 18604 10696
rect 18656 10684 18662 10736
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10656 8171 10659
rect 8202 10656 8208 10668
rect 8159 10628 8208 10656
rect 8159 10625 8171 10628
rect 8113 10619 8171 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9364 10628 9781 10656
rect 9364 10616 9370 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 11238 10656 11244 10668
rect 11199 10628 11244 10656
rect 9769 10619 9827 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11425 10659 11483 10665
rect 11425 10625 11437 10659
rect 11471 10656 11483 10659
rect 11606 10656 11612 10668
rect 11471 10628 11612 10656
rect 11471 10625 11483 10628
rect 11425 10619 11483 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12176 10656 12204 10684
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 12176 10628 12449 10656
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 18708 10665 18736 10764
rect 19518 10752 19524 10764
rect 19576 10792 19582 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19576 10764 19625 10792
rect 19576 10752 19582 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 20070 10792 20076 10804
rect 20031 10764 20076 10792
rect 19613 10755 19671 10761
rect 20070 10752 20076 10764
rect 20128 10752 20134 10804
rect 22002 10792 22008 10804
rect 21100 10764 22008 10792
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15068 10628 15485 10656
rect 15068 10616 15074 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 19334 10656 19340 10668
rect 18831 10628 19340 10656
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9582 10588 9588 10600
rect 9171 10560 9588 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16684 10560 16865 10588
rect 10134 10480 10140 10532
rect 10192 10520 10198 10532
rect 10597 10523 10655 10529
rect 10597 10520 10609 10523
rect 10192 10492 10609 10520
rect 10192 10480 10198 10492
rect 10597 10489 10609 10492
rect 10643 10520 10655 10523
rect 11149 10523 11207 10529
rect 11149 10520 11161 10523
rect 10643 10492 11161 10520
rect 10643 10489 10655 10492
rect 10597 10483 10655 10489
rect 11149 10489 11161 10492
rect 11195 10489 11207 10523
rect 11149 10483 11207 10489
rect 12704 10523 12762 10529
rect 12704 10489 12716 10523
rect 12750 10520 12762 10523
rect 12802 10520 12808 10532
rect 12750 10492 12808 10520
rect 12750 10489 12762 10492
rect 12704 10483 12762 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 15381 10523 15439 10529
rect 15381 10520 15393 10523
rect 14384 10492 15393 10520
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 10321 10455 10379 10461
rect 9732 10424 9777 10452
rect 9732 10412 9738 10424
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 11422 10452 11428 10464
rect 10367 10424 11428 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 11790 10452 11796 10464
rect 11751 10424 11796 10452
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14384 10461 14412 10492
rect 15381 10489 15393 10492
rect 15427 10489 15439 10523
rect 15381 10483 15439 10489
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 13872 10424 14381 10452
rect 13872 10412 13878 10424
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 14369 10415 14427 10421
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 14829 10455 14887 10461
rect 14829 10452 14841 10455
rect 14516 10424 14841 10452
rect 14516 10412 14522 10424
rect 14829 10421 14841 10424
rect 14875 10452 14887 10455
rect 15286 10452 15292 10464
rect 14875 10424 15292 10452
rect 14875 10421 14887 10424
rect 14829 10415 14887 10421
rect 15286 10412 15292 10424
rect 15344 10452 15350 10464
rect 15470 10452 15476 10464
rect 15344 10424 15476 10452
rect 15344 10412 15350 10424
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16684 10461 16712 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 16853 10551 16911 10557
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18598 10588 18604 10600
rect 18012 10560 18604 10588
rect 18012 10548 18018 10560
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 17865 10523 17923 10529
rect 17865 10489 17877 10523
rect 17911 10520 17923 10523
rect 18800 10520 18828 10619
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10588 19947 10591
rect 20622 10588 20628 10600
rect 19935 10560 20628 10588
rect 19935 10557 19947 10560
rect 19889 10551 19947 10557
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 21100 10597 21128 10764
rect 22002 10752 22008 10764
rect 22060 10792 22066 10804
rect 22094 10792 22100 10804
rect 22060 10764 22100 10792
rect 22060 10752 22066 10764
rect 22094 10752 22100 10764
rect 22152 10792 22158 10804
rect 23017 10795 23075 10801
rect 23017 10792 23029 10795
rect 22152 10764 23029 10792
rect 22152 10752 22158 10764
rect 23017 10761 23029 10764
rect 23063 10761 23075 10795
rect 23474 10792 23480 10804
rect 23435 10764 23480 10792
rect 23017 10755 23075 10761
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 23661 10795 23719 10801
rect 23661 10761 23673 10795
rect 23707 10792 23719 10795
rect 24026 10792 24032 10804
rect 23707 10764 24032 10792
rect 23707 10761 23719 10764
rect 23661 10755 23719 10761
rect 24026 10752 24032 10764
rect 24084 10752 24090 10804
rect 25133 10795 25191 10801
rect 25133 10761 25145 10795
rect 25179 10792 25191 10795
rect 25222 10792 25228 10804
rect 25179 10764 25228 10792
rect 25179 10761 25191 10764
rect 25133 10755 25191 10761
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 25409 10795 25467 10801
rect 25409 10761 25421 10795
rect 25455 10792 25467 10795
rect 25774 10792 25780 10804
rect 25455 10764 25780 10792
rect 25455 10761 25467 10764
rect 25409 10755 25467 10761
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 25866 10752 25872 10804
rect 25924 10792 25930 10804
rect 25924 10764 25969 10792
rect 25924 10752 25930 10764
rect 23492 10656 23520 10752
rect 24670 10684 24676 10736
rect 24728 10724 24734 10736
rect 26050 10724 26056 10736
rect 24728 10696 26056 10724
rect 24728 10684 24734 10696
rect 26050 10684 26056 10696
rect 26108 10684 26114 10736
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23492 10628 24225 10656
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10588 21051 10591
rect 21085 10591 21143 10597
rect 21085 10588 21097 10591
rect 21039 10560 21097 10588
rect 21039 10557 21051 10560
rect 20993 10551 21051 10557
rect 21085 10557 21097 10560
rect 21131 10557 21143 10591
rect 21085 10551 21143 10557
rect 23474 10548 23480 10600
rect 23532 10588 23538 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 23532 10560 24685 10588
rect 23532 10548 23538 10560
rect 24673 10557 24685 10560
rect 24719 10588 24731 10591
rect 25038 10588 25044 10600
rect 24719 10560 25044 10588
rect 24719 10557 24731 10560
rect 24673 10551 24731 10557
rect 25038 10548 25044 10560
rect 25096 10548 25102 10600
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10588 25283 10591
rect 25866 10588 25872 10600
rect 25271 10560 25872 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25866 10548 25872 10560
rect 25924 10548 25930 10600
rect 17911 10492 18828 10520
rect 21352 10523 21410 10529
rect 17911 10489 17923 10492
rect 17865 10483 17923 10489
rect 21352 10489 21364 10523
rect 21398 10489 21410 10523
rect 21352 10483 21410 10489
rect 24029 10523 24087 10529
rect 24029 10489 24041 10523
rect 24075 10520 24087 10523
rect 24210 10520 24216 10532
rect 24075 10492 24216 10520
rect 24075 10489 24087 10492
rect 24029 10483 24087 10489
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16632 10424 16681 10452
rect 16632 10412 16638 10424
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 19334 10452 19340 10464
rect 19295 10424 19340 10452
rect 16669 10415 16727 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 20625 10455 20683 10461
rect 20625 10421 20637 10455
rect 20671 10452 20683 10455
rect 21376 10452 21404 10483
rect 24210 10480 24216 10492
rect 24268 10480 24274 10532
rect 21450 10452 21456 10464
rect 20671 10424 21456 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 22336 10424 22477 10452
rect 22336 10412 22342 10424
rect 22465 10421 22477 10424
rect 22511 10421 22523 10455
rect 22465 10415 22523 10421
rect 23842 10412 23848 10464
rect 23900 10452 23906 10464
rect 24121 10455 24179 10461
rect 24121 10452 24133 10455
rect 23900 10424 24133 10452
rect 23900 10412 23906 10424
rect 24121 10421 24133 10424
rect 24167 10421 24179 10455
rect 24121 10415 24179 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 9306 10248 9312 10260
rect 9267 10220 9312 10248
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10100 10220 10609 10248
rect 10100 10208 10106 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 10962 10208 10968 10260
rect 11020 10208 11026 10260
rect 11606 10248 11612 10260
rect 11567 10220 11612 10248
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 15010 10248 15016 10260
rect 14971 10220 15016 10248
rect 15010 10208 15016 10220
rect 15068 10248 15074 10260
rect 15286 10248 15292 10260
rect 15068 10220 15292 10248
rect 15068 10208 15074 10220
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15562 10248 15568 10260
rect 15523 10220 15568 10248
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18656 10220 18797 10248
rect 18656 10208 18662 10220
rect 18785 10217 18797 10220
rect 18831 10217 18843 10251
rect 19150 10248 19156 10260
rect 19111 10220 19156 10248
rect 18785 10211 18843 10217
rect 19150 10208 19156 10220
rect 19208 10248 19214 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19208 10220 19809 10248
rect 19208 10208 19214 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 20898 10248 20904 10260
rect 20859 10220 20904 10248
rect 19797 10211 19855 10217
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 24210 10248 24216 10260
rect 24171 10220 24216 10248
rect 24210 10208 24216 10220
rect 24268 10208 24274 10260
rect 10137 10183 10195 10189
rect 10137 10149 10149 10183
rect 10183 10180 10195 10183
rect 10686 10180 10692 10192
rect 10183 10152 10692 10180
rect 10183 10149 10195 10152
rect 10137 10143 10195 10149
rect 10686 10140 10692 10152
rect 10744 10180 10750 10192
rect 10980 10180 11008 10208
rect 16298 10189 16304 10192
rect 16292 10180 16304 10189
rect 10744 10152 11008 10180
rect 16259 10152 16304 10180
rect 10744 10140 10750 10152
rect 16292 10143 16304 10152
rect 16298 10140 16304 10143
rect 16356 10140 16362 10192
rect 19245 10183 19303 10189
rect 19245 10149 19257 10183
rect 19291 10180 19303 10183
rect 19334 10180 19340 10192
rect 19291 10152 19340 10180
rect 19291 10149 19303 10152
rect 19245 10143 19303 10149
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 21729 10183 21787 10189
rect 21729 10149 21741 10183
rect 21775 10180 21787 10183
rect 22180 10183 22238 10189
rect 22180 10180 22192 10183
rect 21775 10152 22192 10180
rect 21775 10149 21787 10152
rect 21729 10143 21787 10149
rect 22180 10149 22192 10152
rect 22226 10180 22238 10183
rect 22278 10180 22284 10192
rect 22226 10152 22284 10180
rect 22226 10149 22238 10152
rect 22180 10143 22238 10149
rect 22278 10140 22284 10152
rect 22336 10140 22342 10192
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9582 10112 9588 10124
rect 8987 10084 9588 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 10962 10112 10968 10124
rect 10923 10084 10968 10112
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 12158 10112 12164 10124
rect 12119 10084 12164 10112
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12434 10121 12440 10124
rect 12428 10075 12440 10121
rect 12492 10112 12498 10124
rect 16022 10112 16028 10124
rect 12492 10084 12528 10112
rect 15983 10084 16028 10112
rect 12434 10072 12440 10075
rect 12492 10072 12498 10084
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 21913 10115 21971 10121
rect 21913 10081 21925 10115
rect 21959 10112 21971 10115
rect 22002 10112 22008 10124
rect 21959 10084 22008 10112
rect 21959 10081 21971 10084
rect 21913 10075 21971 10081
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 23014 10072 23020 10124
rect 23072 10112 23078 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 23072 10084 24593 10112
rect 23072 10072 23078 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10044 10563 10047
rect 10870 10044 10876 10056
rect 10551 10016 10876 10044
rect 10551 10013 10563 10016
rect 10505 10007 10563 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 11054 10044 11060 10056
rect 11015 10016 11060 10044
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11146 10004 11152 10056
rect 11204 10044 11210 10056
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 11204 10016 11989 10044
rect 11204 10004 11210 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 11992 9908 12020 10007
rect 18690 10004 18696 10056
rect 18748 10044 18754 10056
rect 19337 10047 19395 10053
rect 19337 10044 19349 10047
rect 18748 10016 19349 10044
rect 18748 10004 18754 10016
rect 19337 10013 19349 10016
rect 19383 10044 19395 10047
rect 19426 10044 19432 10056
rect 19383 10016 19432 10044
rect 19383 10013 19395 10016
rect 19337 10007 19395 10013
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 18049 9979 18107 9985
rect 18049 9945 18061 9979
rect 18095 9976 18107 9979
rect 18506 9976 18512 9988
rect 18095 9948 18512 9976
rect 18095 9945 18107 9948
rect 18049 9939 18107 9945
rect 18506 9936 18512 9948
rect 18564 9936 18570 9988
rect 23934 9936 23940 9988
rect 23992 9976 23998 9988
rect 24765 9979 24823 9985
rect 24765 9976 24777 9979
rect 23992 9948 24777 9976
rect 23992 9936 23998 9948
rect 24765 9945 24777 9948
rect 24811 9945 24823 9979
rect 24765 9939 24823 9945
rect 12802 9908 12808 9920
rect 11992 9880 12808 9908
rect 12802 9868 12808 9880
rect 12860 9908 12866 9920
rect 13538 9908 13544 9920
rect 12860 9880 13544 9908
rect 12860 9868 12866 9880
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 17405 9911 17463 9917
rect 17405 9877 17417 9911
rect 17451 9908 17463 9911
rect 17586 9908 17592 9920
rect 17451 9880 17592 9908
rect 17451 9877 17463 9880
rect 17405 9871 17463 9877
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 18322 9908 18328 9920
rect 18283 9880 18328 9908
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 20257 9911 20315 9917
rect 20257 9877 20269 9911
rect 20303 9908 20315 9911
rect 20622 9908 20628 9920
rect 20303 9880 20628 9908
rect 20303 9877 20315 9880
rect 20257 9871 20315 9877
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 21818 9868 21824 9920
rect 21876 9908 21882 9920
rect 23293 9911 23351 9917
rect 23293 9908 23305 9911
rect 21876 9880 23305 9908
rect 21876 9868 21882 9880
rect 23293 9877 23305 9880
rect 23339 9877 23351 9911
rect 23842 9908 23848 9920
rect 23803 9880 23848 9908
rect 23293 9871 23351 9877
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 25130 9908 25136 9920
rect 25091 9880 25136 9908
rect 25130 9868 25136 9880
rect 25188 9868 25194 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 11146 9704 11152 9716
rect 11107 9676 11152 9704
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 12158 9704 12164 9716
rect 12119 9676 12164 9704
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 12434 9704 12440 9716
rect 12400 9676 12440 9704
rect 12400 9664 12406 9676
rect 12434 9664 12440 9676
rect 12492 9704 12498 9716
rect 12618 9704 12624 9716
rect 12492 9676 12624 9704
rect 12492 9664 12498 9676
rect 12618 9664 12624 9676
rect 12676 9704 12682 9716
rect 14642 9704 14648 9716
rect 12676 9676 14648 9704
rect 12676 9664 12682 9676
rect 14642 9664 14648 9676
rect 14700 9704 14706 9716
rect 15105 9707 15163 9713
rect 15105 9704 15117 9707
rect 14700 9676 15117 9704
rect 14700 9664 14706 9676
rect 15105 9673 15117 9676
rect 15151 9704 15163 9707
rect 15286 9704 15292 9716
rect 15151 9676 15292 9704
rect 15151 9673 15163 9676
rect 15105 9667 15163 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 16356 9676 16528 9704
rect 16356 9664 16362 9676
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 10045 9639 10103 9645
rect 10045 9636 10057 9639
rect 9732 9608 10057 9636
rect 9732 9596 9738 9608
rect 10045 9605 10057 9608
rect 10091 9605 10103 9639
rect 10045 9599 10103 9605
rect 10686 9568 10692 9580
rect 10647 9540 10692 9568
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 12176 9568 12204 9664
rect 16206 9636 16212 9648
rect 16167 9608 16212 9636
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 16500 9636 16528 9676
rect 22002 9664 22008 9716
rect 22060 9704 22066 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 22060 9676 22661 9704
rect 22060 9664 22066 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 22649 9667 22707 9673
rect 23014 9664 23020 9716
rect 23072 9704 23078 9716
rect 23290 9704 23296 9716
rect 23072 9676 23296 9704
rect 23072 9664 23078 9676
rect 23290 9664 23296 9676
rect 23348 9704 23354 9716
rect 24397 9707 24455 9713
rect 24397 9704 24409 9707
rect 23348 9676 24409 9704
rect 23348 9664 23354 9676
rect 24397 9673 24409 9676
rect 24443 9673 24455 9707
rect 24397 9667 24455 9673
rect 17221 9639 17279 9645
rect 17221 9636 17233 9639
rect 16500 9608 17233 9636
rect 17221 9605 17233 9608
rect 17267 9605 17279 9639
rect 17221 9599 17279 9605
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 20257 9639 20315 9645
rect 20257 9636 20269 9639
rect 19484 9608 20269 9636
rect 19484 9596 19490 9608
rect 20257 9605 20269 9608
rect 20303 9605 20315 9639
rect 20257 9599 20315 9605
rect 24670 9596 24676 9648
rect 24728 9636 24734 9648
rect 24765 9639 24823 9645
rect 24765 9636 24777 9639
rect 24728 9608 24777 9636
rect 24728 9596 24734 9608
rect 24765 9605 24777 9608
rect 24811 9605 24823 9639
rect 24765 9599 24823 9605
rect 12434 9568 12440 9580
rect 12176 9540 12440 9568
rect 12434 9528 12440 9540
rect 12492 9568 12498 9580
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 12492 9540 13553 9568
rect 12492 9528 12498 9540
rect 13541 9537 13553 9540
rect 13587 9568 13599 9571
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13587 9540 13737 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13725 9537 13737 9540
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16816 9540 16865 9568
rect 16816 9528 16822 9540
rect 16853 9537 16865 9540
rect 16899 9568 16911 9571
rect 16942 9568 16948 9580
rect 16899 9540 16948 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 22278 9568 22284 9580
rect 22239 9540 22284 9568
rect 22278 9528 22284 9540
rect 22336 9528 22342 9580
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 10100 9472 10517 9500
rect 10100 9460 10106 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 12342 9500 12348 9512
rect 11931 9472 12348 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 18322 9500 18328 9512
rect 17788 9472 18328 9500
rect 13265 9435 13323 9441
rect 13265 9401 13277 9435
rect 13311 9432 13323 9435
rect 13992 9435 14050 9441
rect 13992 9432 14004 9435
rect 13311 9404 14004 9432
rect 13311 9401 13323 9404
rect 13265 9395 13323 9401
rect 13992 9401 14004 9404
rect 14038 9432 14050 9435
rect 14274 9432 14280 9444
rect 14038 9404 14280 9432
rect 14038 9401 14050 9404
rect 13992 9395 14050 9401
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 16117 9435 16175 9441
rect 16117 9401 16129 9435
rect 16163 9432 16175 9435
rect 16666 9432 16672 9444
rect 16163 9404 16672 9432
rect 16163 9401 16175 9404
rect 16117 9395 16175 9401
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 17788 9376 17816 9472
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 20898 9460 20904 9512
rect 20956 9500 20962 9512
rect 21177 9503 21235 9509
rect 21177 9500 21189 9503
rect 20956 9472 21189 9500
rect 20956 9460 20962 9472
rect 21177 9469 21189 9472
rect 21223 9500 21235 9503
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21223 9472 22109 9500
rect 21223 9469 21235 9472
rect 21177 9463 21235 9469
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 24578 9500 24584 9512
rect 24539 9472 24584 9500
rect 22097 9463 22155 9469
rect 24578 9460 24584 9472
rect 24636 9500 24642 9512
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 24636 9472 25145 9500
rect 24636 9460 24642 9472
rect 25133 9469 25145 9472
rect 25179 9469 25191 9503
rect 25133 9463 25191 9469
rect 18506 9392 18512 9444
rect 18564 9441 18570 9444
rect 18564 9435 18628 9441
rect 18564 9401 18582 9435
rect 18616 9401 18628 9435
rect 18564 9395 18628 9401
rect 21545 9435 21603 9441
rect 21545 9401 21557 9435
rect 21591 9432 21603 9435
rect 22002 9432 22008 9444
rect 21591 9404 22008 9432
rect 21591 9401 21603 9404
rect 21545 9395 21603 9401
rect 18564 9392 18570 9395
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 9858 9364 9864 9376
rect 9819 9336 9864 9364
rect 9858 9324 9864 9336
rect 9916 9364 9922 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9916 9336 10425 9364
rect 9916 9324 9922 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11204 9336 11529 9364
rect 11204 9324 11210 9336
rect 11517 9333 11529 9336
rect 11563 9364 11575 9367
rect 11882 9364 11888 9376
rect 11563 9336 11888 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 12308 9336 12541 9364
rect 12308 9324 12314 9336
rect 12529 9333 12541 9336
rect 12575 9333 12587 9367
rect 15746 9364 15752 9376
rect 15659 9336 15752 9364
rect 12529 9327 12587 9333
rect 15746 9324 15752 9336
rect 15804 9364 15810 9376
rect 16577 9367 16635 9373
rect 16577 9364 16589 9367
rect 15804 9336 16589 9364
rect 15804 9324 15810 9336
rect 16577 9333 16589 9336
rect 16623 9364 16635 9367
rect 16850 9364 16856 9376
rect 16623 9336 16856 9364
rect 16623 9333 16635 9336
rect 16577 9327 16635 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 19705 9367 19763 9373
rect 19705 9364 19717 9367
rect 18932 9336 19717 9364
rect 18932 9324 18938 9336
rect 19705 9333 19717 9336
rect 19751 9364 19763 9367
rect 20438 9364 20444 9376
rect 19751 9336 20444 9364
rect 19751 9333 19763 9336
rect 19705 9327 19763 9333
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 21637 9367 21695 9373
rect 21637 9333 21649 9367
rect 21683 9364 21695 9367
rect 21726 9364 21732 9376
rect 21683 9336 21732 9364
rect 21683 9333 21695 9336
rect 21637 9327 21695 9333
rect 21726 9324 21732 9336
rect 21784 9324 21790 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 10042 9160 10048 9172
rect 10003 9132 10048 9160
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10689 9163 10747 9169
rect 10689 9129 10701 9163
rect 10735 9160 10747 9163
rect 10962 9160 10968 9172
rect 10735 9132 10968 9160
rect 10735 9129 10747 9132
rect 10689 9123 10747 9129
rect 10962 9120 10968 9132
rect 11020 9160 11026 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11020 9132 11897 9160
rect 11020 9120 11026 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 13449 9163 13507 9169
rect 13449 9129 13461 9163
rect 13495 9160 13507 9163
rect 13722 9160 13728 9172
rect 13495 9132 13728 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 13909 9163 13967 9169
rect 13909 9129 13921 9163
rect 13955 9160 13967 9163
rect 13998 9160 14004 9172
rect 13955 9132 14004 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14553 9163 14611 9169
rect 14553 9129 14565 9163
rect 14599 9160 14611 9163
rect 14642 9160 14648 9172
rect 14599 9132 14648 9160
rect 14599 9129 14611 9132
rect 14553 9123 14611 9129
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 16482 9160 16488 9172
rect 15611 9132 16488 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16942 9160 16948 9172
rect 16903 9132 16948 9160
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 19426 9160 19432 9172
rect 19387 9132 19432 9160
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 19981 9163 20039 9169
rect 19981 9160 19993 9163
rect 19576 9132 19993 9160
rect 19576 9120 19582 9132
rect 19981 9129 19993 9132
rect 20027 9129 20039 9163
rect 20898 9160 20904 9172
rect 20859 9132 20904 9160
rect 19981 9123 20039 9129
rect 20898 9120 20904 9132
rect 20956 9120 20962 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 22830 9160 22836 9172
rect 22152 9132 22836 9160
rect 22152 9120 22158 9132
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 24762 9160 24768 9172
rect 24723 9132 24768 9160
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 13262 9052 13268 9104
rect 13320 9092 13326 9104
rect 13817 9095 13875 9101
rect 13817 9092 13829 9095
rect 13320 9064 13829 9092
rect 13320 9052 13326 9064
rect 13817 9061 13829 9064
rect 13863 9092 13875 9095
rect 14366 9092 14372 9104
rect 13863 9064 14372 9092
rect 13863 9061 13875 9064
rect 13817 9055 13875 9061
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 16022 9052 16028 9104
rect 16080 9092 16086 9104
rect 16390 9092 16396 9104
rect 16080 9064 16396 9092
rect 16080 9052 16086 9064
rect 16390 9052 16396 9064
rect 16448 9092 16454 9104
rect 16577 9095 16635 9101
rect 16577 9092 16589 9095
rect 16448 9064 16589 9092
rect 16448 9052 16454 9064
rect 16577 9061 16589 9064
rect 16623 9092 16635 9095
rect 17770 9092 17776 9104
rect 16623 9064 17776 9092
rect 16623 9061 16635 9064
rect 16577 9055 16635 9061
rect 12250 9024 12256 9036
rect 12211 8996 12256 9024
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 9024 13047 9027
rect 13354 9024 13360 9036
rect 13035 8996 13360 9024
rect 13035 8993 13047 8996
rect 12989 8987 13047 8993
rect 13354 8984 13360 8996
rect 13412 9024 13418 9036
rect 13722 9024 13728 9036
rect 13412 8996 13728 9024
rect 13412 8984 13418 8996
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 15746 8984 15752 9036
rect 15804 9024 15810 9036
rect 17144 9033 17172 9064
rect 17770 9052 17776 9064
rect 17828 9052 17834 9104
rect 22005 9095 22063 9101
rect 22005 9061 22017 9095
rect 22051 9092 22063 9095
rect 22278 9092 22284 9104
rect 22051 9064 22284 9092
rect 22051 9061 22063 9064
rect 22005 9055 22063 9061
rect 22278 9052 22284 9064
rect 22336 9092 22342 9104
rect 22336 9064 23152 9092
rect 22336 9052 22342 9064
rect 17402 9033 17408 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15804 8996 15945 9024
rect 15804 8984 15810 8996
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 8993 17187 9027
rect 17396 9024 17408 9033
rect 17363 8996 17408 9024
rect 17129 8987 17187 8993
rect 17396 8987 17408 8996
rect 17402 8984 17408 8987
rect 17460 8984 17466 9036
rect 19797 9027 19855 9033
rect 19797 8993 19809 9027
rect 19843 9024 19855 9027
rect 20346 9024 20352 9036
rect 19843 8996 20352 9024
rect 19843 8993 19855 8996
rect 19797 8987 19855 8993
rect 20346 8984 20352 8996
rect 20404 8984 20410 9036
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20956 8996 21281 9024
rect 20956 8984 20962 8996
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 22462 8984 22468 9036
rect 22520 9024 22526 9036
rect 22738 9024 22744 9036
rect 22520 8996 22744 9024
rect 22520 8984 22526 8996
rect 22738 8984 22744 8996
rect 22796 9024 22802 9036
rect 22925 9027 22983 9033
rect 22925 9024 22937 9027
rect 22796 8996 22937 9024
rect 22796 8984 22802 8996
rect 22925 8993 22937 8996
rect 22971 8993 22983 9027
rect 22925 8987 22983 8993
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 12342 8956 12348 8968
rect 11756 8928 12348 8956
rect 11756 8916 11762 8928
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12529 8959 12587 8965
rect 12529 8925 12541 8959
rect 12575 8956 12587 8959
rect 12618 8956 12624 8968
rect 12575 8928 12624 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 14274 8956 14280 8968
rect 14139 8928 14280 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8956 15163 8959
rect 16022 8956 16028 8968
rect 15151 8928 16028 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16114 8916 16120 8968
rect 16172 8956 16178 8968
rect 16172 8928 16217 8956
rect 16172 8916 16178 8928
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21361 8959 21419 8965
rect 21361 8956 21373 8959
rect 20680 8928 21373 8956
rect 20680 8916 20686 8928
rect 21361 8925 21373 8928
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 23124 8965 23152 9064
rect 24581 9027 24639 9033
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 24670 9024 24676 9036
rect 24627 8996 24676 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 24670 8984 24676 8996
rect 24728 8984 24734 9036
rect 23109 8959 23167 8965
rect 21508 8928 21553 8956
rect 21508 8916 21514 8928
rect 23109 8925 23121 8959
rect 23155 8956 23167 8959
rect 23198 8956 23204 8968
rect 23155 8928 23204 8956
rect 23155 8925 23167 8928
rect 23109 8919 23167 8925
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 18506 8888 18512 8900
rect 18467 8860 18512 8888
rect 18506 8848 18512 8860
rect 18564 8848 18570 8900
rect 22465 8891 22523 8897
rect 22465 8888 22477 8891
rect 20732 8860 22477 8888
rect 20732 8832 20760 8860
rect 22465 8857 22477 8860
rect 22511 8857 22523 8891
rect 22465 8851 22523 8857
rect 20714 8820 20720 8832
rect 20675 8792 20720 8820
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 11609 8619 11667 8625
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 12250 8616 12256 8628
rect 11655 8588 12256 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 12897 8619 12955 8625
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 12986 8616 12992 8628
rect 12943 8588 12992 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13262 8616 13268 8628
rect 13188 8588 13268 8616
rect 12805 8551 12863 8557
rect 12805 8517 12817 8551
rect 12851 8548 12863 8551
rect 13188 8548 13216 8588
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13998 8616 14004 8628
rect 13959 8588 14004 8616
rect 13998 8576 14004 8588
rect 14056 8616 14062 8628
rect 15378 8616 15384 8628
rect 14056 8588 15384 8616
rect 14056 8576 14062 8588
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15657 8619 15715 8625
rect 15657 8585 15669 8619
rect 15703 8616 15715 8619
rect 16114 8616 16120 8628
rect 15703 8588 16120 8616
rect 15703 8585 15715 8588
rect 15657 8579 15715 8585
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 17497 8619 17555 8625
rect 17497 8585 17509 8619
rect 17543 8616 17555 8619
rect 17770 8616 17776 8628
rect 17543 8588 17776 8616
rect 17543 8585 17555 8588
rect 17497 8579 17555 8585
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18874 8616 18880 8628
rect 18835 8588 18880 8616
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 20806 8576 20812 8628
rect 20864 8616 20870 8628
rect 21269 8619 21327 8625
rect 21269 8616 21281 8619
rect 20864 8588 21281 8616
rect 20864 8576 20870 8588
rect 21269 8585 21281 8588
rect 21315 8585 21327 8619
rect 22830 8616 22836 8628
rect 22791 8588 22836 8616
rect 21269 8579 21327 8585
rect 22830 8576 22836 8588
rect 22888 8576 22894 8628
rect 23198 8616 23204 8628
rect 23159 8588 23204 8616
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 25225 8619 25283 8625
rect 25225 8585 25237 8619
rect 25271 8616 25283 8619
rect 25406 8616 25412 8628
rect 25271 8588 25412 8616
rect 25271 8585 25283 8588
rect 25225 8579 25283 8585
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 12851 8520 13216 8548
rect 13280 8520 14473 8548
rect 12851 8517 12863 8520
rect 12805 8511 12863 8517
rect 13280 8424 13308 8520
rect 14461 8517 14473 8520
rect 14507 8517 14519 8551
rect 18892 8548 18920 8576
rect 20898 8548 20904 8560
rect 18892 8520 19932 8548
rect 20859 8520 20904 8548
rect 14461 8511 14519 8517
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13538 8480 13544 8492
rect 13412 8452 13457 8480
rect 13499 8452 13544 8480
rect 13412 8440 13418 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14700 8452 15025 8480
rect 14700 8440 14706 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16942 8480 16948 8492
rect 16347 8452 16948 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16942 8440 16948 8452
rect 17000 8480 17006 8492
rect 17402 8480 17408 8492
rect 17000 8452 17408 8480
rect 17000 8440 17006 8452
rect 17402 8440 17408 8452
rect 17460 8480 17466 8492
rect 17865 8483 17923 8489
rect 17865 8480 17877 8483
rect 17460 8452 17877 8480
rect 17460 8440 17466 8452
rect 17865 8449 17877 8452
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19904 8489 19932 8520
rect 20898 8508 20904 8520
rect 20956 8508 20962 8560
rect 19797 8483 19855 8489
rect 19797 8480 19809 8483
rect 19484 8452 19809 8480
rect 19484 8440 19490 8452
rect 19797 8449 19809 8452
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8449 19947 8483
rect 21726 8480 21732 8492
rect 21687 8452 21732 8480
rect 19889 8443 19947 8449
rect 21726 8440 21732 8452
rect 21784 8440 21790 8492
rect 21818 8440 21824 8492
rect 21876 8480 21882 8492
rect 24029 8483 24087 8489
rect 21876 8452 21921 8480
rect 21876 8440 21882 8452
rect 24029 8449 24041 8483
rect 24075 8480 24087 8483
rect 24118 8480 24124 8492
rect 24075 8452 24124 8480
rect 24075 8449 24087 8452
rect 24029 8443 24087 8449
rect 24118 8440 24124 8452
rect 24176 8440 24182 8492
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8412 11299 8415
rect 12618 8412 12624 8424
rect 11287 8384 12624 8412
rect 11287 8381 11299 8384
rect 11241 8375 11299 8381
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 13262 8412 13268 8424
rect 13175 8384 13268 8412
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 16632 8384 16865 8412
rect 16632 8372 16638 8384
rect 16853 8381 16865 8384
rect 16899 8412 16911 8415
rect 17770 8412 17776 8424
rect 16899 8384 17776 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 19245 8415 19303 8421
rect 19245 8381 19257 8415
rect 19291 8412 19303 8415
rect 19702 8412 19708 8424
rect 19291 8384 19708 8412
rect 19291 8381 19303 8384
rect 19245 8375 19303 8381
rect 19702 8372 19708 8384
rect 19760 8372 19766 8424
rect 20530 8412 20536 8424
rect 20491 8384 20536 8412
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 20772 8384 21649 8412
rect 20772 8372 20778 8384
rect 21637 8381 21649 8384
rect 21683 8381 21695 8415
rect 21744 8412 21772 8440
rect 22094 8412 22100 8424
rect 21744 8384 22100 8412
rect 21637 8375 21695 8381
rect 22094 8372 22100 8384
rect 22152 8372 22158 8424
rect 25038 8412 25044 8424
rect 24999 8384 25044 8412
rect 25038 8372 25044 8384
rect 25096 8412 25102 8424
rect 25501 8415 25559 8421
rect 25501 8412 25513 8415
rect 25096 8384 25513 8412
rect 25096 8372 25102 8384
rect 25501 8381 25513 8384
rect 25547 8381 25559 8415
rect 25501 8375 25559 8381
rect 11698 8304 11704 8356
rect 11756 8344 11762 8356
rect 11885 8347 11943 8353
rect 11885 8344 11897 8347
rect 11756 8316 11897 8344
rect 11756 8304 11762 8316
rect 11885 8313 11897 8316
rect 11931 8313 11943 8347
rect 11885 8307 11943 8313
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8344 14427 8347
rect 14642 8344 14648 8356
rect 14415 8316 14648 8344
rect 14415 8313 14427 8316
rect 14369 8307 14427 8313
rect 14642 8304 14648 8316
rect 14700 8344 14706 8356
rect 14829 8347 14887 8353
rect 14829 8344 14841 8347
rect 14700 8316 14841 8344
rect 14700 8304 14706 8316
rect 14829 8313 14841 8316
rect 14875 8313 14887 8347
rect 16758 8344 16764 8356
rect 16719 8316 16764 8344
rect 14829 8307 14887 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 18049 8347 18107 8353
rect 18049 8344 18061 8347
rect 17880 8316 18061 8344
rect 17880 8288 17908 8316
rect 18049 8313 18061 8316
rect 18095 8313 18107 8347
rect 18049 8307 18107 8313
rect 14458 8236 14464 8288
rect 14516 8276 14522 8288
rect 14921 8279 14979 8285
rect 14921 8276 14933 8279
rect 14516 8248 14933 8276
rect 14516 8236 14522 8248
rect 14921 8245 14933 8248
rect 14967 8245 14979 8279
rect 14921 8239 14979 8245
rect 15746 8236 15752 8288
rect 15804 8276 15810 8288
rect 16393 8279 16451 8285
rect 16393 8276 16405 8279
rect 15804 8248 16405 8276
rect 15804 8236 15810 8248
rect 16393 8245 16405 8248
rect 16439 8245 16451 8279
rect 16393 8239 16451 8245
rect 17862 8236 17868 8288
rect 17920 8236 17926 8288
rect 22462 8276 22468 8288
rect 22423 8248 22468 8276
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 23842 8236 23848 8288
rect 23900 8276 23906 8288
rect 24581 8279 24639 8285
rect 24581 8276 24593 8279
rect 23900 8248 24593 8276
rect 23900 8236 23906 8248
rect 24581 8245 24593 8248
rect 24627 8276 24639 8279
rect 24670 8276 24676 8288
rect 24627 8248 24676 8276
rect 24627 8245 24639 8248
rect 24581 8239 24639 8245
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 11882 8072 11888 8084
rect 11843 8044 11888 8072
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 13262 8072 13268 8084
rect 13223 8044 13268 8072
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 14550 8072 14556 8084
rect 13679 8044 14556 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15654 8072 15660 8084
rect 15615 8044 15660 8072
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 16025 8075 16083 8081
rect 16025 8041 16037 8075
rect 16071 8072 16083 8075
rect 16482 8072 16488 8084
rect 16071 8044 16488 8072
rect 16071 8041 16083 8044
rect 16025 8035 16083 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 17000 8044 17877 8072
rect 17000 8032 17006 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 20073 8075 20131 8081
rect 20073 8041 20085 8075
rect 20119 8072 20131 8075
rect 20346 8072 20352 8084
rect 20119 8044 20352 8072
rect 20119 8041 20131 8044
rect 20073 8035 20131 8041
rect 20346 8032 20352 8044
rect 20404 8032 20410 8084
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 22833 8075 22891 8081
rect 22152 8044 22197 8072
rect 22152 8032 22158 8044
rect 22833 8041 22845 8075
rect 22879 8072 22891 8075
rect 23106 8072 23112 8084
rect 22879 8044 23112 8072
rect 22879 8041 22891 8044
rect 22833 8035 22891 8041
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 23845 8075 23903 8081
rect 23845 8041 23857 8075
rect 23891 8072 23903 8075
rect 23934 8072 23940 8084
rect 23891 8044 23940 8072
rect 23891 8041 23903 8044
rect 23845 8035 23903 8041
rect 23934 8032 23940 8044
rect 23992 8032 23998 8084
rect 24857 8075 24915 8081
rect 24857 8041 24869 8075
rect 24903 8072 24915 8075
rect 25958 8072 25964 8084
rect 24903 8044 25964 8072
rect 24903 8041 24915 8044
rect 24857 8035 24915 8041
rect 25958 8032 25964 8044
rect 26016 8032 26022 8084
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 12345 8007 12403 8013
rect 12345 8004 12357 8007
rect 10008 7976 12357 8004
rect 10008 7964 10014 7976
rect 12345 7973 12357 7976
rect 12391 8004 12403 8007
rect 12802 8004 12808 8016
rect 12391 7976 12808 8004
rect 12391 7973 12403 7976
rect 12345 7967 12403 7973
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 12989 8007 13047 8013
rect 12989 7973 13001 8007
rect 13035 8004 13047 8007
rect 13538 8004 13544 8016
rect 13035 7976 13544 8004
rect 13035 7973 13047 7976
rect 12989 7967 13047 7973
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 20717 8007 20775 8013
rect 20717 7973 20729 8007
rect 20763 8004 20775 8007
rect 21450 8004 21456 8016
rect 20763 7976 21456 8004
rect 20763 7973 20775 7976
rect 20717 7967 20775 7973
rect 21450 7964 21456 7976
rect 21508 7964 21514 8016
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12253 7939 12311 7945
rect 12253 7936 12265 7939
rect 11940 7908 12265 7936
rect 11940 7896 11946 7908
rect 12253 7905 12265 7908
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 13446 7936 13452 7948
rect 12584 7908 13452 7936
rect 12584 7896 12590 7908
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 14826 7896 14832 7948
rect 14884 7936 14890 7948
rect 15470 7936 15476 7948
rect 14884 7908 15476 7936
rect 14884 7896 14890 7908
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 16485 7939 16543 7945
rect 16485 7936 16497 7939
rect 16448 7908 16497 7936
rect 16448 7896 16454 7908
rect 16485 7905 16497 7908
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 16752 7939 16810 7945
rect 16752 7905 16764 7939
rect 16798 7936 16810 7939
rect 17586 7936 17592 7948
rect 16798 7908 17592 7936
rect 16798 7905 16810 7908
rect 16752 7899 16810 7905
rect 17586 7896 17592 7908
rect 17644 7896 17650 7948
rect 19334 7936 19340 7948
rect 19295 7908 19340 7936
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 21361 7939 21419 7945
rect 21361 7905 21373 7939
rect 21407 7936 21419 7939
rect 21818 7936 21824 7948
rect 21407 7908 21824 7936
rect 21407 7905 21419 7908
rect 21361 7899 21419 7905
rect 21818 7896 21824 7908
rect 21876 7896 21882 7948
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22646 7936 22652 7948
rect 22152 7908 22652 7936
rect 22152 7896 22158 7908
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 23661 7939 23719 7945
rect 23661 7905 23673 7939
rect 23707 7936 23719 7939
rect 23750 7936 23756 7948
rect 23707 7908 23756 7936
rect 23707 7905 23719 7908
rect 23661 7899 23719 7905
rect 23750 7896 23756 7908
rect 23808 7936 23814 7948
rect 24118 7936 24124 7948
rect 23808 7908 24124 7936
rect 23808 7896 23814 7908
rect 24118 7896 24124 7908
rect 24176 7896 24182 7948
rect 24670 7936 24676 7948
rect 24631 7908 24676 7936
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 12618 7868 12624 7880
rect 12483 7840 12624 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 19208 7840 19441 7868
rect 19208 7828 19214 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19610 7868 19616 7880
rect 19523 7840 19616 7868
rect 19429 7831 19487 7837
rect 19610 7828 19616 7840
rect 19668 7868 19674 7880
rect 20622 7868 20628 7880
rect 19668 7840 20628 7868
rect 19668 7828 19674 7840
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 23658 7760 23664 7812
rect 23716 7800 23722 7812
rect 23934 7800 23940 7812
rect 23716 7772 23940 7800
rect 23716 7760 23722 7772
rect 23934 7760 23940 7772
rect 23992 7760 23998 7812
rect 14001 7735 14059 7741
rect 14001 7701 14013 7735
rect 14047 7732 14059 7735
rect 14274 7732 14280 7744
rect 14047 7704 14280 7732
rect 14047 7701 14059 7704
rect 14001 7695 14059 7701
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 14550 7732 14556 7744
rect 14511 7704 14556 7732
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 16390 7732 16396 7744
rect 16351 7704 16396 7732
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 18966 7732 18972 7744
rect 18927 7704 18972 7732
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 11609 7531 11667 7537
rect 11609 7497 11621 7531
rect 11655 7528 11667 7531
rect 12618 7528 12624 7540
rect 11655 7500 12624 7528
rect 11655 7497 11667 7500
rect 11609 7491 11667 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 15013 7531 15071 7537
rect 15013 7497 15025 7531
rect 15059 7528 15071 7531
rect 15746 7528 15752 7540
rect 15059 7500 15752 7528
rect 15059 7497 15071 7500
rect 15013 7491 15071 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16393 7531 16451 7537
rect 16393 7528 16405 7531
rect 16080 7500 16405 7528
rect 16080 7488 16086 7500
rect 16393 7497 16405 7500
rect 16439 7497 16451 7531
rect 16393 7491 16451 7497
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 17828 7500 18061 7528
rect 17828 7488 17834 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 19150 7528 19156 7540
rect 19111 7500 19156 7528
rect 18049 7491 18107 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7528 19671 7531
rect 19978 7528 19984 7540
rect 19659 7500 19984 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 20622 7528 20628 7540
rect 20583 7500 20628 7528
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 22646 7488 22652 7540
rect 22704 7528 22710 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22704 7500 23029 7528
rect 22704 7488 22710 7500
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23842 7528 23848 7540
rect 23803 7500 23848 7528
rect 23017 7491 23075 7497
rect 23842 7488 23848 7500
rect 23900 7488 23906 7540
rect 24118 7528 24124 7540
rect 24079 7500 24124 7528
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 25501 7531 25559 7537
rect 25501 7528 25513 7531
rect 24728 7500 25513 7528
rect 24728 7488 24734 7500
rect 25501 7497 25513 7500
rect 25547 7497 25559 7531
rect 25501 7491 25559 7497
rect 15933 7463 15991 7469
rect 15933 7429 15945 7463
rect 15979 7460 15991 7463
rect 24857 7463 24915 7469
rect 15979 7432 17540 7460
rect 15979 7429 15991 7432
rect 15933 7423 15991 7429
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 14792 7364 15117 7392
rect 14792 7352 14798 7364
rect 15105 7361 15117 7364
rect 15151 7361 15163 7395
rect 16298 7392 16304 7404
rect 16259 7364 16304 7392
rect 15105 7355 15163 7361
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16448 7364 16865 7392
rect 16448 7352 16454 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17512 7401 17540 7432
rect 24857 7429 24869 7463
rect 24903 7460 24915 7463
rect 25314 7460 25320 7472
rect 24903 7432 25320 7460
rect 24903 7429 24915 7432
rect 24857 7423 24915 7429
rect 25314 7420 25320 7432
rect 25372 7420 25378 7472
rect 17497 7395 17555 7401
rect 17000 7364 17045 7392
rect 17000 7352 17006 7364
rect 17497 7361 17509 7395
rect 17543 7392 17555 7395
rect 17586 7392 17592 7404
rect 17543 7364 17592 7392
rect 17543 7361 17555 7364
rect 17497 7355 17555 7361
rect 17586 7352 17592 7364
rect 17644 7392 17650 7404
rect 18693 7395 18751 7401
rect 18693 7392 18705 7395
rect 17644 7364 18705 7392
rect 17644 7352 17650 7364
rect 18693 7361 18705 7364
rect 18739 7392 18751 7395
rect 19610 7392 19616 7404
rect 18739 7364 19616 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19610 7352 19616 7364
rect 19668 7352 19674 7404
rect 20254 7392 20260 7404
rect 20215 7364 20260 7392
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 20990 7352 20996 7404
rect 21048 7392 21054 7404
rect 21177 7395 21235 7401
rect 21177 7392 21189 7395
rect 21048 7364 21189 7392
rect 21048 7352 21054 7364
rect 21177 7361 21189 7364
rect 21223 7361 21235 7395
rect 22554 7392 22560 7404
rect 22515 7364 22560 7392
rect 21177 7355 21235 7361
rect 22554 7352 22560 7364
rect 22612 7352 22618 7404
rect 23934 7352 23940 7404
rect 23992 7392 23998 7404
rect 24118 7392 24124 7404
rect 23992 7364 24124 7392
rect 23992 7352 23998 7364
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 12802 7324 12808 7336
rect 12759 7296 12808 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 16482 7284 16488 7336
rect 16540 7324 16546 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 16540 7296 16773 7324
rect 16540 7284 16546 7296
rect 16761 7293 16773 7296
rect 16807 7324 16819 7327
rect 18966 7324 18972 7336
rect 16807 7296 18972 7324
rect 16807 7293 16819 7296
rect 16761 7287 16819 7293
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 20073 7327 20131 7333
rect 20073 7324 20085 7327
rect 19484 7296 20085 7324
rect 19484 7284 19490 7296
rect 20073 7293 20085 7296
rect 20119 7293 20131 7327
rect 23658 7324 23664 7336
rect 23619 7296 23664 7324
rect 20073 7287 20131 7293
rect 23658 7284 23664 7296
rect 23716 7324 23722 7336
rect 24489 7327 24547 7333
rect 24489 7324 24501 7327
rect 23716 7296 24501 7324
rect 23716 7284 23722 7296
rect 24489 7293 24501 7296
rect 24535 7293 24547 7327
rect 24670 7324 24676 7336
rect 24631 7296 24676 7324
rect 24489 7287 24547 7293
rect 24670 7284 24676 7296
rect 24728 7324 24734 7336
rect 25133 7327 25191 7333
rect 25133 7324 25145 7327
rect 24728 7296 25145 7324
rect 24728 7284 24734 7296
rect 25133 7293 25145 7296
rect 25179 7293 25191 7327
rect 25133 7287 25191 7293
rect 17678 7216 17684 7268
rect 17736 7256 17742 7268
rect 17865 7259 17923 7265
rect 17865 7256 17877 7259
rect 17736 7228 17877 7256
rect 17736 7216 17742 7228
rect 17865 7225 17877 7228
rect 17911 7256 17923 7259
rect 19521 7259 19579 7265
rect 17911 7228 18552 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 18524 7200 18552 7228
rect 19521 7225 19533 7259
rect 19567 7256 19579 7259
rect 19567 7228 20024 7256
rect 19567 7225 19579 7228
rect 19521 7219 19579 7225
rect 19996 7200 20024 7228
rect 11882 7188 11888 7200
rect 11843 7160 11888 7188
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 18138 7148 18144 7200
rect 18196 7188 18202 7200
rect 18417 7191 18475 7197
rect 18417 7188 18429 7191
rect 18196 7160 18429 7188
rect 18196 7148 18202 7160
rect 18417 7157 18429 7160
rect 18463 7157 18475 7191
rect 18417 7151 18475 7157
rect 18506 7148 18512 7200
rect 18564 7188 18570 7200
rect 19978 7188 19984 7200
rect 18564 7160 18609 7188
rect 19939 7160 19984 7188
rect 18564 7148 18570 7160
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 23382 7148 23388 7200
rect 23440 7188 23446 7200
rect 23658 7188 23664 7200
rect 23440 7160 23664 7188
rect 23440 7148 23446 7160
rect 23658 7148 23664 7160
rect 23716 7148 23722 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 15470 6984 15476 6996
rect 15431 6956 15476 6984
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 16853 6987 16911 6993
rect 16853 6953 16865 6987
rect 16899 6984 16911 6987
rect 16942 6984 16948 6996
rect 16899 6956 16948 6984
rect 16899 6953 16911 6956
rect 16853 6947 16911 6953
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17405 6987 17463 6993
rect 17405 6953 17417 6987
rect 17451 6984 17463 6987
rect 17862 6984 17868 6996
rect 17451 6956 17868 6984
rect 17451 6953 17463 6956
rect 17405 6947 17463 6953
rect 17862 6944 17868 6956
rect 17920 6944 17926 6996
rect 19061 6987 19119 6993
rect 19061 6953 19073 6987
rect 19107 6984 19119 6987
rect 19242 6984 19248 6996
rect 19107 6956 19248 6984
rect 19107 6953 19119 6956
rect 19061 6947 19119 6953
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 19613 6987 19671 6993
rect 19613 6984 19625 6987
rect 19484 6956 19625 6984
rect 19484 6944 19490 6956
rect 19613 6953 19625 6956
rect 19659 6953 19671 6987
rect 19613 6947 19671 6953
rect 20073 6987 20131 6993
rect 20073 6953 20085 6987
rect 20119 6984 20131 6987
rect 20254 6984 20260 6996
rect 20119 6956 20260 6984
rect 20119 6953 20131 6956
rect 20073 6947 20131 6953
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 16117 6851 16175 6857
rect 16117 6817 16129 6851
rect 16163 6848 16175 6851
rect 16482 6848 16488 6860
rect 16163 6820 16488 6848
rect 16163 6817 16175 6820
rect 16117 6811 16175 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 23750 6848 23756 6860
rect 23711 6820 23756 6848
rect 23750 6808 23756 6820
rect 23808 6808 23814 6860
rect 24762 6848 24768 6860
rect 24723 6820 24768 6848
rect 24762 6808 24768 6820
rect 24820 6808 24826 6860
rect 16758 6740 16764 6792
rect 16816 6780 16822 6792
rect 16816 6752 17080 6780
rect 16816 6740 16822 6752
rect 17052 6721 17080 6752
rect 17402 6740 17408 6792
rect 17460 6780 17466 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 17460 6752 17509 6780
rect 17460 6740 17466 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 17644 6752 17689 6780
rect 17644 6740 17650 6752
rect 17037 6715 17095 6721
rect 17037 6681 17049 6715
rect 17083 6681 17095 6715
rect 17037 6675 17095 6681
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 16942 6644 16948 6656
rect 16531 6616 16948 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 16942 6604 16948 6616
rect 17000 6644 17006 6656
rect 17604 6644 17632 6740
rect 23934 6712 23940 6724
rect 23895 6684 23940 6712
rect 23934 6672 23940 6684
rect 23992 6672 23998 6724
rect 18138 6644 18144 6656
rect 17000 6616 17632 6644
rect 18099 6616 18144 6644
rect 17000 6604 17006 6616
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 15436 6412 16221 6440
rect 15436 6400 15442 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 16390 6440 16396 6452
rect 16351 6412 16396 6440
rect 16209 6403 16267 6409
rect 16224 6236 16252 6403
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17862 6440 17868 6452
rect 17823 6412 17868 6440
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 23750 6400 23756 6452
rect 23808 6440 23814 6452
rect 23845 6443 23903 6449
rect 23845 6440 23857 6443
rect 23808 6412 23857 6440
rect 23808 6400 23814 6412
rect 23845 6409 23857 6412
rect 23891 6409 23903 6443
rect 23845 6403 23903 6409
rect 16942 6304 16948 6316
rect 16903 6276 16948 6304
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 16853 6239 16911 6245
rect 16853 6236 16865 6239
rect 16224 6208 16865 6236
rect 16853 6205 16865 6208
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 16448 6072 16773 6100
rect 16448 6060 16454 6072
rect 16761 6069 16773 6072
rect 16807 6069 16819 6103
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 16761 6063 16819 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 16390 5896 16396 5908
rect 16351 5868 16396 5896
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 17037 5899 17095 5905
rect 17037 5896 17049 5899
rect 17000 5868 17049 5896
rect 17000 5856 17006 5868
rect 17037 5865 17049 5868
rect 17083 5865 17095 5899
rect 17037 5859 17095 5865
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 12437 2499 12495 2505
rect 12437 2465 12449 2499
rect 12483 2496 12495 2499
rect 13164 2499 13222 2505
rect 13164 2496 13176 2499
rect 12483 2468 13176 2496
rect 12483 2465 12495 2468
rect 12437 2459 12495 2465
rect 13164 2465 13176 2468
rect 13210 2496 13222 2499
rect 13722 2496 13728 2508
rect 13210 2468 13728 2496
rect 13210 2465 13222 2468
rect 13164 2459 13222 2465
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2428 12038 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12032 2400 12909 2428
rect 12032 2388 12038 2400
rect 12452 2372 12480 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 12434 2320 12440 2372
rect 12492 2320 12498 2372
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 10048 25984 10100 26036
rect 14832 25984 14884 26036
rect 8024 25916 8076 25968
rect 18604 25916 18656 25968
rect 13268 25848 13320 25900
rect 21548 25848 21600 25900
rect 9588 25780 9640 25832
rect 18052 25780 18104 25832
rect 10968 25712 11020 25764
rect 16304 25712 16356 25764
rect 1400 25644 1452 25696
rect 11704 25644 11756 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 1400 25483 1452 25492
rect 1400 25449 1409 25483
rect 1409 25449 1443 25483
rect 1443 25449 1452 25483
rect 1400 25440 1452 25449
rect 2872 25440 2924 25492
rect 2964 25440 3016 25492
rect 5080 25440 5132 25492
rect 7288 25440 7340 25492
rect 8024 25483 8076 25492
rect 8024 25449 8033 25483
rect 8033 25449 8067 25483
rect 8067 25449 8076 25483
rect 8024 25440 8076 25449
rect 10968 25440 11020 25492
rect 3976 25304 4028 25356
rect 8760 25304 8812 25356
rect 9588 25304 9640 25356
rect 10692 25304 10744 25356
rect 17132 25440 17184 25492
rect 20076 25440 20128 25492
rect 21824 25440 21876 25492
rect 22836 25440 22888 25492
rect 24768 25440 24820 25492
rect 2872 25279 2924 25288
rect 2872 25245 2881 25279
rect 2881 25245 2915 25279
rect 2915 25245 2924 25279
rect 2872 25236 2924 25245
rect 3056 25279 3108 25288
rect 3056 25245 3065 25279
rect 3065 25245 3099 25279
rect 3099 25245 3108 25279
rect 3056 25236 3108 25245
rect 5540 25236 5592 25288
rect 4068 25168 4120 25220
rect 5448 25168 5500 25220
rect 8300 25236 8352 25288
rect 9128 25236 9180 25288
rect 11796 25304 11848 25356
rect 11612 25279 11664 25288
rect 11612 25245 11621 25279
rect 11621 25245 11655 25279
rect 11655 25245 11664 25279
rect 11612 25236 11664 25245
rect 12992 25347 13044 25356
rect 12992 25313 13001 25347
rect 13001 25313 13035 25347
rect 13035 25313 13044 25347
rect 12992 25304 13044 25313
rect 10600 25168 10652 25220
rect 10968 25211 11020 25220
rect 10968 25177 10977 25211
rect 10977 25177 11011 25211
rect 11011 25177 11020 25211
rect 10968 25168 11020 25177
rect 1952 25143 2004 25152
rect 1952 25109 1961 25143
rect 1961 25109 1995 25143
rect 1995 25109 2004 25143
rect 1952 25100 2004 25109
rect 2320 25143 2372 25152
rect 2320 25109 2329 25143
rect 2329 25109 2363 25143
rect 2363 25109 2372 25143
rect 2320 25100 2372 25109
rect 2412 25143 2464 25152
rect 2412 25109 2421 25143
rect 2421 25109 2455 25143
rect 2455 25109 2464 25143
rect 3424 25143 3476 25152
rect 2412 25100 2464 25109
rect 3424 25109 3433 25143
rect 3433 25109 3467 25143
rect 3467 25109 3476 25143
rect 3424 25100 3476 25109
rect 3516 25100 3568 25152
rect 5080 25143 5132 25152
rect 5080 25109 5089 25143
rect 5089 25109 5123 25143
rect 5123 25109 5132 25143
rect 5080 25100 5132 25109
rect 6644 25143 6696 25152
rect 6644 25109 6653 25143
rect 6653 25109 6687 25143
rect 6687 25109 6696 25143
rect 6644 25100 6696 25109
rect 8944 25100 8996 25152
rect 9128 25143 9180 25152
rect 9128 25109 9137 25143
rect 9137 25109 9171 25143
rect 9171 25109 9180 25143
rect 9128 25100 9180 25109
rect 12716 25236 12768 25288
rect 13176 25236 13228 25288
rect 16120 25372 16172 25424
rect 21548 25415 21600 25424
rect 21548 25381 21557 25415
rect 21557 25381 21591 25415
rect 21591 25381 21600 25415
rect 23756 25415 23808 25424
rect 21548 25372 21600 25381
rect 14464 25304 14516 25356
rect 15568 25304 15620 25356
rect 16212 25304 16264 25356
rect 17040 25304 17092 25356
rect 23756 25381 23765 25415
rect 23765 25381 23799 25415
rect 23799 25381 23808 25415
rect 23756 25372 23808 25381
rect 24400 25415 24452 25424
rect 24400 25381 24409 25415
rect 24409 25381 24443 25415
rect 24443 25381 24452 25415
rect 24400 25372 24452 25381
rect 24492 25347 24544 25356
rect 16120 25279 16172 25288
rect 11980 25143 12032 25152
rect 11980 25109 11989 25143
rect 11989 25109 12023 25143
rect 12023 25109 12032 25143
rect 11980 25100 12032 25109
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 24492 25313 24501 25347
rect 24501 25313 24535 25347
rect 24535 25313 24544 25347
rect 24492 25304 24544 25313
rect 25596 25347 25648 25356
rect 25596 25313 25605 25347
rect 25605 25313 25639 25347
rect 25639 25313 25648 25347
rect 25596 25304 25648 25313
rect 20076 25236 20128 25288
rect 18512 25168 18564 25220
rect 20628 25168 20680 25220
rect 24124 25168 24176 25220
rect 24860 25236 24912 25288
rect 15292 25100 15344 25152
rect 16580 25143 16632 25152
rect 16580 25109 16589 25143
rect 16589 25109 16623 25143
rect 16623 25109 16632 25143
rect 16580 25100 16632 25109
rect 18144 25143 18196 25152
rect 18144 25109 18153 25143
rect 18153 25109 18187 25143
rect 18187 25109 18196 25143
rect 18144 25100 18196 25109
rect 22560 25100 22612 25152
rect 24032 25143 24084 25152
rect 24032 25109 24041 25143
rect 24041 25109 24075 25143
rect 24075 25109 24084 25143
rect 24032 25100 24084 25109
rect 25228 25143 25280 25152
rect 25228 25109 25237 25143
rect 25237 25109 25271 25143
rect 25271 25109 25280 25143
rect 25228 25100 25280 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1400 24896 1452 24948
rect 3516 24896 3568 24948
rect 4344 24896 4396 24948
rect 8852 24896 8904 24948
rect 10692 24939 10744 24948
rect 10692 24905 10701 24939
rect 10701 24905 10735 24939
rect 10735 24905 10744 24939
rect 10692 24896 10744 24905
rect 12992 24939 13044 24948
rect 12992 24905 13001 24939
rect 13001 24905 13035 24939
rect 13035 24905 13044 24939
rect 12992 24896 13044 24905
rect 13360 24896 13412 24948
rect 16120 24939 16172 24948
rect 5448 24828 5500 24880
rect 1676 24760 1728 24812
rect 2504 24760 2556 24812
rect 2688 24803 2740 24812
rect 2688 24769 2697 24803
rect 2697 24769 2731 24803
rect 2731 24769 2740 24803
rect 2688 24760 2740 24769
rect 12716 24828 12768 24880
rect 7104 24760 7156 24812
rect 7288 24803 7340 24812
rect 7288 24769 7297 24803
rect 7297 24769 7331 24803
rect 7331 24769 7340 24803
rect 7288 24760 7340 24769
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 13176 24760 13228 24812
rect 13820 24828 13872 24880
rect 15292 24828 15344 24880
rect 16120 24905 16129 24939
rect 16129 24905 16163 24939
rect 16163 24905 16172 24939
rect 16120 24896 16172 24905
rect 17040 24896 17092 24948
rect 18512 24939 18564 24948
rect 18512 24905 18521 24939
rect 18521 24905 18555 24939
rect 18555 24905 18564 24939
rect 18512 24896 18564 24905
rect 20628 24896 20680 24948
rect 23756 24896 23808 24948
rect 24768 24939 24820 24948
rect 24768 24905 24777 24939
rect 24777 24905 24811 24939
rect 24811 24905 24820 24939
rect 24768 24896 24820 24905
rect 21456 24871 21508 24880
rect 21456 24837 21465 24871
rect 21465 24837 21499 24871
rect 21499 24837 21508 24871
rect 21456 24828 21508 24837
rect 2412 24692 2464 24744
rect 3240 24692 3292 24744
rect 3424 24735 3476 24744
rect 3424 24701 3458 24735
rect 3458 24701 3476 24735
rect 3424 24692 3476 24701
rect 4436 24692 4488 24744
rect 5448 24692 5500 24744
rect 6552 24692 6604 24744
rect 7012 24692 7064 24744
rect 8300 24692 8352 24744
rect 8484 24735 8536 24744
rect 8484 24701 8493 24735
rect 8493 24701 8527 24735
rect 8527 24701 8536 24735
rect 8484 24692 8536 24701
rect 11980 24692 12032 24744
rect 2228 24624 2280 24676
rect 1952 24556 2004 24608
rect 2688 24624 2740 24676
rect 8116 24624 8168 24676
rect 9128 24624 9180 24676
rect 9588 24624 9640 24676
rect 11612 24624 11664 24676
rect 12164 24624 12216 24676
rect 2872 24556 2924 24608
rect 3332 24556 3384 24608
rect 3884 24556 3936 24608
rect 4804 24556 4856 24608
rect 6736 24556 6788 24608
rect 7196 24599 7248 24608
rect 7196 24565 7205 24599
rect 7205 24565 7239 24599
rect 7239 24565 7248 24599
rect 7196 24556 7248 24565
rect 9864 24599 9916 24608
rect 9864 24565 9873 24599
rect 9873 24565 9907 24599
rect 9907 24565 9916 24599
rect 9864 24556 9916 24565
rect 11520 24599 11572 24608
rect 11520 24565 11529 24599
rect 11529 24565 11563 24599
rect 11563 24565 11572 24599
rect 11520 24556 11572 24565
rect 12900 24667 12952 24676
rect 12900 24633 12909 24667
rect 12909 24633 12943 24667
rect 12943 24633 12952 24667
rect 12900 24624 12952 24633
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 18972 24760 19024 24812
rect 22560 24803 22612 24812
rect 22560 24769 22569 24803
rect 22569 24769 22603 24803
rect 22603 24769 22612 24803
rect 22560 24760 22612 24769
rect 14740 24624 14792 24676
rect 16212 24692 16264 24744
rect 16580 24735 16632 24744
rect 16580 24701 16589 24735
rect 16589 24701 16623 24735
rect 16623 24701 16632 24735
rect 16580 24692 16632 24701
rect 18144 24692 18196 24744
rect 13728 24556 13780 24608
rect 14004 24599 14056 24608
rect 14004 24565 14013 24599
rect 14013 24565 14047 24599
rect 14047 24565 14056 24599
rect 14004 24556 14056 24565
rect 14832 24556 14884 24608
rect 15476 24599 15528 24608
rect 15476 24565 15485 24599
rect 15485 24565 15519 24599
rect 15519 24565 15528 24599
rect 15476 24556 15528 24565
rect 16764 24599 16816 24608
rect 16764 24565 16773 24599
rect 16773 24565 16807 24599
rect 16807 24565 16816 24599
rect 16764 24556 16816 24565
rect 17040 24556 17092 24608
rect 21456 24692 21508 24744
rect 22284 24692 22336 24744
rect 22652 24692 22704 24744
rect 23756 24760 23808 24812
rect 24860 24760 24912 24812
rect 25228 24735 25280 24744
rect 18880 24599 18932 24608
rect 18880 24565 18889 24599
rect 18889 24565 18923 24599
rect 18923 24565 18932 24599
rect 18880 24556 18932 24565
rect 19248 24599 19300 24608
rect 19248 24565 19257 24599
rect 19257 24565 19291 24599
rect 19291 24565 19300 24599
rect 19248 24556 19300 24565
rect 19432 24556 19484 24608
rect 21916 24667 21968 24676
rect 21916 24633 21925 24667
rect 21925 24633 21959 24667
rect 21959 24633 21968 24667
rect 21916 24624 21968 24633
rect 25228 24701 25237 24735
rect 25237 24701 25271 24735
rect 25271 24701 25280 24735
rect 25228 24692 25280 24701
rect 23940 24624 23992 24676
rect 25136 24624 25188 24676
rect 25596 24624 25648 24676
rect 20444 24599 20496 24608
rect 20444 24565 20453 24599
rect 20453 24565 20487 24599
rect 20487 24565 20496 24599
rect 20444 24556 20496 24565
rect 20536 24556 20588 24608
rect 22008 24599 22060 24608
rect 22008 24565 22017 24599
rect 22017 24565 22051 24599
rect 22051 24565 22060 24599
rect 22008 24556 22060 24565
rect 23204 24556 23256 24608
rect 23664 24599 23716 24608
rect 23664 24565 23673 24599
rect 23673 24565 23707 24599
rect 23707 24565 23716 24599
rect 23664 24556 23716 24565
rect 25412 24599 25464 24608
rect 25412 24565 25421 24599
rect 25421 24565 25455 24599
rect 25455 24565 25464 24599
rect 25412 24556 25464 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1676 24352 1728 24404
rect 3056 24352 3108 24404
rect 3884 24395 3936 24404
rect 3884 24361 3893 24395
rect 3893 24361 3927 24395
rect 3927 24361 3936 24395
rect 3884 24352 3936 24361
rect 4160 24352 4212 24404
rect 4712 24352 4764 24404
rect 6920 24352 6972 24404
rect 7472 24352 7524 24404
rect 8116 24395 8168 24404
rect 8116 24361 8125 24395
rect 8125 24361 8159 24395
rect 8159 24361 8168 24395
rect 8116 24352 8168 24361
rect 8760 24395 8812 24404
rect 8760 24361 8769 24395
rect 8769 24361 8803 24395
rect 8803 24361 8812 24395
rect 8760 24352 8812 24361
rect 9864 24352 9916 24404
rect 10692 24395 10744 24404
rect 10692 24361 10701 24395
rect 10701 24361 10735 24395
rect 10735 24361 10744 24395
rect 10692 24352 10744 24361
rect 11152 24395 11204 24404
rect 11152 24361 11161 24395
rect 11161 24361 11195 24395
rect 11195 24361 11204 24395
rect 11152 24352 11204 24361
rect 11796 24395 11848 24404
rect 11796 24361 11805 24395
rect 11805 24361 11839 24395
rect 11839 24361 11848 24395
rect 11796 24352 11848 24361
rect 14648 24352 14700 24404
rect 18052 24352 18104 24404
rect 19340 24395 19392 24404
rect 19340 24361 19349 24395
rect 19349 24361 19383 24395
rect 19383 24361 19392 24395
rect 19340 24352 19392 24361
rect 20076 24395 20128 24404
rect 20076 24361 20085 24395
rect 20085 24361 20119 24395
rect 20119 24361 20128 24395
rect 20076 24352 20128 24361
rect 22008 24352 22060 24404
rect 24124 24352 24176 24404
rect 24216 24352 24268 24404
rect 25320 24352 25372 24404
rect 2504 24284 2556 24336
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 1952 24216 2004 24268
rect 6092 24284 6144 24336
rect 10876 24284 10928 24336
rect 11244 24284 11296 24336
rect 12072 24284 12124 24336
rect 17592 24284 17644 24336
rect 24032 24284 24084 24336
rect 3332 24148 3384 24200
rect 6368 24216 6420 24268
rect 8116 24216 8168 24268
rect 12716 24259 12768 24268
rect 12716 24225 12725 24259
rect 12725 24225 12759 24259
rect 12759 24225 12768 24259
rect 12716 24216 12768 24225
rect 14648 24216 14700 24268
rect 16120 24259 16172 24268
rect 16120 24225 16129 24259
rect 16129 24225 16163 24259
rect 16163 24225 16172 24259
rect 16120 24216 16172 24225
rect 17408 24216 17460 24268
rect 19064 24216 19116 24268
rect 22468 24216 22520 24268
rect 23296 24216 23348 24268
rect 24860 24216 24912 24268
rect 4620 24191 4672 24200
rect 4620 24157 4629 24191
rect 4629 24157 4663 24191
rect 4663 24157 4672 24191
rect 4620 24148 4672 24157
rect 5356 24148 5408 24200
rect 5540 24123 5592 24132
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 5540 24089 5549 24123
rect 5549 24089 5583 24123
rect 5583 24089 5592 24123
rect 5540 24080 5592 24089
rect 3240 24012 3292 24064
rect 3976 24012 4028 24064
rect 4160 24055 4212 24064
rect 4160 24021 4169 24055
rect 4169 24021 4203 24055
rect 4203 24021 4212 24055
rect 4160 24012 4212 24021
rect 5356 24012 5408 24064
rect 9312 24148 9364 24200
rect 11796 24148 11848 24200
rect 13728 24148 13780 24200
rect 15752 24148 15804 24200
rect 16212 24191 16264 24200
rect 16212 24157 16221 24191
rect 16221 24157 16255 24191
rect 16255 24157 16264 24191
rect 16212 24148 16264 24157
rect 16304 24191 16356 24200
rect 16304 24157 16313 24191
rect 16313 24157 16347 24191
rect 16347 24157 16356 24191
rect 17224 24191 17276 24200
rect 16304 24148 16356 24157
rect 17224 24157 17233 24191
rect 17233 24157 17267 24191
rect 17267 24157 17276 24191
rect 17224 24148 17276 24157
rect 21456 24148 21508 24200
rect 7104 24123 7156 24132
rect 7104 24089 7113 24123
rect 7113 24089 7147 24123
rect 7147 24089 7156 24123
rect 7104 24080 7156 24089
rect 10784 24080 10836 24132
rect 17408 24080 17460 24132
rect 21640 24123 21692 24132
rect 21640 24089 21649 24123
rect 21649 24089 21683 24123
rect 21683 24089 21692 24123
rect 23572 24148 23624 24200
rect 21640 24080 21692 24089
rect 23204 24080 23256 24132
rect 25780 24148 25832 24200
rect 6000 24012 6052 24064
rect 8300 24012 8352 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 12256 24055 12308 24064
rect 12256 24021 12265 24055
rect 12265 24021 12299 24055
rect 12299 24021 12308 24055
rect 12256 24012 12308 24021
rect 12992 24012 13044 24064
rect 14464 24012 14516 24064
rect 14740 24012 14792 24064
rect 16488 24012 16540 24064
rect 17316 24055 17368 24064
rect 17316 24021 17325 24055
rect 17325 24021 17359 24055
rect 17359 24021 17368 24055
rect 17316 24012 17368 24021
rect 19064 24055 19116 24064
rect 19064 24021 19073 24055
rect 19073 24021 19107 24055
rect 19107 24021 19116 24055
rect 19064 24012 19116 24021
rect 20536 24055 20588 24064
rect 20536 24021 20545 24055
rect 20545 24021 20579 24055
rect 20579 24021 20588 24055
rect 20536 24012 20588 24021
rect 21732 24055 21784 24064
rect 21732 24021 21741 24055
rect 21741 24021 21775 24055
rect 21775 24021 21784 24055
rect 21732 24012 21784 24021
rect 23848 24012 23900 24064
rect 24860 24055 24912 24064
rect 24860 24021 24869 24055
rect 24869 24021 24903 24055
rect 24903 24021 24912 24055
rect 24860 24012 24912 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1768 23808 1820 23860
rect 1952 23851 2004 23860
rect 1952 23817 1961 23851
rect 1961 23817 1995 23851
rect 1995 23817 2004 23851
rect 1952 23808 2004 23817
rect 8116 23808 8168 23860
rect 9312 23851 9364 23860
rect 9312 23817 9321 23851
rect 9321 23817 9355 23851
rect 9355 23817 9364 23851
rect 9312 23808 9364 23817
rect 11796 23851 11848 23860
rect 11796 23817 11805 23851
rect 11805 23817 11839 23851
rect 11839 23817 11848 23851
rect 11796 23808 11848 23817
rect 5356 23783 5408 23792
rect 5356 23749 5365 23783
rect 5365 23749 5399 23783
rect 5399 23749 5408 23783
rect 5356 23740 5408 23749
rect 8024 23740 8076 23792
rect 8484 23740 8536 23792
rect 9128 23740 9180 23792
rect 11520 23740 11572 23792
rect 12716 23808 12768 23860
rect 14004 23808 14056 23860
rect 14556 23808 14608 23860
rect 16212 23808 16264 23860
rect 16396 23808 16448 23860
rect 16580 23808 16632 23860
rect 17408 23851 17460 23860
rect 17408 23817 17417 23851
rect 17417 23817 17451 23851
rect 17451 23817 17460 23851
rect 17408 23808 17460 23817
rect 17592 23808 17644 23860
rect 19064 23808 19116 23860
rect 22468 23808 22520 23860
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 25412 23851 25464 23860
rect 25412 23817 25421 23851
rect 25421 23817 25455 23851
rect 25455 23817 25464 23851
rect 25412 23808 25464 23817
rect 25780 23851 25832 23860
rect 25780 23817 25789 23851
rect 25789 23817 25823 23851
rect 25823 23817 25832 23851
rect 25780 23808 25832 23817
rect 12072 23740 12124 23792
rect 19340 23783 19392 23792
rect 19340 23749 19349 23783
rect 19349 23749 19383 23783
rect 19383 23749 19392 23783
rect 19340 23740 19392 23749
rect 19984 23740 20036 23792
rect 20444 23740 20496 23792
rect 3240 23672 3292 23724
rect 3976 23715 4028 23724
rect 3976 23681 3985 23715
rect 3985 23681 4019 23715
rect 4019 23681 4028 23715
rect 3976 23672 4028 23681
rect 6368 23715 6420 23724
rect 6368 23681 6377 23715
rect 6377 23681 6411 23715
rect 6411 23681 6420 23715
rect 6368 23672 6420 23681
rect 8760 23672 8812 23724
rect 12992 23715 13044 23724
rect 2136 23604 2188 23656
rect 2504 23604 2556 23656
rect 2780 23647 2832 23656
rect 2780 23613 2789 23647
rect 2789 23613 2823 23647
rect 2823 23613 2832 23647
rect 2780 23604 2832 23613
rect 3424 23604 3476 23656
rect 3884 23604 3936 23656
rect 4528 23536 4580 23588
rect 9312 23604 9364 23656
rect 8116 23579 8168 23588
rect 8116 23545 8125 23579
rect 8125 23545 8159 23579
rect 8159 23545 8168 23579
rect 8116 23536 8168 23545
rect 9864 23604 9916 23656
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 18236 23672 18288 23724
rect 18972 23715 19024 23724
rect 18972 23681 18981 23715
rect 18981 23681 19015 23715
rect 19015 23681 19024 23715
rect 18972 23672 19024 23681
rect 24124 23715 24176 23724
rect 24124 23681 24133 23715
rect 24133 23681 24167 23715
rect 24167 23681 24176 23715
rect 24124 23672 24176 23681
rect 24308 23715 24360 23724
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 15384 23604 15436 23656
rect 15752 23647 15804 23656
rect 15752 23613 15786 23647
rect 15786 23613 15804 23647
rect 15752 23604 15804 23613
rect 18052 23604 18104 23656
rect 20260 23604 20312 23656
rect 11520 23536 11572 23588
rect 13544 23536 13596 23588
rect 2780 23468 2832 23520
rect 3056 23468 3108 23520
rect 4804 23468 4856 23520
rect 6000 23511 6052 23520
rect 6000 23477 6009 23511
rect 6009 23477 6043 23511
rect 6043 23477 6052 23511
rect 6000 23468 6052 23477
rect 6184 23468 6236 23520
rect 7012 23511 7064 23520
rect 7012 23477 7021 23511
rect 7021 23477 7055 23511
rect 7055 23477 7064 23511
rect 7012 23468 7064 23477
rect 7104 23468 7156 23520
rect 8208 23511 8260 23520
rect 8208 23477 8217 23511
rect 8217 23477 8251 23511
rect 8251 23477 8260 23511
rect 8208 23468 8260 23477
rect 8668 23511 8720 23520
rect 8668 23477 8677 23511
rect 8677 23477 8711 23511
rect 8711 23477 8720 23511
rect 8668 23468 8720 23477
rect 11152 23511 11204 23520
rect 11152 23477 11161 23511
rect 11161 23477 11195 23511
rect 11195 23477 11204 23511
rect 11152 23468 11204 23477
rect 11888 23468 11940 23520
rect 14924 23468 14976 23520
rect 16120 23468 16172 23520
rect 20996 23604 21048 23656
rect 24032 23647 24084 23656
rect 23572 23536 23624 23588
rect 24032 23613 24041 23647
rect 24041 23613 24075 23647
rect 24075 23613 24084 23647
rect 24032 23604 24084 23613
rect 25596 23604 25648 23656
rect 24308 23536 24360 23588
rect 21548 23468 21600 23520
rect 21640 23468 21692 23520
rect 23296 23511 23348 23520
rect 23296 23477 23305 23511
rect 23305 23477 23339 23511
rect 23339 23477 23348 23511
rect 23296 23468 23348 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 3608 23264 3660 23316
rect 1308 23196 1360 23248
rect 4620 23264 4672 23316
rect 4712 23307 4764 23316
rect 4712 23273 4721 23307
rect 4721 23273 4755 23307
rect 4755 23273 4764 23307
rect 4712 23264 4764 23273
rect 6828 23264 6880 23316
rect 8208 23264 8260 23316
rect 8576 23264 8628 23316
rect 10876 23264 10928 23316
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 13176 23264 13228 23316
rect 18236 23264 18288 23316
rect 18972 23264 19024 23316
rect 19340 23264 19392 23316
rect 21456 23307 21508 23316
rect 21456 23273 21465 23307
rect 21465 23273 21499 23307
rect 21499 23273 21508 23307
rect 21456 23264 21508 23273
rect 22928 23307 22980 23316
rect 22928 23273 22937 23307
rect 22937 23273 22971 23307
rect 22971 23273 22980 23307
rect 22928 23264 22980 23273
rect 23664 23264 23716 23316
rect 7748 23196 7800 23248
rect 8944 23196 8996 23248
rect 11796 23239 11848 23248
rect 11796 23205 11830 23239
rect 11830 23205 11848 23239
rect 11796 23196 11848 23205
rect 16212 23196 16264 23248
rect 16396 23239 16448 23248
rect 16396 23205 16430 23239
rect 16430 23205 16448 23239
rect 16396 23196 16448 23205
rect 19984 23196 20036 23248
rect 21640 23196 21692 23248
rect 24860 23264 24912 23316
rect 25320 23264 25372 23316
rect 25688 23264 25740 23316
rect 24768 23196 24820 23248
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 2780 23128 2832 23137
rect 3240 23128 3292 23180
rect 3884 23128 3936 23180
rect 3976 23128 4028 23180
rect 1952 23035 2004 23044
rect 1952 23001 1961 23035
rect 1961 23001 1995 23035
rect 1995 23001 2004 23035
rect 1952 22992 2004 23001
rect 3240 22992 3292 23044
rect 5172 23171 5224 23180
rect 5172 23137 5206 23171
rect 5206 23137 5224 23171
rect 10048 23171 10100 23180
rect 5172 23128 5224 23137
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 11336 23128 11388 23180
rect 11520 23171 11572 23180
rect 11520 23137 11529 23171
rect 11529 23137 11563 23171
rect 11563 23137 11572 23171
rect 11520 23128 11572 23137
rect 13912 23128 13964 23180
rect 4160 23060 4212 23112
rect 4804 23060 4856 23112
rect 8668 23103 8720 23112
rect 8668 23069 8677 23103
rect 8677 23069 8711 23103
rect 8711 23069 8720 23103
rect 8668 23060 8720 23069
rect 15108 23103 15160 23112
rect 6644 22992 6696 23044
rect 9496 22992 9548 23044
rect 9864 22992 9916 23044
rect 15108 23069 15117 23103
rect 15117 23069 15151 23103
rect 15151 23069 15160 23103
rect 15108 23060 15160 23069
rect 2320 22967 2372 22976
rect 2320 22933 2329 22967
rect 2329 22933 2363 22967
rect 2363 22933 2372 22967
rect 2320 22924 2372 22933
rect 2504 22924 2556 22976
rect 3792 22967 3844 22976
rect 3792 22933 3801 22967
rect 3801 22933 3835 22967
rect 3835 22933 3844 22967
rect 3792 22924 3844 22933
rect 3884 22924 3936 22976
rect 6920 22967 6972 22976
rect 6920 22933 6929 22967
rect 6929 22933 6963 22967
rect 6963 22933 6972 22967
rect 6920 22924 6972 22933
rect 13544 22967 13596 22976
rect 13544 22933 13553 22967
rect 13553 22933 13587 22967
rect 13587 22933 13596 22967
rect 13544 22924 13596 22933
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 15384 22924 15436 22976
rect 20996 23060 21048 23112
rect 21548 23103 21600 23112
rect 21548 23069 21557 23103
rect 21557 23069 21591 23103
rect 21591 23069 21600 23103
rect 21548 23060 21600 23069
rect 17500 23035 17552 23044
rect 17500 23001 17509 23035
rect 17509 23001 17543 23035
rect 17543 23001 17552 23035
rect 17500 22992 17552 23001
rect 21456 22992 21508 23044
rect 24308 22992 24360 23044
rect 24676 22992 24728 23044
rect 16304 22924 16356 22976
rect 20260 22967 20312 22976
rect 20260 22933 20269 22967
rect 20269 22933 20303 22967
rect 20303 22933 20312 22967
rect 20260 22924 20312 22933
rect 23204 22924 23256 22976
rect 24124 22924 24176 22976
rect 25596 22924 25648 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2780 22720 2832 22772
rect 3516 22720 3568 22772
rect 4436 22763 4488 22772
rect 4436 22729 4445 22763
rect 4445 22729 4479 22763
rect 4479 22729 4488 22763
rect 4436 22720 4488 22729
rect 6460 22720 6512 22772
rect 2320 22584 2372 22636
rect 2504 22584 2556 22636
rect 1768 22516 1820 22568
rect 1952 22516 2004 22568
rect 3608 22652 3660 22704
rect 2780 22584 2832 22636
rect 2964 22584 3016 22636
rect 4988 22652 5040 22704
rect 3884 22627 3936 22636
rect 3884 22593 3893 22627
rect 3893 22593 3927 22627
rect 3927 22593 3936 22627
rect 3884 22584 3936 22593
rect 5356 22627 5408 22636
rect 5356 22593 5365 22627
rect 5365 22593 5399 22627
rect 5399 22593 5408 22627
rect 5356 22584 5408 22593
rect 4068 22516 4120 22568
rect 5080 22516 5132 22568
rect 5264 22559 5316 22568
rect 5264 22525 5273 22559
rect 5273 22525 5307 22559
rect 5307 22525 5316 22559
rect 5264 22516 5316 22525
rect 4436 22448 4488 22500
rect 8668 22720 8720 22772
rect 8760 22720 8812 22772
rect 11336 22720 11388 22772
rect 11796 22720 11848 22772
rect 14648 22720 14700 22772
rect 16396 22763 16448 22772
rect 16396 22729 16405 22763
rect 16405 22729 16439 22763
rect 16439 22729 16448 22763
rect 16396 22720 16448 22729
rect 18972 22720 19024 22772
rect 19800 22720 19852 22772
rect 20996 22763 21048 22772
rect 20996 22729 21005 22763
rect 21005 22729 21039 22763
rect 21039 22729 21048 22763
rect 20996 22720 21048 22729
rect 22744 22720 22796 22772
rect 24860 22720 24912 22772
rect 26148 22720 26200 22772
rect 10048 22652 10100 22704
rect 15200 22652 15252 22704
rect 16028 22652 16080 22704
rect 16488 22652 16540 22704
rect 22192 22652 22244 22704
rect 8024 22627 8076 22636
rect 8024 22593 8033 22627
rect 8033 22593 8067 22627
rect 8067 22593 8076 22627
rect 8024 22584 8076 22593
rect 10968 22627 11020 22636
rect 10968 22593 10977 22627
rect 10977 22593 11011 22627
rect 11011 22593 11020 22627
rect 10968 22584 11020 22593
rect 9772 22516 9824 22568
rect 16580 22584 16632 22636
rect 21640 22584 21692 22636
rect 8116 22448 8168 22500
rect 10784 22448 10836 22500
rect 10968 22448 11020 22500
rect 1308 22380 1360 22432
rect 1860 22380 1912 22432
rect 3792 22380 3844 22432
rect 4804 22423 4856 22432
rect 4804 22389 4813 22423
rect 4813 22389 4847 22423
rect 4847 22389 4856 22423
rect 4804 22380 4856 22389
rect 6184 22380 6236 22432
rect 7012 22423 7064 22432
rect 7012 22389 7021 22423
rect 7021 22389 7055 22423
rect 7055 22389 7064 22423
rect 7012 22380 7064 22389
rect 9772 22380 9824 22432
rect 9864 22380 9916 22432
rect 12348 22380 12400 22432
rect 12716 22423 12768 22432
rect 12716 22389 12725 22423
rect 12725 22389 12759 22423
rect 12759 22389 12768 22423
rect 12716 22380 12768 22389
rect 13452 22423 13504 22432
rect 13452 22389 13461 22423
rect 13461 22389 13495 22423
rect 13495 22389 13504 22423
rect 13452 22380 13504 22389
rect 13544 22380 13596 22432
rect 15384 22516 15436 22568
rect 16396 22516 16448 22568
rect 17776 22516 17828 22568
rect 18420 22559 18472 22568
rect 18420 22525 18429 22559
rect 18429 22525 18463 22559
rect 18463 22525 18472 22559
rect 18420 22516 18472 22525
rect 13820 22448 13872 22500
rect 16764 22491 16816 22500
rect 16764 22457 16773 22491
rect 16773 22457 16807 22491
rect 16807 22457 16816 22491
rect 16764 22448 16816 22457
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 18880 22380 18932 22432
rect 19340 22380 19392 22432
rect 21548 22559 21600 22568
rect 21548 22525 21557 22559
rect 21557 22525 21591 22559
rect 21591 22525 21600 22559
rect 21548 22516 21600 22525
rect 19800 22448 19852 22500
rect 24124 22559 24176 22568
rect 24124 22525 24133 22559
rect 24133 22525 24167 22559
rect 24167 22525 24176 22559
rect 24124 22516 24176 22525
rect 25228 22559 25280 22568
rect 25228 22525 25237 22559
rect 25237 22525 25271 22559
rect 25271 22525 25280 22559
rect 25228 22516 25280 22525
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 23112 22423 23164 22432
rect 23112 22389 23121 22423
rect 23121 22389 23155 22423
rect 23155 22389 23164 22423
rect 23112 22380 23164 22389
rect 24676 22423 24728 22432
rect 24676 22389 24685 22423
rect 24685 22389 24719 22423
rect 24719 22389 24728 22423
rect 24676 22380 24728 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1676 22176 1728 22228
rect 2504 22176 2556 22228
rect 3240 22176 3292 22228
rect 3884 22176 3936 22228
rect 5172 22219 5224 22228
rect 5172 22185 5181 22219
rect 5181 22185 5215 22219
rect 5215 22185 5224 22219
rect 5172 22176 5224 22185
rect 5264 22176 5316 22228
rect 8576 22219 8628 22228
rect 8576 22185 8585 22219
rect 8585 22185 8619 22219
rect 8619 22185 8628 22219
rect 8576 22176 8628 22185
rect 9496 22219 9548 22228
rect 9496 22185 9505 22219
rect 9505 22185 9539 22219
rect 9539 22185 9548 22219
rect 9496 22176 9548 22185
rect 9956 22176 10008 22228
rect 10140 22176 10192 22228
rect 10968 22219 11020 22228
rect 10968 22185 10977 22219
rect 10977 22185 11011 22219
rect 11011 22185 11020 22219
rect 10968 22176 11020 22185
rect 16212 22219 16264 22228
rect 16212 22185 16221 22219
rect 16221 22185 16255 22219
rect 16255 22185 16264 22219
rect 16212 22176 16264 22185
rect 16764 22219 16816 22228
rect 16764 22185 16773 22219
rect 16773 22185 16807 22219
rect 16807 22185 16816 22219
rect 16764 22176 16816 22185
rect 22192 22219 22244 22228
rect 22192 22185 22201 22219
rect 22201 22185 22235 22219
rect 22235 22185 22244 22219
rect 22192 22176 22244 22185
rect 23112 22176 23164 22228
rect 4436 22151 4488 22160
rect 4436 22117 4445 22151
rect 4445 22117 4479 22151
rect 4479 22117 4488 22151
rect 4436 22108 4488 22117
rect 6000 22108 6052 22160
rect 6828 22108 6880 22160
rect 10048 22108 10100 22160
rect 10600 22108 10652 22160
rect 12256 22108 12308 22160
rect 13176 22108 13228 22160
rect 16672 22108 16724 22160
rect 1860 22040 1912 22092
rect 3424 22040 3476 22092
rect 3792 22040 3844 22092
rect 6092 22040 6144 22092
rect 11336 22083 11388 22092
rect 11336 22049 11345 22083
rect 11345 22049 11379 22083
rect 11379 22049 11388 22083
rect 11336 22040 11388 22049
rect 14556 22040 14608 22092
rect 15568 22040 15620 22092
rect 17776 22083 17828 22092
rect 17776 22049 17785 22083
rect 17785 22049 17819 22083
rect 17819 22049 17828 22083
rect 17776 22040 17828 22049
rect 17868 22040 17920 22092
rect 24124 22176 24176 22228
rect 24768 22219 24820 22228
rect 24768 22185 24777 22219
rect 24777 22185 24811 22219
rect 24811 22185 24820 22219
rect 24768 22176 24820 22185
rect 23848 22151 23900 22160
rect 23848 22117 23857 22151
rect 23857 22117 23891 22151
rect 23891 22117 23900 22151
rect 23848 22108 23900 22117
rect 1952 21972 2004 22024
rect 2228 21972 2280 22024
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 5172 21972 5224 22024
rect 6184 22015 6236 22024
rect 6184 21981 6193 22015
rect 6193 21981 6227 22015
rect 6227 21981 6236 22015
rect 6184 21972 6236 21981
rect 8392 21972 8444 22024
rect 9036 21972 9088 22024
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 11152 21972 11204 22024
rect 13912 21972 13964 22024
rect 15476 21972 15528 22024
rect 15752 21972 15804 22024
rect 17132 21972 17184 22024
rect 17592 21972 17644 22024
rect 18052 21972 18104 22024
rect 21732 21972 21784 22024
rect 22008 21972 22060 22024
rect 22560 21972 22612 22024
rect 22928 21972 22980 22024
rect 23480 21972 23532 22024
rect 24676 22108 24728 22160
rect 24216 22040 24268 22092
rect 24860 22040 24912 22092
rect 25228 22040 25280 22092
rect 1400 21904 1452 21956
rect 3424 21904 3476 21956
rect 12440 21904 12492 21956
rect 14372 21904 14424 21956
rect 15384 21904 15436 21956
rect 15844 21947 15896 21956
rect 15844 21913 15853 21947
rect 15853 21913 15887 21947
rect 15887 21913 15896 21947
rect 15844 21904 15896 21913
rect 19708 21947 19760 21956
rect 19708 21913 19717 21947
rect 19717 21913 19751 21947
rect 19751 21913 19760 21947
rect 19708 21904 19760 21913
rect 21548 21947 21600 21956
rect 21548 21913 21557 21947
rect 21557 21913 21591 21947
rect 21591 21913 21600 21947
rect 21548 21904 21600 21913
rect 25872 21904 25924 21956
rect 2228 21836 2280 21888
rect 2504 21836 2556 21888
rect 3608 21836 3660 21888
rect 7564 21879 7616 21888
rect 7564 21845 7573 21879
rect 7573 21845 7607 21879
rect 7607 21845 7616 21879
rect 7564 21836 7616 21845
rect 8116 21879 8168 21888
rect 8116 21845 8125 21879
rect 8125 21845 8159 21879
rect 8159 21845 8168 21879
rect 8116 21836 8168 21845
rect 10876 21836 10928 21888
rect 12164 21836 12216 21888
rect 12532 21836 12584 21888
rect 13820 21836 13872 21888
rect 15476 21879 15528 21888
rect 15476 21845 15485 21879
rect 15485 21845 15519 21879
rect 15519 21845 15528 21879
rect 15476 21836 15528 21845
rect 16580 21836 16632 21888
rect 17776 21836 17828 21888
rect 18696 21836 18748 21888
rect 19524 21836 19576 21888
rect 21180 21836 21232 21888
rect 23664 21836 23716 21888
rect 23940 21836 23992 21888
rect 24768 21836 24820 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1676 21632 1728 21684
rect 2688 21632 2740 21684
rect 5172 21632 5224 21684
rect 6000 21632 6052 21684
rect 8300 21675 8352 21684
rect 8300 21641 8309 21675
rect 8309 21641 8343 21675
rect 8343 21641 8352 21675
rect 8300 21632 8352 21641
rect 10232 21675 10284 21684
rect 10232 21641 10241 21675
rect 10241 21641 10275 21675
rect 10275 21641 10284 21675
rect 10232 21632 10284 21641
rect 10600 21675 10652 21684
rect 10600 21641 10609 21675
rect 10609 21641 10643 21675
rect 10643 21641 10652 21675
rect 10600 21632 10652 21641
rect 11152 21632 11204 21684
rect 12256 21675 12308 21684
rect 1952 21564 2004 21616
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 12164 21564 12216 21616
rect 6184 21496 6236 21548
rect 7564 21496 7616 21548
rect 7748 21496 7800 21548
rect 9404 21496 9456 21548
rect 1400 21428 1452 21480
rect 2504 21428 2556 21480
rect 1768 21292 1820 21344
rect 3608 21403 3660 21412
rect 3608 21369 3642 21403
rect 3642 21369 3660 21403
rect 3608 21360 3660 21369
rect 3700 21292 3752 21344
rect 7196 21471 7248 21480
rect 7196 21437 7205 21471
rect 7205 21437 7239 21471
rect 7239 21437 7248 21471
rect 7196 21428 7248 21437
rect 7288 21471 7340 21480
rect 7288 21437 7297 21471
rect 7297 21437 7331 21471
rect 7331 21437 7340 21471
rect 7288 21428 7340 21437
rect 9956 21496 10008 21548
rect 10508 21496 10560 21548
rect 11336 21539 11388 21548
rect 11336 21505 11345 21539
rect 11345 21505 11379 21539
rect 11379 21505 11388 21539
rect 11336 21496 11388 21505
rect 13544 21632 13596 21684
rect 15384 21632 15436 21684
rect 16396 21675 16448 21684
rect 16396 21641 16405 21675
rect 16405 21641 16439 21675
rect 16439 21641 16448 21675
rect 16396 21632 16448 21641
rect 17868 21675 17920 21684
rect 17868 21641 17877 21675
rect 17877 21641 17911 21675
rect 17911 21641 17920 21675
rect 17868 21632 17920 21641
rect 21456 21675 21508 21684
rect 21456 21641 21465 21675
rect 21465 21641 21499 21675
rect 21499 21641 21508 21675
rect 21456 21632 21508 21641
rect 22560 21675 22612 21684
rect 22560 21641 22569 21675
rect 22569 21641 22603 21675
rect 22603 21641 22612 21675
rect 22560 21632 22612 21641
rect 23480 21632 23532 21684
rect 23940 21632 23992 21684
rect 24676 21632 24728 21684
rect 25504 21675 25556 21684
rect 25504 21641 25513 21675
rect 25513 21641 25547 21675
rect 25547 21641 25556 21675
rect 25504 21632 25556 21641
rect 15476 21496 15528 21548
rect 17040 21539 17092 21548
rect 17040 21505 17049 21539
rect 17049 21505 17083 21539
rect 17083 21505 17092 21539
rect 17040 21496 17092 21505
rect 17592 21496 17644 21548
rect 20904 21539 20956 21548
rect 20904 21505 20913 21539
rect 20913 21505 20947 21539
rect 20947 21505 20956 21539
rect 20904 21496 20956 21505
rect 22100 21496 22152 21548
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 24768 21496 24820 21548
rect 11244 21471 11296 21480
rect 11244 21437 11253 21471
rect 11253 21437 11287 21471
rect 11287 21437 11296 21471
rect 11244 21428 11296 21437
rect 12440 21428 12492 21480
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 13360 21428 13412 21480
rect 16672 21428 16724 21480
rect 9588 21403 9640 21412
rect 9588 21369 9597 21403
rect 9597 21369 9631 21403
rect 9631 21369 9640 21403
rect 9588 21360 9640 21369
rect 12348 21360 12400 21412
rect 16396 21360 16448 21412
rect 6368 21292 6420 21344
rect 6460 21292 6512 21344
rect 9220 21335 9272 21344
rect 9220 21301 9229 21335
rect 9229 21301 9263 21335
rect 9263 21301 9272 21335
rect 9220 21292 9272 21301
rect 9772 21292 9824 21344
rect 13820 21292 13872 21344
rect 16948 21292 17000 21344
rect 17132 21292 17184 21344
rect 18052 21292 18104 21344
rect 19064 21428 19116 21480
rect 20536 21428 20588 21480
rect 21916 21428 21968 21480
rect 18696 21360 18748 21412
rect 19432 21360 19484 21412
rect 21548 21360 21600 21412
rect 20352 21335 20404 21344
rect 20352 21301 20361 21335
rect 20361 21301 20395 21335
rect 20395 21301 20404 21335
rect 20352 21292 20404 21301
rect 21640 21292 21692 21344
rect 23388 21428 23440 21480
rect 23480 21360 23532 21412
rect 24860 21428 24912 21480
rect 25320 21471 25372 21480
rect 25320 21437 25329 21471
rect 25329 21437 25363 21471
rect 25363 21437 25372 21471
rect 25320 21428 25372 21437
rect 23848 21360 23900 21412
rect 25780 21292 25832 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1400 21131 1452 21140
rect 1400 21097 1409 21131
rect 1409 21097 1443 21131
rect 1443 21097 1452 21131
rect 1400 21088 1452 21097
rect 1860 21131 1912 21140
rect 1860 21097 1869 21131
rect 1869 21097 1903 21131
rect 1903 21097 1912 21131
rect 1860 21088 1912 21097
rect 2044 21088 2096 21140
rect 2412 21131 2464 21140
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 3332 21088 3384 21140
rect 6184 21088 6236 21140
rect 6276 21088 6328 21140
rect 7380 21131 7432 21140
rect 7380 21097 7389 21131
rect 7389 21097 7423 21131
rect 7423 21097 7432 21131
rect 7932 21131 7984 21140
rect 7380 21088 7432 21097
rect 4068 21020 4120 21072
rect 6000 21063 6052 21072
rect 6000 21029 6009 21063
rect 6009 21029 6043 21063
rect 6043 21029 6052 21063
rect 6000 21020 6052 21029
rect 7472 21020 7524 21072
rect 7932 21097 7941 21131
rect 7941 21097 7975 21131
rect 7975 21097 7984 21131
rect 7932 21088 7984 21097
rect 9404 21088 9456 21140
rect 9956 21131 10008 21140
rect 9956 21097 9965 21131
rect 9965 21097 9999 21131
rect 9999 21097 10008 21131
rect 9956 21088 10008 21097
rect 10048 21088 10100 21140
rect 11244 21088 11296 21140
rect 11796 21088 11848 21140
rect 12072 21131 12124 21140
rect 7840 21020 7892 21072
rect 10968 21020 11020 21072
rect 12072 21097 12081 21131
rect 12081 21097 12115 21131
rect 12115 21097 12124 21131
rect 12072 21088 12124 21097
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13360 21088 13412 21097
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 15936 21088 15988 21140
rect 16396 21131 16448 21140
rect 16396 21097 16405 21131
rect 16405 21097 16439 21131
rect 16439 21097 16448 21131
rect 16396 21088 16448 21097
rect 17868 21088 17920 21140
rect 19248 21131 19300 21140
rect 2872 20927 2924 20936
rect 2872 20893 2881 20927
rect 2881 20893 2915 20927
rect 2915 20893 2924 20927
rect 2872 20884 2924 20893
rect 3608 20952 3660 21004
rect 4160 20952 4212 21004
rect 6920 20952 6972 21004
rect 8576 20952 8628 21004
rect 10876 20995 10928 21004
rect 10876 20961 10885 20995
rect 10885 20961 10919 20995
rect 10919 20961 10928 20995
rect 10876 20952 10928 20961
rect 3700 20884 3752 20936
rect 7840 20884 7892 20936
rect 9220 20884 9272 20936
rect 11704 20952 11756 21004
rect 1860 20816 1912 20868
rect 3056 20816 3108 20868
rect 2596 20748 2648 20800
rect 7288 20816 7340 20868
rect 8668 20859 8720 20868
rect 8668 20825 8677 20859
rect 8677 20825 8711 20859
rect 8711 20825 8720 20859
rect 8668 20816 8720 20825
rect 12072 20884 12124 20936
rect 14372 21020 14424 21072
rect 15752 21020 15804 21072
rect 16580 21020 16632 21072
rect 17040 21063 17092 21072
rect 17040 21029 17074 21063
rect 17074 21029 17092 21063
rect 17040 21020 17092 21029
rect 18696 21063 18748 21072
rect 18696 21029 18705 21063
rect 18705 21029 18739 21063
rect 18739 21029 18748 21063
rect 18696 21020 18748 21029
rect 19248 21097 19257 21131
rect 19257 21097 19291 21131
rect 19291 21097 19300 21131
rect 19248 21088 19300 21097
rect 21548 21088 21600 21140
rect 22008 21131 22060 21140
rect 22008 21097 22017 21131
rect 22017 21097 22051 21131
rect 22051 21097 22060 21131
rect 22008 21088 22060 21097
rect 22192 21088 22244 21140
rect 23664 21088 23716 21140
rect 19800 21020 19852 21072
rect 20352 21020 20404 21072
rect 21364 21063 21416 21072
rect 21364 21029 21373 21063
rect 21373 21029 21407 21063
rect 21407 21029 21416 21063
rect 21364 21020 21416 21029
rect 14832 20952 14884 21004
rect 16396 20952 16448 21004
rect 19248 20952 19300 21004
rect 23296 20952 23348 21004
rect 24676 20952 24728 21004
rect 16764 20927 16816 20936
rect 11152 20816 11204 20868
rect 13544 20816 13596 20868
rect 16764 20893 16773 20927
rect 16773 20893 16807 20927
rect 16807 20893 16816 20927
rect 16764 20884 16816 20893
rect 19340 20884 19392 20936
rect 15568 20816 15620 20868
rect 17776 20816 17828 20868
rect 19800 20927 19852 20936
rect 19800 20893 19809 20927
rect 19809 20893 19843 20927
rect 19843 20893 19852 20927
rect 19800 20884 19852 20893
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 22928 20859 22980 20868
rect 22928 20825 22937 20859
rect 22937 20825 22971 20859
rect 22971 20825 22980 20859
rect 22928 20816 22980 20825
rect 23940 20816 23992 20868
rect 24216 20816 24268 20868
rect 24860 20884 24912 20936
rect 5448 20791 5500 20800
rect 5448 20757 5457 20791
rect 5457 20757 5491 20791
rect 5491 20757 5500 20791
rect 5448 20748 5500 20757
rect 5540 20748 5592 20800
rect 6736 20791 6788 20800
rect 6736 20757 6745 20791
rect 6745 20757 6779 20791
rect 6779 20757 6788 20791
rect 6736 20748 6788 20757
rect 8300 20791 8352 20800
rect 8300 20757 8309 20791
rect 8309 20757 8343 20791
rect 8343 20757 8352 20791
rect 8300 20748 8352 20757
rect 11520 20791 11572 20800
rect 11520 20757 11529 20791
rect 11529 20757 11563 20791
rect 11563 20757 11572 20791
rect 11520 20748 11572 20757
rect 14556 20748 14608 20800
rect 21272 20748 21324 20800
rect 23848 20791 23900 20800
rect 23848 20757 23857 20791
rect 23857 20757 23891 20791
rect 23891 20757 23900 20791
rect 23848 20748 23900 20757
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 25320 20791 25372 20800
rect 25320 20757 25329 20791
rect 25329 20757 25363 20791
rect 25363 20757 25372 20791
rect 25320 20748 25372 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1400 20383 1452 20392
rect 1400 20349 1434 20383
rect 1434 20349 1452 20383
rect 2320 20544 2372 20596
rect 3148 20544 3200 20596
rect 3516 20544 3568 20596
rect 4528 20544 4580 20596
rect 5448 20544 5500 20596
rect 6276 20587 6328 20596
rect 6276 20553 6285 20587
rect 6285 20553 6319 20587
rect 6319 20553 6328 20587
rect 6276 20544 6328 20553
rect 6828 20587 6880 20596
rect 6828 20553 6837 20587
rect 6837 20553 6871 20587
rect 6871 20553 6880 20587
rect 6828 20544 6880 20553
rect 8116 20544 8168 20596
rect 10968 20544 11020 20596
rect 11704 20587 11756 20596
rect 11704 20553 11713 20587
rect 11713 20553 11747 20587
rect 11747 20553 11756 20587
rect 11704 20544 11756 20553
rect 14372 20587 14424 20596
rect 14372 20553 14381 20587
rect 14381 20553 14415 20587
rect 14415 20553 14424 20587
rect 14372 20544 14424 20553
rect 18328 20544 18380 20596
rect 19248 20544 19300 20596
rect 19524 20544 19576 20596
rect 20536 20587 20588 20596
rect 20536 20553 20545 20587
rect 20545 20553 20579 20587
rect 20579 20553 20588 20587
rect 20536 20544 20588 20553
rect 21364 20544 21416 20596
rect 22100 20544 22152 20596
rect 3976 20476 4028 20528
rect 1400 20340 1452 20349
rect 2780 20340 2832 20392
rect 4160 20408 4212 20460
rect 6736 20476 6788 20528
rect 7288 20451 7340 20460
rect 7288 20417 7297 20451
rect 7297 20417 7331 20451
rect 7331 20417 7340 20451
rect 7288 20408 7340 20417
rect 12164 20408 12216 20460
rect 3240 20383 3292 20392
rect 3240 20349 3249 20383
rect 3249 20349 3283 20383
rect 3283 20349 3292 20383
rect 3240 20340 3292 20349
rect 3516 20340 3568 20392
rect 3976 20340 4028 20392
rect 6828 20340 6880 20392
rect 8668 20340 8720 20392
rect 10876 20383 10928 20392
rect 10876 20349 10885 20383
rect 10885 20349 10919 20383
rect 10919 20349 10928 20383
rect 10876 20340 10928 20349
rect 3332 20315 3384 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 1860 20204 1912 20256
rect 3332 20281 3341 20315
rect 3341 20281 3375 20315
rect 3375 20281 3384 20315
rect 3332 20272 3384 20281
rect 3700 20272 3752 20324
rect 4252 20272 4304 20324
rect 6368 20272 6420 20324
rect 8760 20272 8812 20324
rect 12624 20272 12676 20324
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 3516 20204 3568 20256
rect 5172 20204 5224 20256
rect 5448 20247 5500 20256
rect 5448 20213 5457 20247
rect 5457 20213 5491 20247
rect 5491 20213 5500 20247
rect 5448 20204 5500 20213
rect 6828 20204 6880 20256
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 8576 20204 8628 20256
rect 11060 20247 11112 20256
rect 11060 20213 11069 20247
rect 11069 20213 11103 20247
rect 11103 20213 11112 20247
rect 11060 20204 11112 20213
rect 12072 20247 12124 20256
rect 12072 20213 12081 20247
rect 12081 20213 12115 20247
rect 12115 20213 12124 20247
rect 12072 20204 12124 20213
rect 13912 20204 13964 20256
rect 14832 20247 14884 20256
rect 14832 20213 14841 20247
rect 14841 20213 14875 20247
rect 14875 20213 14884 20247
rect 14832 20204 14884 20213
rect 14924 20204 14976 20256
rect 16764 20340 16816 20392
rect 17316 20383 17368 20392
rect 17316 20349 17325 20383
rect 17325 20349 17359 20383
rect 17359 20349 17368 20383
rect 17316 20340 17368 20349
rect 17960 20340 18012 20392
rect 19432 20408 19484 20460
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 20904 20340 20956 20392
rect 23296 20544 23348 20596
rect 23664 20544 23716 20596
rect 24032 20544 24084 20596
rect 25412 20587 25464 20596
rect 25412 20553 25421 20587
rect 25421 20553 25455 20587
rect 25455 20553 25464 20587
rect 25412 20544 25464 20553
rect 23848 20408 23900 20460
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 15752 20272 15804 20324
rect 25228 20383 25280 20392
rect 25228 20349 25237 20383
rect 25237 20349 25271 20383
rect 25271 20349 25280 20383
rect 25228 20340 25280 20349
rect 16764 20247 16816 20256
rect 16764 20213 16773 20247
rect 16773 20213 16807 20247
rect 16807 20213 16816 20247
rect 16764 20204 16816 20213
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 17776 20204 17828 20213
rect 18972 20247 19024 20256
rect 18972 20213 18981 20247
rect 18981 20213 19015 20247
rect 19015 20213 19024 20247
rect 21916 20272 21968 20324
rect 24768 20272 24820 20324
rect 18972 20204 19024 20213
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 23756 20204 23808 20256
rect 24676 20247 24728 20256
rect 24676 20213 24685 20247
rect 24685 20213 24719 20247
rect 24719 20213 24728 20247
rect 24676 20204 24728 20213
rect 25872 20204 25924 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2412 20043 2464 20052
rect 2412 20009 2421 20043
rect 2421 20009 2455 20043
rect 2455 20009 2464 20043
rect 2412 20000 2464 20009
rect 3056 20000 3108 20052
rect 4068 20043 4120 20052
rect 4068 20009 4077 20043
rect 4077 20009 4111 20043
rect 4111 20009 4120 20043
rect 4068 20000 4120 20009
rect 7196 20000 7248 20052
rect 8760 20000 8812 20052
rect 12624 20000 12676 20052
rect 13544 20043 13596 20052
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 13636 20043 13688 20052
rect 13636 20009 13645 20043
rect 13645 20009 13679 20043
rect 13679 20009 13688 20043
rect 14648 20043 14700 20052
rect 13636 20000 13688 20009
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 17040 20000 17092 20052
rect 17408 20043 17460 20052
rect 17408 20009 17417 20043
rect 17417 20009 17451 20043
rect 17451 20009 17460 20043
rect 17408 20000 17460 20009
rect 19432 20000 19484 20052
rect 21088 20043 21140 20052
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 21548 20043 21600 20052
rect 21548 20009 21557 20043
rect 21557 20009 21591 20043
rect 21591 20009 21600 20043
rect 21548 20000 21600 20009
rect 23388 20000 23440 20052
rect 2136 19932 2188 19984
rect 3332 19932 3384 19984
rect 4620 19932 4672 19984
rect 7840 19975 7892 19984
rect 7840 19941 7849 19975
rect 7849 19941 7883 19975
rect 7883 19941 7892 19975
rect 7840 19932 7892 19941
rect 9680 19932 9732 19984
rect 12072 19932 12124 19984
rect 2596 19864 2648 19916
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 4160 19864 4212 19916
rect 2872 19796 2924 19848
rect 4528 19839 4580 19848
rect 2412 19728 2464 19780
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 5448 19864 5500 19916
rect 6368 19864 6420 19916
rect 8852 19864 8904 19916
rect 9220 19864 9272 19916
rect 21456 19932 21508 19984
rect 25044 20000 25096 20052
rect 12164 19864 12216 19916
rect 13636 19864 13688 19916
rect 14004 19907 14056 19916
rect 14004 19873 14013 19907
rect 14013 19873 14047 19907
rect 14047 19873 14056 19907
rect 14004 19864 14056 19873
rect 8668 19796 8720 19848
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 11612 19839 11664 19848
rect 9680 19796 9732 19805
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 12624 19839 12676 19848
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 12624 19796 12676 19805
rect 13820 19796 13872 19848
rect 15292 19864 15344 19916
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 15476 19796 15528 19848
rect 15844 19864 15896 19916
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 18604 19907 18656 19916
rect 18604 19873 18638 19907
rect 18638 19873 18656 19907
rect 18604 19864 18656 19873
rect 20812 19864 20864 19916
rect 23020 19864 23072 19916
rect 23296 19864 23348 19916
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16764 19796 16816 19848
rect 6828 19728 6880 19780
rect 8760 19728 8812 19780
rect 19340 19796 19392 19848
rect 19984 19796 20036 19848
rect 20904 19728 20956 19780
rect 24308 19796 24360 19848
rect 25136 19839 25188 19848
rect 25136 19805 25145 19839
rect 25145 19805 25179 19839
rect 25179 19805 25188 19839
rect 25136 19796 25188 19805
rect 23664 19728 23716 19780
rect 1492 19660 1544 19712
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 2044 19660 2096 19712
rect 3700 19703 3752 19712
rect 3700 19669 3709 19703
rect 3709 19669 3743 19703
rect 3743 19669 3752 19703
rect 3700 19660 3752 19669
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 6736 19660 6788 19712
rect 7288 19660 7340 19712
rect 9312 19703 9364 19712
rect 9312 19669 9321 19703
rect 9321 19669 9355 19703
rect 9355 19669 9364 19703
rect 9312 19660 9364 19669
rect 13176 19703 13228 19712
rect 13176 19669 13185 19703
rect 13185 19669 13219 19703
rect 13219 19669 13228 19703
rect 13176 19660 13228 19669
rect 13452 19660 13504 19712
rect 14004 19660 14056 19712
rect 16396 19703 16448 19712
rect 16396 19669 16405 19703
rect 16405 19669 16439 19703
rect 16439 19669 16448 19703
rect 16396 19660 16448 19669
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 19984 19660 20036 19712
rect 21916 19703 21968 19712
rect 21916 19669 21925 19703
rect 21925 19669 21959 19703
rect 21959 19669 21968 19703
rect 21916 19660 21968 19669
rect 23296 19660 23348 19712
rect 24216 19660 24268 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 3056 19456 3108 19508
rect 5172 19499 5224 19508
rect 1124 19388 1176 19440
rect 3792 19388 3844 19440
rect 4068 19388 4120 19440
rect 5172 19465 5181 19499
rect 5181 19465 5215 19499
rect 5215 19465 5224 19499
rect 5172 19456 5224 19465
rect 6368 19456 6420 19508
rect 8668 19456 8720 19508
rect 9680 19456 9732 19508
rect 13636 19456 13688 19508
rect 7288 19388 7340 19440
rect 7840 19388 7892 19440
rect 9312 19388 9364 19440
rect 2044 19320 2096 19372
rect 3700 19320 3752 19372
rect 1860 19252 1912 19304
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 3884 19252 3936 19304
rect 5356 19320 5408 19372
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 9588 19320 9640 19372
rect 9864 19320 9916 19372
rect 5540 19295 5592 19304
rect 1676 19184 1728 19236
rect 2228 19227 2280 19236
rect 2228 19193 2237 19227
rect 2237 19193 2271 19227
rect 2271 19193 2280 19227
rect 2228 19184 2280 19193
rect 3792 19184 3844 19236
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 7288 19252 7340 19304
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 9220 19252 9272 19304
rect 9496 19252 9548 19304
rect 12348 19320 12400 19372
rect 11152 19252 11204 19304
rect 14832 19456 14884 19508
rect 15292 19456 15344 19508
rect 16764 19456 16816 19508
rect 17224 19499 17276 19508
rect 17224 19465 17233 19499
rect 17233 19465 17267 19499
rect 17267 19465 17276 19499
rect 17224 19456 17276 19465
rect 17316 19456 17368 19508
rect 13084 19252 13136 19304
rect 13452 19295 13504 19304
rect 13452 19261 13461 19295
rect 13461 19261 13495 19295
rect 13495 19261 13504 19295
rect 13452 19252 13504 19261
rect 14832 19295 14884 19304
rect 14832 19261 14866 19295
rect 14866 19261 14884 19295
rect 15936 19320 15988 19372
rect 25044 19456 25096 19508
rect 25136 19388 25188 19440
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 14832 19252 14884 19261
rect 20904 19295 20956 19304
rect 20904 19261 20913 19295
rect 20913 19261 20947 19295
rect 20947 19261 20956 19295
rect 20904 19252 20956 19261
rect 1952 19116 2004 19168
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 5080 19159 5132 19168
rect 5080 19125 5089 19159
rect 5089 19125 5123 19159
rect 5123 19125 5132 19159
rect 5080 19116 5132 19125
rect 7012 19116 7064 19168
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7288 19116 7340 19125
rect 8208 19116 8260 19168
rect 8852 19116 8904 19168
rect 12164 19184 12216 19236
rect 9404 19116 9456 19168
rect 10692 19116 10744 19168
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 13728 19184 13780 19236
rect 14280 19184 14332 19236
rect 13084 19116 13136 19168
rect 14556 19116 14608 19168
rect 18512 19184 18564 19236
rect 20444 19184 20496 19236
rect 21180 19227 21232 19236
rect 21180 19193 21214 19227
rect 21214 19193 21232 19227
rect 21180 19184 21232 19193
rect 18604 19116 18656 19168
rect 20812 19159 20864 19168
rect 20812 19125 20821 19159
rect 20821 19125 20855 19159
rect 20855 19125 20864 19159
rect 20812 19116 20864 19125
rect 23204 19184 23256 19236
rect 23020 19116 23072 19168
rect 25136 19252 25188 19304
rect 23848 19116 23900 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2136 18912 2188 18964
rect 2872 18955 2924 18964
rect 2872 18921 2881 18955
rect 2881 18921 2915 18955
rect 2915 18921 2924 18955
rect 2872 18912 2924 18921
rect 4620 18912 4672 18964
rect 5356 18912 5408 18964
rect 5540 18912 5592 18964
rect 6184 18912 6236 18964
rect 7012 18912 7064 18964
rect 7196 18912 7248 18964
rect 7840 18955 7892 18964
rect 7840 18921 7849 18955
rect 7849 18921 7883 18955
rect 7883 18921 7892 18955
rect 7840 18912 7892 18921
rect 11152 18912 11204 18964
rect 13360 18955 13412 18964
rect 13360 18921 13369 18955
rect 13369 18921 13403 18955
rect 13403 18921 13412 18955
rect 13360 18912 13412 18921
rect 14832 18912 14884 18964
rect 15016 18955 15068 18964
rect 15016 18921 15025 18955
rect 15025 18921 15059 18955
rect 15059 18921 15068 18955
rect 15016 18912 15068 18921
rect 17500 18955 17552 18964
rect 17500 18921 17509 18955
rect 17509 18921 17543 18955
rect 17543 18921 17552 18955
rect 17500 18912 17552 18921
rect 17776 18912 17828 18964
rect 18604 18955 18656 18964
rect 18604 18921 18613 18955
rect 18613 18921 18647 18955
rect 18647 18921 18656 18955
rect 18604 18912 18656 18921
rect 19248 18912 19300 18964
rect 21732 18912 21784 18964
rect 22008 18912 22060 18964
rect 24768 18955 24820 18964
rect 24768 18921 24777 18955
rect 24777 18921 24811 18955
rect 24811 18921 24820 18955
rect 24768 18912 24820 18921
rect 25228 18955 25280 18964
rect 25228 18921 25237 18955
rect 25237 18921 25271 18955
rect 25271 18921 25280 18955
rect 25228 18912 25280 18921
rect 3884 18844 3936 18896
rect 4344 18844 4396 18896
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 2688 18776 2740 18828
rect 2964 18776 3016 18828
rect 6184 18819 6236 18828
rect 6184 18785 6193 18819
rect 6193 18785 6227 18819
rect 6227 18785 6236 18819
rect 6184 18776 6236 18785
rect 6552 18776 6604 18828
rect 2044 18751 2096 18760
rect 2044 18717 2053 18751
rect 2053 18717 2087 18751
rect 2087 18717 2096 18751
rect 2044 18708 2096 18717
rect 4436 18708 4488 18760
rect 3240 18640 3292 18692
rect 5080 18640 5132 18692
rect 7104 18708 7156 18760
rect 7472 18844 7524 18896
rect 8760 18887 8812 18896
rect 8760 18853 8769 18887
rect 8769 18853 8803 18887
rect 8803 18853 8812 18887
rect 8760 18844 8812 18853
rect 9680 18844 9732 18896
rect 15292 18844 15344 18896
rect 10968 18776 11020 18828
rect 11152 18776 11204 18828
rect 13912 18776 13964 18828
rect 16304 18819 16356 18828
rect 16304 18785 16313 18819
rect 16313 18785 16347 18819
rect 16347 18785 16356 18819
rect 16304 18776 16356 18785
rect 9680 18708 9732 18760
rect 9864 18708 9916 18760
rect 11060 18708 11112 18760
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 16212 18708 16264 18760
rect 16580 18708 16632 18760
rect 19064 18776 19116 18828
rect 21364 18776 21416 18828
rect 21824 18776 21876 18828
rect 23756 18844 23808 18896
rect 8024 18640 8076 18692
rect 9496 18683 9548 18692
rect 9496 18649 9505 18683
rect 9505 18649 9539 18683
rect 9539 18649 9548 18683
rect 9496 18640 9548 18649
rect 18604 18708 18656 18760
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 21180 18751 21232 18760
rect 19432 18640 19484 18692
rect 21180 18717 21189 18751
rect 21189 18717 21223 18751
rect 21223 18717 21232 18751
rect 21180 18708 21232 18717
rect 21916 18708 21968 18760
rect 23296 18776 23348 18828
rect 23664 18751 23716 18760
rect 23664 18717 23673 18751
rect 23673 18717 23707 18751
rect 23707 18717 23716 18751
rect 23664 18708 23716 18717
rect 23848 18751 23900 18760
rect 23848 18717 23857 18751
rect 23857 18717 23891 18751
rect 23891 18717 23900 18751
rect 23848 18708 23900 18717
rect 24952 18776 25004 18828
rect 25780 18708 25832 18760
rect 21640 18683 21692 18692
rect 21640 18649 21649 18683
rect 21649 18649 21683 18683
rect 21683 18649 21692 18683
rect 21640 18640 21692 18649
rect 22744 18640 22796 18692
rect 23388 18640 23440 18692
rect 2136 18572 2188 18624
rect 7012 18572 7064 18624
rect 7288 18572 7340 18624
rect 8668 18572 8720 18624
rect 12072 18572 12124 18624
rect 13820 18615 13872 18624
rect 13820 18581 13829 18615
rect 13829 18581 13863 18615
rect 13863 18581 13872 18615
rect 13820 18572 13872 18581
rect 15476 18615 15528 18624
rect 15476 18581 15485 18615
rect 15485 18581 15519 18615
rect 15519 18581 15528 18615
rect 15476 18572 15528 18581
rect 18604 18572 18656 18624
rect 20168 18615 20220 18624
rect 20168 18581 20177 18615
rect 20177 18581 20211 18615
rect 20211 18581 20220 18615
rect 20168 18572 20220 18581
rect 22560 18572 22612 18624
rect 23848 18572 23900 18624
rect 24308 18640 24360 18692
rect 25136 18640 25188 18692
rect 24216 18615 24268 18624
rect 24216 18581 24225 18615
rect 24225 18581 24259 18615
rect 24259 18581 24268 18615
rect 24216 18572 24268 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 4068 18368 4120 18420
rect 5080 18368 5132 18420
rect 9588 18368 9640 18420
rect 12532 18368 12584 18420
rect 13636 18368 13688 18420
rect 17408 18411 17460 18420
rect 6552 18300 6604 18352
rect 12716 18300 12768 18352
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 1952 18096 2004 18148
rect 2136 18028 2188 18080
rect 2780 18028 2832 18080
rect 4160 18232 4212 18284
rect 6184 18232 6236 18284
rect 7840 18232 7892 18284
rect 8668 18232 8720 18284
rect 13728 18232 13780 18284
rect 17408 18377 17417 18411
rect 17417 18377 17451 18411
rect 17451 18377 17460 18411
rect 17408 18368 17460 18377
rect 17776 18368 17828 18420
rect 21732 18411 21784 18420
rect 21732 18377 21741 18411
rect 21741 18377 21775 18411
rect 21775 18377 21784 18411
rect 21732 18368 21784 18377
rect 23480 18411 23532 18420
rect 23480 18377 23489 18411
rect 23489 18377 23523 18411
rect 23523 18377 23532 18411
rect 23480 18368 23532 18377
rect 16672 18232 16724 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 20168 18232 20220 18284
rect 21824 18300 21876 18352
rect 3424 18207 3476 18216
rect 3424 18173 3447 18207
rect 3447 18173 3476 18207
rect 3424 18164 3476 18173
rect 6000 18164 6052 18216
rect 5816 18071 5868 18080
rect 5816 18037 5825 18071
rect 5825 18037 5859 18071
rect 5859 18037 5868 18071
rect 5816 18028 5868 18037
rect 7380 18164 7432 18216
rect 6920 18096 6972 18148
rect 6368 18028 6420 18080
rect 6644 18028 6696 18080
rect 8024 18028 8076 18080
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 8208 18028 8260 18037
rect 8576 18028 8628 18080
rect 9496 18164 9548 18216
rect 10140 18164 10192 18216
rect 9036 18096 9088 18148
rect 12716 18164 12768 18216
rect 14556 18207 14608 18216
rect 14556 18173 14590 18207
rect 14590 18173 14608 18207
rect 14556 18164 14608 18173
rect 15660 18164 15712 18216
rect 17408 18164 17460 18216
rect 21180 18232 21232 18284
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 22560 18275 22612 18284
rect 22560 18241 22569 18275
rect 22569 18241 22603 18275
rect 22603 18241 22612 18275
rect 22560 18232 22612 18241
rect 25228 18368 25280 18420
rect 25504 18368 25556 18420
rect 25780 18411 25832 18420
rect 25780 18377 25789 18411
rect 25789 18377 25823 18411
rect 25823 18377 25832 18411
rect 25780 18368 25832 18377
rect 26240 18411 26292 18420
rect 26240 18377 26249 18411
rect 26249 18377 26283 18411
rect 26283 18377 26292 18411
rect 26240 18368 26292 18377
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24216 18232 24268 18241
rect 20720 18164 20772 18216
rect 21640 18164 21692 18216
rect 23112 18164 23164 18216
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 10048 18028 10100 18080
rect 11520 18071 11572 18080
rect 11520 18037 11529 18071
rect 11529 18037 11563 18071
rect 11563 18037 11572 18071
rect 11520 18028 11572 18037
rect 15292 18096 15344 18148
rect 16212 18096 16264 18148
rect 18328 18096 18380 18148
rect 19064 18139 19116 18148
rect 19064 18105 19073 18139
rect 19073 18105 19107 18139
rect 19107 18105 19116 18139
rect 19064 18096 19116 18105
rect 20168 18096 20220 18148
rect 22928 18096 22980 18148
rect 23848 18096 23900 18148
rect 13912 18028 13964 18080
rect 16304 18071 16356 18080
rect 16304 18037 16313 18071
rect 16313 18037 16347 18071
rect 16347 18037 16356 18071
rect 16304 18028 16356 18037
rect 17316 18028 17368 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 20260 18028 20312 18080
rect 20444 18071 20496 18080
rect 20444 18037 20453 18071
rect 20453 18037 20487 18071
rect 20487 18037 20496 18071
rect 20444 18028 20496 18037
rect 21364 18028 21416 18080
rect 21640 18028 21692 18080
rect 22008 18028 22060 18080
rect 23664 18071 23716 18080
rect 23664 18037 23673 18071
rect 23673 18037 23707 18071
rect 23707 18037 23716 18071
rect 23664 18028 23716 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2044 17824 2096 17876
rect 2872 17824 2924 17876
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 4068 17824 4120 17876
rect 4344 17824 4396 17876
rect 6736 17867 6788 17876
rect 6736 17833 6745 17867
rect 6745 17833 6779 17867
rect 6779 17833 6788 17867
rect 6736 17824 6788 17833
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 8208 17824 8260 17876
rect 9312 17824 9364 17876
rect 10784 17867 10836 17876
rect 10784 17833 10793 17867
rect 10793 17833 10827 17867
rect 10827 17833 10836 17867
rect 10784 17824 10836 17833
rect 12440 17824 12492 17876
rect 14004 17824 14056 17876
rect 14556 17824 14608 17876
rect 16580 17824 16632 17876
rect 18604 17824 18656 17876
rect 19432 17824 19484 17876
rect 20076 17824 20128 17876
rect 22192 17824 22244 17876
rect 22376 17824 22428 17876
rect 23388 17824 23440 17876
rect 1492 17756 1544 17808
rect 7288 17756 7340 17808
rect 11060 17756 11112 17808
rect 12072 17756 12124 17808
rect 12164 17756 12216 17808
rect 14188 17756 14240 17808
rect 2228 17688 2280 17740
rect 5080 17731 5132 17740
rect 5080 17697 5114 17731
rect 5114 17697 5132 17731
rect 5080 17688 5132 17697
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 9128 17688 9180 17740
rect 11520 17688 11572 17740
rect 15660 17688 15712 17740
rect 16120 17688 16172 17740
rect 17040 17756 17092 17808
rect 21456 17756 21508 17808
rect 22468 17756 22520 17808
rect 18144 17688 18196 17740
rect 19432 17688 19484 17740
rect 19984 17688 20036 17740
rect 22560 17688 22612 17740
rect 23664 17688 23716 17740
rect 25320 17688 25372 17740
rect 1492 17663 1544 17672
rect 1492 17629 1501 17663
rect 1501 17629 1535 17663
rect 1535 17629 1544 17663
rect 1492 17620 1544 17629
rect 4804 17663 4856 17672
rect 4804 17629 4813 17663
rect 4813 17629 4847 17663
rect 4847 17629 4856 17663
rect 4804 17620 4856 17629
rect 6828 17620 6880 17672
rect 7748 17620 7800 17672
rect 10232 17620 10284 17672
rect 11336 17620 11388 17672
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 16580 17620 16632 17672
rect 20904 17663 20956 17672
rect 15752 17552 15804 17604
rect 16856 17552 16908 17604
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 22100 17620 22152 17672
rect 22928 17620 22980 17672
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 4436 17484 4488 17536
rect 6184 17527 6236 17536
rect 6184 17493 6193 17527
rect 6193 17493 6227 17527
rect 6227 17493 6236 17527
rect 6184 17484 6236 17493
rect 6920 17484 6972 17536
rect 8576 17484 8628 17536
rect 9404 17527 9456 17536
rect 9404 17493 9413 17527
rect 9413 17493 9447 17527
rect 9447 17493 9456 17527
rect 9404 17484 9456 17493
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 11152 17484 11204 17536
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 23204 17484 23256 17536
rect 24216 17484 24268 17536
rect 24952 17484 25004 17536
rect 25136 17527 25188 17536
rect 25136 17493 25145 17527
rect 25145 17493 25179 17527
rect 25179 17493 25188 17527
rect 25136 17484 25188 17493
rect 25228 17484 25280 17536
rect 25964 17484 26016 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1492 17280 1544 17332
rect 2780 17280 2832 17332
rect 3424 17323 3476 17332
rect 3424 17289 3433 17323
rect 3433 17289 3467 17323
rect 3467 17289 3476 17323
rect 3424 17280 3476 17289
rect 4712 17323 4764 17332
rect 4712 17289 4721 17323
rect 4721 17289 4755 17323
rect 4755 17289 4764 17323
rect 4712 17280 4764 17289
rect 5356 17280 5408 17332
rect 6276 17280 6328 17332
rect 6828 17280 6880 17332
rect 7012 17323 7064 17332
rect 7012 17289 7021 17323
rect 7021 17289 7055 17323
rect 7055 17289 7064 17323
rect 7012 17280 7064 17289
rect 7380 17323 7432 17332
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 11520 17280 11572 17332
rect 12072 17280 12124 17332
rect 13268 17280 13320 17332
rect 13544 17323 13596 17332
rect 13544 17289 13553 17323
rect 13553 17289 13587 17323
rect 13587 17289 13596 17323
rect 13544 17280 13596 17289
rect 16488 17280 16540 17332
rect 16856 17280 16908 17332
rect 4252 17212 4304 17264
rect 4804 17212 4856 17264
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 11428 17187 11480 17196
rect 5448 17144 5500 17153
rect 11428 17153 11437 17187
rect 11437 17153 11471 17187
rect 11471 17153 11480 17187
rect 11428 17144 11480 17153
rect 15384 17144 15436 17196
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 17684 17144 17736 17196
rect 21364 17280 21416 17332
rect 22468 17323 22520 17332
rect 22468 17289 22477 17323
rect 22477 17289 22511 17323
rect 22511 17289 22520 17323
rect 22468 17280 22520 17289
rect 20904 17255 20956 17264
rect 20904 17221 20913 17255
rect 20913 17221 20947 17255
rect 20947 17221 20956 17255
rect 20904 17212 20956 17221
rect 2872 17076 2924 17128
rect 4344 17076 4396 17128
rect 7380 17076 7432 17128
rect 7564 17076 7616 17128
rect 8576 17076 8628 17128
rect 9404 17076 9456 17128
rect 9956 17076 10008 17128
rect 3148 17008 3200 17060
rect 5080 17008 5132 17060
rect 5172 17008 5224 17060
rect 7288 17008 7340 17060
rect 7840 17008 7892 17060
rect 10048 17008 10100 17060
rect 10232 17008 10284 17060
rect 10784 17076 10836 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 14004 17119 14056 17128
rect 14004 17085 14038 17119
rect 14038 17085 14056 17119
rect 14004 17076 14056 17085
rect 16488 17076 16540 17128
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 18696 17076 18748 17128
rect 12808 17008 12860 17060
rect 15660 17051 15712 17060
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 5540 16940 5592 16992
rect 8576 16940 8628 16992
rect 9680 16940 9732 16992
rect 15660 17017 15669 17051
rect 15669 17017 15703 17051
rect 15703 17017 15712 17051
rect 15660 17008 15712 17017
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 12900 16940 12952 16992
rect 14556 16940 14608 16992
rect 15936 16940 15988 16992
rect 16120 16983 16172 16992
rect 16120 16949 16129 16983
rect 16129 16949 16163 16983
rect 16163 16949 16172 16983
rect 16120 16940 16172 16949
rect 21364 17119 21416 17128
rect 21364 17085 21398 17119
rect 21398 17085 21416 17119
rect 21364 17076 21416 17085
rect 24216 17008 24268 17060
rect 22100 16940 22152 16992
rect 23020 16940 23072 16992
rect 25044 16983 25096 16992
rect 25044 16949 25053 16983
rect 25053 16949 25087 16983
rect 25087 16949 25096 16983
rect 25044 16940 25096 16949
rect 25320 16940 25372 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1584 16736 1636 16788
rect 2044 16736 2096 16788
rect 2872 16736 2924 16788
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 4344 16736 4396 16788
rect 5080 16736 5132 16788
rect 5264 16736 5316 16788
rect 7656 16736 7708 16788
rect 7932 16779 7984 16788
rect 7932 16745 7941 16779
rect 7941 16745 7975 16779
rect 7975 16745 7984 16779
rect 7932 16736 7984 16745
rect 8300 16779 8352 16788
rect 8300 16745 8309 16779
rect 8309 16745 8343 16779
rect 8343 16745 8352 16779
rect 8300 16736 8352 16745
rect 11428 16736 11480 16788
rect 15384 16736 15436 16788
rect 17684 16779 17736 16788
rect 17684 16745 17693 16779
rect 17693 16745 17727 16779
rect 17727 16745 17736 16779
rect 17684 16736 17736 16745
rect 18696 16779 18748 16788
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 19156 16779 19208 16788
rect 1216 16668 1268 16720
rect 4528 16668 4580 16720
rect 5448 16668 5500 16720
rect 7840 16711 7892 16720
rect 7840 16677 7849 16711
rect 7849 16677 7883 16711
rect 7883 16677 7892 16711
rect 7840 16668 7892 16677
rect 2596 16600 2648 16652
rect 3884 16643 3936 16652
rect 3884 16609 3893 16643
rect 3893 16609 3927 16643
rect 3927 16609 3936 16643
rect 3884 16600 3936 16609
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 6184 16600 6236 16652
rect 2688 16532 2740 16584
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 3148 16532 3200 16584
rect 4804 16532 4856 16584
rect 5356 16532 5408 16584
rect 7656 16600 7708 16652
rect 9036 16600 9088 16652
rect 9128 16600 9180 16652
rect 10876 16668 10928 16720
rect 19156 16745 19165 16779
rect 19165 16745 19199 16779
rect 19199 16745 19208 16779
rect 19156 16736 19208 16745
rect 20720 16736 20772 16788
rect 21272 16779 21324 16788
rect 21272 16745 21281 16779
rect 21281 16745 21315 16779
rect 21315 16745 21324 16779
rect 21272 16736 21324 16745
rect 22560 16779 22612 16788
rect 22560 16745 22569 16779
rect 22569 16745 22603 16779
rect 22603 16745 22612 16779
rect 22560 16736 22612 16745
rect 22928 16779 22980 16788
rect 22928 16745 22937 16779
rect 22937 16745 22971 16779
rect 22971 16745 22980 16779
rect 22928 16736 22980 16745
rect 24400 16779 24452 16788
rect 24400 16745 24409 16779
rect 24409 16745 24443 16779
rect 24443 16745 24452 16779
rect 24400 16736 24452 16745
rect 20812 16668 20864 16720
rect 23296 16711 23348 16720
rect 23296 16677 23330 16711
rect 23330 16677 23348 16711
rect 23296 16668 23348 16677
rect 7104 16532 7156 16584
rect 8576 16575 8628 16584
rect 296 16464 348 16516
rect 1400 16396 1452 16448
rect 2228 16439 2280 16448
rect 2228 16405 2237 16439
rect 2237 16405 2271 16439
rect 2271 16405 2280 16439
rect 2228 16396 2280 16405
rect 2412 16439 2464 16448
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 8300 16464 8352 16516
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 9496 16532 9548 16584
rect 9864 16600 9916 16652
rect 11060 16600 11112 16652
rect 11336 16600 11388 16652
rect 11704 16643 11756 16652
rect 11704 16609 11738 16643
rect 11738 16609 11756 16643
rect 11704 16600 11756 16609
rect 13820 16600 13872 16652
rect 15660 16600 15712 16652
rect 15752 16600 15804 16652
rect 16580 16643 16632 16652
rect 16580 16609 16614 16643
rect 16614 16609 16632 16643
rect 16580 16600 16632 16609
rect 19248 16643 19300 16652
rect 19248 16609 19257 16643
rect 19257 16609 19291 16643
rect 19291 16609 19300 16643
rect 19248 16600 19300 16609
rect 21272 16600 21324 16652
rect 10232 16532 10284 16584
rect 10968 16532 11020 16584
rect 11428 16575 11480 16584
rect 11428 16541 11437 16575
rect 11437 16541 11471 16575
rect 11471 16541 11480 16575
rect 11428 16532 11480 16541
rect 21456 16575 21508 16584
rect 19156 16464 19208 16516
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 21364 16464 21416 16516
rect 22008 16464 22060 16516
rect 7288 16396 7340 16448
rect 12072 16396 12124 16448
rect 14004 16396 14056 16448
rect 14372 16439 14424 16448
rect 14372 16405 14381 16439
rect 14381 16405 14415 16439
rect 14415 16405 14424 16439
rect 14372 16396 14424 16405
rect 16580 16396 16632 16448
rect 17040 16396 17092 16448
rect 18604 16396 18656 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2044 16192 2096 16244
rect 5356 16192 5408 16244
rect 6000 16192 6052 16244
rect 5448 16056 5500 16108
rect 7564 16192 7616 16244
rect 8392 16192 8444 16244
rect 10232 16192 10284 16244
rect 12440 16235 12492 16244
rect 12440 16201 12449 16235
rect 12449 16201 12483 16235
rect 12483 16201 12492 16235
rect 13912 16235 13964 16244
rect 12440 16192 12492 16201
rect 13912 16201 13921 16235
rect 13921 16201 13955 16235
rect 13955 16201 13964 16235
rect 13912 16192 13964 16201
rect 14096 16192 14148 16244
rect 15752 16192 15804 16244
rect 16488 16192 16540 16244
rect 19156 16235 19208 16244
rect 19156 16201 19165 16235
rect 19165 16201 19199 16235
rect 19199 16201 19208 16235
rect 19156 16192 19208 16201
rect 20444 16192 20496 16244
rect 21180 16192 21232 16244
rect 21916 16192 21968 16244
rect 22100 16192 22152 16244
rect 23020 16235 23072 16244
rect 23020 16201 23029 16235
rect 23029 16201 23063 16235
rect 23063 16201 23072 16235
rect 23020 16192 23072 16201
rect 3240 15988 3292 16040
rect 7380 15988 7432 16040
rect 12808 16056 12860 16108
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 23296 16124 23348 16176
rect 21456 16056 21508 16108
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 11428 15988 11480 16040
rect 14188 15988 14240 16040
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 20996 15988 21048 16040
rect 21916 16031 21968 16040
rect 2044 15963 2096 15972
rect 2044 15929 2053 15963
rect 2053 15929 2087 15963
rect 2087 15929 2096 15963
rect 2044 15920 2096 15929
rect 3516 15920 3568 15972
rect 7104 15963 7156 15972
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 3976 15895 4028 15904
rect 3976 15861 3985 15895
rect 3985 15861 4019 15895
rect 4019 15861 4028 15895
rect 3976 15852 4028 15861
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 7104 15929 7138 15963
rect 7138 15929 7156 15963
rect 7104 15920 7156 15929
rect 10968 15920 11020 15972
rect 13728 15920 13780 15972
rect 20536 15920 20588 15972
rect 21916 15997 21925 16031
rect 21925 15997 21959 16031
rect 21959 15997 21968 16031
rect 21916 15988 21968 15997
rect 23572 15988 23624 16040
rect 7196 15852 7248 15904
rect 7472 15852 7524 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 13360 15852 13412 15904
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 15476 15895 15528 15904
rect 14464 15852 14516 15861
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 18052 15895 18104 15904
rect 18052 15861 18061 15895
rect 18061 15861 18095 15895
rect 18095 15861 18104 15895
rect 18052 15852 18104 15861
rect 20996 15895 21048 15904
rect 20996 15861 21005 15895
rect 21005 15861 21039 15895
rect 21039 15861 21048 15895
rect 20996 15852 21048 15861
rect 23112 15920 23164 15972
rect 24216 15852 24268 15904
rect 25228 15852 25280 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1676 15648 1728 15700
rect 2504 15648 2556 15700
rect 2780 15648 2832 15700
rect 2872 15648 2924 15700
rect 5172 15648 5224 15700
rect 5448 15648 5500 15700
rect 6092 15648 6144 15700
rect 8576 15648 8628 15700
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 9496 15691 9548 15700
rect 9496 15657 9505 15691
rect 9505 15657 9539 15691
rect 9539 15657 9548 15691
rect 9496 15648 9548 15657
rect 10784 15648 10836 15700
rect 10968 15691 11020 15700
rect 10968 15657 10977 15691
rect 10977 15657 11011 15691
rect 11011 15657 11020 15691
rect 10968 15648 11020 15657
rect 11704 15648 11756 15700
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 14832 15648 14884 15700
rect 16028 15648 16080 15700
rect 17040 15648 17092 15700
rect 19156 15691 19208 15700
rect 19156 15657 19165 15691
rect 19165 15657 19199 15691
rect 19199 15657 19208 15691
rect 19156 15648 19208 15657
rect 20352 15648 20404 15700
rect 20812 15648 20864 15700
rect 21456 15648 21508 15700
rect 23112 15648 23164 15700
rect 2596 15580 2648 15632
rect 3148 15623 3200 15632
rect 3148 15589 3157 15623
rect 3157 15589 3191 15623
rect 3191 15589 3200 15623
rect 3148 15580 3200 15589
rect 4804 15623 4856 15632
rect 4804 15589 4813 15623
rect 4813 15589 4847 15623
rect 4847 15589 4856 15623
rect 4804 15580 4856 15589
rect 1400 15512 1452 15564
rect 3516 15555 3568 15564
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 3516 15521 3525 15555
rect 3525 15521 3559 15555
rect 3559 15521 3568 15555
rect 3516 15512 3568 15521
rect 4712 15555 4764 15564
rect 4712 15521 4721 15555
rect 4721 15521 4755 15555
rect 4755 15521 4764 15555
rect 4712 15512 4764 15521
rect 5080 15512 5132 15564
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 3976 15376 4028 15428
rect 4344 15419 4396 15428
rect 4344 15385 4353 15419
rect 4353 15385 4387 15419
rect 4387 15385 4396 15419
rect 4344 15376 4396 15385
rect 1400 15308 1452 15360
rect 4160 15308 4212 15360
rect 6276 15580 6328 15632
rect 6368 15580 6420 15632
rect 9588 15580 9640 15632
rect 10876 15580 10928 15632
rect 6000 15512 6052 15564
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 8668 15512 8720 15564
rect 10968 15512 11020 15564
rect 11428 15555 11480 15564
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 11520 15512 11572 15564
rect 12072 15512 12124 15564
rect 13912 15555 13964 15564
rect 13912 15521 13921 15555
rect 13921 15521 13955 15555
rect 13955 15521 13964 15555
rect 13912 15512 13964 15521
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 15752 15512 15804 15564
rect 16764 15555 16816 15564
rect 16764 15521 16798 15555
rect 16798 15521 16816 15555
rect 16764 15512 16816 15521
rect 19248 15512 19300 15564
rect 19340 15512 19392 15564
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 10140 15444 10192 15496
rect 9036 15376 9088 15428
rect 9956 15376 10008 15428
rect 15384 15444 15436 15496
rect 21640 15512 21692 15564
rect 24124 15580 24176 15632
rect 22100 15512 22152 15564
rect 23848 15512 23900 15564
rect 24768 15512 24820 15564
rect 21548 15487 21600 15496
rect 13820 15376 13872 15428
rect 14464 15376 14516 15428
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 23664 15444 23716 15496
rect 24032 15444 24084 15496
rect 25228 15444 25280 15496
rect 20628 15376 20680 15428
rect 23020 15376 23072 15428
rect 23480 15376 23532 15428
rect 24216 15376 24268 15428
rect 7012 15308 7064 15360
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 20076 15308 20128 15360
rect 24032 15351 24084 15360
rect 24032 15317 24041 15351
rect 24041 15317 24075 15351
rect 24075 15317 24084 15351
rect 24032 15308 24084 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 2504 15104 2556 15156
rect 4160 15104 4212 15156
rect 4344 15104 4396 15156
rect 4804 15104 4856 15156
rect 6276 15104 6328 15156
rect 10140 15104 10192 15156
rect 10784 15147 10836 15156
rect 10784 15113 10793 15147
rect 10793 15113 10827 15147
rect 10827 15113 10836 15147
rect 10784 15104 10836 15113
rect 11428 15104 11480 15156
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 1860 15036 1912 15088
rect 4712 15079 4764 15088
rect 4712 15045 4721 15079
rect 4721 15045 4755 15079
rect 4755 15045 4764 15079
rect 4712 15036 4764 15045
rect 11336 15036 11388 15088
rect 3976 14968 4028 15020
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 6368 14968 6420 15020
rect 11520 14968 11572 15020
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 13544 14968 13596 15020
rect 15384 15104 15436 15156
rect 16212 15104 16264 15156
rect 16764 15104 16816 15156
rect 18052 15104 18104 15156
rect 21640 15104 21692 15156
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 23848 15147 23900 15156
rect 23848 15113 23857 15147
rect 23857 15113 23891 15147
rect 23891 15113 23900 15147
rect 23848 15104 23900 15113
rect 24676 15104 24728 15156
rect 17592 15036 17644 15088
rect 23388 15036 23440 15088
rect 24124 15036 24176 15088
rect 25228 15079 25280 15088
rect 25228 15045 25237 15079
rect 25237 15045 25271 15079
rect 25271 15045 25280 15079
rect 25228 15036 25280 15045
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 4712 14900 4764 14952
rect 5172 14900 5224 14952
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 13452 14900 13504 14952
rect 16672 14900 16724 14952
rect 18052 14900 18104 14952
rect 22468 14943 22520 14952
rect 3884 14832 3936 14884
rect 7104 14832 7156 14884
rect 10600 14875 10652 14884
rect 10600 14841 10609 14875
rect 10609 14841 10643 14875
rect 10643 14841 10652 14875
rect 10600 14832 10652 14841
rect 3700 14764 3752 14816
rect 5080 14764 5132 14816
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 5632 14764 5684 14773
rect 7748 14764 7800 14816
rect 9220 14764 9272 14816
rect 10140 14764 10192 14816
rect 11428 14764 11480 14816
rect 12624 14764 12676 14816
rect 14188 14832 14240 14884
rect 14832 14832 14884 14884
rect 20076 14832 20128 14884
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 16396 14764 16448 14816
rect 18420 14764 18472 14816
rect 18696 14764 18748 14816
rect 19340 14807 19392 14816
rect 19340 14773 19349 14807
rect 19349 14773 19383 14807
rect 19383 14773 19392 14807
rect 19340 14764 19392 14773
rect 20904 14764 20956 14816
rect 21548 14807 21600 14816
rect 21548 14773 21557 14807
rect 21557 14773 21591 14807
rect 21591 14773 21600 14807
rect 21548 14764 21600 14773
rect 24216 14807 24268 14816
rect 24216 14773 24225 14807
rect 24225 14773 24259 14807
rect 24259 14773 24268 14807
rect 24216 14764 24268 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2596 14560 2648 14612
rect 3976 14560 4028 14612
rect 4068 14560 4120 14612
rect 5632 14560 5684 14612
rect 6920 14560 6972 14612
rect 9588 14560 9640 14612
rect 11520 14560 11572 14612
rect 13268 14560 13320 14612
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 13820 14560 13872 14612
rect 17592 14603 17644 14612
rect 17592 14569 17601 14603
rect 17601 14569 17635 14603
rect 17635 14569 17644 14603
rect 17592 14560 17644 14569
rect 18696 14603 18748 14612
rect 18696 14569 18705 14603
rect 18705 14569 18739 14603
rect 18739 14569 18748 14603
rect 18696 14560 18748 14569
rect 19248 14560 19300 14612
rect 20536 14603 20588 14612
rect 1492 14492 1544 14544
rect 1860 14492 1912 14544
rect 5816 14492 5868 14544
rect 7012 14492 7064 14544
rect 11796 14492 11848 14544
rect 18328 14492 18380 14544
rect 20536 14569 20545 14603
rect 20545 14569 20579 14603
rect 20579 14569 20588 14603
rect 20536 14560 20588 14569
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 24768 14560 24820 14612
rect 25596 14603 25648 14612
rect 25596 14569 25605 14603
rect 25605 14569 25639 14603
rect 25639 14569 25648 14603
rect 25596 14560 25648 14569
rect 20628 14492 20680 14544
rect 23664 14492 23716 14544
rect 3148 14424 3200 14476
rect 4620 14424 4672 14476
rect 5080 14424 5132 14476
rect 5448 14424 5500 14476
rect 6368 14467 6420 14476
rect 6368 14433 6377 14467
rect 6377 14433 6411 14467
rect 6411 14433 6420 14467
rect 6368 14424 6420 14433
rect 8668 14424 8720 14476
rect 11244 14424 11296 14476
rect 12072 14424 12124 14476
rect 12992 14424 13044 14476
rect 13452 14424 13504 14476
rect 15384 14424 15436 14476
rect 16212 14467 16264 14476
rect 16212 14433 16221 14467
rect 16221 14433 16255 14467
rect 16255 14433 16264 14467
rect 16212 14424 16264 14433
rect 16304 14424 16356 14476
rect 21180 14467 21232 14476
rect 21180 14433 21214 14467
rect 21214 14433 21232 14467
rect 21180 14424 21232 14433
rect 23848 14424 23900 14476
rect 24676 14424 24728 14476
rect 25136 14424 25188 14476
rect 2872 14356 2924 14408
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 9496 14356 9548 14408
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 19156 14399 19208 14408
rect 14188 14356 14240 14365
rect 19156 14365 19165 14399
rect 19165 14365 19199 14399
rect 19199 14365 19208 14399
rect 19156 14356 19208 14365
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 24124 14356 24176 14408
rect 3240 14288 3292 14340
rect 7748 14331 7800 14340
rect 7748 14297 7757 14331
rect 7757 14297 7791 14331
rect 7791 14297 7800 14331
rect 7748 14288 7800 14297
rect 12348 14331 12400 14340
rect 12348 14297 12357 14331
rect 12357 14297 12391 14331
rect 12391 14297 12400 14331
rect 12348 14288 12400 14297
rect 1400 14220 1452 14272
rect 2688 14220 2740 14272
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 9588 14220 9640 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 12624 14220 12676 14272
rect 14464 14220 14516 14272
rect 14832 14220 14884 14272
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 18788 14220 18840 14272
rect 23296 14220 23348 14272
rect 23756 14263 23808 14272
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1584 14059 1636 14068
rect 1584 14025 1593 14059
rect 1593 14025 1627 14059
rect 1627 14025 1636 14059
rect 1584 14016 1636 14025
rect 1860 14016 1912 14068
rect 2228 14016 2280 14068
rect 3424 14016 3476 14068
rect 3792 14016 3844 14068
rect 6368 14059 6420 14068
rect 2872 13948 2924 14000
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7380 14016 7432 14068
rect 5172 13991 5224 14000
rect 5172 13957 5181 13991
rect 5181 13957 5215 13991
rect 5215 13957 5224 13991
rect 5172 13948 5224 13957
rect 9496 14016 9548 14068
rect 11244 14016 11296 14068
rect 12164 14016 12216 14068
rect 14096 14016 14148 14068
rect 16304 14016 16356 14068
rect 18604 14016 18656 14068
rect 19248 14016 19300 14068
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 23296 14016 23348 14068
rect 24860 14016 24912 14068
rect 8208 13948 8260 14000
rect 13452 13948 13504 14000
rect 14464 13948 14516 14000
rect 16212 13948 16264 14000
rect 16764 13948 16816 14000
rect 1676 13880 1728 13932
rect 2228 13880 2280 13932
rect 3884 13880 3936 13932
rect 4988 13880 5040 13932
rect 5816 13923 5868 13932
rect 5816 13889 5825 13923
rect 5825 13889 5859 13923
rect 5859 13889 5868 13923
rect 5816 13880 5868 13889
rect 6276 13880 6328 13932
rect 8116 13880 8168 13932
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 8760 13880 8812 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3608 13812 3660 13864
rect 3516 13744 3568 13796
rect 3608 13719 3660 13728
rect 3608 13685 3617 13719
rect 3617 13685 3651 13719
rect 3651 13685 3660 13719
rect 3608 13676 3660 13685
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 9496 13812 9548 13864
rect 16028 13880 16080 13932
rect 10140 13812 10192 13864
rect 11060 13812 11112 13864
rect 13452 13855 13504 13864
rect 13452 13821 13461 13855
rect 13461 13821 13495 13855
rect 13495 13821 13504 13855
rect 13452 13812 13504 13821
rect 15384 13855 15436 13864
rect 15384 13821 15393 13855
rect 15393 13821 15427 13855
rect 15427 13821 15436 13855
rect 15384 13812 15436 13821
rect 18328 13948 18380 14000
rect 20076 13948 20128 14000
rect 24124 13948 24176 14000
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 23388 13880 23440 13932
rect 23756 13880 23808 13932
rect 25136 13880 25188 13932
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 18696 13812 18748 13864
rect 6920 13676 6972 13728
rect 7380 13676 7432 13728
rect 11152 13744 11204 13796
rect 13820 13744 13872 13796
rect 18788 13744 18840 13796
rect 19248 13744 19300 13796
rect 19524 13744 19576 13796
rect 21272 13812 21324 13864
rect 22468 13812 22520 13864
rect 23664 13812 23716 13864
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 25228 13855 25280 13864
rect 25228 13821 25237 13855
rect 25237 13821 25271 13855
rect 25271 13821 25280 13855
rect 25228 13812 25280 13821
rect 21548 13744 21600 13796
rect 22100 13744 22152 13796
rect 10968 13719 11020 13728
rect 10968 13685 10977 13719
rect 10977 13685 11011 13719
rect 11011 13685 11020 13719
rect 10968 13676 11020 13685
rect 12256 13719 12308 13728
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 12532 13676 12584 13728
rect 15936 13719 15988 13728
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 16304 13719 16356 13728
rect 16304 13685 16313 13719
rect 16313 13685 16347 13719
rect 16347 13685 16356 13719
rect 16304 13676 16356 13685
rect 20904 13676 20956 13728
rect 21272 13676 21324 13728
rect 22008 13676 22060 13728
rect 23296 13744 23348 13796
rect 24676 13719 24728 13728
rect 24676 13685 24685 13719
rect 24685 13685 24719 13719
rect 24719 13685 24728 13719
rect 24676 13676 24728 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 1768 13472 1820 13524
rect 2136 13472 2188 13524
rect 2780 13472 2832 13524
rect 3516 13472 3568 13524
rect 3976 13472 4028 13524
rect 4896 13515 4948 13524
rect 4896 13481 4905 13515
rect 4905 13481 4939 13515
rect 4939 13481 4948 13515
rect 4896 13472 4948 13481
rect 5356 13472 5408 13524
rect 5540 13472 5592 13524
rect 6460 13515 6512 13524
rect 6460 13481 6469 13515
rect 6469 13481 6503 13515
rect 6503 13481 6512 13515
rect 6460 13472 6512 13481
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 8116 13472 8168 13524
rect 8484 13472 8536 13524
rect 9036 13472 9088 13524
rect 9404 13515 9456 13524
rect 9404 13481 9413 13515
rect 9413 13481 9447 13515
rect 9447 13481 9456 13515
rect 9404 13472 9456 13481
rect 10692 13472 10744 13524
rect 11060 13472 11112 13524
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 14188 13472 14240 13524
rect 18604 13472 18656 13524
rect 19156 13515 19208 13524
rect 19156 13481 19165 13515
rect 19165 13481 19199 13515
rect 19199 13481 19208 13515
rect 19156 13472 19208 13481
rect 21180 13515 21232 13524
rect 21180 13481 21189 13515
rect 21189 13481 21223 13515
rect 21223 13481 21232 13515
rect 21180 13472 21232 13481
rect 23388 13472 23440 13524
rect 24032 13472 24084 13524
rect 5816 13447 5868 13456
rect 5816 13413 5825 13447
rect 5825 13413 5859 13447
rect 5859 13413 5868 13447
rect 5816 13404 5868 13413
rect 16396 13404 16448 13456
rect 19708 13447 19760 13456
rect 19708 13413 19717 13447
rect 19717 13413 19751 13447
rect 19751 13413 19760 13447
rect 19708 13404 19760 13413
rect 2136 13336 2188 13388
rect 2780 13336 2832 13388
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 6920 13336 6972 13388
rect 8116 13336 8168 13388
rect 8300 13336 8352 13388
rect 10968 13336 11020 13388
rect 12716 13379 12768 13388
rect 12716 13345 12750 13379
rect 12750 13345 12768 13379
rect 15752 13379 15804 13388
rect 12716 13336 12768 13345
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 20628 13336 20680 13388
rect 22008 13336 22060 13388
rect 5264 13268 5316 13320
rect 6552 13268 6604 13320
rect 7012 13268 7064 13320
rect 8760 13268 8812 13320
rect 9404 13268 9456 13320
rect 9956 13311 10008 13320
rect 9956 13277 9965 13311
rect 9965 13277 9999 13311
rect 9999 13277 10008 13311
rect 9956 13268 10008 13277
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 20444 13268 20496 13320
rect 21272 13311 21324 13320
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 7196 13200 7248 13252
rect 18788 13200 18840 13252
rect 23204 13404 23256 13456
rect 25044 13404 25096 13456
rect 23572 13336 23624 13388
rect 24032 13336 24084 13388
rect 25228 13336 25280 13388
rect 25872 13200 25924 13252
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 11336 13175 11388 13184
rect 11336 13141 11345 13175
rect 11345 13141 11379 13175
rect 11379 13141 11388 13175
rect 11336 13132 11388 13141
rect 12072 13132 12124 13184
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 19156 13132 19208 13184
rect 20260 13175 20312 13184
rect 20260 13141 20269 13175
rect 20269 13141 20303 13175
rect 20303 13141 20312 13175
rect 20260 13132 20312 13141
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 25504 13175 25556 13184
rect 25504 13141 25513 13175
rect 25513 13141 25547 13175
rect 25547 13141 25556 13175
rect 25504 13132 25556 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1492 12928 1544 12980
rect 3608 12928 3660 12980
rect 4804 12928 4856 12980
rect 6276 12971 6328 12980
rect 6276 12937 6285 12971
rect 6285 12937 6319 12971
rect 6319 12937 6328 12971
rect 6276 12928 6328 12937
rect 6368 12928 6420 12980
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 8300 12928 8352 12980
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 8852 12928 8904 12980
rect 9956 12928 10008 12980
rect 10692 12928 10744 12980
rect 10968 12928 11020 12980
rect 12440 12928 12492 12980
rect 12992 12971 13044 12980
rect 12992 12937 13001 12971
rect 13001 12937 13035 12971
rect 13035 12937 13044 12971
rect 12992 12928 13044 12937
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 2688 12903 2740 12912
rect 2688 12869 2697 12903
rect 2697 12869 2731 12903
rect 2731 12869 2740 12903
rect 2688 12860 2740 12869
rect 2780 12860 2832 12912
rect 4344 12860 4396 12912
rect 4988 12903 5040 12912
rect 4988 12869 4997 12903
rect 4997 12869 5031 12903
rect 5031 12869 5040 12903
rect 4988 12860 5040 12869
rect 6092 12792 6144 12844
rect 6184 12792 6236 12844
rect 2044 12699 2096 12708
rect 2044 12665 2053 12699
rect 2053 12665 2087 12699
rect 2087 12665 2096 12699
rect 2044 12656 2096 12665
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 5264 12724 5316 12776
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 6644 12724 6696 12776
rect 6920 12792 6972 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 14832 12860 14884 12912
rect 16212 12928 16264 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 16764 12971 16816 12980
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 17868 12928 17920 12980
rect 18052 12971 18104 12980
rect 18052 12937 18061 12971
rect 18061 12937 18095 12971
rect 18095 12937 18104 12971
rect 18052 12928 18104 12937
rect 19708 12928 19760 12980
rect 20168 12928 20220 12980
rect 20628 12971 20680 12980
rect 20628 12937 20637 12971
rect 20637 12937 20671 12971
rect 20671 12937 20680 12971
rect 20628 12928 20680 12937
rect 20904 12928 20956 12980
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 9404 12792 9456 12844
rect 13728 12792 13780 12844
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 20352 12860 20404 12912
rect 22100 12860 22152 12912
rect 8116 12724 8168 12776
rect 9956 12724 10008 12776
rect 13452 12767 13504 12776
rect 13452 12733 13461 12767
rect 13461 12733 13495 12767
rect 13495 12733 13504 12767
rect 14004 12767 14056 12776
rect 13452 12724 13504 12733
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 15476 12767 15528 12776
rect 15476 12733 15485 12767
rect 15485 12733 15519 12767
rect 15519 12733 15528 12767
rect 15476 12724 15528 12733
rect 16304 12792 16356 12844
rect 18236 12792 18288 12844
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 22284 12792 22336 12844
rect 23296 12928 23348 12980
rect 24032 12928 24084 12980
rect 25044 12971 25096 12980
rect 25044 12937 25053 12971
rect 25053 12937 25087 12971
rect 25087 12937 25096 12971
rect 25044 12928 25096 12937
rect 25228 12928 25280 12980
rect 22744 12860 22796 12912
rect 22928 12860 22980 12912
rect 15936 12724 15988 12776
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 20628 12724 20680 12776
rect 22008 12724 22060 12776
rect 23388 12792 23440 12844
rect 24492 12860 24544 12912
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 25044 12724 25096 12776
rect 2596 12656 2648 12708
rect 2320 12631 2372 12640
rect 2320 12597 2329 12631
rect 2329 12597 2363 12631
rect 2363 12597 2372 12631
rect 2320 12588 2372 12597
rect 6092 12656 6144 12708
rect 9128 12699 9180 12708
rect 9128 12665 9137 12699
rect 9137 12665 9171 12699
rect 9171 12665 9180 12699
rect 9128 12656 9180 12665
rect 9588 12656 9640 12708
rect 11152 12656 11204 12708
rect 9864 12588 9916 12640
rect 11612 12588 11664 12640
rect 12440 12588 12492 12640
rect 12716 12588 12768 12640
rect 18328 12656 18380 12708
rect 20720 12656 20772 12708
rect 22284 12699 22336 12708
rect 22284 12665 22293 12699
rect 22293 12665 22327 12699
rect 22327 12665 22336 12699
rect 22284 12656 22336 12665
rect 22376 12656 22428 12708
rect 13820 12588 13872 12640
rect 16120 12588 16172 12640
rect 17408 12588 17460 12640
rect 18512 12631 18564 12640
rect 18512 12597 18521 12631
rect 18521 12597 18555 12631
rect 18555 12597 18564 12631
rect 18512 12588 18564 12597
rect 19524 12588 19576 12640
rect 21272 12588 21324 12640
rect 21916 12588 21968 12640
rect 25412 12631 25464 12640
rect 25412 12597 25421 12631
rect 25421 12597 25455 12631
rect 25455 12597 25464 12631
rect 25412 12588 25464 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1768 12427 1820 12436
rect 1768 12393 1777 12427
rect 1777 12393 1811 12427
rect 1811 12393 1820 12427
rect 1768 12384 1820 12393
rect 2136 12427 2188 12436
rect 2136 12393 2145 12427
rect 2145 12393 2179 12427
rect 2179 12393 2188 12427
rect 2136 12384 2188 12393
rect 3240 12427 3292 12436
rect 3240 12393 3249 12427
rect 3249 12393 3283 12427
rect 3283 12393 3292 12427
rect 3240 12384 3292 12393
rect 4620 12384 4672 12436
rect 4804 12427 4856 12436
rect 4804 12393 4813 12427
rect 4813 12393 4847 12427
rect 4847 12393 4856 12427
rect 4804 12384 4856 12393
rect 5632 12427 5684 12436
rect 5632 12393 5641 12427
rect 5641 12393 5675 12427
rect 5675 12393 5684 12427
rect 5632 12384 5684 12393
rect 7104 12384 7156 12436
rect 8300 12384 8352 12436
rect 1400 12316 1452 12368
rect 4896 12316 4948 12368
rect 9864 12384 9916 12436
rect 12440 12384 12492 12436
rect 16672 12384 16724 12436
rect 18328 12384 18380 12436
rect 18604 12384 18656 12436
rect 20260 12384 20312 12436
rect 21456 12427 21508 12436
rect 21456 12393 21465 12427
rect 21465 12393 21499 12427
rect 21499 12393 21508 12427
rect 21456 12384 21508 12393
rect 11336 12316 11388 12368
rect 1860 12248 1912 12300
rect 2596 12248 2648 12300
rect 2780 12248 2832 12300
rect 3332 12248 3384 12300
rect 5448 12248 5500 12300
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 6368 12248 6420 12300
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10692 12248 10744 12300
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 14648 12316 14700 12368
rect 11796 12291 11848 12300
rect 11796 12257 11830 12291
rect 11830 12257 11848 12291
rect 11796 12248 11848 12257
rect 14096 12248 14148 12300
rect 15384 12248 15436 12300
rect 18880 12316 18932 12368
rect 16856 12248 16908 12300
rect 17776 12248 17828 12300
rect 20444 12248 20496 12300
rect 20720 12291 20772 12300
rect 20720 12257 20729 12291
rect 20729 12257 20763 12291
rect 20763 12257 20772 12291
rect 20720 12248 20772 12257
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 6736 12180 6788 12232
rect 7288 12180 7340 12232
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 6644 12112 6696 12164
rect 7472 12112 7524 12164
rect 10140 12180 10192 12232
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 18328 12223 18380 12232
rect 18328 12189 18337 12223
rect 18337 12189 18371 12223
rect 18371 12189 18380 12223
rect 18328 12180 18380 12189
rect 22008 12384 22060 12436
rect 23388 12384 23440 12436
rect 24308 12427 24360 12436
rect 24308 12393 24317 12427
rect 24317 12393 24351 12427
rect 24351 12393 24360 12427
rect 24308 12384 24360 12393
rect 24676 12384 24728 12436
rect 23204 12316 23256 12368
rect 25596 12248 25648 12300
rect 22100 12180 22152 12232
rect 25044 12180 25096 12232
rect 25412 12223 25464 12232
rect 25412 12189 25421 12223
rect 25421 12189 25455 12223
rect 25455 12189 25464 12223
rect 25412 12180 25464 12189
rect 8576 12112 8628 12164
rect 11428 12112 11480 12164
rect 24400 12112 24452 12164
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 13820 12044 13872 12096
rect 16212 12044 16264 12096
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 16948 12044 17000 12096
rect 17868 12044 17920 12096
rect 20444 12044 20496 12096
rect 21364 12044 21416 12096
rect 22744 12044 22796 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2320 11840 2372 11892
rect 2780 11883 2832 11892
rect 2780 11849 2789 11883
rect 2789 11849 2823 11883
rect 2823 11849 2832 11883
rect 2780 11840 2832 11849
rect 5172 11840 5224 11892
rect 6460 11840 6512 11892
rect 6644 11883 6696 11892
rect 6644 11849 6653 11883
rect 6653 11849 6687 11883
rect 6687 11849 6696 11883
rect 6644 11840 6696 11849
rect 7564 11840 7616 11892
rect 9036 11840 9088 11892
rect 10048 11840 10100 11892
rect 10784 11883 10836 11892
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 11520 11840 11572 11892
rect 12164 11840 12216 11892
rect 12992 11840 13044 11892
rect 14648 11883 14700 11892
rect 1860 11815 1912 11824
rect 1860 11781 1869 11815
rect 1869 11781 1903 11815
rect 1903 11781 1912 11815
rect 1860 11772 1912 11781
rect 1952 11772 2004 11824
rect 5356 11772 5408 11824
rect 6276 11772 6328 11824
rect 6368 11772 6420 11824
rect 7748 11704 7800 11756
rect 8576 11704 8628 11756
rect 9220 11704 9272 11756
rect 9312 11704 9364 11756
rect 12256 11772 12308 11824
rect 10784 11704 10836 11756
rect 11060 11704 11112 11756
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 11428 11747 11480 11756
rect 11428 11713 11437 11747
rect 11437 11713 11471 11747
rect 11471 11713 11480 11747
rect 11428 11704 11480 11713
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 15476 11840 15528 11892
rect 22652 11883 22704 11892
rect 22652 11849 22661 11883
rect 22661 11849 22695 11883
rect 22695 11849 22704 11883
rect 22652 11840 22704 11849
rect 23480 11883 23532 11892
rect 23480 11849 23489 11883
rect 23489 11849 23523 11883
rect 23523 11849 23532 11883
rect 23480 11840 23532 11849
rect 23664 11883 23716 11892
rect 23664 11849 23673 11883
rect 23673 11849 23707 11883
rect 23707 11849 23716 11883
rect 23664 11840 23716 11849
rect 25044 11840 25096 11892
rect 25688 11840 25740 11892
rect 16028 11772 16080 11824
rect 16212 11747 16264 11756
rect 7932 11636 7984 11688
rect 9496 11636 9548 11688
rect 11152 11679 11204 11688
rect 11152 11645 11161 11679
rect 11161 11645 11195 11679
rect 11195 11645 11204 11679
rect 11152 11636 11204 11645
rect 16212 11713 16221 11747
rect 16221 11713 16255 11747
rect 16255 11713 16264 11747
rect 16212 11704 16264 11713
rect 17960 11772 18012 11824
rect 16672 11704 16724 11756
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 18236 11704 18288 11756
rect 23204 11704 23256 11756
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 24308 11704 24360 11713
rect 25412 11704 25464 11756
rect 15384 11636 15436 11688
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 17960 11636 18012 11688
rect 22468 11679 22520 11688
rect 8300 11568 8352 11620
rect 9680 11611 9732 11620
rect 9680 11577 9689 11611
rect 9689 11577 9723 11611
rect 9723 11577 9732 11611
rect 9680 11568 9732 11577
rect 11796 11568 11848 11620
rect 13728 11568 13780 11620
rect 18328 11568 18380 11620
rect 22468 11645 22477 11679
rect 22477 11645 22511 11679
rect 22511 11645 22520 11679
rect 22468 11636 22520 11645
rect 24032 11679 24084 11688
rect 24032 11645 24041 11679
rect 24041 11645 24075 11679
rect 24075 11645 24084 11679
rect 24032 11636 24084 11645
rect 20168 11611 20220 11620
rect 20168 11577 20202 11611
rect 20202 11577 20220 11611
rect 20168 11568 20220 11577
rect 22744 11568 22796 11620
rect 11336 11500 11388 11552
rect 17408 11500 17460 11552
rect 17500 11500 17552 11552
rect 19340 11500 19392 11552
rect 21456 11500 21508 11552
rect 22100 11500 22152 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 6828 11296 6880 11348
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 7932 11296 7984 11348
rect 8484 11296 8536 11348
rect 8944 11296 8996 11348
rect 9312 11339 9364 11348
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 11244 11296 11296 11348
rect 14372 11296 14424 11348
rect 16304 11296 16356 11348
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 17960 11296 18012 11348
rect 18512 11296 18564 11348
rect 18788 11296 18840 11348
rect 21272 11296 21324 11348
rect 23204 11296 23256 11348
rect 24032 11339 24084 11348
rect 24032 11305 24041 11339
rect 24041 11305 24075 11339
rect 24075 11305 24084 11339
rect 24032 11296 24084 11305
rect 24308 11296 24360 11348
rect 25228 11296 25280 11348
rect 10048 11228 10100 11280
rect 11428 11228 11480 11280
rect 11888 11228 11940 11280
rect 15568 11271 15620 11280
rect 15568 11237 15602 11271
rect 15602 11237 15620 11271
rect 15568 11228 15620 11237
rect 16028 11228 16080 11280
rect 18604 11271 18656 11280
rect 18604 11237 18638 11271
rect 18638 11237 18656 11271
rect 18604 11228 18656 11237
rect 25136 11228 25188 11280
rect 25596 11271 25648 11280
rect 25596 11237 25605 11271
rect 25605 11237 25639 11271
rect 25639 11237 25648 11271
rect 25596 11228 25648 11237
rect 8392 11160 8444 11212
rect 8668 11160 8720 11212
rect 11244 11160 11296 11212
rect 11796 11160 11848 11212
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 15384 11160 15436 11212
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 11428 11135 11480 11144
rect 8576 11092 8628 11101
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 6000 11024 6052 11076
rect 8116 11024 8168 11076
rect 11704 11092 11756 11144
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 10876 10956 10928 11008
rect 13728 11092 13780 11144
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 21916 11092 21968 11144
rect 17960 11024 18012 11076
rect 19340 11024 19392 11076
rect 20168 11024 20220 11076
rect 21824 11024 21876 11076
rect 22100 11135 22152 11144
rect 22100 11101 22109 11135
rect 22109 11101 22143 11135
rect 22143 11101 22152 11135
rect 22100 11092 22152 11101
rect 24216 11024 24268 11076
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 12532 10956 12584 10965
rect 24032 10956 24084 11008
rect 24952 10956 25004 11008
rect 25136 10956 25188 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 8116 10752 8168 10804
rect 8484 10795 8536 10804
rect 8484 10761 8493 10795
rect 8493 10761 8527 10795
rect 8527 10761 8536 10795
rect 8484 10752 8536 10761
rect 9220 10795 9272 10804
rect 9220 10761 9229 10795
rect 9229 10761 9263 10795
rect 9263 10761 9272 10795
rect 9220 10752 9272 10761
rect 9680 10752 9732 10804
rect 13820 10795 13872 10804
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 15384 10752 15436 10804
rect 16028 10752 16080 10804
rect 16120 10752 16172 10804
rect 16580 10752 16632 10804
rect 18052 10752 18104 10804
rect 12164 10727 12216 10736
rect 12164 10693 12173 10727
rect 12173 10693 12207 10727
rect 12207 10693 12216 10727
rect 12164 10684 12216 10693
rect 13912 10684 13964 10736
rect 18604 10684 18656 10736
rect 8208 10616 8260 10668
rect 9312 10616 9364 10668
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 11612 10616 11664 10668
rect 15016 10616 15068 10668
rect 19524 10752 19576 10804
rect 20076 10795 20128 10804
rect 20076 10761 20085 10795
rect 20085 10761 20119 10795
rect 20119 10761 20128 10795
rect 20076 10752 20128 10761
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 10140 10480 10192 10532
rect 12808 10480 12860 10532
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 11428 10412 11480 10464
rect 11796 10455 11848 10464
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 13820 10412 13872 10464
rect 14464 10412 14516 10464
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 15476 10412 15528 10464
rect 16580 10412 16632 10464
rect 17960 10548 18012 10600
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 19340 10616 19392 10668
rect 20628 10548 20680 10600
rect 22008 10752 22060 10804
rect 22100 10752 22152 10804
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 23480 10752 23532 10761
rect 24032 10752 24084 10804
rect 25228 10752 25280 10804
rect 25780 10752 25832 10804
rect 25872 10795 25924 10804
rect 25872 10761 25881 10795
rect 25881 10761 25915 10795
rect 25915 10761 25924 10795
rect 25872 10752 25924 10761
rect 24676 10684 24728 10736
rect 26056 10684 26108 10736
rect 23480 10548 23532 10600
rect 25044 10548 25096 10600
rect 25872 10548 25924 10600
rect 19340 10455 19392 10464
rect 19340 10421 19349 10455
rect 19349 10421 19383 10455
rect 19383 10421 19392 10455
rect 19340 10412 19392 10421
rect 24216 10480 24268 10532
rect 21456 10412 21508 10464
rect 22284 10412 22336 10464
rect 23848 10412 23900 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 10048 10208 10100 10260
rect 10968 10208 11020 10260
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 15016 10251 15068 10260
rect 15016 10217 15025 10251
rect 15025 10217 15059 10251
rect 15059 10217 15068 10251
rect 15016 10208 15068 10217
rect 15292 10208 15344 10260
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 18604 10208 18656 10260
rect 19156 10251 19208 10260
rect 19156 10217 19165 10251
rect 19165 10217 19199 10251
rect 19199 10217 19208 10251
rect 19156 10208 19208 10217
rect 20904 10251 20956 10260
rect 20904 10217 20913 10251
rect 20913 10217 20947 10251
rect 20947 10217 20956 10251
rect 20904 10208 20956 10217
rect 24216 10251 24268 10260
rect 24216 10217 24225 10251
rect 24225 10217 24259 10251
rect 24259 10217 24268 10251
rect 24216 10208 24268 10217
rect 10692 10140 10744 10192
rect 16304 10183 16356 10192
rect 16304 10149 16338 10183
rect 16338 10149 16356 10183
rect 16304 10140 16356 10149
rect 19340 10140 19392 10192
rect 22284 10140 22336 10192
rect 9588 10072 9640 10124
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12440 10115 12492 10124
rect 12440 10081 12474 10115
rect 12474 10081 12492 10115
rect 16028 10115 16080 10124
rect 12440 10072 12492 10081
rect 16028 10081 16037 10115
rect 16037 10081 16071 10115
rect 16071 10081 16080 10115
rect 16028 10072 16080 10081
rect 22008 10072 22060 10124
rect 23020 10072 23072 10124
rect 10876 10004 10928 10056
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 18696 10004 18748 10056
rect 19432 10004 19484 10056
rect 18512 9936 18564 9988
rect 23940 9936 23992 9988
rect 12808 9868 12860 9920
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 13544 9868 13596 9877
rect 17592 9868 17644 9920
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 18328 9868 18380 9877
rect 20628 9868 20680 9920
rect 21824 9868 21876 9920
rect 23848 9911 23900 9920
rect 23848 9877 23857 9911
rect 23857 9877 23891 9911
rect 23891 9877 23900 9911
rect 23848 9868 23900 9877
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 11152 9707 11204 9716
rect 11152 9673 11161 9707
rect 11161 9673 11195 9707
rect 11195 9673 11204 9707
rect 11152 9664 11204 9673
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 12348 9664 12400 9716
rect 12440 9664 12492 9716
rect 12624 9664 12676 9716
rect 14648 9664 14700 9716
rect 15292 9664 15344 9716
rect 16304 9664 16356 9716
rect 9680 9596 9732 9648
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 16212 9639 16264 9648
rect 16212 9605 16221 9639
rect 16221 9605 16255 9639
rect 16255 9605 16264 9639
rect 16212 9596 16264 9605
rect 22008 9664 22060 9716
rect 23020 9664 23072 9716
rect 23296 9664 23348 9716
rect 19432 9596 19484 9648
rect 24676 9596 24728 9648
rect 12440 9528 12492 9580
rect 16764 9528 16816 9580
rect 16948 9528 17000 9580
rect 22284 9571 22336 9580
rect 22284 9537 22293 9571
rect 22293 9537 22327 9571
rect 22327 9537 22336 9571
rect 22284 9528 22336 9537
rect 10048 9460 10100 9512
rect 12348 9460 12400 9512
rect 18328 9503 18380 9512
rect 14280 9392 14332 9444
rect 16672 9435 16724 9444
rect 16672 9401 16681 9435
rect 16681 9401 16715 9435
rect 16715 9401 16724 9435
rect 16672 9392 16724 9401
rect 18328 9469 18337 9503
rect 18337 9469 18371 9503
rect 18371 9469 18380 9503
rect 18328 9460 18380 9469
rect 20904 9460 20956 9512
rect 24584 9503 24636 9512
rect 24584 9469 24593 9503
rect 24593 9469 24627 9503
rect 24627 9469 24636 9503
rect 24584 9460 24636 9469
rect 18512 9392 18564 9444
rect 22008 9435 22060 9444
rect 22008 9401 22017 9435
rect 22017 9401 22051 9435
rect 22051 9401 22060 9435
rect 22008 9392 22060 9401
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 11152 9324 11204 9376
rect 11888 9324 11940 9376
rect 12256 9324 12308 9376
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 16856 9324 16908 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 18880 9324 18932 9376
rect 20444 9324 20496 9376
rect 21732 9324 21784 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 10968 9120 11020 9172
rect 13728 9120 13780 9172
rect 14004 9120 14056 9172
rect 14648 9120 14700 9172
rect 16488 9120 16540 9172
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 19432 9163 19484 9172
rect 19432 9129 19441 9163
rect 19441 9129 19475 9163
rect 19475 9129 19484 9163
rect 19432 9120 19484 9129
rect 19524 9120 19576 9172
rect 20904 9163 20956 9172
rect 20904 9129 20913 9163
rect 20913 9129 20947 9163
rect 20947 9129 20956 9163
rect 20904 9120 20956 9129
rect 22100 9120 22152 9172
rect 22836 9163 22888 9172
rect 22836 9129 22845 9163
rect 22845 9129 22879 9163
rect 22879 9129 22888 9163
rect 22836 9120 22888 9129
rect 24768 9163 24820 9172
rect 24768 9129 24777 9163
rect 24777 9129 24811 9163
rect 24811 9129 24820 9163
rect 24768 9120 24820 9129
rect 13268 9052 13320 9104
rect 14372 9052 14424 9104
rect 16028 9052 16080 9104
rect 16396 9052 16448 9104
rect 12256 9027 12308 9036
rect 12256 8993 12265 9027
rect 12265 8993 12299 9027
rect 12299 8993 12308 9027
rect 12256 8984 12308 8993
rect 13360 8984 13412 9036
rect 13728 8984 13780 9036
rect 15752 8984 15804 9036
rect 17776 9052 17828 9104
rect 22284 9052 22336 9104
rect 17408 9027 17460 9036
rect 17408 8993 17442 9027
rect 17442 8993 17460 9027
rect 17408 8984 17460 8993
rect 20352 8984 20404 9036
rect 20904 8984 20956 9036
rect 22468 8984 22520 9036
rect 22744 8984 22796 9036
rect 11704 8916 11756 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 12624 8916 12676 8968
rect 14280 8916 14332 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 16120 8959 16172 8968
rect 16120 8925 16129 8959
rect 16129 8925 16163 8959
rect 16163 8925 16172 8959
rect 16120 8916 16172 8925
rect 20628 8916 20680 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 24676 8984 24728 9036
rect 21456 8916 21508 8925
rect 23204 8916 23256 8968
rect 18512 8891 18564 8900
rect 18512 8857 18521 8891
rect 18521 8857 18555 8891
rect 18555 8857 18564 8891
rect 18512 8848 18564 8857
rect 20720 8823 20772 8832
rect 20720 8789 20729 8823
rect 20729 8789 20763 8823
rect 20763 8789 20772 8823
rect 20720 8780 20772 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 12256 8576 12308 8628
rect 12992 8576 13044 8628
rect 13268 8576 13320 8628
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 15384 8576 15436 8628
rect 16120 8576 16172 8628
rect 17776 8576 17828 8628
rect 18880 8619 18932 8628
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 20812 8576 20864 8628
rect 22836 8619 22888 8628
rect 22836 8585 22845 8619
rect 22845 8585 22879 8619
rect 22879 8585 22888 8619
rect 22836 8576 22888 8585
rect 23204 8619 23256 8628
rect 23204 8585 23213 8619
rect 23213 8585 23247 8619
rect 23247 8585 23256 8619
rect 23204 8576 23256 8585
rect 25412 8576 25464 8628
rect 20904 8551 20956 8560
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13544 8483 13596 8492
rect 13360 8440 13412 8449
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 14648 8440 14700 8492
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17408 8440 17460 8492
rect 19432 8440 19484 8492
rect 20904 8517 20913 8551
rect 20913 8517 20947 8551
rect 20947 8517 20956 8551
rect 20904 8508 20956 8517
rect 21732 8483 21784 8492
rect 21732 8449 21741 8483
rect 21741 8449 21775 8483
rect 21775 8449 21784 8483
rect 21732 8440 21784 8449
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 24124 8440 24176 8492
rect 12624 8372 12676 8424
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 16580 8372 16632 8424
rect 17776 8372 17828 8424
rect 19708 8415 19760 8424
rect 19708 8381 19717 8415
rect 19717 8381 19751 8415
rect 19751 8381 19760 8415
rect 19708 8372 19760 8381
rect 20536 8415 20588 8424
rect 20536 8381 20545 8415
rect 20545 8381 20579 8415
rect 20579 8381 20588 8415
rect 20536 8372 20588 8381
rect 20720 8372 20772 8424
rect 22100 8372 22152 8424
rect 25044 8415 25096 8424
rect 25044 8381 25053 8415
rect 25053 8381 25087 8415
rect 25087 8381 25096 8415
rect 25044 8372 25096 8381
rect 11704 8304 11756 8356
rect 14648 8304 14700 8356
rect 16764 8347 16816 8356
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 14464 8236 14516 8288
rect 15752 8236 15804 8288
rect 17868 8236 17920 8288
rect 22468 8279 22520 8288
rect 22468 8245 22477 8279
rect 22477 8245 22511 8279
rect 22511 8245 22520 8279
rect 22468 8236 22520 8245
rect 23848 8236 23900 8288
rect 24676 8236 24728 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 11888 8075 11940 8084
rect 11888 8041 11897 8075
rect 11897 8041 11931 8075
rect 11931 8041 11940 8075
rect 11888 8032 11940 8041
rect 13268 8075 13320 8084
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 14556 8032 14608 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 15660 8075 15712 8084
rect 15660 8041 15669 8075
rect 15669 8041 15703 8075
rect 15703 8041 15712 8075
rect 15660 8032 15712 8041
rect 16488 8032 16540 8084
rect 16948 8032 17000 8084
rect 20352 8032 20404 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 22100 8075 22152 8084
rect 22100 8041 22109 8075
rect 22109 8041 22143 8075
rect 22143 8041 22152 8075
rect 22100 8032 22152 8041
rect 23112 8032 23164 8084
rect 23940 8032 23992 8084
rect 25964 8032 26016 8084
rect 9956 7964 10008 8016
rect 12808 7964 12860 8016
rect 13544 7964 13596 8016
rect 21456 7964 21508 8016
rect 11888 7896 11940 7948
rect 12532 7896 12584 7948
rect 13452 7939 13504 7948
rect 13452 7905 13461 7939
rect 13461 7905 13495 7939
rect 13495 7905 13504 7939
rect 13452 7896 13504 7905
rect 14832 7896 14884 7948
rect 15476 7939 15528 7948
rect 15476 7905 15485 7939
rect 15485 7905 15519 7939
rect 15519 7905 15528 7939
rect 15476 7896 15528 7905
rect 16396 7896 16448 7948
rect 17592 7896 17644 7948
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 21824 7896 21876 7948
rect 22100 7896 22152 7948
rect 22652 7939 22704 7948
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 23756 7896 23808 7948
rect 24124 7896 24176 7948
rect 24676 7939 24728 7948
rect 24676 7905 24685 7939
rect 24685 7905 24719 7939
rect 24719 7905 24728 7939
rect 24676 7896 24728 7905
rect 12624 7828 12676 7880
rect 19156 7828 19208 7880
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 20628 7828 20680 7880
rect 23664 7760 23716 7812
rect 23940 7760 23992 7812
rect 14280 7692 14332 7744
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 16396 7735 16448 7744
rect 16396 7701 16405 7735
rect 16405 7701 16439 7735
rect 16439 7701 16448 7735
rect 16396 7692 16448 7701
rect 18972 7735 19024 7744
rect 18972 7701 18981 7735
rect 18981 7701 19015 7735
rect 19015 7701 19024 7735
rect 18972 7692 19024 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 12624 7488 12676 7540
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 15752 7488 15804 7540
rect 16028 7488 16080 7540
rect 17776 7488 17828 7540
rect 19156 7531 19208 7540
rect 19156 7497 19165 7531
rect 19165 7497 19199 7531
rect 19199 7497 19208 7531
rect 19156 7488 19208 7497
rect 19984 7488 20036 7540
rect 20628 7531 20680 7540
rect 20628 7497 20637 7531
rect 20637 7497 20671 7531
rect 20671 7497 20680 7531
rect 20628 7488 20680 7497
rect 22652 7488 22704 7540
rect 23848 7531 23900 7540
rect 23848 7497 23857 7531
rect 23857 7497 23891 7531
rect 23891 7497 23900 7531
rect 23848 7488 23900 7497
rect 24124 7531 24176 7540
rect 24124 7497 24133 7531
rect 24133 7497 24167 7531
rect 24167 7497 24176 7531
rect 24124 7488 24176 7497
rect 24676 7488 24728 7540
rect 14740 7352 14792 7404
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 16396 7352 16448 7404
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 25320 7420 25372 7472
rect 16948 7352 17000 7361
rect 17592 7352 17644 7404
rect 19616 7352 19668 7404
rect 20260 7395 20312 7404
rect 20260 7361 20269 7395
rect 20269 7361 20303 7395
rect 20303 7361 20312 7395
rect 20260 7352 20312 7361
rect 20996 7352 21048 7404
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 23940 7352 23992 7404
rect 24124 7352 24176 7404
rect 12808 7284 12860 7336
rect 16488 7284 16540 7336
rect 18972 7284 19024 7336
rect 19432 7284 19484 7336
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 17684 7216 17736 7268
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 18144 7148 18196 7200
rect 18512 7191 18564 7200
rect 18512 7157 18521 7191
rect 18521 7157 18555 7191
rect 18555 7157 18564 7191
rect 19984 7191 20036 7200
rect 18512 7148 18564 7157
rect 19984 7157 19993 7191
rect 19993 7157 20027 7191
rect 20027 7157 20036 7191
rect 19984 7148 20036 7157
rect 23388 7148 23440 7200
rect 23664 7148 23716 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 15476 6987 15528 6996
rect 15476 6953 15485 6987
rect 15485 6953 15519 6987
rect 15519 6953 15528 6987
rect 15476 6944 15528 6953
rect 16948 6944 17000 6996
rect 17868 6944 17920 6996
rect 19248 6944 19300 6996
rect 19432 6944 19484 6996
rect 20260 6944 20312 6996
rect 16488 6808 16540 6860
rect 23756 6851 23808 6860
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 24768 6851 24820 6860
rect 24768 6817 24777 6851
rect 24777 6817 24811 6851
rect 24811 6817 24820 6851
rect 24768 6808 24820 6817
rect 16764 6740 16816 6792
rect 17408 6740 17460 6792
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 16948 6604 17000 6656
rect 23940 6715 23992 6724
rect 23940 6681 23949 6715
rect 23949 6681 23983 6715
rect 23983 6681 23992 6715
rect 23940 6672 23992 6681
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 15384 6400 15436 6452
rect 16396 6443 16448 6452
rect 16396 6409 16405 6443
rect 16405 6409 16439 6443
rect 16439 6409 16448 6443
rect 16396 6400 16448 6409
rect 17868 6443 17920 6452
rect 17868 6409 17877 6443
rect 17877 6409 17911 6443
rect 17911 6409 17920 6443
rect 17868 6400 17920 6409
rect 23756 6400 23808 6452
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 16396 6060 16448 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 16396 5899 16448 5908
rect 16396 5865 16405 5899
rect 16405 5865 16439 5899
rect 16439 5865 16448 5899
rect 16396 5856 16448 5865
rect 16948 5856 17000 5908
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 13728 2456 13780 2508
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12440 2320 12492 2372
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 2042 27520 2098 28000
rect 2594 27520 2650 28000
rect 3146 27520 3202 28000
rect 3790 27520 3846 28000
rect 4158 27704 4214 27713
rect 4158 27639 4214 27648
rect 308 16522 336 27520
rect 860 19009 888 27520
rect 1412 25786 1440 27520
rect 1858 26616 1914 26625
rect 1858 26551 1914 26560
rect 1228 25758 1440 25786
rect 1122 20360 1178 20369
rect 1122 20295 1178 20304
rect 1136 19446 1164 20295
rect 1124 19440 1176 19446
rect 1124 19382 1176 19388
rect 846 19000 902 19009
rect 846 18935 902 18944
rect 1228 16726 1256 25758
rect 1400 25696 1452 25702
rect 1400 25638 1452 25644
rect 1412 25498 1440 25638
rect 1400 25492 1452 25498
rect 1400 25434 1452 25440
rect 1306 25392 1362 25401
rect 1306 25327 1362 25336
rect 1320 23254 1348 25327
rect 1766 25256 1822 25265
rect 1766 25191 1822 25200
rect 1400 24948 1452 24954
rect 1400 24890 1452 24896
rect 1412 24274 1440 24890
rect 1676 24812 1728 24818
rect 1676 24754 1728 24760
rect 1688 24410 1716 24754
rect 1676 24404 1728 24410
rect 1504 24364 1676 24392
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1308 23248 1360 23254
rect 1308 23190 1360 23196
rect 1320 22438 1348 23190
rect 1308 22432 1360 22438
rect 1308 22374 1360 22380
rect 1400 21956 1452 21962
rect 1400 21898 1452 21904
rect 1412 21570 1440 21898
rect 1320 21542 1440 21570
rect 1216 16720 1268 16726
rect 1216 16662 1268 16668
rect 296 16516 348 16522
rect 296 16458 348 16464
rect 1320 15450 1348 21542
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 21146 1440 21422
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 17218 1440 20334
rect 1504 20097 1532 24364
rect 1676 24346 1728 24352
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 1596 23361 1624 24006
rect 1780 23866 1808 25191
rect 1768 23860 1820 23866
rect 1768 23802 1820 23808
rect 1582 23352 1638 23361
rect 1582 23287 1638 23296
rect 1872 23100 1900 26551
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 1964 24614 1992 25094
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1952 24268 2004 24274
rect 1952 24210 2004 24216
rect 1964 23866 1992 24210
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1688 23072 1900 23100
rect 1950 23080 2006 23089
rect 1688 22234 1716 23072
rect 1950 23015 1952 23024
rect 2004 23015 2006 23024
rect 1952 22986 2004 22992
rect 1964 22574 1992 22986
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1952 22568 2004 22574
rect 1952 22510 2004 22516
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1688 21690 1716 22170
rect 1676 21684 1728 21690
rect 1676 21626 1728 21632
rect 1780 21434 1808 22510
rect 1860 22432 1912 22438
rect 1860 22374 1912 22380
rect 1872 22098 1900 22374
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1688 21406 1808 21434
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1490 20088 1546 20097
rect 1490 20023 1546 20032
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 17814 1532 19654
rect 1492 17808 1544 17814
rect 1492 17750 1544 17756
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1504 17338 1532 17614
rect 1596 17513 1624 20198
rect 1688 19961 1716 21406
rect 1768 21344 1820 21350
rect 1768 21286 1820 21292
rect 1674 19952 1730 19961
rect 1674 19887 1730 19896
rect 1676 19236 1728 19242
rect 1676 19178 1728 19184
rect 1582 17504 1638 17513
rect 1582 17439 1638 17448
rect 1492 17332 1544 17338
rect 1492 17274 1544 17280
rect 1582 17232 1638 17241
rect 1412 17190 1532 17218
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 1412 15570 1440 16390
rect 1504 15586 1532 17190
rect 1582 17167 1638 17176
rect 1596 16794 1624 17167
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1596 15745 1624 15846
rect 1582 15736 1638 15745
rect 1688 15706 1716 19178
rect 1780 18834 1808 21286
rect 1872 21146 1900 22034
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1964 21622 1992 21966
rect 2056 21706 2084 27520
rect 2320 25152 2372 25158
rect 2320 25094 2372 25100
rect 2412 25152 2464 25158
rect 2412 25094 2464 25100
rect 2134 24712 2190 24721
rect 2134 24647 2190 24656
rect 2228 24676 2280 24682
rect 2148 23662 2176 24647
rect 2228 24618 2280 24624
rect 2136 23656 2188 23662
rect 2136 23598 2188 23604
rect 2240 22030 2268 24618
rect 2332 22982 2360 25094
rect 2424 24750 2452 25094
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2516 24426 2544 24754
rect 2424 24398 2544 24426
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22642 2360 22918
rect 2320 22636 2372 22642
rect 2320 22578 2372 22584
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 2424 21944 2452 24398
rect 2504 24336 2556 24342
rect 2504 24278 2556 24284
rect 2516 23662 2544 24278
rect 2504 23656 2556 23662
rect 2504 23598 2556 23604
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 2516 22817 2544 22918
rect 2502 22808 2558 22817
rect 2502 22743 2558 22752
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2516 22234 2544 22578
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 2332 21916 2452 21944
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2056 21678 2176 21706
rect 1952 21616 2004 21622
rect 1952 21558 2004 21564
rect 2042 21584 2098 21593
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 1872 20874 1900 21082
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 1860 20256 1912 20262
rect 1964 20244 1992 21558
rect 2042 21519 2044 21528
rect 2096 21519 2098 21528
rect 2044 21490 2096 21496
rect 2056 21146 2084 21490
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 1912 20216 1992 20244
rect 1860 20198 1912 20204
rect 1872 19718 1900 20198
rect 2148 19990 2176 21678
rect 2136 19984 2188 19990
rect 2136 19926 2188 19932
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 2056 19378 2084 19654
rect 2044 19372 2096 19378
rect 2240 19360 2268 21830
rect 2332 20602 2360 21916
rect 2504 21888 2556 21894
rect 2410 21856 2466 21865
rect 2504 21830 2556 21836
rect 2410 21791 2466 21800
rect 2424 21146 2452 21791
rect 2516 21486 2544 21830
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 2608 20890 2636 27520
rect 2872 25492 2924 25498
rect 2700 25452 2872 25480
rect 2700 24818 2728 25452
rect 2872 25434 2924 25440
rect 2964 25492 3016 25498
rect 2964 25434 3016 25440
rect 2872 25288 2924 25294
rect 2872 25230 2924 25236
rect 2778 24848 2834 24857
rect 2688 24812 2740 24818
rect 2778 24783 2834 24792
rect 2688 24754 2740 24760
rect 2688 24676 2740 24682
rect 2688 24618 2740 24624
rect 2700 22273 2728 24618
rect 2792 23662 2820 24783
rect 2884 24614 2912 25230
rect 2872 24608 2924 24614
rect 2872 24550 2924 24556
rect 2870 24304 2926 24313
rect 2870 24239 2926 24248
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2780 23520 2832 23526
rect 2778 23488 2780 23497
rect 2832 23488 2834 23497
rect 2778 23423 2834 23432
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 22778 2820 23122
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2686 22264 2742 22273
rect 2686 22199 2742 22208
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2516 20862 2636 20890
rect 2700 20890 2728 21626
rect 2792 21457 2820 22578
rect 2778 21448 2834 21457
rect 2778 21383 2834 21392
rect 2884 21026 2912 24239
rect 2976 22642 3004 25434
rect 3054 25392 3110 25401
rect 3054 25327 3110 25336
rect 3068 25294 3096 25327
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3068 24410 3096 25230
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3056 23520 3108 23526
rect 3056 23462 3108 23468
rect 2964 22636 3016 22642
rect 2964 22578 3016 22584
rect 3068 22001 3096 23462
rect 3054 21992 3110 22001
rect 3054 21927 3110 21936
rect 2884 20998 3004 21026
rect 2872 20936 2924 20942
rect 2700 20862 2820 20890
rect 2872 20878 2924 20884
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 2410 20496 2466 20505
rect 2410 20431 2466 20440
rect 2424 20058 2452 20431
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2318 19544 2374 19553
rect 2318 19479 2374 19488
rect 2044 19314 2096 19320
rect 2148 19332 2268 19360
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1582 15671 1638 15680
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1400 15564 1452 15570
rect 1504 15558 1716 15586
rect 1400 15506 1452 15512
rect 1320 15422 1532 15450
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1412 14958 1440 15302
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1504 14550 1532 15422
rect 1582 15192 1638 15201
rect 1582 15127 1584 15136
rect 1636 15127 1638 15136
rect 1584 15098 1636 15104
rect 1582 14648 1638 14657
rect 1582 14583 1638 14592
rect 1492 14544 1544 14550
rect 1492 14486 1544 14492
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 13870 1440 14214
rect 1596 14074 1624 14583
rect 1584 14068 1636 14074
rect 1584 14010 1636 14016
rect 1490 13968 1546 13977
rect 1688 13938 1716 15558
rect 1490 13903 1546 13912
rect 1676 13932 1728 13938
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 12374 1440 13806
rect 1504 12986 1532 13903
rect 1676 13874 1728 13880
rect 1780 13530 1808 18770
rect 1872 15094 1900 19246
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1964 18873 1992 19110
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 1964 18290 1992 18799
rect 2056 18766 2084 19314
rect 2148 18970 2176 19332
rect 2332 19310 2360 19479
rect 2320 19304 2372 19310
rect 2226 19272 2282 19281
rect 2320 19246 2372 19252
rect 2226 19207 2228 19216
rect 2280 19207 2282 19216
rect 2228 19178 2280 19184
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 2148 18714 2176 18906
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1860 15088 1912 15094
rect 1860 15030 1912 15036
rect 1860 14544 1912 14550
rect 1860 14486 1912 14492
rect 1872 14074 1900 14486
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1596 13433 1624 13466
rect 1582 13424 1638 13433
rect 1582 13359 1638 13368
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1400 12368 1452 12374
rect 1780 12345 1808 12378
rect 1400 12310 1452 12316
rect 1766 12336 1822 12345
rect 1766 12271 1822 12280
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1872 11830 1900 12242
rect 1964 11830 1992 18090
rect 2056 17882 2084 18702
rect 2148 18686 2268 18714
rect 2136 18624 2188 18630
rect 2136 18566 2188 18572
rect 2148 18086 2176 18566
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16794 2084 17138
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2056 16250 2084 16730
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2042 16008 2098 16017
rect 2042 15943 2044 15952
rect 2096 15943 2098 15952
rect 2044 15914 2096 15920
rect 2148 13530 2176 18022
rect 2240 17921 2268 18686
rect 2226 17912 2282 17921
rect 2226 17847 2282 17856
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 16454 2268 17682
rect 2424 16969 2452 19722
rect 2410 16960 2466 16969
rect 2410 16895 2466 16904
rect 2516 16810 2544 20862
rect 2596 20800 2648 20806
rect 2596 20742 2648 20748
rect 2608 19922 2636 20742
rect 2792 20641 2820 20862
rect 2778 20632 2834 20641
rect 2778 20567 2834 20576
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2792 19922 2820 20334
rect 2884 20262 2912 20878
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2332 16782 2544 16810
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2226 16280 2282 16289
rect 2226 16215 2282 16224
rect 2240 14074 2268 16215
rect 2332 14396 2360 16782
rect 2608 16658 2636 19858
rect 2792 19802 2820 19858
rect 2700 19774 2820 19802
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2700 18834 2728 19774
rect 2778 19680 2834 19689
rect 2778 19615 2834 19624
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2792 18170 2820 19615
rect 2884 18970 2912 19790
rect 2976 19394 3004 20998
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 3068 20058 3096 20810
rect 3160 20602 3188 27520
rect 3606 27160 3662 27169
rect 3606 27095 3662 27104
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3436 24750 3464 25094
rect 3528 24954 3556 25094
rect 3516 24948 3568 24954
rect 3516 24890 3568 24896
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3252 24070 3280 24686
rect 3332 24608 3384 24614
rect 3330 24576 3332 24585
rect 3384 24576 3386 24585
rect 3330 24511 3386 24520
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3344 23848 3372 24142
rect 3252 23820 3372 23848
rect 3252 23730 3280 23820
rect 3330 23760 3386 23769
rect 3240 23724 3292 23730
rect 3330 23695 3386 23704
rect 3240 23666 3292 23672
rect 3252 23186 3280 23666
rect 3240 23180 3292 23186
rect 3240 23122 3292 23128
rect 3252 23050 3280 23122
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3252 22234 3280 22986
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3238 21312 3294 21321
rect 3238 21247 3294 21256
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3146 20496 3202 20505
rect 3146 20431 3202 20440
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3068 19514 3096 19994
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 2976 19366 3096 19394
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2700 18142 2820 18170
rect 2700 16674 2728 18142
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2792 17338 2820 18022
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 2884 17542 2912 17818
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2884 17134 2912 17478
rect 2976 17377 3004 18770
rect 2962 17368 3018 17377
rect 2962 17303 3018 17312
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 16794 2912 17070
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2596 16652 2648 16658
rect 2700 16646 3004 16674
rect 2596 16594 2648 16600
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2424 14521 2452 16390
rect 2594 16144 2650 16153
rect 2594 16079 2650 16088
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2516 15502 2544 15642
rect 2608 15638 2636 16079
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 15162 2544 15438
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2608 14618 2636 15574
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2410 14512 2466 14521
rect 2410 14447 2466 14456
rect 2332 14368 2452 14396
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2042 12744 2098 12753
rect 2042 12679 2044 12688
rect 2096 12679 2098 12688
rect 2044 12650 2096 12656
rect 2148 12442 2176 13330
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 1860 11824 1912 11830
rect 1860 11766 1912 11772
rect 1952 11824 2004 11830
rect 1952 11766 2004 11772
rect 2240 9081 2268 13874
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2332 11898 2360 12582
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2424 10441 2452 14368
rect 2700 14278 2728 16526
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 2792 15706 2820 15807
rect 2884 15706 2912 16526
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2976 15008 3004 16646
rect 3068 16153 3096 19366
rect 3160 19145 3188 20431
rect 3252 20398 3280 21247
rect 3344 21146 3372 23695
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3436 22098 3464 23598
rect 3528 22778 3556 24890
rect 3620 23322 3648 27095
rect 3804 24834 3832 27520
rect 3882 26072 3938 26081
rect 3882 26007 3938 26016
rect 3712 24806 3832 24834
rect 3608 23316 3660 23322
rect 3608 23258 3660 23264
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3620 22710 3648 23258
rect 3608 22704 3660 22710
rect 3608 22646 3660 22652
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3620 22001 3648 22646
rect 3606 21992 3662 22001
rect 3424 21956 3476 21962
rect 3606 21927 3662 21936
rect 3424 21898 3476 21904
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3436 20890 3464 21898
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3620 21418 3648 21830
rect 3712 21457 3740 24806
rect 3896 24732 3924 26007
rect 3976 25356 4028 25362
rect 3976 25298 4028 25304
rect 3988 25265 4016 25298
rect 3974 25256 4030 25265
rect 3974 25191 4030 25200
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 3804 24704 3924 24732
rect 3804 23066 3832 24704
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3896 24410 3924 24550
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3896 23662 3924 24346
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3988 23730 4016 24006
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3896 23186 3924 23598
rect 3988 23186 4016 23666
rect 3884 23180 3936 23186
rect 3884 23122 3936 23128
rect 3976 23180 4028 23186
rect 3976 23122 4028 23128
rect 3804 23038 4016 23066
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3884 22976 3936 22982
rect 3884 22918 3936 22924
rect 3804 22438 3832 22918
rect 3896 22642 3924 22918
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3896 22234 3924 22578
rect 3884 22228 3936 22234
rect 3884 22170 3936 22176
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3698 21448 3754 21457
rect 3608 21412 3660 21418
rect 3698 21383 3754 21392
rect 3608 21354 3660 21360
rect 3620 21010 3648 21354
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3608 21004 3660 21010
rect 3608 20946 3660 20952
rect 3712 20942 3740 21286
rect 3344 20862 3464 20890
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3344 20448 3372 20862
rect 3516 20596 3568 20602
rect 3516 20538 3568 20544
rect 3344 20420 3464 20448
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 3330 20360 3386 20369
rect 3146 19136 3202 19145
rect 3146 19071 3202 19080
rect 3252 18698 3280 20334
rect 3330 20295 3332 20304
rect 3384 20295 3386 20304
rect 3332 20266 3384 20272
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3344 18408 3372 19926
rect 3252 18380 3372 18408
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3160 16590 3188 17002
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3054 16144 3110 16153
rect 3054 16079 3110 16088
rect 3160 15638 3188 16526
rect 3252 16046 3280 18380
rect 3436 18306 3464 20420
rect 3528 20398 3556 20538
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3712 20330 3740 20878
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3528 18737 3556 20198
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 3712 19378 3740 19654
rect 3804 19446 3832 22034
rect 3882 21584 3938 21593
rect 3882 21519 3938 21528
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3896 19310 3924 21519
rect 3988 20534 4016 23038
rect 4080 22574 4108 25162
rect 4172 24410 4200 27639
rect 4342 27520 4398 28000
rect 4894 27520 4950 28000
rect 5538 27520 5594 28000
rect 6090 27520 6146 28000
rect 6642 27520 6698 28000
rect 7286 27520 7342 28000
rect 7838 27520 7894 28000
rect 8390 27520 8446 28000
rect 9034 27520 9090 28000
rect 9586 27520 9642 28000
rect 10138 27520 10194 28000
rect 10782 27520 10838 28000
rect 11334 27520 11390 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 16026 27520 16082 28000
rect 16578 27520 16634 28000
rect 17130 27520 17186 28000
rect 17774 27520 17830 28000
rect 18326 27520 18382 28000
rect 18878 27520 18934 28000
rect 19522 27520 19578 28000
rect 20074 27520 20130 28000
rect 20626 27520 20682 28000
rect 21270 27520 21326 28000
rect 21822 27520 21878 28000
rect 22374 27520 22430 28000
rect 23018 27520 23074 28000
rect 23570 27520 23626 28000
rect 23754 27704 23810 27713
rect 23754 27639 23810 27648
rect 4356 24954 4384 27520
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4436 24744 4488 24750
rect 4436 24686 4488 24692
rect 4160 24404 4212 24410
rect 4160 24346 4212 24352
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 4172 23497 4200 24006
rect 4158 23488 4214 23497
rect 4158 23423 4214 23432
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4068 22568 4120 22574
rect 4068 22510 4120 22516
rect 4080 22409 4108 22510
rect 4066 22400 4122 22409
rect 4066 22335 4122 22344
rect 4172 21593 4200 23054
rect 4448 22778 4476 24686
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4526 23760 4582 23769
rect 4526 23695 4582 23704
rect 4540 23594 4568 23695
rect 4528 23588 4580 23594
rect 4528 23530 4580 23536
rect 4632 23322 4660 24142
rect 4724 23322 4752 24346
rect 4816 23526 4844 24550
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4804 23112 4856 23118
rect 4804 23054 4856 23060
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4448 22506 4476 22714
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 4816 22438 4844 23054
rect 4908 22556 4936 27520
rect 5552 25514 5580 27520
rect 5080 25492 5132 25498
rect 5552 25486 6040 25514
rect 5080 25434 5132 25440
rect 5092 25158 5120 25434
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5448 25220 5500 25226
rect 5448 25162 5500 25168
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 4988 22704 5040 22710
rect 4986 22672 4988 22681
rect 5040 22672 5042 22681
rect 4986 22607 5042 22616
rect 5092 22574 5120 25094
rect 5460 24886 5488 25162
rect 5448 24880 5500 24886
rect 5448 24822 5500 24828
rect 5460 24750 5488 24822
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 5354 24440 5410 24449
rect 5354 24375 5410 24384
rect 5368 24206 5396 24375
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5368 24070 5396 24142
rect 5552 24138 5580 25230
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24857 6040 25486
rect 5998 24848 6054 24857
rect 5998 24783 6054 24792
rect 6104 24342 6132 27520
rect 6656 25945 6684 27520
rect 6642 25936 6698 25945
rect 6642 25871 6698 25880
rect 7300 25498 7328 27520
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6552 24744 6604 24750
rect 6656 24721 6684 25094
rect 7300 24857 7328 25434
rect 7010 24848 7066 24857
rect 7286 24848 7342 24857
rect 7010 24783 7066 24792
rect 7104 24812 7156 24818
rect 7024 24750 7052 24783
rect 7286 24783 7288 24792
rect 7104 24754 7156 24760
rect 7340 24783 7342 24792
rect 7472 24812 7524 24818
rect 7288 24754 7340 24760
rect 7472 24754 7524 24760
rect 7012 24744 7064 24750
rect 6552 24686 6604 24692
rect 6642 24712 6698 24721
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 5540 24132 5592 24138
rect 5540 24074 5592 24080
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 6000 24064 6052 24070
rect 6104 24041 6132 24278
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6000 24006 6052 24012
rect 6090 24032 6146 24041
rect 5368 23798 5396 24006
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5354 23624 5410 23633
rect 5354 23559 5410 23568
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 5080 22568 5132 22574
rect 4908 22528 5028 22556
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4436 22160 4488 22166
rect 4436 22102 4488 22108
rect 4342 21992 4398 22001
rect 4342 21927 4398 21936
rect 4158 21584 4214 21593
rect 4158 21519 4214 21528
rect 4080 21078 4108 21109
rect 4068 21072 4120 21078
rect 4066 21040 4068 21049
rect 4120 21040 4122 21049
rect 4066 20975 4122 20984
rect 4160 21004 4212 21010
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3792 19236 3844 19242
rect 3792 19178 3844 19184
rect 3608 19168 3660 19174
rect 3606 19136 3608 19145
rect 3660 19136 3662 19145
rect 3606 19071 3662 19080
rect 3606 19000 3662 19009
rect 3606 18935 3662 18944
rect 3514 18728 3570 18737
rect 3514 18663 3570 18672
rect 3344 18278 3464 18306
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 2792 14980 3004 15008
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2792 13530 2820 14980
rect 2962 14920 3018 14929
rect 2962 14855 3018 14864
rect 2870 14784 2926 14793
rect 2870 14719 2926 14728
rect 2884 14414 2912 14719
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2884 14006 2912 14350
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 12918 2820 13330
rect 2688 12912 2740 12918
rect 2686 12880 2688 12889
rect 2780 12912 2832 12918
rect 2740 12880 2742 12889
rect 2780 12854 2832 12860
rect 2686 12815 2742 12824
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2608 12306 2636 12650
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11898 2820 12242
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2976 11801 3004 14855
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3068 13297 3096 13806
rect 3054 13288 3110 13297
rect 3054 13223 3110 13232
rect 3160 13190 3188 14418
rect 3240 14340 3292 14346
rect 3240 14282 3292 14288
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12889 3188 13126
rect 3146 12880 3202 12889
rect 3146 12815 3202 12824
rect 3146 12608 3202 12617
rect 3146 12543 3202 12552
rect 2962 11792 3018 11801
rect 2962 11727 3018 11736
rect 2410 10432 2466 10441
rect 2410 10367 2466 10376
rect 3160 9489 3188 12543
rect 3252 12442 3280 14282
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3344 12306 3372 18278
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3436 17882 3464 18158
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3436 17338 3464 17818
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3528 15745 3556 15914
rect 3514 15736 3570 15745
rect 3514 15671 3570 15680
rect 3528 15570 3556 15671
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3514 14512 3570 14521
rect 3514 14447 3570 14456
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3146 9480 3202 9489
rect 3146 9415 3202 9424
rect 2226 9072 2282 9081
rect 2226 9007 2282 9016
rect 3436 7562 3464 14010
rect 3528 13802 3556 14447
rect 3620 13870 3648 18935
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3528 13530 3556 13738
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3620 12986 3648 13670
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3620 12782 3648 12922
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3712 12628 3740 14758
rect 3804 14074 3832 19178
rect 3896 18902 3924 19246
rect 3884 18896 3936 18902
rect 3884 18838 3936 18844
rect 3882 18592 3938 18601
rect 3882 18527 3938 18536
rect 3896 17785 3924 18527
rect 3882 17776 3938 17785
rect 3882 17711 3938 17720
rect 3988 17105 4016 20334
rect 4080 20058 4108 20975
rect 4160 20946 4212 20952
rect 4172 20466 4200 20946
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4172 19922 4200 20402
rect 4252 20324 4304 20330
rect 4252 20266 4304 20272
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 4080 18578 4108 19382
rect 4080 18550 4200 18578
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4080 17882 4108 18362
rect 4172 18290 4200 18550
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4264 17270 4292 20266
rect 4356 18902 4384 21927
rect 4448 21865 4476 22102
rect 4528 22024 4580 22030
rect 4526 21992 4528 22001
rect 4580 21992 4582 22001
rect 4526 21927 4582 21936
rect 4434 21856 4490 21865
rect 4434 21791 4490 21800
rect 4448 21593 4476 21791
rect 4434 21584 4490 21593
rect 4434 21519 4490 21528
rect 4434 20632 4490 20641
rect 4540 20602 4568 21927
rect 4434 20567 4490 20576
rect 4528 20596 4580 20602
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4356 17882 4384 18838
rect 4448 18766 4476 20567
rect 4528 20538 4580 20544
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4540 19145 4568 19790
rect 4632 19174 4660 19926
rect 4620 19168 4672 19174
rect 4526 19136 4582 19145
rect 4620 19110 4672 19116
rect 4526 19071 4582 19080
rect 4632 18970 4660 19110
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4252 17264 4304 17270
rect 4252 17206 4304 17212
rect 4356 17134 4384 17818
rect 4448 17542 4476 18702
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4344 17128 4396 17134
rect 3974 17096 4030 17105
rect 4344 17070 4396 17076
rect 3974 17031 4030 17040
rect 4066 16960 4122 16969
rect 4066 16895 4122 16904
rect 3882 16688 3938 16697
rect 4080 16658 4108 16895
rect 4250 16824 4306 16833
rect 4356 16794 4384 17070
rect 4250 16759 4252 16768
rect 4304 16759 4306 16768
rect 4344 16788 4396 16794
rect 4252 16730 4304 16736
rect 4344 16730 4396 16736
rect 3882 16623 3884 16632
rect 3936 16623 3938 16632
rect 4068 16652 4120 16658
rect 3884 16594 3936 16600
rect 4068 16594 4120 16600
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3988 15434 4016 15846
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 3988 15026 4016 15370
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3896 13938 3924 14826
rect 3988 14618 4016 14962
rect 4080 14618 4108 16594
rect 4342 15464 4398 15473
rect 4342 15399 4344 15408
rect 4396 15399 4398 15408
rect 4344 15370 4396 15376
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4172 15162 4200 15302
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13530 4016 13670
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4356 12918 4384 15098
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 3620 12600 3740 12628
rect 3620 9489 3648 12600
rect 4448 11393 4476 17478
rect 4710 17368 4766 17377
rect 4710 17303 4712 17312
rect 4764 17303 4766 17312
rect 4712 17274 4764 17280
rect 4816 17270 4844 17614
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4540 14521 4568 16662
rect 4816 16590 4844 17206
rect 4896 16992 4948 16998
rect 5000 16969 5028 22528
rect 5080 22510 5132 22516
rect 5184 22234 5212 23122
rect 5262 22808 5318 22817
rect 5262 22743 5318 22752
rect 5276 22574 5304 22743
rect 5368 22642 5396 23559
rect 6012 23526 6040 24006
rect 6090 23967 6146 23976
rect 6380 23730 6408 24210
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5264 22568 5316 22574
rect 5264 22510 5316 22516
rect 5276 22234 5304 22510
rect 6196 22438 6224 23462
rect 6458 23352 6514 23361
rect 6458 23287 6514 23296
rect 6472 22778 6500 23287
rect 6460 22772 6512 22778
rect 6460 22714 6512 22720
rect 6184 22432 6236 22438
rect 6090 22400 6146 22409
rect 6184 22374 6236 22380
rect 6090 22335 6146 22344
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5184 22030 5212 22170
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5184 21690 5212 21966
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21690 6040 22102
rect 6104 22098 6132 22335
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6196 22030 6224 22374
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6090 21720 6146 21729
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 6000 21684 6052 21690
rect 6090 21655 6146 21664
rect 6000 21626 6052 21632
rect 6104 21570 6132 21655
rect 6012 21542 6132 21570
rect 6196 21554 6224 21966
rect 6184 21548 6236 21554
rect 6012 21457 6040 21542
rect 6184 21490 6236 21496
rect 5998 21448 6054 21457
rect 6564 21434 6592 24686
rect 7012 24686 7064 24692
rect 6642 24647 6698 24656
rect 6656 23050 6684 24647
rect 6736 24608 6788 24614
rect 6736 24550 6788 24556
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6748 21457 6776 24550
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6828 23316 6880 23322
rect 6932 23304 6960 24346
rect 7116 24138 7144 24754
rect 7300 24723 7328 24754
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7208 24177 7236 24550
rect 7484 24410 7512 24754
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7194 24168 7250 24177
rect 7104 24132 7156 24138
rect 7194 24103 7250 24112
rect 7104 24074 7156 24080
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7746 23488 7802 23497
rect 6880 23276 6960 23304
rect 6828 23258 6880 23264
rect 6840 22166 6868 23258
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 6932 22681 6960 22918
rect 6918 22672 6974 22681
rect 6918 22607 6974 22616
rect 7024 22545 7052 23462
rect 7010 22536 7066 22545
rect 7010 22471 7066 22480
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 5998 21383 6054 21392
rect 6104 21406 6592 21434
rect 6734 21448 6790 21457
rect 6000 21072 6052 21078
rect 5998 21040 6000 21049
rect 6052 21040 6054 21049
rect 5998 20975 6054 20984
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5460 20602 5488 20742
rect 5448 20596 5500 20602
rect 5448 20538 5500 20544
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5448 20256 5500 20262
rect 5552 20244 5580 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5500 20216 5580 20244
rect 5448 20198 5500 20204
rect 5184 19825 5212 20198
rect 5460 19922 5488 20198
rect 5998 19952 6054 19961
rect 5448 19916 5500 19922
rect 5368 19876 5448 19904
rect 5170 19816 5226 19825
rect 5170 19751 5226 19760
rect 5184 19514 5212 19751
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5368 19378 5396 19876
rect 5998 19887 6054 19896
rect 5448 19858 5500 19864
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5446 19544 5502 19553
rect 5552 19530 5580 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5502 19502 5580 19530
rect 5446 19479 5502 19488
rect 5538 19408 5594 19417
rect 5356 19372 5408 19378
rect 5538 19343 5594 19352
rect 5356 19314 5408 19320
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 5092 18698 5120 19110
rect 5368 18970 5396 19314
rect 5552 19310 5580 19343
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5552 18970 5580 19246
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 5092 18426 5120 18634
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 6012 18222 6040 19887
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 5816 18080 5868 18086
rect 5814 18048 5816 18057
rect 5868 18048 5870 18057
rect 5814 17983 5870 17992
rect 5080 17740 5132 17746
rect 5080 17682 5132 17688
rect 5092 17066 5120 17682
rect 5354 17640 5410 17649
rect 5354 17575 5410 17584
rect 5368 17338 5396 17575
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 4896 16934 4948 16940
rect 4986 16960 5042 16969
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4724 15094 4752 15506
rect 4816 15162 4844 15574
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4712 15088 4764 15094
rect 4712 15030 4764 15036
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4526 14512 4582 14521
rect 4526 14447 4582 14456
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4632 12442 4660 14418
rect 4724 14278 4752 14894
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4724 13977 4752 14214
rect 4710 13968 4766 13977
rect 4710 13903 4766 13912
rect 4908 13530 4936 16934
rect 4986 16895 5042 16904
rect 5092 16794 5120 17002
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5184 16674 5212 17002
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5092 16646 5212 16674
rect 4986 16552 5042 16561
rect 4986 16487 5042 16496
rect 5000 15502 5028 16487
rect 5092 15570 5120 16646
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15706 5212 15846
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5092 14482 5120 14758
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5184 14006 5212 14894
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 4988 13932 5040 13938
rect 4988 13874 5040 13880
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4816 12986 4844 13330
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4710 12472 4766 12481
rect 4620 12436 4672 12442
rect 4816 12442 4844 12922
rect 4710 12407 4766 12416
rect 4804 12436 4856 12442
rect 4620 12378 4672 12384
rect 4434 11384 4490 11393
rect 4434 11319 4490 11328
rect 4724 11121 4752 12407
rect 4804 12378 4856 12384
rect 4908 12374 4936 13466
rect 5000 12918 5028 13874
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 5184 11898 5212 13942
rect 5276 13326 5304 16730
rect 5460 16726 5488 17138
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5368 16250 5396 16526
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5460 16114 5488 16662
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15706 5488 16050
rect 5552 15910 5580 16934
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5552 15065 5580 15846
rect 6012 15570 6040 16186
rect 6104 15858 6132 21406
rect 6734 21383 6790 21392
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6196 18970 6224 21082
rect 6288 20602 6316 21082
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6380 20330 6408 21286
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6380 19922 6408 20266
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6380 19514 6408 19858
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6196 18290 6224 18770
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 6196 18057 6224 18226
rect 6368 18080 6420 18086
rect 6182 18048 6238 18057
rect 6368 18022 6420 18028
rect 6182 17983 6238 17992
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6196 16658 6224 17478
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6104 15830 6224 15858
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5538 15056 5594 15065
rect 5538 14991 5594 15000
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14618 5672 14758
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5828 14550 5856 14962
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5356 14408 5408 14414
rect 5354 14376 5356 14385
rect 5408 14376 5410 14385
rect 5354 14311 5410 14320
rect 5368 13530 5396 14311
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5460 13512 5488 14418
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5540 13524 5592 13530
rect 5460 13484 5540 13512
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12782 5304 13262
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5460 12424 5488 13484
rect 5540 13466 5592 13472
rect 5828 13462 5856 13874
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5630 12880 5686 12889
rect 6104 12850 6132 15642
rect 6196 12850 6224 15830
rect 6288 15638 6316 17274
rect 6380 16153 6408 18022
rect 6366 16144 6422 16153
rect 6366 16079 6422 16088
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6288 15162 6316 15574
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6288 13938 6316 15098
rect 6380 15026 6408 15574
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6380 14482 6408 14962
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6380 14074 6408 14418
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6288 12986 6316 13874
rect 6472 13530 6500 21286
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6826 20768 6882 20777
rect 6748 20534 6776 20742
rect 6826 20703 6882 20712
rect 6840 20602 6868 20703
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 6748 19718 6776 20470
rect 6840 20398 6868 20538
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6828 20256 6880 20262
rect 6932 20244 6960 20946
rect 7024 20505 7052 22374
rect 7010 20496 7066 20505
rect 7010 20431 7066 20440
rect 6880 20216 6960 20244
rect 6828 20198 6880 20204
rect 6826 20088 6882 20097
rect 6826 20023 6882 20032
rect 6840 19786 6868 20023
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6564 18358 6592 18770
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6564 16289 6592 18294
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6550 16280 6606 16289
rect 6550 16215 6606 16224
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6380 12986 6408 13330
rect 6552 13320 6604 13326
rect 6472 13280 6552 13308
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 5630 12815 5686 12824
rect 6092 12844 6144 12850
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5368 12396 5488 12424
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5368 11830 5396 12396
rect 5448 12300 5500 12306
rect 5552 12288 5580 12718
rect 5644 12442 5672 12815
rect 6092 12786 6144 12792
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6104 12714 6132 12786
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5500 12260 5580 12288
rect 6000 12300 6052 12306
rect 5448 12242 5500 12248
rect 6000 12242 6052 12248
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 4710 11112 4766 11121
rect 6012 11082 6040 12242
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11830 6316 12174
rect 6380 11830 6408 12242
rect 6472 11898 6500 13280
rect 6552 13262 6604 13268
rect 6656 12782 6684 18022
rect 6734 17912 6790 17921
rect 6734 17847 6736 17856
rect 6788 17847 6790 17856
rect 6736 17818 6788 17824
rect 6840 17762 6868 19722
rect 6932 18154 6960 20216
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7024 18970 7052 19110
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7024 18630 7052 18906
rect 7116 18850 7144 23462
rect 7746 23423 7802 23432
rect 7760 23254 7788 23423
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 7470 22944 7526 22953
rect 7470 22879 7526 22888
rect 7194 22808 7250 22817
rect 7194 22743 7250 22752
rect 7208 21486 7236 22743
rect 7196 21480 7248 21486
rect 7288 21480 7340 21486
rect 7196 21422 7248 21428
rect 7286 21448 7288 21457
rect 7340 21448 7342 21457
rect 7286 21383 7342 21392
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7300 20466 7328 20810
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7208 20058 7236 20198
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7208 18970 7236 19994
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19446 7328 19654
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7300 19174 7328 19246
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7116 18822 7236 18850
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 7116 17882 7144 18702
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 6748 17734 6868 17762
rect 7010 17776 7066 17785
rect 6748 15688 6776 17734
rect 7010 17711 7066 17720
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17338 6868 17614
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6748 15660 6868 15688
rect 6840 13954 6868 15660
rect 6932 14618 6960 17478
rect 7024 17338 7052 17711
rect 7208 17377 7236 18822
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 17814 7328 18566
rect 7392 18222 7420 21082
rect 7484 21078 7512 22879
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7576 21554 7604 21830
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7472 21072 7524 21078
rect 7472 21014 7524 21020
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7484 18902 7512 19314
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7470 18456 7526 18465
rect 7470 18391 7526 18400
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7288 17808 7340 17814
rect 7288 17750 7340 17756
rect 7378 17776 7434 17785
rect 7194 17368 7250 17377
rect 7012 17332 7064 17338
rect 7194 17303 7250 17312
rect 7012 17274 7064 17280
rect 7300 17066 7328 17750
rect 7378 17711 7434 17720
rect 7392 17338 7420 17711
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7392 17134 7420 17274
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 7010 16008 7066 16017
rect 7116 15978 7144 16526
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7010 15943 7066 15952
rect 7104 15972 7156 15978
rect 7024 15609 7052 15943
rect 7104 15914 7156 15920
rect 7010 15600 7066 15609
rect 7010 15535 7066 15544
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7024 14550 7052 15302
rect 7116 14890 7144 15914
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 6748 13926 6868 13954
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6748 12238 6776 13926
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13394 6960 13670
rect 7024 13530 7052 14486
rect 7102 13968 7158 13977
rect 7102 13903 7158 13912
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 7024 13326 7052 13466
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6644 12164 6696 12170
rect 6644 12106 6696 12112
rect 6656 11898 6684 12106
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6840 11354 6868 12922
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 12102 6960 12786
rect 7116 12442 7144 13903
rect 7208 13258 7236 15846
rect 7300 14249 7328 16390
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7484 15994 7512 18391
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7668 17649 7696 17682
rect 7760 17678 7788 21490
rect 7852 21078 7880 27520
rect 8024 25968 8076 25974
rect 8024 25910 8076 25916
rect 8036 25498 8064 25910
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8312 24750 8340 25230
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8116 24676 8168 24682
rect 8116 24618 8168 24624
rect 8128 24449 8156 24618
rect 8114 24440 8170 24449
rect 8114 24375 8116 24384
rect 8168 24375 8170 24384
rect 8116 24346 8168 24352
rect 8128 24315 8156 24346
rect 8312 24313 8340 24686
rect 8298 24304 8354 24313
rect 8116 24268 8168 24274
rect 8298 24239 8354 24248
rect 8116 24210 8168 24216
rect 8128 23866 8156 24210
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8024 23792 8076 23798
rect 8024 23734 8076 23740
rect 8036 22642 8064 23734
rect 8128 23594 8156 23802
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8128 23361 8156 23530
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8114 23352 8170 23361
rect 8220 23322 8248 23462
rect 8114 23287 8170 23296
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8312 23225 8340 24006
rect 8298 23216 8354 23225
rect 8298 23151 8354 23160
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 8116 22500 8168 22506
rect 8116 22442 8168 22448
rect 8128 21894 8156 22442
rect 8404 22030 8432 27520
rect 8760 25356 8812 25362
rect 8760 25298 8812 25304
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 8496 23798 8524 24686
rect 8772 24410 8800 25298
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 8852 24948 8904 24954
rect 8852 24890 8904 24896
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 8484 23792 8536 23798
rect 8484 23734 8536 23740
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8668 23520 8720 23526
rect 8666 23488 8668 23497
rect 8720 23488 8722 23497
rect 8666 23423 8722 23432
rect 8576 23316 8628 23322
rect 8576 23258 8628 23264
rect 8588 22234 8616 23258
rect 8666 23216 8722 23225
rect 8666 23151 8722 23160
rect 8680 23118 8708 23151
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8680 22778 8708 23054
rect 8772 22778 8800 23666
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8760 22772 8812 22778
rect 8760 22714 8812 22720
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8392 22024 8444 22030
rect 8298 21992 8354 22001
rect 8392 21966 8444 21972
rect 8298 21927 8354 21936
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 7930 21584 7986 21593
rect 7930 21519 7986 21528
rect 7944 21146 7972 21519
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7852 19990 7880 20878
rect 8128 20602 8156 21830
rect 8312 21690 8340 21927
rect 8300 21684 8352 21690
rect 8300 21626 8352 21632
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7852 19446 7880 19926
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7840 19304 7892 19310
rect 7838 19272 7840 19281
rect 7892 19272 7894 19281
rect 7838 19207 7894 19216
rect 7838 19000 7894 19009
rect 7838 18935 7840 18944
rect 7892 18935 7894 18944
rect 7840 18906 7892 18912
rect 7852 18290 7880 18906
rect 8024 18692 8076 18698
rect 8024 18634 8076 18640
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 8036 18086 8064 18634
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7748 17672 7800 17678
rect 7654 17640 7710 17649
rect 7748 17614 7800 17620
rect 7654 17575 7710 17584
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 16250 7604 17070
rect 7668 16794 7696 17575
rect 7746 17368 7802 17377
rect 7746 17303 7802 17312
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7286 14240 7342 14249
rect 7286 14175 7342 14184
rect 7392 14074 7420 15982
rect 7484 15966 7604 15994
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15745 7512 15846
rect 7470 15736 7526 15745
rect 7470 15671 7526 15680
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7392 13734 7420 14010
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7286 13288 7342 13297
rect 7196 13252 7248 13258
rect 7286 13223 7342 13232
rect 7196 13194 7248 13200
rect 7300 12850 7328 13223
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 4710 11047 4766 11056
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 3882 10432 3938 10441
rect 3882 10367 3938 10376
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3160 7534 3464 7562
rect 2962 6896 3018 6905
rect 2962 6831 3018 6840
rect 2976 6089 3004 6831
rect 2962 6080 3018 6089
rect 2962 6015 3018 6024
rect 3160 377 3188 7534
rect 3896 4865 3924 10367
rect 4080 10033 4108 10639
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 3974 9616 4030 9625
rect 3974 9551 4030 9560
rect 3988 8945 4016 9551
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 3974 8936 4030 8945
rect 3974 8871 4030 8880
rect 4080 7177 4108 9279
rect 6932 9217 6960 12038
rect 7300 11354 7328 12174
rect 7484 12170 7512 15671
rect 7576 12306 7604 15966
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7472 12164 7524 12170
rect 7472 12106 7524 12112
rect 7576 11898 7604 12242
rect 7668 12238 7696 16594
rect 7760 16436 7788 17303
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7852 16726 7880 17002
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7840 16720 7892 16726
rect 7944 16697 7972 16730
rect 7840 16662 7892 16668
rect 7930 16688 7986 16697
rect 7852 16561 7880 16662
rect 7930 16623 7986 16632
rect 7838 16552 7894 16561
rect 7838 16487 7894 16496
rect 7760 16408 7880 16436
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14385 7788 14758
rect 7746 14376 7802 14385
rect 7746 14311 7748 14320
rect 7800 14311 7802 14320
rect 7748 14282 7800 14288
rect 7852 13954 7880 16408
rect 7930 16280 7986 16289
rect 7930 16215 7986 16224
rect 7760 13926 7880 13954
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7760 11762 7788 13926
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 12617 7880 13806
rect 7838 12608 7894 12617
rect 7838 12543 7894 12552
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7944 11694 7972 16215
rect 8036 15609 8064 18022
rect 8022 15600 8078 15609
rect 8022 15535 8078 15544
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7944 11354 7972 11630
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 6918 9208 6974 9217
rect 6918 9143 6974 9152
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 8036 8265 8064 15535
rect 8128 14793 8156 20538
rect 8312 19417 8340 20742
rect 8588 20262 8616 20946
rect 8864 20913 8892 24890
rect 8956 23254 8984 25094
rect 9048 23474 9076 27520
rect 9402 25936 9458 25945
rect 9402 25871 9458 25880
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 9140 25158 9168 25230
rect 9128 25152 9180 25158
rect 9128 25094 9180 25100
rect 9140 24682 9168 25094
rect 9128 24676 9180 24682
rect 9128 24618 9180 24624
rect 9312 24200 9364 24206
rect 9312 24142 9364 24148
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23798 9168 24006
rect 9324 23866 9352 24142
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9324 23662 9352 23802
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9048 23446 9168 23474
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 8666 20904 8722 20913
rect 8666 20839 8668 20848
rect 8720 20839 8722 20848
rect 8850 20904 8906 20913
rect 8850 20839 8906 20848
rect 8668 20810 8720 20816
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8298 19408 8354 19417
rect 8298 19343 8354 19352
rect 8208 19168 8260 19174
rect 8588 19122 8616 20198
rect 8680 19854 8708 20334
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8772 20058 8800 20266
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8680 19514 8708 19790
rect 8772 19786 8800 19994
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8760 19780 8812 19786
rect 8760 19722 8812 19728
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8864 19174 8892 19858
rect 8942 19408 8998 19417
rect 8942 19343 8998 19352
rect 8260 19116 8616 19122
rect 8208 19110 8616 19116
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8220 19094 8616 19110
rect 8588 18193 8616 19094
rect 8760 18896 8812 18902
rect 8758 18864 8760 18873
rect 8812 18864 8814 18873
rect 8758 18799 8814 18808
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8680 18290 8708 18566
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8574 18184 8630 18193
rect 8574 18119 8630 18128
rect 8208 18080 8260 18086
rect 8576 18080 8628 18086
rect 8208 18022 8260 18028
rect 8298 18048 8354 18057
rect 8220 17882 8248 18022
rect 8576 18022 8628 18028
rect 8298 17983 8354 17992
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8206 16960 8262 16969
rect 8206 16895 8262 16904
rect 8114 14784 8170 14793
rect 8114 14719 8170 14728
rect 8220 14090 8248 16895
rect 8312 16794 8340 17983
rect 8588 17542 8616 18022
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 17134 8616 17478
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8300 16788 8352 16794
rect 8352 16748 8432 16776
rect 8300 16730 8352 16736
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8312 15502 8340 16458
rect 8404 16250 8432 16748
rect 8588 16590 8616 16934
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8588 15706 8616 16526
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8680 15570 8708 18226
rect 8864 16561 8892 19110
rect 8850 16552 8906 16561
rect 8850 16487 8906 16496
rect 8864 15881 8892 16487
rect 8850 15872 8906 15881
rect 8850 15807 8906 15816
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8772 15609 8800 15642
rect 8758 15600 8814 15609
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8668 15564 8720 15570
rect 8758 15535 8814 15544
rect 8668 15506 8720 15512
rect 8300 15496 8352 15502
rect 8298 15464 8300 15473
rect 8352 15464 8354 15473
rect 8298 15399 8354 15408
rect 8220 14062 8340 14090
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8128 13530 8156 13874
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8114 13424 8170 13433
rect 8114 13359 8116 13368
rect 8168 13359 8170 13368
rect 8116 13330 8168 13336
rect 8114 13254 8170 13263
rect 8114 13189 8170 13198
rect 8128 12782 8156 13189
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8220 12424 8248 13942
rect 8312 13394 8340 14062
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8312 12986 8340 13330
rect 8496 12986 8524 13466
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8300 12436 8352 12442
rect 8220 12396 8300 12424
rect 8300 12378 8352 12384
rect 8588 12170 8616 15506
rect 8850 15056 8906 15065
rect 8850 14991 8906 15000
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8680 13938 8708 14418
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13938 8800 14214
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8666 13560 8722 13569
rect 8666 13495 8722 13504
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11626 8340 12038
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8390 11384 8446 11393
rect 8390 11319 8446 11328
rect 8484 11348 8536 11354
rect 8404 11218 8432 11319
rect 8484 11290 8536 11296
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8404 11098 8432 11154
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8220 11070 8432 11098
rect 8128 10810 8156 11018
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8220 10674 8248 11070
rect 8496 10810 8524 11290
rect 8588 11150 8616 11698
rect 8680 11218 8708 13495
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8772 12986 8800 13262
rect 8864 12986 8892 14991
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8956 11354 8984 19343
rect 9048 18154 9076 21966
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 9048 16658 9076 18090
rect 9140 17746 9168 23446
rect 9416 21554 9444 25871
rect 9600 25838 9628 27520
rect 10048 26036 10100 26042
rect 10048 25978 10100 25984
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9600 25362 9628 25774
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9600 24562 9628 24618
rect 9864 24608 9916 24614
rect 9600 24534 9812 24562
rect 10060 24585 10088 25978
rect 10046 24576 10102 24585
rect 9864 24550 9916 24556
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9508 22234 9536 22986
rect 9784 22574 9812 24534
rect 9876 24410 9904 24550
rect 9968 24534 10046 24562
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9876 23662 9904 24346
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9876 23050 9904 23598
rect 9864 23044 9916 23050
rect 9864 22986 9916 22992
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9784 22001 9812 22374
rect 9586 21992 9642 22001
rect 9586 21927 9642 21936
rect 9770 21992 9826 22001
rect 9770 21927 9826 21936
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9220 21344 9272 21350
rect 9220 21286 9272 21292
rect 9232 20942 9260 21286
rect 9416 21146 9444 21490
rect 9600 21418 9628 21927
rect 9588 21412 9640 21418
rect 9588 21354 9640 21360
rect 9772 21344 9824 21350
rect 9772 21286 9824 21292
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9678 20088 9734 20097
rect 9678 20023 9734 20032
rect 9692 19990 9720 20023
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9232 19310 9260 19858
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9324 19446 9352 19654
rect 9692 19514 9720 19790
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 16658 9168 17682
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 9048 15065 9076 15370
rect 9034 15056 9090 15065
rect 9034 14991 9090 15000
rect 9140 14362 9168 16594
rect 9232 14822 9260 19246
rect 9324 17882 9352 19382
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9496 19304 9548 19310
rect 9600 19281 9628 19314
rect 9496 19246 9548 19252
rect 9586 19272 9642 19281
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9416 18601 9444 19110
rect 9508 18698 9536 19246
rect 9586 19207 9642 19216
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9402 18592 9458 18601
rect 9402 18527 9458 18536
rect 9508 18222 9536 18634
rect 9600 18426 9628 19207
rect 9678 19136 9734 19145
rect 9678 19071 9734 19080
rect 9692 18902 9720 19071
rect 9680 18896 9732 18902
rect 9680 18838 9732 18844
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9692 17898 9720 18702
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9416 17870 9720 17898
rect 9416 17542 9444 17870
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9416 17241 9444 17478
rect 9402 17232 9458 17241
rect 9402 17167 9458 17176
rect 9404 17128 9456 17134
rect 9692 17105 9720 17478
rect 9404 17070 9456 17076
rect 9678 17096 9734 17105
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9048 14334 9168 14362
rect 9048 13530 9076 14334
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9034 13152 9090 13161
rect 9034 13087 9090 13096
rect 9048 11898 9076 13087
rect 9126 12744 9182 12753
rect 9126 12679 9128 12688
rect 9180 12679 9182 12688
rect 9128 12650 9180 12656
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9232 11762 9260 14758
rect 9416 13530 9444 17070
rect 9678 17031 9734 17040
rect 9680 16992 9732 16998
rect 9678 16960 9680 16969
rect 9732 16960 9734 16969
rect 9678 16895 9734 16904
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9508 15706 9536 16526
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9600 14618 9628 15574
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9508 14074 9536 14350
rect 9588 14272 9640 14278
rect 9586 14240 9588 14249
rect 9640 14240 9642 14249
rect 9586 14175 9642 14184
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9508 13870 9536 14010
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9416 13326 9444 13466
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12850 9444 13262
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9494 12744 9550 12753
rect 9494 12679 9550 12688
rect 9588 12708 9640 12714
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11354 9352 11698
rect 9508 11694 9536 12679
rect 9588 12650 9640 12656
rect 9496 11688 9548 11694
rect 9402 11656 9458 11665
rect 9496 11630 9548 11636
rect 9402 11591 9458 11600
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9218 11248 9274 11257
rect 8668 11212 8720 11218
rect 9416 11234 9444 11591
rect 9218 11183 9274 11192
rect 9324 11206 9444 11234
rect 8668 11154 8720 11160
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 9232 10810 9260 11183
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9324 10674 9352 11206
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 10266 9352 10610
rect 9600 10606 9628 12650
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 10810 9720 11562
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9588 10124 9640 10130
rect 9692 10112 9720 10406
rect 9640 10084 9720 10112
rect 9588 10066 9640 10072
rect 9692 9654 9720 10084
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 7562 8256 7618 8265
rect 7562 8191 7618 8200
rect 8022 8256 8078 8265
rect 8022 8191 8078 8200
rect 7576 7721 7604 8191
rect 7562 7712 7618 7721
rect 5622 7644 5918 7664
rect 7562 7647 7618 7656
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 9784 7449 9812 21286
rect 9876 21026 9904 22374
rect 9968 22234 9996 24534
rect 10046 24511 10102 24520
rect 10152 23769 10180 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10690 25528 10746 25537
rect 10612 25472 10690 25480
rect 10612 25463 10746 25472
rect 10612 25452 10732 25463
rect 10612 25226 10640 25452
rect 10692 25356 10744 25362
rect 10692 25298 10744 25304
rect 10600 25220 10652 25226
rect 10600 25162 10652 25168
rect 10704 24954 10732 25298
rect 10692 24948 10744 24954
rect 10692 24890 10744 24896
rect 10690 24712 10746 24721
rect 10690 24647 10746 24656
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 24410 10732 24647
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10796 24138 10824 27520
rect 10968 25764 11020 25770
rect 10968 25706 11020 25712
rect 10980 25498 11008 25706
rect 11348 25514 11376 27520
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 11256 25486 11376 25514
rect 10966 25256 11022 25265
rect 10966 25191 10968 25200
rect 11020 25191 11022 25200
rect 10968 25162 11020 25168
rect 11150 24848 11206 24857
rect 11150 24783 11206 24792
rect 11164 24410 11192 24783
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 10876 24336 10928 24342
rect 10876 24278 10928 24284
rect 10888 24177 10916 24278
rect 10874 24168 10930 24177
rect 10784 24132 10836 24138
rect 10874 24103 10930 24112
rect 10784 24074 10836 24080
rect 10138 23760 10194 23769
rect 10138 23695 10194 23704
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10060 22710 10088 23122
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 10060 22166 10088 22646
rect 10796 22506 10824 24074
rect 10888 23322 10916 24103
rect 11164 23848 11192 24346
rect 11256 24342 11284 25486
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11426 24848 11482 24857
rect 11426 24783 11482 24792
rect 11244 24336 11296 24342
rect 11440 24313 11468 24783
rect 11624 24682 11652 25230
rect 11612 24676 11664 24682
rect 11612 24618 11664 24624
rect 11520 24608 11572 24614
rect 11518 24576 11520 24585
rect 11572 24576 11574 24585
rect 11518 24511 11574 24520
rect 11716 24392 11744 25638
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11808 24410 11836 25298
rect 11624 24364 11744 24392
rect 11796 24404 11848 24410
rect 11244 24278 11296 24284
rect 11426 24304 11482 24313
rect 11426 24239 11482 24248
rect 11518 24032 11574 24041
rect 11518 23967 11574 23976
rect 11072 23820 11192 23848
rect 10966 23488 11022 23497
rect 10966 23423 11022 23432
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10980 22642 11008 23423
rect 11072 23322 11100 23820
rect 11532 23798 11560 23967
rect 11520 23792 11572 23798
rect 11520 23734 11572 23740
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11164 23225 11192 23462
rect 11150 23216 11206 23225
rect 11426 23216 11482 23225
rect 11150 23151 11206 23160
rect 11336 23180 11388 23186
rect 11532 23186 11560 23530
rect 11426 23151 11482 23160
rect 11520 23180 11572 23186
rect 11336 23122 11388 23128
rect 11348 22778 11376 23122
rect 11336 22772 11388 22778
rect 11164 22732 11336 22760
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10968 22500 11020 22506
rect 10968 22442 11020 22448
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10980 22234 11008 22442
rect 10140 22228 10192 22234
rect 10968 22228 11020 22234
rect 10192 22188 10272 22216
rect 10140 22170 10192 22176
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 10244 21690 10272 22188
rect 10612 22166 10640 22197
rect 10968 22170 11020 22176
rect 10600 22160 10652 22166
rect 10598 22128 10600 22137
rect 10652 22128 10654 22137
rect 10598 22063 10654 22072
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10520 21593 10548 21966
rect 10612 21690 10640 22063
rect 11164 22030 11192 22732
rect 11336 22714 11388 22720
rect 11334 22672 11390 22681
rect 11334 22607 11390 22616
rect 11348 22098 11376 22607
rect 11440 22545 11468 23151
rect 11520 23122 11572 23128
rect 11426 22536 11482 22545
rect 11426 22471 11482 22480
rect 11624 22114 11652 24364
rect 11796 24346 11848 24352
rect 11900 24290 11928 27520
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11992 24750 12020 25094
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11716 24262 11928 24290
rect 11716 22953 11744 24262
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11808 24041 11836 24142
rect 11794 24032 11850 24041
rect 11794 23967 11850 23976
rect 11808 23866 11836 23967
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11808 23254 11836 23802
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 11796 23248 11848 23254
rect 11796 23190 11848 23196
rect 11702 22944 11758 22953
rect 11702 22879 11758 22888
rect 11808 22778 11836 23190
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11336 22092 11388 22098
rect 11624 22086 11735 22114
rect 11707 22080 11735 22086
rect 11707 22052 11744 22080
rect 11336 22034 11388 22040
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10600 21684 10652 21690
rect 10652 21644 10824 21672
rect 10600 21626 10652 21632
rect 10506 21584 10562 21593
rect 9956 21548 10008 21554
rect 10506 21519 10508 21528
rect 9956 21490 10008 21496
rect 10560 21519 10562 21528
rect 10508 21490 10560 21496
rect 9968 21146 9996 21490
rect 10520 21459 10548 21490
rect 10046 21312 10102 21321
rect 10046 21247 10102 21256
rect 10060 21146 10088 21247
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 9876 20998 9996 21026
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9876 18766 9904 19314
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9862 18592 9918 18601
rect 9862 18527 9918 18536
rect 9876 16658 9904 18527
rect 9968 17785 9996 20998
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10138 19000 10194 19009
rect 10289 18992 10585 19012
rect 10138 18935 10194 18944
rect 10152 18222 10180 18935
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9954 17776 10010 17785
rect 9954 17711 10010 17720
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9968 16538 9996 17070
rect 10060 17066 10088 18022
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10152 16572 10180 18158
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10244 17066 10272 17614
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10232 16584 10284 16590
rect 10152 16544 10232 16572
rect 9876 16510 9996 16538
rect 10232 16526 10284 16532
rect 9876 12646 9904 16510
rect 10244 16250 10272 16526
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10138 15736 10194 15745
rect 10289 15728 10585 15748
rect 10138 15671 10194 15680
rect 10152 15502 10180 15671
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9956 15428 10008 15434
rect 9956 15370 10008 15376
rect 9968 14249 9996 15370
rect 10152 15162 10180 15438
rect 10140 15156 10192 15162
rect 10060 15116 10140 15144
rect 9954 14240 10010 14249
rect 9954 14175 10010 14184
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9968 12986 9996 13262
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9876 12442 9904 12582
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9864 9376 9916 9382
rect 9862 9344 9864 9353
rect 9916 9344 9918 9353
rect 9862 9279 9918 9288
rect 9968 8022 9996 12718
rect 10060 12481 10088 15116
rect 10140 15098 10192 15104
rect 10598 14920 10654 14929
rect 10598 14855 10600 14864
rect 10652 14855 10654 14864
rect 10600 14826 10652 14832
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10152 14521 10180 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10138 14512 10194 14521
rect 10138 14447 10194 14456
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10046 12472 10102 12481
rect 10046 12407 10102 12416
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11898 10088 12242
rect 10152 12238 10180 13806
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 19110
rect 10796 17882 10824 21644
rect 10888 21010 10916 21830
rect 11058 21720 11114 21729
rect 11164 21690 11192 21966
rect 11058 21655 11114 21664
rect 11152 21684 11204 21690
rect 11072 21321 11100 21655
rect 11152 21626 11204 21632
rect 11348 21554 11376 22034
rect 11336 21548 11388 21554
rect 11336 21490 11388 21496
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11058 21312 11114 21321
rect 11058 21247 11114 21256
rect 11256 21146 11284 21422
rect 11610 21312 11666 21321
rect 11610 21247 11666 21256
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 10968 21072 11020 21078
rect 10966 21040 10968 21049
rect 11020 21040 11022 21049
rect 10876 21004 10928 21010
rect 10966 20975 11022 20984
rect 10876 20946 10928 20952
rect 10888 20641 10916 20946
rect 10874 20632 10930 20641
rect 10980 20602 11008 20975
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 10874 20567 10930 20576
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10876 20392 10928 20398
rect 10874 20360 10876 20369
rect 10928 20360 10930 20369
rect 10874 20295 10930 20304
rect 11060 20256 11112 20262
rect 10874 20224 10930 20233
rect 11060 20198 11112 20204
rect 10874 20159 10930 20168
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10796 17134 10824 17818
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10796 16833 10824 16934
rect 10782 16824 10838 16833
rect 10782 16759 10838 16768
rect 10888 16726 10916 20159
rect 11072 19417 11100 20198
rect 11058 19408 11114 19417
rect 11058 19343 11114 19352
rect 11164 19310 11192 20810
rect 11520 20800 11572 20806
rect 11518 20768 11520 20777
rect 11572 20768 11574 20777
rect 11518 20703 11574 20712
rect 11624 19938 11652 21247
rect 11716 21010 11744 22052
rect 11808 21146 11836 22714
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 11704 21004 11756 21010
rect 11704 20946 11756 20952
rect 11716 20602 11744 20946
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11624 19910 11836 19938
rect 11612 19848 11664 19854
rect 11610 19816 11612 19825
rect 11664 19816 11666 19825
rect 11610 19751 11666 19760
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11152 19168 11204 19174
rect 11150 19136 11152 19145
rect 11204 19136 11206 19145
rect 11150 19071 11206 19080
rect 11164 18970 11192 19071
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 10980 16810 11008 18770
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 17814 11100 18702
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 11164 17542 11192 18770
rect 11244 18760 11296 18766
rect 11242 18728 11244 18737
rect 11428 18760 11480 18766
rect 11296 18728 11298 18737
rect 11428 18702 11480 18708
rect 11242 18663 11298 18672
rect 11440 18068 11468 18702
rect 11520 18080 11572 18086
rect 11440 18040 11520 18068
rect 11520 18022 11572 18028
rect 11532 17746 11560 18022
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 10980 16782 11100 16810
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 11072 16658 11100 16782
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10968 16584 11020 16590
rect 11164 16538 11192 17478
rect 11348 17218 11376 17614
rect 11532 17338 11560 17682
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11426 17232 11482 17241
rect 11348 17190 11426 17218
rect 11426 17167 11428 17176
rect 11480 17167 11482 17176
rect 11428 17138 11480 17144
rect 11440 16794 11468 17138
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11532 16674 11560 17274
rect 11808 17116 11836 19910
rect 11900 17218 11928 23462
rect 11992 20505 12020 24686
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12072 24336 12124 24342
rect 12072 24278 12124 24284
rect 12084 23798 12112 24278
rect 12072 23792 12124 23798
rect 12070 23760 12072 23769
rect 12124 23760 12126 23769
rect 12070 23695 12126 23704
rect 12070 22536 12126 22545
rect 12070 22471 12126 22480
rect 12084 21146 12112 22471
rect 12176 21894 12204 24618
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23905 12296 24006
rect 12254 23896 12310 23905
rect 12254 23831 12310 23840
rect 12438 22944 12494 22953
rect 12438 22879 12494 22888
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12268 21690 12296 22102
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 11978 20496 12034 20505
rect 11978 20431 12034 20440
rect 12084 20262 12112 20878
rect 12176 20466 12204 21558
rect 12360 21418 12388 22374
rect 12452 22273 12480 22879
rect 12438 22264 12494 22273
rect 12438 22199 12494 22208
rect 12544 22114 12572 27520
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12728 24886 12756 25230
rect 13004 24954 13032 25298
rect 12992 24948 13044 24954
rect 12992 24890 13044 24896
rect 12716 24880 12768 24886
rect 13096 24834 13124 27520
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 12716 24822 12768 24828
rect 12728 24721 12756 24822
rect 12820 24806 13124 24834
rect 13188 24818 13216 25230
rect 13176 24812 13228 24818
rect 12714 24712 12770 24721
rect 12714 24647 12770 24656
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12728 23866 12756 24210
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12716 22432 12768 22438
rect 12714 22400 12716 22409
rect 12768 22400 12770 22409
rect 12714 22335 12770 22344
rect 12544 22086 12664 22114
rect 12636 22080 12664 22086
rect 12636 22052 12756 22080
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12452 21486 12480 21898
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12544 21298 12572 21830
rect 12624 21480 12676 21486
rect 12622 21448 12624 21457
rect 12676 21448 12678 21457
rect 12622 21383 12678 21392
rect 12544 21270 12664 21298
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12084 19990 12112 20198
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 12084 19689 12112 19926
rect 12176 19922 12204 20402
rect 12636 20330 12664 21270
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12636 20058 12664 20266
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12070 19680 12126 19689
rect 12070 19615 12126 19624
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 17814 12112 18566
rect 12176 17814 12204 19178
rect 12360 18306 12388 19314
rect 12636 18737 12664 19790
rect 12622 18728 12678 18737
rect 12622 18663 12678 18672
rect 12622 18456 12678 18465
rect 12532 18420 12584 18426
rect 12728 18442 12756 22052
rect 12678 18414 12756 18442
rect 12622 18391 12678 18400
rect 12532 18362 12584 18368
rect 12544 18329 12572 18362
rect 12728 18358 12756 18414
rect 12716 18352 12768 18358
rect 12530 18320 12586 18329
rect 12360 18278 12480 18306
rect 12452 17882 12480 18278
rect 12716 18294 12768 18300
rect 12530 18255 12586 18264
rect 12728 18222 12756 18294
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 12084 17338 12112 17750
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 11900 17190 12020 17218
rect 11808 17088 11928 17116
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11440 16646 11560 16674
rect 11702 16688 11758 16697
rect 11020 16532 11192 16538
rect 10968 16526 11192 16532
rect 10980 16510 11192 16526
rect 10874 16280 10930 16289
rect 10874 16215 10930 16224
rect 10782 15872 10838 15881
rect 10782 15807 10838 15816
rect 10796 15706 10824 15807
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10888 15638 10916 16215
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10980 15745 11008 15914
rect 10966 15736 11022 15745
rect 10966 15671 10968 15680
rect 11020 15671 11022 15680
rect 10968 15642 11020 15648
rect 10876 15632 10928 15638
rect 11072 15586 11100 16510
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 10876 15574 10928 15580
rect 10980 15570 11100 15586
rect 10968 15564 11100 15570
rect 11020 15558 11100 15564
rect 10968 15506 11020 15512
rect 11072 15473 11100 15558
rect 11058 15464 11114 15473
rect 11058 15399 11114 15408
rect 10782 15328 10838 15337
rect 10782 15263 10838 15272
rect 10796 15162 10824 15263
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 11256 14482 11284 15846
rect 11348 15094 11376 16594
rect 11440 16590 11468 16646
rect 11702 16623 11704 16632
rect 11756 16623 11758 16632
rect 11704 16594 11756 16600
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11440 16046 11468 16526
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11440 15570 11468 15982
rect 11716 15706 11744 16594
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11440 15162 11468 15506
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11532 15026 11560 15506
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13870 11100 14214
rect 11256 14074 11284 14418
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10782 13560 10838 13569
rect 10692 13524 10744 13530
rect 10782 13495 10838 13504
rect 10692 13466 10744 13472
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12306 10732 12922
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10060 11286 10088 11834
rect 10152 11354 10180 12174
rect 10796 11898 10824 13495
rect 10980 13394 11008 13670
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10980 12986 11008 13330
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10046 11112 10102 11121
rect 10046 11047 10102 11056
rect 10060 10266 10088 11047
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10152 10441 10180 10474
rect 10138 10432 10194 10441
rect 10138 10367 10194 10376
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10692 10192 10744 10198
rect 10046 10160 10102 10169
rect 10692 10134 10744 10140
rect 10046 10095 10102 10104
rect 10060 9518 10088 10095
rect 10704 9586 10732 10134
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 9178 10088 9454
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 9956 8016 10008 8022
rect 10796 7993 10824 11698
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10062 10916 10950
rect 10980 10266 11008 12922
rect 11072 11762 11100 13466
rect 11164 12714 11192 13738
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11348 12374 11376 13126
rect 11440 12889 11468 14758
rect 11532 14618 11560 14962
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11808 14550 11836 15098
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11426 12880 11482 12889
rect 11426 12815 11482 12824
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11426 12200 11482 12209
rect 11426 12135 11428 12144
rect 11480 12135 11482 12144
rect 11428 12106 11480 12112
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11150 11792 11206 11801
rect 11060 11756 11112 11762
rect 11256 11762 11284 12038
rect 11440 11762 11468 12106
rect 11532 11898 11560 12242
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11150 11727 11206 11736
rect 11244 11756 11296 11762
rect 11060 11698 11112 11704
rect 11164 11694 11192 11727
rect 11244 11698 11296 11704
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11256 11354 11284 11698
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11244 11212 11296 11218
rect 11348 11200 11376 11494
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11296 11172 11376 11200
rect 11244 11154 11296 11160
rect 11256 10674 11284 11154
rect 11440 11150 11468 11222
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11440 10470 11468 11086
rect 11624 10674 11652 12582
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11702 12064 11758 12073
rect 11702 11999 11758 12008
rect 11716 11150 11744 11999
rect 11808 11665 11836 12242
rect 11794 11656 11850 11665
rect 11794 11591 11796 11600
rect 11848 11591 11850 11600
rect 11796 11562 11848 11568
rect 11900 11286 11928 17088
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10980 9178 11008 10066
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11072 9466 11100 9998
rect 11164 9722 11192 9998
rect 11440 9761 11468 10406
rect 11624 10266 11652 10610
rect 11808 10470 11836 11154
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11426 9752 11482 9761
rect 11152 9716 11204 9722
rect 11426 9687 11482 9696
rect 11152 9658 11204 9664
rect 11072 9438 11192 9466
rect 11164 9382 11192 9438
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11716 8362 11744 8910
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 9956 7958 10008 7964
rect 10782 7984 10838 7993
rect 10782 7919 10838 7928
rect 9770 7440 9826 7449
rect 9770 7375 9826 7384
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 4066 5400 4122 5409
rect 5622 5392 5918 5412
rect 4066 5335 4122 5344
rect 3882 4856 3938 4865
rect 3882 4791 3938 4800
rect 4080 4593 4108 5335
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 3974 4040 4030 4049
rect 3974 3975 4030 3984
rect 3330 3632 3386 3641
rect 3330 3567 3386 3576
rect 3344 921 3372 3567
rect 3988 3233 4016 3975
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 4066 3768 4122 3777
rect 10289 3760 10585 3780
rect 4066 3703 4122 3712
rect 3974 3224 4030 3233
rect 3974 3159 4030 3168
rect 4080 3097 4108 3703
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 4066 3088 4122 3097
rect 4066 3023 4122 3032
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 3514 2680 3570 2689
rect 10289 2672 10585 2692
rect 3514 2615 3570 2624
rect 3528 1601 3556 2615
rect 11716 2553 11744 8298
rect 11702 2544 11758 2553
rect 11702 2479 11758 2488
rect 4618 2408 4674 2417
rect 4618 2343 4674 2352
rect 3514 1592 3570 1601
rect 3514 1527 3570 1536
rect 3330 912 3386 921
rect 3330 847 3386 856
rect 4632 480 4660 2343
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 11808 1601 11836 10406
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 8090 11928 9318
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7206 11928 7890
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 3641 11928 7142
rect 11886 3632 11942 3641
rect 11886 3567 11942 3576
rect 11992 3505 12020 17190
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 15570 12112 16390
rect 12452 16250 12480 17070
rect 12820 17066 12848 24806
rect 13176 24754 13228 24760
rect 12900 24676 12952 24682
rect 12900 24618 12952 24624
rect 12912 22817 12940 24618
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 13004 23730 13032 24006
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12990 23352 13046 23361
rect 13188 23322 13216 24754
rect 12990 23287 13046 23296
rect 13176 23316 13228 23322
rect 12898 22808 12954 22817
rect 12898 22743 12954 22752
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15745 12848 16050
rect 12806 15736 12862 15745
rect 12806 15671 12808 15680
rect 12860 15671 12862 15680
rect 12808 15642 12860 15648
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 12912 15065 12940 16934
rect 12898 15056 12954 15065
rect 12898 14991 12954 15000
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12084 13190 12112 14418
rect 12162 14376 12218 14385
rect 12162 14311 12218 14320
rect 12346 14376 12402 14385
rect 12346 14311 12348 14320
rect 12176 14074 12204 14311
rect 12400 14311 12402 14320
rect 12348 14282 12400 14288
rect 12636 14278 12664 14758
rect 13004 14482 13032 23287
rect 13176 23258 13228 23264
rect 13188 22166 13216 23258
rect 13176 22160 13228 22166
rect 13176 22102 13228 22108
rect 13174 20904 13230 20913
rect 13174 20839 13230 20848
rect 13188 19718 13216 20839
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13096 19174 13124 19246
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13096 17377 13124 19110
rect 13082 17368 13138 17377
rect 13280 17338 13308 25842
rect 13648 25106 13676 27520
rect 14292 25650 14320 27520
rect 14844 26042 14872 27520
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14922 25800 14978 25809
rect 14922 25735 14978 25744
rect 13556 25078 13676 25106
rect 14108 25622 14320 25650
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13372 24614 13400 24890
rect 13360 24608 13412 24614
rect 13556 24562 13584 25078
rect 13820 24880 13872 24886
rect 13360 24550 13412 24556
rect 13464 24534 13584 24562
rect 13648 24828 13820 24834
rect 13648 24822 13872 24828
rect 13910 24848 13966 24857
rect 13648 24806 13860 24822
rect 13464 23497 13492 24534
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13450 23488 13506 23497
rect 13450 23423 13506 23432
rect 13556 22982 13584 23530
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22681 13584 22918
rect 13542 22672 13598 22681
rect 13542 22607 13598 22616
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13358 21584 13414 21593
rect 13358 21519 13414 21528
rect 13372 21486 13400 21519
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13372 21146 13400 21422
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13464 20777 13492 22374
rect 13556 21690 13584 22374
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 13648 21146 13676 24806
rect 13910 24783 13966 24792
rect 13726 24712 13782 24721
rect 13726 24647 13782 24656
rect 13740 24614 13768 24647
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13924 24449 13952 24783
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 13910 24440 13966 24449
rect 13910 24375 13966 24384
rect 13728 24200 13780 24206
rect 13726 24168 13728 24177
rect 13780 24168 13782 24177
rect 13726 24103 13782 24112
rect 14016 24041 14044 24550
rect 14002 24032 14058 24041
rect 14002 23967 14058 23976
rect 14016 23866 14044 23967
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13820 22500 13872 22506
rect 13820 22442 13872 22448
rect 13832 21894 13860 22442
rect 13924 22030 13952 23122
rect 14108 23089 14136 25622
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14370 24848 14426 24857
rect 14370 24783 14426 24792
rect 14094 23080 14150 23089
rect 14094 23015 14150 23024
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22545 14320 22918
rect 14278 22536 14334 22545
rect 14278 22471 14334 22480
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13832 21350 13860 21830
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13832 21049 13860 21286
rect 13818 21040 13874 21049
rect 13818 20975 13874 20984
rect 13634 20904 13690 20913
rect 13544 20868 13596 20874
rect 13924 20890 13952 21966
rect 14384 21962 14412 24783
rect 14476 24070 14504 25298
rect 14936 25140 14964 25735
rect 14660 25112 14964 25140
rect 15292 25152 15344 25158
rect 14660 24410 14688 25112
rect 15292 25094 15344 25100
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15304 24886 15332 25094
rect 15292 24880 15344 24886
rect 15292 24822 15344 24828
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 13924 20862 14228 20890
rect 13634 20839 13690 20848
rect 13544 20810 13596 20816
rect 13450 20768 13506 20777
rect 13450 20703 13506 20712
rect 13556 20058 13584 20810
rect 13648 20058 13676 20839
rect 14094 20768 14150 20777
rect 14094 20703 14150 20712
rect 13912 20256 13964 20262
rect 13912 20198 13964 20204
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13464 19310 13492 19654
rect 13648 19514 13676 19858
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13452 19304 13504 19310
rect 13358 19272 13414 19281
rect 13452 19246 13504 19252
rect 13358 19207 13414 19216
rect 13372 18970 13400 19207
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13082 17303 13138 17312
rect 13268 17332 13320 17338
rect 13096 14532 13124 17303
rect 13268 17274 13320 17280
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13266 15464 13322 15473
rect 13266 15399 13322 15408
rect 13280 15026 13308 15399
rect 13372 15366 13400 15846
rect 13360 15360 13412 15366
rect 13358 15328 13360 15337
rect 13412 15328 13414 15337
rect 13358 15263 13414 15272
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13188 14657 13216 14894
rect 13174 14648 13230 14657
rect 13280 14618 13308 14962
rect 13464 14958 13492 19246
rect 13648 18426 13676 19450
rect 13832 19258 13860 19790
rect 13740 19242 13860 19258
rect 13728 19236 13860 19242
rect 13780 19230 13860 19236
rect 13728 19178 13780 19184
rect 13726 18864 13782 18873
rect 13924 18834 13952 20198
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 14016 19718 14044 19858
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13726 18799 13782 18808
rect 13912 18828 13964 18834
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13648 17626 13676 18362
rect 13740 18290 13768 18799
rect 13912 18770 13964 18776
rect 13820 18624 13872 18630
rect 13818 18592 13820 18601
rect 13872 18592 13874 18601
rect 13818 18527 13874 18536
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13556 17598 13676 17626
rect 13556 17338 13584 17598
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13556 16969 13584 17274
rect 13924 17116 13952 18022
rect 14016 17882 14044 19654
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14004 17128 14056 17134
rect 13924 17088 14004 17116
rect 14004 17070 14056 17076
rect 13542 16960 13598 16969
rect 13542 16895 13598 16904
rect 13910 16688 13966 16697
rect 13820 16652 13872 16658
rect 13910 16623 13966 16632
rect 13820 16594 13872 16600
rect 13542 16008 13598 16017
rect 13832 15994 13860 16594
rect 13924 16250 13952 16623
rect 14016 16454 14044 17070
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13740 15978 13860 15994
rect 13542 15943 13598 15952
rect 13728 15972 13860 15978
rect 13556 15858 13584 15943
rect 13780 15966 13860 15972
rect 13728 15914 13780 15920
rect 13556 15830 13676 15858
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13556 14618 13584 14962
rect 13174 14583 13230 14592
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13096 14504 13216 14532
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 11257 12112 13126
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12070 11248 12126 11257
rect 12070 11183 12126 11192
rect 12176 10742 12204 11834
rect 12268 11830 12296 13670
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12452 12986 12480 13262
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12544 12753 12572 13670
rect 12530 12744 12586 12753
rect 12530 12679 12586 12688
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12442 12480 12582
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12636 12356 12664 14214
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12728 12646 12756 13330
rect 13082 13288 13138 13297
rect 13082 13223 13138 13232
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12636 12328 12756 12356
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12176 10130 12204 10678
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12176 9722 12204 10066
rect 12452 9722 12480 10066
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12360 9518 12388 9658
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 9042 12296 9318
rect 12346 9208 12402 9217
rect 12346 9143 12402 9152
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12268 8634 12296 8978
rect 12360 8974 12388 9143
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 11978 3496 12034 3505
rect 11978 3431 12034 3440
rect 11980 2440 12032 2446
rect 11978 2408 11980 2417
rect 12032 2408 12034 2417
rect 12452 2378 12480 9522
rect 12544 7954 12572 10950
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12636 8974 12664 9658
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8430 12664 8910
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12636 7886 12664 8366
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7546 12664 7822
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12728 6769 12756 12328
rect 13004 11898 13032 12922
rect 13096 12753 13124 13223
rect 13082 12744 13138 12753
rect 13082 12679 13138 12688
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12912 11121 12940 11154
rect 12992 11144 13044 11150
rect 12898 11112 12954 11121
rect 12992 11086 13044 11092
rect 12898 11047 12954 11056
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 9926 12848 10474
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 13004 8634 13032 11086
rect 13188 10305 13216 14504
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 14006 13492 14418
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13452 13864 13504 13870
rect 13556 13852 13584 14554
rect 13504 13824 13584 13852
rect 13452 13806 13504 13812
rect 13542 13696 13598 13705
rect 13542 13631 13598 13640
rect 13450 13424 13506 13433
rect 13450 13359 13506 13368
rect 13266 13288 13322 13297
rect 13266 13223 13322 13232
rect 13280 12889 13308 13223
rect 13266 12880 13322 12889
rect 13266 12815 13322 12824
rect 13174 10296 13230 10305
rect 13174 10231 13230 10240
rect 13280 9110 13308 12815
rect 13464 12782 13492 13359
rect 13556 12986 13584 13631
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13648 10577 13676 15830
rect 13726 15736 13782 15745
rect 13726 15671 13782 15680
rect 13740 12850 13768 15671
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 14618 13860 15370
rect 13924 14822 13952 15506
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 14016 14770 14044 16390
rect 14108 16250 14136 20703
rect 14200 17814 14228 20862
rect 14384 20602 14412 21014
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19242 14320 19790
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14188 17808 14240 17814
rect 14188 17750 14240 17756
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14200 16289 14228 17614
rect 14384 17377 14412 20538
rect 14370 17368 14426 17377
rect 14370 17303 14426 17312
rect 14476 17218 14504 24006
rect 14554 23896 14610 23905
rect 14554 23831 14556 23840
rect 14608 23831 14610 23840
rect 14556 23802 14608 23808
rect 14554 23624 14610 23633
rect 14554 23559 14610 23568
rect 14568 22953 14596 23559
rect 14660 22982 14688 24210
rect 14752 24070 14780 24618
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14648 22976 14700 22982
rect 14554 22944 14610 22953
rect 14648 22918 14700 22924
rect 14554 22879 14610 22888
rect 14660 22778 14688 22918
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14556 22092 14608 22098
rect 14556 22034 14608 22040
rect 14568 20806 14596 22034
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14568 19258 14596 20742
rect 14646 20632 14702 20641
rect 14646 20567 14702 20576
rect 14660 20058 14688 20567
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14568 19230 14688 19258
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18222 14596 19110
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14568 17882 14596 18158
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14292 17190 14504 17218
rect 14186 16280 14242 16289
rect 14096 16244 14148 16250
rect 14186 16215 14242 16224
rect 14096 16186 14148 16192
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14200 14890 14228 15982
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13832 13530 13860 13738
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13924 13161 13952 14758
rect 14016 14742 14228 14770
rect 14200 14414 14228 14742
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14108 14074 14136 14350
rect 14200 14249 14228 14350
rect 14186 14240 14242 14249
rect 14186 14175 14242 14184
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 13910 13152 13966 13161
rect 13910 13087 13966 13096
rect 14108 12968 14136 14010
rect 14200 13530 14228 14175
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 13924 12940 14136 12968
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13820 12640 13872 12646
rect 13924 12628 13952 12940
rect 14002 12880 14058 12889
rect 14002 12815 14058 12824
rect 14096 12844 14148 12850
rect 14016 12782 14044 12815
rect 14096 12786 14148 12792
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13924 12600 14044 12628
rect 13820 12582 13872 12588
rect 13832 12102 13860 12582
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 11150 13768 11562
rect 13832 11257 13860 12038
rect 13818 11248 13874 11257
rect 13818 11183 13874 11192
rect 13728 11144 13780 11150
rect 13780 11104 13860 11132
rect 13728 11086 13780 11092
rect 13832 10810 13860 11104
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13634 10568 13690 10577
rect 13634 10503 13690 10512
rect 13820 10464 13872 10470
rect 13634 10432 13690 10441
rect 13634 10367 13690 10376
rect 13740 10424 13820 10452
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13280 8634 13308 9046
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8498 13400 8978
rect 13556 8498 13584 9862
rect 13648 9625 13676 10367
rect 13634 9616 13690 9625
rect 13634 9551 13690 9560
rect 13740 9178 13768 10424
rect 13820 10406 13872 10412
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13924 9058 13952 10678
rect 14016 9178 14044 12600
rect 14108 12306 14136 12786
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14094 11928 14150 11937
rect 14094 11863 14150 11872
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 13740 9042 13952 9058
rect 13728 9036 13952 9042
rect 13780 9030 13952 9036
rect 13728 8978 13780 8984
rect 14016 8634 14044 9114
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 8090 13308 8366
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13556 8022 13584 8434
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 12820 7342 12848 7958
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7546 13492 7890
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 12808 7336 12860 7342
rect 12806 7304 12808 7313
rect 12860 7304 12862 7313
rect 12806 7239 12862 7248
rect 14108 6905 14136 11863
rect 14200 11393 14228 12174
rect 14186 11384 14242 11393
rect 14186 11319 14242 11328
rect 14186 10024 14242 10033
rect 14186 9959 14242 9968
rect 14200 7721 14228 9959
rect 14292 9625 14320 17190
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 15910 14412 16390
rect 14568 16114 14596 16934
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14372 15904 14424 15910
rect 14370 15872 14372 15881
rect 14464 15904 14516 15910
rect 14424 15872 14426 15881
rect 14464 15846 14516 15852
rect 14370 15807 14426 15816
rect 14370 15600 14426 15609
rect 14370 15535 14426 15544
rect 14384 11354 14412 15535
rect 14476 15434 14504 15846
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14476 14006 14504 14214
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14476 12073 14504 13942
rect 14660 13410 14688 19230
rect 14568 13382 14688 13410
rect 14568 12481 14596 13382
rect 14554 12472 14610 12481
rect 14554 12407 14610 12416
rect 14648 12368 14700 12374
rect 14554 12336 14610 12345
rect 14648 12310 14700 12316
rect 14554 12271 14610 12280
rect 14462 12064 14518 12073
rect 14462 11999 14518 12008
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10169 14504 10406
rect 14462 10160 14518 10169
rect 14462 10095 14518 10104
rect 14462 9752 14518 9761
rect 14462 9687 14518 9696
rect 14278 9616 14334 9625
rect 14278 9551 14334 9560
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14292 8974 14320 9386
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 7750 14320 8910
rect 14280 7744 14332 7750
rect 14186 7712 14242 7721
rect 14280 7686 14332 7692
rect 14186 7647 14242 7656
rect 14094 6896 14150 6905
rect 14094 6831 14150 6840
rect 12714 6760 12770 6769
rect 12714 6695 12770 6704
rect 14292 2650 14320 7686
rect 14384 5953 14412 9046
rect 14476 8294 14504 9687
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 7732 14504 8230
rect 14568 8090 14596 12271
rect 14660 11898 14688 12310
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14660 9178 14688 9658
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14660 8498 14688 9114
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14556 7744 14608 7750
rect 14476 7704 14556 7732
rect 14556 7686 14608 7692
rect 14568 7177 14596 7686
rect 14554 7168 14610 7177
rect 14554 7103 14610 7112
rect 14660 6769 14688 8298
rect 14752 7410 14780 24006
rect 14844 23361 14872 24550
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 14830 23352 14886 23361
rect 14830 23287 14886 23296
rect 14936 23089 14964 23462
rect 15108 23112 15160 23118
rect 14922 23080 14978 23089
rect 14922 23015 14978 23024
rect 15106 23080 15108 23089
rect 15160 23080 15162 23089
rect 15106 23015 15162 23024
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15200 22704 15252 22710
rect 15198 22672 15200 22681
rect 15252 22672 15254 22681
rect 15198 22607 15254 22616
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21593 15332 24822
rect 15396 24721 15424 27520
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15382 24712 15438 24721
rect 15382 24647 15438 24656
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15396 22982 15424 23598
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15396 22574 15424 22918
rect 15384 22568 15436 22574
rect 15384 22510 15436 22516
rect 15488 22030 15516 24550
rect 15580 24041 15608 25298
rect 16040 24800 16068 27520
rect 16304 25764 16356 25770
rect 16304 25706 16356 25712
rect 16120 25424 16172 25430
rect 16120 25366 16172 25372
rect 16132 25294 16160 25366
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 16132 24954 16160 25230
rect 16120 24948 16172 24954
rect 16120 24890 16172 24896
rect 15672 24772 16068 24800
rect 15566 24032 15622 24041
rect 15566 23967 15622 23976
rect 15580 22273 15608 23967
rect 15566 22264 15622 22273
rect 15566 22199 15622 22208
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15396 21690 15424 21898
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15290 21584 15346 21593
rect 15488 21554 15516 21830
rect 15290 21519 15346 21528
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14844 20262 14872 20946
rect 15580 20874 15608 22034
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14844 20097 14872 20198
rect 14830 20088 14886 20097
rect 14830 20023 14886 20032
rect 14936 19972 14964 20198
rect 14844 19944 14964 19972
rect 14844 19514 14872 19944
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19514 15332 19858
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 14844 18970 14872 19246
rect 15014 19136 15070 19145
rect 15014 19071 15070 19080
rect 15028 18970 15056 19071
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15304 18902 15332 19450
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15488 18630 15516 19790
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 15108 17672 15160 17678
rect 15106 17640 15108 17649
rect 15160 17640 15162 17649
rect 15106 17575 15162 17584
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14830 15872 14886 15881
rect 14830 15807 14886 15816
rect 14844 15706 14872 15807
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14278 14872 14826
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14844 7954 14872 12854
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15028 10266 15056 10610
rect 15304 10470 15332 18090
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15396 17202 15424 17478
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15396 16794 15424 17138
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15488 16017 15516 18566
rect 15474 16008 15530 16017
rect 15474 15943 15530 15952
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15745 15516 15846
rect 15474 15736 15530 15745
rect 15474 15671 15530 15680
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15396 15162 15424 15438
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 14249 15424 14418
rect 15488 14278 15516 15506
rect 15476 14272 15528 14278
rect 15382 14240 15438 14249
rect 15476 14214 15528 14220
rect 15382 14175 15438 14184
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15396 13705 15424 13806
rect 15382 13696 15438 13705
rect 15382 13631 15438 13640
rect 15488 13569 15516 14214
rect 15474 13560 15530 13569
rect 15474 13495 15530 13504
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15488 12782 15516 13126
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15396 11694 15424 12242
rect 15488 11898 15516 12718
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11218 15424 11630
rect 15580 11529 15608 20810
rect 15672 18222 15700 24772
rect 16224 24750 16252 25298
rect 16212 24744 16264 24750
rect 15934 24712 15990 24721
rect 16212 24686 16264 24692
rect 15934 24647 15990 24656
rect 15842 24304 15898 24313
rect 15842 24239 15898 24248
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15764 23905 15792 24142
rect 15750 23896 15806 23905
rect 15750 23831 15806 23840
rect 15764 23662 15792 23831
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15764 21842 15792 21966
rect 15856 21962 15884 24239
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15764 21814 15884 21842
rect 15856 21457 15884 21814
rect 15842 21448 15898 21457
rect 15842 21383 15898 21392
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15764 20330 15792 21014
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 15856 19922 15884 21383
rect 15948 21146 15976 24647
rect 16316 24562 16344 25706
rect 16592 25242 16620 27520
rect 17038 25528 17094 25537
rect 17144 25498 17172 27520
rect 17590 25936 17646 25945
rect 17590 25871 17646 25880
rect 17038 25463 17094 25472
rect 17132 25492 17184 25498
rect 17052 25362 17080 25463
rect 17132 25434 17184 25440
rect 17222 25392 17278 25401
rect 17040 25356 17092 25362
rect 17222 25327 17278 25336
rect 17040 25298 17092 25304
rect 16592 25214 16712 25242
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24750 16620 25094
rect 16684 24857 16712 25214
rect 17052 24954 17080 25298
rect 17040 24948 17092 24954
rect 17040 24890 17092 24896
rect 16670 24848 16726 24857
rect 16670 24783 16726 24792
rect 16580 24744 16632 24750
rect 16580 24686 16632 24692
rect 16040 24534 16344 24562
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 16040 22710 16068 24534
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 16132 23526 16160 24210
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16304 24200 16356 24206
rect 16776 24177 16804 24550
rect 16304 24142 16356 24148
rect 16578 24168 16634 24177
rect 16224 23866 16252 24142
rect 16212 23860 16264 23866
rect 16212 23802 16264 23808
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 16212 23248 16264 23254
rect 16212 23190 16264 23196
rect 16028 22704 16080 22710
rect 16028 22646 16080 22652
rect 16224 22234 16252 23190
rect 16316 22982 16344 24142
rect 16578 24103 16634 24112
rect 16762 24168 16818 24177
rect 16762 24103 16818 24112
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16408 23254 16436 23802
rect 16396 23248 16448 23254
rect 16396 23190 16448 23196
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16394 22944 16450 22953
rect 16394 22879 16450 22888
rect 16408 22778 16436 22879
rect 16500 22817 16528 24006
rect 16592 23866 16620 24103
rect 17052 24041 17080 24550
rect 17236 24206 17264 25327
rect 17604 24342 17632 25871
rect 17788 24721 17816 27520
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 17774 24712 17830 24721
rect 17774 24647 17830 24656
rect 18064 24410 18092 25774
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18156 24750 18184 25094
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 18052 24404 18104 24410
rect 18052 24346 18104 24352
rect 17592 24336 17644 24342
rect 17592 24278 17644 24284
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17420 24138 17448 24210
rect 17408 24132 17460 24138
rect 17408 24074 17460 24080
rect 17316 24064 17368 24070
rect 17038 24032 17094 24041
rect 17316 24006 17368 24012
rect 17038 23967 17094 23976
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 17328 23225 17356 24006
rect 17420 23866 17448 24074
rect 17604 23866 17632 24278
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 18064 23662 18092 24346
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17314 23216 17370 23225
rect 17314 23151 17370 23160
rect 16762 23080 16818 23089
rect 16762 23015 16818 23024
rect 17498 23080 17554 23089
rect 17498 23015 17500 23024
rect 16486 22808 16542 22817
rect 16396 22772 16448 22778
rect 16486 22743 16542 22752
rect 16396 22714 16448 22720
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16396 22568 16448 22574
rect 16396 22510 16448 22516
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 16408 21690 16436 22510
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16396 21412 16448 21418
rect 16396 21354 16448 21360
rect 16408 21321 16436 21354
rect 16394 21312 16450 21321
rect 16394 21247 16450 21256
rect 16408 21146 16436 21247
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15948 19378 15976 19790
rect 16408 19718 16436 20946
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 16224 18154 16252 18702
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16316 18086 16344 18770
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 15672 17066 15700 17682
rect 15752 17604 15804 17610
rect 15752 17546 15804 17552
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15764 16969 15792 17546
rect 16132 16998 16160 17682
rect 15936 16992 15988 16998
rect 15750 16960 15806 16969
rect 15936 16934 15988 16940
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 15750 16895 15806 16904
rect 15764 16658 15792 16895
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15672 11801 15700 16594
rect 15764 16250 15792 16594
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15764 15570 15792 16186
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15750 15328 15806 15337
rect 15750 15263 15806 15272
rect 15764 13682 15792 15263
rect 15948 15201 15976 16934
rect 16026 16008 16082 16017
rect 16026 15943 16082 15952
rect 16040 15706 16068 15943
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15934 15192 15990 15201
rect 15934 15127 15990 15136
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 16040 13938 16068 14214
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 15936 13728 15988 13734
rect 15764 13654 15884 13682
rect 15936 13670 15988 13676
rect 15750 13424 15806 13433
rect 15750 13359 15752 13368
rect 15804 13359 15806 13368
rect 15752 13330 15804 13336
rect 15658 11792 15714 11801
rect 15658 11727 15714 11736
rect 15566 11520 15622 11529
rect 15566 11455 15622 11464
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15396 10810 15424 11154
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9722 15332 10202
rect 15488 9897 15516 10406
rect 15580 10266 15608 11222
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15474 9888 15530 9897
rect 15474 9823 15530 9832
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15658 9616 15714 9625
rect 15658 9551 15714 9560
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15396 8401 15424 8570
rect 15382 8392 15438 8401
rect 15382 8327 15438 8336
rect 15106 8256 15162 8265
rect 15106 8191 15162 8200
rect 15120 8090 15148 8191
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14646 6760 14702 6769
rect 14646 6695 14702 6704
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15396 6458 15424 8327
rect 15672 8090 15700 9551
rect 15750 9480 15806 9489
rect 15750 9415 15806 9424
rect 15764 9382 15792 9415
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15764 8294 15792 8978
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15488 7002 15516 7890
rect 15764 7546 15792 8230
rect 15856 7857 15884 13654
rect 15948 12782 15976 13670
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 16040 11830 16068 13874
rect 16132 12646 16160 16934
rect 16316 16425 16344 18022
rect 16302 16416 16358 16425
rect 16302 16351 16358 16360
rect 16408 16130 16436 19654
rect 16500 17338 16528 22646
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16592 21894 16620 22578
rect 16776 22506 16804 23015
rect 17552 23015 17554 23024
rect 17500 22986 17552 22992
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16776 22234 16804 22442
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16672 22160 16724 22166
rect 16672 22102 16724 22108
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 21078 16620 21830
rect 16684 21486 16712 22102
rect 17788 22098 17816 22510
rect 18052 22432 18104 22438
rect 18050 22400 18052 22409
rect 18104 22400 18106 22409
rect 18050 22335 18106 22344
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17132 22024 17184 22030
rect 17592 22024 17644 22030
rect 17132 21966 17184 21972
rect 17590 21992 17592 22001
rect 17644 21992 17646 22001
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16592 17882 16620 18702
rect 16684 18290 16712 21422
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16776 20398 16804 20878
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 19854 16804 20198
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16776 19514 16804 19790
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16762 17640 16818 17649
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16500 16250 16528 17070
rect 16592 16658 16620 17614
rect 16762 17575 16818 17584
rect 16856 17604 16908 17610
rect 16776 17134 16804 17575
rect 16856 17546 16908 17552
rect 16868 17338 16896 17546
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16592 16454 16620 16594
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16408 16102 16528 16130
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16224 14482 16252 15098
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16224 14006 16252 14418
rect 16316 14074 16344 14418
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16316 13190 16344 13670
rect 16408 13462 16436 14758
rect 16396 13456 16448 13462
rect 16396 13398 16448 13404
rect 16304 13184 16356 13190
rect 16302 13152 16304 13161
rect 16356 13152 16358 13161
rect 16302 13087 16358 13096
rect 16408 12986 16436 13398
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16224 12209 16252 12922
rect 16500 12866 16528 16102
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16764 15564 16816 15570
rect 16764 15506 16816 15512
rect 16776 15162 16804 15506
rect 16868 15337 16896 15846
rect 16960 15586 16988 21286
rect 17052 21078 17080 21490
rect 17144 21350 17172 21966
rect 17590 21927 17646 21936
rect 17604 21554 17632 21927
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 17052 20058 17080 21014
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17144 19258 17172 21286
rect 17788 20874 17816 21830
rect 17880 21690 17908 22034
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17880 21146 17908 21626
rect 18064 21350 18092 21966
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17776 20868 17828 20874
rect 17776 20810 17828 20816
rect 17406 20632 17462 20641
rect 17406 20567 17462 20576
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17236 19514 17264 19858
rect 17328 19514 17356 20334
rect 17420 20058 17448 20567
rect 17498 20496 17554 20505
rect 17498 20431 17554 20440
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17222 19272 17278 19281
rect 17144 19230 17222 19258
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 17052 17202 17080 17750
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16114 17080 16390
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17052 15706 17080 16050
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 16960 15558 17080 15586
rect 16854 15328 16910 15337
rect 16854 15263 16910 15272
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16408 12838 16528 12866
rect 16210 12200 16266 12209
rect 16210 12135 16266 12144
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 16118 11792 16174 11801
rect 16040 11286 16068 11766
rect 16224 11762 16252 12038
rect 16118 11727 16174 11736
rect 16212 11756 16264 11762
rect 16132 11694 16160 11727
rect 16212 11698 16264 11704
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 16132 10810 16160 11630
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16040 10130 16068 10746
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16040 9110 16068 10066
rect 16224 9654 16252 11698
rect 16316 11354 16344 12786
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16316 10198 16344 11290
rect 16408 10792 16436 12838
rect 16684 12442 16712 14894
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16776 13394 16804 13942
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16776 12986 16804 13330
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16948 12776 17000 12782
rect 17052 12753 17080 15558
rect 16948 12718 17000 12724
rect 17038 12744 17094 12753
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11762 16712 12038
rect 16868 11762 16896 12242
rect 16960 12102 16988 12718
rect 17038 12679 17094 12688
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16672 11756 16724 11762
rect 16856 11756 16908 11762
rect 16672 11698 16724 11704
rect 16776 11716 16856 11744
rect 16580 10804 16632 10810
rect 16408 10764 16580 10792
rect 16580 10746 16632 10752
rect 16580 10464 16632 10470
rect 16500 10424 16580 10452
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16316 9722 16344 10134
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16500 9178 16528 10424
rect 16580 10406 16632 10412
rect 16776 9586 16804 11716
rect 16856 11698 16908 11704
rect 17144 10713 17172 19230
rect 17222 19207 17278 19216
rect 17512 18970 17540 20431
rect 17960 20392 18012 20398
rect 17880 20340 17960 20346
rect 17880 20334 18012 20340
rect 17880 20318 18000 20334
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17788 18970 17816 20198
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17406 18728 17462 18737
rect 17406 18663 17462 18672
rect 17420 18426 17448 18663
rect 17788 18426 17816 18906
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17420 18222 17448 18362
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17222 17640 17278 17649
rect 17222 17575 17278 17584
rect 17236 15473 17264 17575
rect 17222 15464 17278 15473
rect 17222 15399 17278 15408
rect 17130 10704 17186 10713
rect 17130 10639 17186 10648
rect 17328 10033 17356 18022
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17696 16794 17724 17138
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15609 17448 15846
rect 17406 15600 17462 15609
rect 17406 15535 17462 15544
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17604 14618 17632 15030
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17880 12986 17908 20318
rect 18064 19718 18092 21286
rect 18156 20913 18184 24686
rect 18234 24440 18290 24449
rect 18234 24375 18290 24384
rect 18248 23730 18276 24375
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18248 23322 18276 23666
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 18142 20904 18198 20913
rect 18142 20839 18198 20848
rect 18340 20602 18368 27520
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18512 25220 18564 25226
rect 18512 25162 18564 25168
rect 18524 24954 18552 25162
rect 18512 24948 18564 24954
rect 18512 24890 18564 24896
rect 18418 23352 18474 23361
rect 18418 23287 18474 23296
rect 18432 22574 18460 23287
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18616 22250 18644 25910
rect 18892 24834 18920 27520
rect 18800 24806 18920 24834
rect 19246 24848 19302 24857
rect 18972 24812 19024 24818
rect 18800 22545 18828 24806
rect 19246 24783 19302 24792
rect 18972 24754 19024 24760
rect 18880 24608 18932 24614
rect 18878 24576 18880 24585
rect 18932 24576 18934 24585
rect 18878 24511 18934 24520
rect 18984 23730 19012 24754
rect 19260 24614 19288 24783
rect 19338 24712 19394 24721
rect 19338 24647 19394 24656
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19352 24410 19380 24647
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19076 24070 19104 24210
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 19076 23866 19104 24006
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18984 23322 19012 23666
rect 19352 23322 19380 23734
rect 19444 23497 19472 24550
rect 19536 24313 19564 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20088 25498 20116 27520
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20088 24410 20116 25230
rect 20640 25226 20668 27520
rect 20628 25220 20680 25226
rect 20628 25162 20680 25168
rect 20628 24948 20680 24954
rect 20628 24890 20680 24896
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19522 24304 19578 24313
rect 19522 24239 19578 24248
rect 20456 23798 20484 24550
rect 20548 24070 20576 24550
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 20444 23792 20496 23798
rect 20444 23734 20496 23740
rect 19430 23488 19486 23497
rect 19430 23423 19486 23432
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 18972 23316 19024 23322
rect 18972 23258 19024 23264
rect 19340 23316 19392 23322
rect 19340 23258 19392 23264
rect 18984 22778 19012 23258
rect 19996 23254 20024 23734
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 19984 23248 20036 23254
rect 19984 23190 20036 23196
rect 20272 22982 20300 23598
rect 20260 22976 20312 22982
rect 20258 22944 20260 22953
rect 20312 22944 20314 22953
rect 20258 22879 20314 22888
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 18786 22536 18842 22545
rect 19812 22506 19840 22714
rect 19982 22536 20038 22545
rect 18786 22471 18842 22480
rect 19800 22500 19852 22506
rect 19982 22471 20038 22480
rect 19800 22442 19852 22448
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 18432 22222 18644 22250
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19378 18092 19654
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 18326 18184 18382 18193
rect 18326 18119 18328 18128
rect 18380 18119 18382 18128
rect 18328 18090 18380 18096
rect 18326 17776 18382 17785
rect 18144 17740 18196 17746
rect 18326 17711 18382 17720
rect 18144 17682 18196 17688
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 18064 15162 18092 15846
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18064 14958 18092 15098
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18050 13152 18106 13161
rect 18050 13087 18106 13096
rect 18064 12986 18092 13087
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 17682 12744 17738 12753
rect 17682 12679 17738 12688
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 11558 17448 12582
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17314 10024 17370 10033
rect 17314 9959 17370 9968
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16670 9480 16726 9489
rect 16670 9415 16672 9424
rect 16724 9415 16726 9424
rect 16672 9386 16724 9392
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16028 9104 16080 9110
rect 16028 9046 16080 9052
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16028 8968 16080 8974
rect 16120 8968 16172 8974
rect 16028 8910 16080 8916
rect 16118 8936 16120 8945
rect 16172 8936 16174 8945
rect 15842 7848 15898 7857
rect 15842 7783 15898 7792
rect 16040 7546 16068 8910
rect 16118 8871 16174 8880
rect 16132 8634 16160 8871
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16408 7954 16436 9046
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 8084 16540 8090
rect 16592 8072 16620 8366
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16776 8265 16804 8298
rect 16762 8256 16818 8265
rect 16762 8191 16818 8200
rect 16540 8044 16620 8072
rect 16488 8026 16540 8032
rect 16396 7948 16448 7954
rect 16316 7908 16396 7936
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16316 7410 16344 7908
rect 16396 7890 16448 7896
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16408 7410 16436 7686
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 16408 6458 16436 7346
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16500 6866 16528 7278
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16776 6798 16804 8191
rect 16764 6792 16816 6798
rect 16486 6760 16542 6769
rect 16764 6734 16816 6740
rect 16486 6695 16542 6704
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5953 16436 6054
rect 14370 5944 14426 5953
rect 14370 5879 14426 5888
rect 16394 5944 16450 5953
rect 16394 5879 16396 5888
rect 16448 5879 16450 5888
rect 16396 5850 16448 5856
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13740 2394 13768 2450
rect 11978 2343 12034 2352
rect 12440 2372 12492 2378
rect 13740 2366 13952 2394
rect 12440 2314 12492 2320
rect 11794 1592 11850 1601
rect 11794 1527 11850 1536
rect 13924 480 13952 2366
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 16500 1601 16528 6695
rect 16868 5273 16896 9318
rect 16960 9178 16988 9522
rect 17038 9344 17094 9353
rect 17038 9279 17094 9288
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17052 9081 17080 9279
rect 17038 9072 17094 9081
rect 17038 9007 17094 9016
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17420 8498 17448 8978
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 16960 8090 16988 8434
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16960 7410 16988 8026
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16960 7002 16988 7346
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17406 6896 17462 6905
rect 17406 6831 17462 6840
rect 17420 6798 17448 6831
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16960 6322 16988 6598
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16960 5914 16988 6258
rect 17420 6118 17448 6734
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16854 5264 16910 5273
rect 16854 5199 16910 5208
rect 17420 3097 17448 6054
rect 17512 4049 17540 11494
rect 17696 10713 17724 12679
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17788 11354 17816 12242
rect 17868 12096 17920 12102
rect 17920 12044 18092 12050
rect 17868 12038 18092 12044
rect 17880 12022 18092 12038
rect 17960 11824 18012 11830
rect 17958 11792 17960 11801
rect 18012 11792 18014 11801
rect 17958 11727 18014 11736
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17866 11520 17922 11529
rect 17866 11455 17922 11464
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17682 10704 17738 10713
rect 17682 10639 17738 10648
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 7954 17632 9862
rect 17880 9625 17908 11455
rect 17972 11393 18000 11630
rect 17958 11384 18014 11393
rect 17958 11319 17960 11328
rect 18012 11319 18014 11328
rect 17960 11290 18012 11296
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17972 10606 18000 11018
rect 18064 10810 18092 12022
rect 18156 10985 18184 17682
rect 18340 14550 18368 17711
rect 18432 14822 18460 22222
rect 18892 22137 18920 22374
rect 18878 22128 18934 22137
rect 19352 22114 19380 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 18878 22063 18934 22072
rect 19076 22086 19380 22114
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18708 21418 18736 21830
rect 19076 21486 19104 22086
rect 19706 21992 19762 22001
rect 19706 21927 19708 21936
rect 19760 21927 19762 21936
rect 19708 21898 19760 21904
rect 19524 21888 19576 21894
rect 19246 21856 19302 21865
rect 19524 21830 19576 21836
rect 19246 21791 19302 21800
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18696 21412 18748 21418
rect 18696 21354 18748 21360
rect 18708 21078 18736 21354
rect 19260 21146 19288 21791
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 19260 20602 19288 20946
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19352 20482 19380 20878
rect 19260 20454 19380 20482
rect 19444 20466 19472 21354
rect 19536 20602 19564 21830
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19800 21072 19852 21078
rect 19800 21014 19852 21020
rect 19812 20942 19840 21014
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19522 20496 19578 20505
rect 19432 20460 19484 20466
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18524 18612 18552 19178
rect 18616 19174 18644 19858
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18616 18970 18644 19110
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18616 18766 18644 18906
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18604 18624 18656 18630
rect 18524 18584 18604 18612
rect 18604 18566 18656 18572
rect 18616 18290 18644 18566
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18510 18184 18566 18193
rect 18510 18119 18566 18128
rect 18524 18086 18552 18119
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18616 17882 18644 18226
rect 18604 17876 18656 17882
rect 18604 17818 18656 17824
rect 18694 17232 18750 17241
rect 18694 17167 18750 17176
rect 18708 17134 18736 17167
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18708 16794 18736 17070
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18708 16697 18736 16730
rect 18694 16688 18750 16697
rect 18694 16623 18750 16632
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 16114 18644 16390
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18524 14929 18552 15982
rect 18510 14920 18566 14929
rect 18510 14855 18566 14864
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18340 14006 18368 14486
rect 18616 14074 18644 16050
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18708 14618 18736 14758
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18616 13530 18644 13806
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18616 13410 18644 13466
rect 18524 13382 18644 13410
rect 18524 12866 18552 13382
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18432 12838 18552 12866
rect 18248 11762 18276 12786
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18340 12442 18368 12650
rect 18432 12458 18460 12838
rect 18510 12744 18566 12753
rect 18510 12679 18566 12688
rect 18524 12646 18552 12679
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18328 12436 18380 12442
rect 18432 12430 18552 12458
rect 18328 12378 18380 12384
rect 18328 12232 18380 12238
rect 18524 12186 18552 12430
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18380 12180 18552 12186
rect 18328 12174 18552 12180
rect 18340 12158 18552 12174
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18340 11626 18368 12158
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18340 11150 18368 11562
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18142 10976 18198 10985
rect 18142 10911 18198 10920
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 18340 9926 18368 11086
rect 18524 10112 18552 11290
rect 18616 11286 18644 12378
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18616 10742 18644 11222
rect 18708 10792 18736 13806
rect 18800 13802 18828 14214
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18800 13258 18828 13738
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18800 11354 18828 13194
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18892 11937 18920 12310
rect 18878 11928 18934 11937
rect 18878 11863 18934 11872
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18708 10764 18828 10792
rect 18604 10736 18656 10742
rect 18656 10684 18736 10690
rect 18604 10678 18736 10684
rect 18616 10662 18736 10678
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 10266 18644 10542
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18524 10084 18644 10112
rect 18512 9988 18564 9994
rect 18512 9930 18564 9936
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17866 9616 17922 9625
rect 17866 9551 17922 9560
rect 18340 9518 18368 9862
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18524 9450 18552 9930
rect 18616 9761 18644 10084
rect 18708 10062 18736 10662
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18602 9752 18658 9761
rect 18602 9687 18658 9696
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9110 17816 9318
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17788 8634 17816 9046
rect 18524 8945 18552 9386
rect 18510 8936 18566 8945
rect 18510 8871 18512 8880
rect 18564 8871 18566 8880
rect 18512 8842 18564 8848
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17682 8120 17738 8129
rect 17682 8055 17738 8064
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17604 7410 17632 7890
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 6798 17632 7346
rect 17696 7274 17724 8055
rect 17788 7546 17816 8366
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17880 7002 17908 8230
rect 18144 7200 18196 7206
rect 18144 7142 18196 7148
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17880 6458 17908 6938
rect 18156 6662 18184 7142
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18156 5137 18184 6598
rect 18142 5128 18198 5137
rect 18142 5063 18198 5072
rect 18524 4049 18552 7142
rect 18800 6361 18828 10764
rect 18984 10441 19012 20198
rect 19260 18970 19288 20454
rect 19522 20431 19578 20440
rect 19432 20402 19484 20408
rect 19444 20058 19472 20402
rect 19536 20398 19564 20431
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19076 18154 19104 18770
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 19246 17096 19302 17105
rect 19246 17031 19302 17040
rect 19154 16824 19210 16833
rect 19154 16759 19156 16768
rect 19208 16759 19210 16768
rect 19156 16730 19208 16736
rect 19260 16658 19288 17031
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 19168 16250 19196 16458
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19168 15706 19196 16186
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19260 15570 19288 16594
rect 19352 15881 19380 19790
rect 19444 18698 19472 19994
rect 19996 19854 20024 22471
rect 20548 21486 20576 24006
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20364 21078 20392 21286
rect 20352 21072 20404 21078
rect 20352 21014 20404 21020
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 19984 19848 20036 19854
rect 20548 19825 20576 20538
rect 19984 19790 20036 19796
rect 20534 19816 20590 19825
rect 20534 19751 20590 19760
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19444 17882 19472 18634
rect 19536 18086 19564 18702
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19338 15872 19394 15881
rect 19338 15807 19394 15816
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 14822 19380 15506
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19246 14648 19302 14657
rect 19246 14583 19248 14592
rect 19300 14583 19302 14592
rect 19248 14554 19300 14560
rect 19246 14512 19302 14521
rect 19246 14447 19302 14456
rect 19260 14414 19288 14447
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19168 13530 19196 14350
rect 19260 14074 19288 14350
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19248 13796 19300 13802
rect 19248 13738 19300 13744
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19168 13297 19196 13466
rect 19154 13288 19210 13297
rect 19154 13223 19210 13232
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 18970 10432 19026 10441
rect 18970 10367 19026 10376
rect 19168 10266 19196 13126
rect 19260 12753 19288 13738
rect 19246 12744 19302 12753
rect 19246 12679 19302 12688
rect 19246 11928 19302 11937
rect 19246 11863 19302 11872
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19154 9888 19210 9897
rect 19154 9823 19210 9832
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18892 8634 18920 9318
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 19168 7886 19196 9823
rect 19260 8514 19288 11863
rect 19352 11665 19380 14758
rect 19338 11656 19394 11665
rect 19338 11591 19394 11600
rect 19352 11558 19380 11591
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19352 10674 19380 11018
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19340 10464 19392 10470
rect 19444 10452 19472 17682
rect 19536 13802 19564 18022
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17746 20024 19654
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20074 19136 20130 19145
rect 20074 19071 20130 19080
rect 20088 17882 20116 19071
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20180 18290 20208 18566
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19982 15192 20038 15201
rect 19982 15127 20038 15136
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19708 13456 19760 13462
rect 19708 13398 19760 13404
rect 19720 12986 19748 13398
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19536 10810 19564 12582
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19996 10577 20024 15127
rect 20088 14890 20116 15302
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 20088 14006 20116 14826
rect 20180 14793 20208 18090
rect 20456 18086 20484 19178
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20166 14784 20222 14793
rect 20166 14719 20222 14728
rect 20272 14498 20300 18022
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 16114 20392 17478
rect 20456 16250 20484 18022
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20364 15706 20392 16050
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20548 14618 20576 15914
rect 20640 15434 20668 24890
rect 21284 24857 21312 27520
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21560 25430 21588 25842
rect 21836 25498 21864 27520
rect 21824 25492 21876 25498
rect 21824 25434 21876 25440
rect 21548 25424 21600 25430
rect 21362 25392 21418 25401
rect 21548 25366 21600 25372
rect 21362 25327 21418 25336
rect 21270 24848 21326 24857
rect 21270 24783 21326 24792
rect 20718 24304 20774 24313
rect 20718 24239 20774 24248
rect 20732 23633 20760 24239
rect 20996 23656 21048 23662
rect 20718 23624 20774 23633
rect 20996 23598 21048 23604
rect 20718 23559 20774 23568
rect 21008 23118 21036 23598
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21008 22778 21036 23054
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 20902 21584 20958 21593
rect 20902 21519 20904 21528
rect 20956 21519 20958 21528
rect 20904 21490 20956 21496
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 21086 20360 21142 20369
rect 20916 20262 20944 20334
rect 21086 20295 21142 20304
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20824 19174 20852 19858
rect 20916 19786 20944 20198
rect 21100 20058 21128 20295
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20916 19310 20944 19722
rect 21192 19360 21220 21830
rect 21376 21078 21404 25327
rect 21456 24880 21508 24886
rect 21456 24822 21508 24828
rect 21468 24750 21496 24822
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 22284 24744 22336 24750
rect 22388 24721 22416 27520
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22572 24818 22600 25094
rect 22742 24848 22798 24857
rect 22560 24812 22612 24818
rect 22742 24783 22798 24792
rect 22560 24754 22612 24760
rect 22652 24744 22704 24750
rect 22284 24686 22336 24692
rect 22374 24712 22430 24721
rect 21916 24676 21968 24682
rect 21916 24618 21968 24624
rect 21928 24313 21956 24618
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 22020 24410 22048 24550
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 21914 24304 21970 24313
rect 22296 24290 22324 24686
rect 22374 24647 22430 24656
rect 22650 24712 22652 24721
rect 22704 24712 22706 24721
rect 22650 24647 22706 24656
rect 22296 24262 22416 24290
rect 21914 24239 21970 24248
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21468 23322 21496 24142
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21652 23526 21680 24074
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21468 23050 21496 23258
rect 21560 23118 21588 23462
rect 21652 23254 21680 23462
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21560 22574 21588 23054
rect 21652 22642 21680 23190
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21454 22128 21510 22137
rect 21454 22063 21510 22072
rect 21468 21690 21496 22063
rect 21744 22030 21772 24006
rect 22388 23338 22416 24262
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22480 23866 22508 24210
rect 22468 23860 22520 23866
rect 22468 23802 22520 23808
rect 22296 23310 22416 23338
rect 22296 23236 22324 23310
rect 22112 23208 22324 23236
rect 22112 23202 22140 23208
rect 21836 23174 22140 23202
rect 21732 22024 21784 22030
rect 21546 21992 21602 22001
rect 21732 21966 21784 21972
rect 21546 21927 21548 21936
rect 21600 21927 21602 21936
rect 21548 21898 21600 21904
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21560 21418 21588 21898
rect 21548 21412 21600 21418
rect 21548 21354 21600 21360
rect 21560 21146 21588 21354
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21100 19332 21220 19360
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20720 18216 20772 18222
rect 20824 18193 20852 19110
rect 20720 18158 20772 18164
rect 20810 18184 20866 18193
rect 20732 16794 20760 18158
rect 20810 18119 20866 18128
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20916 17270 20944 17614
rect 20904 17264 20956 17270
rect 20904 17206 20956 17212
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20824 15706 20852 16662
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 21008 15910 21036 15982
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20718 15464 20774 15473
rect 20628 15428 20680 15434
rect 20718 15399 20774 15408
rect 20628 15370 20680 15376
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20640 14550 20668 15370
rect 20628 14544 20680 14550
rect 20272 14470 20576 14498
rect 20628 14486 20680 14492
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20088 11393 20116 13942
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20180 11744 20208 12922
rect 20272 12850 20300 13126
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20272 12442 20300 12786
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 20180 11716 20300 11744
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20074 11384 20130 11393
rect 20074 11319 20130 11328
rect 20180 11082 20208 11562
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20074 10976 20130 10985
rect 20272 10962 20300 11716
rect 20074 10911 20130 10920
rect 20180 10934 20300 10962
rect 20088 10810 20116 10911
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 19982 10568 20038 10577
rect 19982 10503 20038 10512
rect 19444 10424 20116 10452
rect 19340 10406 19392 10412
rect 19352 10198 19380 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19352 8634 19380 10134
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19444 9654 19472 9998
rect 19982 9888 20038 9897
rect 19982 9823 20038 9832
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19522 9616 19578 9625
rect 19522 9551 19578 9560
rect 19430 9344 19486 9353
rect 19430 9279 19486 9288
rect 19444 9178 19472 9279
rect 19536 9178 19564 9551
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19444 8673 19472 9114
rect 19430 8664 19486 8673
rect 19340 8628 19392 8634
rect 19430 8599 19486 8608
rect 19340 8570 19392 8576
rect 19260 8486 19380 8514
rect 19444 8498 19472 8599
rect 19706 8528 19762 8537
rect 19352 8072 19380 8486
rect 19432 8492 19484 8498
rect 19706 8463 19762 8472
rect 19432 8434 19484 8440
rect 19720 8430 19748 8463
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19352 8044 19472 8072
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18984 7342 19012 7686
rect 19168 7546 19196 7822
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19352 7177 19380 7890
rect 19444 7342 19472 8044
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19628 7410 19656 7822
rect 19996 7546 20024 9823
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19338 7168 19394 7177
rect 19260 7126 19338 7154
rect 19260 7002 19288 7126
rect 19338 7103 19394 7112
rect 19444 7002 19472 7278
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 18786 6352 18842 6361
rect 18786 6287 18842 6296
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4185 20024 7142
rect 20088 6769 20116 10424
rect 20074 6760 20130 6769
rect 20074 6695 20130 6704
rect 20180 4729 20208 10934
rect 20258 9752 20314 9761
rect 20258 9687 20314 9696
rect 20272 7410 20300 9687
rect 20364 9042 20392 12854
rect 20456 12306 20484 13262
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20456 12102 20484 12242
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11529 20484 12038
rect 20442 11520 20498 11529
rect 20442 11455 20498 11464
rect 20456 9382 20484 11455
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20352 9036 20404 9042
rect 20352 8978 20404 8984
rect 20364 8090 20392 8978
rect 20548 8945 20576 14470
rect 20732 14385 20760 15399
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20916 14414 20944 14758
rect 20904 14408 20956 14414
rect 20718 14376 20774 14385
rect 20904 14350 20956 14356
rect 20718 14311 20774 14320
rect 20916 13734 20944 14350
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20640 12986 20668 13330
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20640 12288 20668 12718
rect 20732 12714 20760 13126
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20732 12617 20760 12650
rect 20718 12608 20774 12617
rect 20718 12543 20774 12552
rect 20720 12300 20772 12306
rect 20640 12260 20720 12288
rect 20640 12209 20668 12260
rect 20720 12242 20772 12248
rect 20626 12200 20682 12209
rect 20626 12135 20682 12144
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20640 9926 20668 10542
rect 20916 10266 20944 12922
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20628 9920 20680 9926
rect 20680 9868 20852 9874
rect 20628 9862 20852 9868
rect 20640 9846 20852 9862
rect 20628 8968 20680 8974
rect 20534 8936 20590 8945
rect 20628 8910 20680 8916
rect 20534 8871 20590 8880
rect 20536 8424 20588 8430
rect 20534 8392 20536 8401
rect 20640 8412 20668 8910
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 8430 20760 8774
rect 20824 8634 20852 9846
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20916 9178 20944 9454
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20916 8809 20944 8978
rect 20902 8800 20958 8809
rect 20902 8735 20958 8744
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20916 8566 20944 8735
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20588 8392 20668 8412
rect 20590 8384 20668 8392
rect 20720 8424 20772 8430
rect 20916 8401 20944 8502
rect 20720 8366 20772 8372
rect 20902 8392 20958 8401
rect 20534 8327 20590 8336
rect 20902 8327 20958 8336
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 7546 20668 7822
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 21008 7410 21036 15846
rect 21100 7585 21128 19332
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21192 18766 21220 19178
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21192 18290 21220 18702
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21178 18184 21234 18193
rect 21178 18119 21234 18128
rect 21192 16250 21220 18119
rect 21284 16794 21312 20742
rect 21376 20602 21404 21014
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21468 19990 21496 20878
rect 21560 20058 21588 21082
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21456 19984 21508 19990
rect 21652 19938 21680 21286
rect 21456 19926 21508 19932
rect 21362 18864 21418 18873
rect 21362 18799 21364 18808
rect 21416 18799 21418 18808
rect 21364 18770 21416 18776
rect 21376 18086 21404 18770
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21468 17898 21496 19926
rect 21376 17870 21496 17898
rect 21560 19910 21680 19938
rect 21376 17338 21404 17870
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21376 17134 21404 17274
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21284 16658 21312 16730
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21376 16522 21404 17070
rect 21468 16590 21496 17750
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21468 16114 21496 16526
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 15706 21496 16050
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21560 15586 21588 19910
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21652 18222 21680 18634
rect 21744 18426 21772 18906
rect 21836 18834 21864 23174
rect 22756 22778 22784 24783
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22204 22234 22232 22646
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21928 21026 21956 21422
rect 22020 21146 22048 21966
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 21928 20998 22048 21026
rect 21916 20324 21968 20330
rect 21916 20266 21968 20272
rect 21928 19718 21956 20266
rect 21916 19712 21968 19718
rect 21916 19654 21968 19660
rect 21928 18873 21956 19654
rect 22020 18970 22048 20998
rect 22112 20602 22140 21490
rect 22204 21146 22232 22170
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 21914 18864 21970 18873
rect 21824 18828 21876 18834
rect 21914 18799 21970 18808
rect 21824 18770 21876 18776
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 21836 18358 21864 18770
rect 21916 18760 21968 18766
rect 21968 18708 22232 18714
rect 21916 18702 22232 18708
rect 21928 18686 22232 18702
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21376 15558 21588 15586
rect 21652 15570 21680 18022
rect 22020 17898 22048 18022
rect 22020 17870 22140 17898
rect 22204 17882 22232 18686
rect 22112 17678 22140 17870
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22100 17672 22152 17678
rect 22296 17649 22324 22374
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22572 21690 22600 21966
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22744 18692 22796 18698
rect 22664 18652 22744 18680
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22374 18320 22430 18329
rect 22572 18290 22600 18566
rect 22374 18255 22376 18264
rect 22428 18255 22430 18264
rect 22560 18284 22612 18290
rect 22376 18226 22428 18232
rect 22560 18226 22612 18232
rect 22388 17882 22416 18226
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22468 17808 22520 17814
rect 22468 17750 22520 17756
rect 22100 17614 22152 17620
rect 22282 17640 22338 17649
rect 22282 17575 22338 17584
rect 22480 17338 22508 17750
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 21916 16244 21968 16250
rect 21916 16186 21968 16192
rect 21928 16046 21956 16186
rect 22020 16114 22048 16458
rect 22112 16250 22140 16934
rect 22572 16794 22600 17682
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22190 16416 22246 16425
rect 22190 16351 22246 16360
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 22112 15570 22140 16186
rect 21640 15564 21692 15570
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21192 13530 21220 14418
rect 21270 14104 21326 14113
rect 21270 14039 21272 14048
rect 21324 14039 21326 14048
rect 21272 14010 21324 14016
rect 21284 13870 21312 14010
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21284 13326 21312 13670
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 12646 21312 13262
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21284 11354 21312 12242
rect 21376 12102 21404 15558
rect 21640 15506 21692 15512
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21560 14822 21588 15438
rect 21652 15162 21680 15506
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21454 14648 21510 14657
rect 21454 14583 21510 14592
rect 21468 12442 21496 14583
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21914 13832 21970 13841
rect 21548 13796 21600 13802
rect 21914 13767 21970 13776
rect 21548 13738 21600 13744
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21284 11121 21312 11290
rect 21270 11112 21326 11121
rect 21270 11047 21326 11056
rect 21468 10470 21496 11494
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21468 8974 21496 10406
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21468 8022 21496 8910
rect 21560 8090 21588 13738
rect 21928 12986 21956 13767
rect 22020 13734 22048 13874
rect 22100 13796 22152 13802
rect 22100 13738 22152 13744
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 22020 13394 22048 13670
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22020 12782 22048 13330
rect 22112 12918 22140 13738
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21928 12322 21956 12582
rect 22020 12442 22048 12718
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21928 12294 22140 12322
rect 22112 12238 22140 12294
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22112 11558 22140 12174
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22112 11150 22140 11494
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21836 9926 21864 11018
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21638 9480 21694 9489
rect 21638 9415 21694 9424
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21086 7576 21142 7585
rect 21086 7511 21142 7520
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 20272 7002 20300 7346
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20166 4720 20222 4729
rect 20166 4655 20222 4664
rect 19982 4176 20038 4185
rect 19982 4111 20038 4120
rect 17498 4040 17554 4049
rect 17498 3975 17554 3984
rect 18510 4040 18566 4049
rect 18510 3975 18566 3984
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 17498 3632 17554 3641
rect 17498 3567 17554 3576
rect 17406 3088 17462 3097
rect 17406 3023 17462 3032
rect 17512 1737 17540 3567
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 21652 2553 21680 9415
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21744 8498 21772 9318
rect 21836 8498 21864 9862
rect 21928 9602 21956 11086
rect 22112 10810 22140 11086
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22020 10130 22048 10746
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22020 9722 22048 10066
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 21928 9574 22140 9602
rect 22006 9480 22062 9489
rect 22006 9415 22008 9424
rect 22060 9415 22062 9424
rect 22008 9386 22060 9392
rect 22112 9178 22140 9574
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 22006 8936 22062 8945
rect 22006 8871 22062 8880
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21836 7954 21864 8434
rect 22020 7970 22048 8871
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22112 8090 22140 8366
rect 22204 8129 22232 16351
rect 22374 16144 22430 16153
rect 22374 16079 22430 16088
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22296 14521 22324 14554
rect 22282 14512 22338 14521
rect 22282 14447 22338 14456
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22296 12714 22324 12786
rect 22388 12714 22416 16079
rect 22664 15552 22692 18652
rect 22744 18634 22796 18640
rect 22848 15858 22876 25434
rect 23032 24177 23060 27520
rect 23584 25809 23612 27520
rect 23570 25800 23626 25809
rect 23570 25735 23626 25744
rect 23768 25430 23796 27639
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25870 27520 25926 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 23756 25424 23808 25430
rect 23756 25366 23808 25372
rect 23768 24954 23796 25366
rect 24136 25226 24164 27520
rect 24674 26616 24730 26625
rect 24674 26551 24730 26560
rect 24398 26072 24454 26081
rect 24398 26007 24454 26016
rect 24412 25430 24440 26007
rect 24400 25424 24452 25430
rect 24228 25384 24400 25412
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 23768 24818 23796 24890
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23940 24676 23992 24682
rect 23940 24618 23992 24624
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23018 24168 23074 24177
rect 23216 24138 23244 24550
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 23018 24103 23074 24112
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 22926 23896 22982 23905
rect 22926 23831 22982 23840
rect 22940 23322 22968 23831
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 22940 22030 22968 23258
rect 23018 23080 23074 23089
rect 23018 23015 23074 23024
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22926 20904 22982 20913
rect 22926 20839 22928 20848
rect 22980 20839 22982 20848
rect 22928 20810 22980 20816
rect 22926 19952 22982 19961
rect 23032 19922 23060 23015
rect 23216 22982 23244 24074
rect 23308 23526 23336 24210
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23584 23594 23612 24142
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 23124 22234 23152 22374
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 22926 19887 22982 19896
rect 23020 19916 23072 19922
rect 22940 18154 22968 19887
rect 23020 19858 23072 19864
rect 23216 19242 23244 22918
rect 23308 21010 23336 23462
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23492 21690 23520 21966
rect 23480 21684 23532 21690
rect 23480 21626 23532 21632
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 23308 20602 23336 20946
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23400 20058 23428 21422
rect 23480 21412 23532 21418
rect 23480 21354 23532 21360
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 23308 19718 23336 19858
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23204 19236 23256 19242
rect 23204 19178 23256 19184
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22928 18148 22980 18154
rect 22928 18090 22980 18096
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 22940 16794 22968 17614
rect 23032 16998 23060 19110
rect 23308 18834 23336 19654
rect 23386 18864 23442 18873
rect 23296 18828 23348 18834
rect 23386 18799 23442 18808
rect 23296 18770 23348 18776
rect 23400 18698 23428 18799
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23112 18216 23164 18222
rect 23112 18158 23164 18164
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 23032 16590 23060 16934
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23032 16250 23060 16526
rect 23020 16244 23072 16250
rect 23020 16186 23072 16192
rect 23124 15978 23152 18158
rect 23400 17882 23428 18634
rect 23492 18426 23520 21354
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23478 18048 23534 18057
rect 23478 17983 23534 17992
rect 23388 17876 23440 17882
rect 23388 17818 23440 17824
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23112 15972 23164 15978
rect 23112 15914 23164 15920
rect 22848 15830 22968 15858
rect 22572 15524 22692 15552
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22480 13870 22508 14894
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22296 11801 22324 12650
rect 22282 11792 22338 11801
rect 22282 11727 22338 11736
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22296 10198 22324 10406
rect 22284 10192 22336 10198
rect 22284 10134 22336 10140
rect 22296 9586 22324 10134
rect 22284 9580 22336 9586
rect 22284 9522 22336 9528
rect 22296 9110 22324 9522
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22190 8120 22246 8129
rect 22100 8084 22152 8090
rect 22190 8055 22246 8064
rect 22100 8026 22152 8032
rect 22020 7954 22140 7970
rect 21824 7948 21876 7954
rect 22020 7948 22152 7954
rect 22020 7942 22100 7948
rect 21824 7890 21876 7896
rect 22100 7890 22152 7896
rect 22388 6089 22416 12650
rect 22468 11688 22520 11694
rect 22466 11656 22468 11665
rect 22520 11656 22522 11665
rect 22466 11591 22522 11600
rect 22572 9081 22600 15524
rect 22650 15056 22706 15065
rect 22650 14991 22706 15000
rect 22664 11898 22692 14991
rect 22940 12918 22968 15830
rect 23124 15706 23152 15914
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23020 15428 23072 15434
rect 23020 15370 23072 15376
rect 22744 12912 22796 12918
rect 22742 12880 22744 12889
rect 22928 12912 22980 12918
rect 22796 12880 22798 12889
rect 22928 12854 22980 12860
rect 22742 12815 22798 12824
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22756 11626 22784 12038
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22558 9072 22614 9081
rect 22468 9036 22520 9042
rect 22756 9042 22784 11562
rect 23032 10130 23060 15370
rect 23216 13462 23244 17478
rect 23294 16960 23350 16969
rect 23294 16895 23350 16904
rect 23308 16726 23336 16895
rect 23296 16720 23348 16726
rect 23492 16674 23520 17983
rect 23296 16662 23348 16668
rect 23308 16182 23336 16662
rect 23400 16646 23520 16674
rect 23296 16176 23348 16182
rect 23296 16118 23348 16124
rect 23400 15094 23428 16646
rect 23584 16130 23612 23530
rect 23676 23322 23704 24550
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23754 23760 23810 23769
rect 23754 23695 23810 23704
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23768 23202 23796 23695
rect 23676 23174 23796 23202
rect 23676 22001 23704 23174
rect 23754 23080 23810 23089
rect 23754 23015 23810 23024
rect 23662 21992 23718 22001
rect 23662 21927 23718 21936
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23676 21146 23704 21830
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23676 20602 23704 21082
rect 23768 20641 23796 23015
rect 23860 22166 23888 24006
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23860 21418 23888 22102
rect 23952 21894 23980 24618
rect 24044 24342 24072 25094
rect 24228 24410 24256 25384
rect 24400 25366 24452 25372
rect 24490 25392 24546 25401
rect 24490 25327 24492 25336
rect 24544 25327 24546 25336
rect 24492 25298 24544 25304
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24688 24426 24716 26551
rect 24780 25498 24808 27520
rect 25332 27282 25360 27520
rect 25148 27254 25360 27282
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24780 24954 24808 25327
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24872 24818 24900 25230
rect 25148 24857 25176 27254
rect 25318 27160 25374 27169
rect 25318 27095 25374 27104
rect 25228 25152 25280 25158
rect 25228 25094 25280 25100
rect 25134 24848 25190 24857
rect 24860 24812 24912 24818
rect 25134 24783 25190 24792
rect 24860 24754 24912 24760
rect 25240 24750 25268 25094
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 25136 24676 25188 24682
rect 25136 24618 25188 24624
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24216 24404 24268 24410
rect 24688 24398 24900 24426
rect 24216 24346 24268 24352
rect 24032 24336 24084 24342
rect 24032 24278 24084 24284
rect 24044 23662 24072 24278
rect 24136 23730 24164 24346
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24032 23656 24084 23662
rect 24032 23598 24084 23604
rect 24030 23488 24086 23497
rect 24030 23423 24086 23432
rect 24044 22114 24072 23423
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24136 22574 24164 22918
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24136 22234 24164 22510
rect 24124 22228 24176 22234
rect 24124 22170 24176 22176
rect 24044 22086 24164 22114
rect 24228 22098 24256 24346
rect 24872 24274 24900 24398
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24872 24154 24900 24210
rect 24872 24126 24992 24154
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24320 23594 24348 23666
rect 24308 23588 24360 23594
rect 24308 23530 24360 23536
rect 24320 23050 24348 23530
rect 24872 23322 24900 24006
rect 24964 23866 24992 24126
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24964 23769 24992 23802
rect 24950 23760 25006 23769
rect 24950 23695 25006 23704
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24308 23044 24360 23050
rect 24308 22986 24360 22992
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22438 24716 22986
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24688 22166 24716 22374
rect 24780 22234 24808 23190
rect 24872 22778 24900 23258
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 25042 22672 25098 22681
rect 25042 22607 25098 22616
rect 24768 22228 24820 22234
rect 24768 22170 24820 22176
rect 24676 22160 24728 22166
rect 24676 22102 24728 22108
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23952 20874 23980 21626
rect 24136 21570 24164 22086
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21690 24716 22102
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24044 21542 24164 21570
rect 24780 21554 24808 21830
rect 24308 21548 24360 21554
rect 24044 21026 24072 21542
rect 24308 21490 24360 21496
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24320 21128 24348 21490
rect 24872 21486 24900 22034
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24228 21100 24348 21128
rect 24044 20998 24164 21026
rect 23940 20868 23992 20874
rect 23940 20810 23992 20816
rect 23848 20800 23900 20806
rect 23848 20742 23900 20748
rect 23754 20632 23810 20641
rect 23664 20596 23716 20602
rect 23754 20567 23810 20576
rect 23664 20538 23716 20544
rect 23860 20466 23888 20742
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23676 18766 23704 19722
rect 23768 18902 23796 20198
rect 23848 19168 23900 19174
rect 23848 19110 23900 19116
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23860 18766 23888 19110
rect 23664 18760 23716 18766
rect 23662 18728 23664 18737
rect 23848 18760 23900 18766
rect 23716 18728 23718 18737
rect 23848 18702 23900 18708
rect 23662 18663 23718 18672
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 18154 23888 18566
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23676 17746 23704 18022
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23492 16102 23612 16130
rect 23492 15434 23520 16102
rect 23572 16040 23624 16046
rect 23572 15982 23624 15988
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23478 15328 23534 15337
rect 23478 15263 23534 15272
rect 23492 15162 23520 15263
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23478 14240 23534 14249
rect 23308 14074 23336 14214
rect 23478 14175 23534 14184
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23308 13802 23336 14010
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 23400 13530 23428 13874
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23204 13456 23256 13462
rect 23204 13398 23256 13404
rect 23110 13288 23166 13297
rect 23110 13223 23166 13232
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 23032 9722 23060 10066
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22558 9007 22614 9016
rect 22744 9036 22796 9042
rect 22468 8978 22520 8984
rect 22744 8978 22796 8984
rect 22480 8294 22508 8978
rect 22848 8634 22876 9114
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22558 8392 22614 8401
rect 22558 8327 22614 8336
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22374 6080 22430 6089
rect 22374 6015 22430 6024
rect 22480 4593 22508 8230
rect 22572 7410 22600 8327
rect 23124 8090 23152 13223
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12986 23336 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23294 12744 23350 12753
rect 23294 12679 23350 12688
rect 23204 12368 23256 12374
rect 23204 12310 23256 12316
rect 23308 12322 23336 12679
rect 23400 12442 23428 12786
rect 23492 12481 23520 14175
rect 23584 13394 23612 15982
rect 23754 15736 23810 15745
rect 23754 15671 23810 15680
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23676 14550 23704 15438
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23676 13870 23704 14486
rect 23768 14362 23796 15671
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23860 15162 23888 15506
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23860 14482 23888 15098
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23768 14334 23888 14362
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13938 23796 14214
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23676 13172 23704 13806
rect 23584 13144 23704 13172
rect 23756 13184 23808 13190
rect 23478 12472 23534 12481
rect 23388 12436 23440 12442
rect 23478 12407 23534 12416
rect 23388 12378 23440 12384
rect 23216 11762 23244 12310
rect 23308 12294 23520 12322
rect 23492 11898 23520 12294
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23216 11354 23244 11698
rect 23478 11384 23534 11393
rect 23204 11348 23256 11354
rect 23478 11319 23534 11328
rect 23204 11290 23256 11296
rect 23492 10810 23520 11319
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23216 8634 23244 8910
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22664 7546 22692 7890
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 23308 6905 23336 9658
rect 23492 8378 23520 10542
rect 23400 8350 23520 8378
rect 23400 7206 23428 8350
rect 23478 8256 23534 8265
rect 23478 8191 23534 8200
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23294 6896 23350 6905
rect 23294 6831 23350 6840
rect 23492 5137 23520 8191
rect 23584 7698 23612 13144
rect 23756 13126 23808 13132
rect 23662 12608 23718 12617
rect 23662 12543 23718 12552
rect 23676 11898 23704 12543
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23662 11656 23718 11665
rect 23662 11591 23718 11600
rect 23676 8945 23704 11591
rect 23662 8936 23718 8945
rect 23662 8871 23718 8880
rect 23662 8664 23718 8673
rect 23662 8599 23718 8608
rect 23676 7818 23704 8599
rect 23768 7954 23796 13126
rect 23860 10554 23888 14334
rect 23952 10690 23980 20810
rect 24032 20596 24084 20602
rect 24032 20538 24084 20544
rect 24044 15502 24072 20538
rect 24136 16153 24164 20998
rect 24228 20874 24256 21100
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24216 20868 24268 20874
rect 24216 20810 24268 20816
rect 24228 19718 24256 20810
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24320 19854 24348 20402
rect 24688 20262 24716 20946
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24872 20505 24900 20878
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24858 20496 24914 20505
rect 24858 20431 24914 20440
rect 24964 20346 24992 20742
rect 24780 20330 24992 20346
rect 24768 20324 24992 20330
rect 24820 20318 24992 20324
rect 24768 20266 24820 20272
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24308 19848 24360 19854
rect 24308 19790 24360 19796
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24674 19680 24730 19689
rect 24289 19612 24585 19632
rect 24674 19615 24730 19624
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24306 19408 24362 19417
rect 24306 19343 24362 19352
rect 24320 18698 24348 19343
rect 24308 18692 24360 18698
rect 24308 18634 24360 18640
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24228 18290 24256 18566
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17066 24256 17478
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17060 24268 17066
rect 24216 17002 24268 17008
rect 24122 16144 24178 16153
rect 24122 16079 24178 16088
rect 24228 15910 24256 17002
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24412 16697 24440 16730
rect 24398 16688 24454 16697
rect 24398 16623 24454 16632
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 15904 24268 15910
rect 24216 15846 24268 15852
rect 24124 15632 24176 15638
rect 24124 15574 24176 15580
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 24044 13530 24072 15302
rect 24136 15094 24164 15574
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24124 15088 24176 15094
rect 24124 15030 24176 15036
rect 24136 14414 24164 15030
rect 24228 14822 24256 15370
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 19615
rect 24780 18970 24808 20266
rect 25056 20058 25084 22607
rect 25148 22001 25176 24618
rect 25240 23497 25268 24686
rect 25332 24410 25360 27095
rect 25596 25356 25648 25362
rect 25596 25298 25648 25304
rect 25410 24848 25466 24857
rect 25410 24783 25466 24792
rect 25424 24614 25452 24783
rect 25608 24682 25636 25298
rect 25596 24676 25648 24682
rect 25596 24618 25648 24624
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 25226 23488 25282 23497
rect 25226 23423 25282 23432
rect 25332 23322 25360 24346
rect 25780 24200 25832 24206
rect 25780 24142 25832 24148
rect 25410 24032 25466 24041
rect 25410 23967 25466 23976
rect 25424 23866 25452 23967
rect 25792 23866 25820 24142
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25780 23860 25832 23866
rect 25780 23802 25832 23808
rect 25778 23760 25834 23769
rect 25778 23695 25834 23704
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25320 23316 25372 23322
rect 25320 23258 25372 23264
rect 25608 22982 25636 23598
rect 25688 23316 25740 23322
rect 25688 23258 25740 23264
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25228 22568 25280 22574
rect 25226 22536 25228 22545
rect 25280 22536 25282 22545
rect 25226 22471 25282 22480
rect 25502 22536 25558 22545
rect 25502 22471 25558 22480
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25134 21992 25190 22001
rect 25134 21927 25190 21936
rect 25240 21332 25268 22034
rect 25410 21992 25466 22001
rect 25410 21927 25466 21936
rect 25320 21480 25372 21486
rect 25318 21448 25320 21457
rect 25372 21448 25374 21457
rect 25318 21383 25374 21392
rect 25240 21304 25360 21332
rect 25332 20806 25360 21304
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25056 19514 25084 19994
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 25148 19446 25176 19790
rect 25136 19440 25188 19446
rect 25136 19382 25188 19388
rect 25148 19310 25176 19382
rect 25136 19304 25188 19310
rect 25240 19281 25268 20334
rect 25332 19394 25360 20742
rect 25424 20602 25452 21927
rect 25516 21690 25544 22471
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25502 21448 25558 21457
rect 25502 21383 25558 21392
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25332 19366 25452 19394
rect 25136 19246 25188 19252
rect 25226 19272 25282 19281
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 24766 18592 24822 18601
rect 24766 18527 24822 18536
rect 24780 15722 24808 18527
rect 24964 17542 24992 18770
rect 25148 18698 25176 19246
rect 25226 19207 25282 19216
rect 25240 18970 25268 19207
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25240 18426 25268 18906
rect 25228 18420 25280 18426
rect 25228 18362 25280 18368
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25240 17542 25268 18158
rect 25320 17740 25372 17746
rect 25320 17682 25372 17688
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 24780 15694 24900 15722
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24136 14006 24164 14350
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24124 13864 24176 13870
rect 24122 13832 24124 13841
rect 24176 13832 24178 13841
rect 24122 13767 24178 13776
rect 24228 13716 24256 14758
rect 24780 14618 24808 15506
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 13734 24716 14418
rect 24872 14074 24900 15694
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24964 13954 24992 17478
rect 25044 16992 25096 16998
rect 25042 16960 25044 16969
rect 25096 16960 25098 16969
rect 25042 16895 25098 16904
rect 25148 16833 25176 17478
rect 25332 16998 25360 17682
rect 25320 16992 25372 16998
rect 25320 16934 25372 16940
rect 25134 16824 25190 16833
rect 25134 16759 25190 16768
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25240 15502 25268 15846
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25240 15094 25268 15438
rect 25228 15088 25280 15094
rect 25228 15030 25280 15036
rect 25226 14920 25282 14929
rect 25226 14855 25282 14864
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 24872 13926 24992 13954
rect 25148 13938 25176 14418
rect 25136 13932 25188 13938
rect 24136 13688 24256 13716
rect 24676 13728 24728 13734
rect 24674 13696 24676 13705
rect 24728 13696 24730 13705
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24044 12986 24072 13330
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 24030 11928 24086 11937
rect 24030 11863 24086 11872
rect 24044 11694 24072 11863
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 24044 11354 24072 11630
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 24044 10810 24072 10950
rect 24032 10804 24084 10810
rect 24032 10746 24084 10752
rect 23952 10662 24072 10690
rect 23860 10526 23980 10554
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 9926 23888 10406
rect 23952 9994 23980 10526
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23848 9920 23900 9926
rect 23846 9888 23848 9897
rect 23900 9888 23902 9897
rect 23846 9823 23902 9832
rect 24044 8401 24072 10662
rect 24136 8498 24164 13688
rect 24674 13631 24730 13640
rect 24766 13424 24822 13433
rect 24766 13359 24822 13368
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24320 12442 24348 12786
rect 24504 12481 24532 12854
rect 24490 12472 24546 12481
rect 24308 12436 24360 12442
rect 24490 12407 24546 12416
rect 24674 12472 24730 12481
rect 24674 12407 24676 12416
rect 24308 12378 24360 12384
rect 24728 12407 24730 12416
rect 24676 12378 24728 12384
rect 24674 12336 24730 12345
rect 24674 12271 24730 12280
rect 24398 12200 24454 12209
rect 24398 12135 24400 12144
rect 24452 12135 24454 12144
rect 24400 12106 24452 12112
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24320 11529 24348 11698
rect 24306 11520 24362 11529
rect 24306 11455 24362 11464
rect 24320 11354 24348 11455
rect 24688 11393 24716 12271
rect 24674 11384 24730 11393
rect 24308 11348 24360 11354
rect 24674 11319 24730 11328
rect 24308 11290 24360 11296
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24228 10538 24256 11018
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24676 10736 24728 10742
rect 24676 10678 24728 10684
rect 24306 10568 24362 10577
rect 24216 10532 24268 10538
rect 24306 10503 24362 10512
rect 24216 10474 24268 10480
rect 24228 10266 24256 10474
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24320 10146 24348 10503
rect 24228 10118 24348 10146
rect 24228 8514 24256 10118
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9654 24716 10678
rect 24676 9648 24728 9654
rect 24676 9590 24728 9596
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24596 9217 24624 9454
rect 24582 9208 24638 9217
rect 24780 9178 24808 13359
rect 24582 9143 24638 9152
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24872 9058 24900 13926
rect 25136 13874 25188 13880
rect 25044 13456 25096 13462
rect 25044 13398 25096 13404
rect 25056 12986 25084 13398
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25056 12345 25084 12718
rect 25042 12336 25098 12345
rect 25042 12271 25098 12280
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25056 11898 25084 12174
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25148 11286 25176 13874
rect 25240 13870 25268 14855
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25240 13297 25268 13330
rect 25226 13288 25282 13297
rect 25226 13223 25282 13232
rect 25240 12986 25268 13223
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25226 12880 25282 12889
rect 25226 12815 25282 12824
rect 25240 11354 25268 12815
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25136 11280 25188 11286
rect 25136 11222 25188 11228
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 25136 11008 25188 11014
rect 25136 10950 25188 10956
rect 24964 10792 24992 10950
rect 24964 10764 25084 10792
rect 24950 10704 25006 10713
rect 24950 10639 25006 10648
rect 24964 10033 24992 10639
rect 25056 10606 25084 10764
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 24950 10024 25006 10033
rect 24950 9959 25006 9968
rect 25148 9926 25176 10950
rect 25240 10810 25268 11290
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 9920 25188 9926
rect 25134 9888 25136 9897
rect 25188 9888 25190 9897
rect 25134 9823 25190 9832
rect 24676 9036 24728 9042
rect 24676 8978 24728 8984
rect 24780 9030 24900 9058
rect 25042 9072 25098 9081
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24124 8492 24176 8498
rect 24228 8486 24348 8514
rect 24124 8434 24176 8440
rect 24030 8392 24086 8401
rect 24030 8327 24086 8336
rect 24214 8392 24270 8401
rect 24214 8327 24270 8336
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23756 7948 23808 7954
rect 23756 7890 23808 7896
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23584 7670 23796 7698
rect 23662 7576 23718 7585
rect 23662 7511 23718 7520
rect 23676 7342 23704 7511
rect 23768 7426 23796 7670
rect 23860 7546 23888 8230
rect 23938 8120 23994 8129
rect 23938 8055 23940 8064
rect 23992 8055 23994 8064
rect 23940 8026 23992 8032
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 23848 7540 23900 7546
rect 23848 7482 23900 7488
rect 23768 7398 23888 7426
rect 23952 7410 23980 7754
rect 24136 7546 24164 7890
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 23664 7336 23716 7342
rect 23570 7304 23626 7313
rect 23664 7278 23716 7284
rect 23570 7239 23626 7248
rect 23478 5128 23534 5137
rect 23478 5063 23534 5072
rect 22466 4584 22522 4593
rect 22466 4519 22522 4528
rect 23478 4176 23534 4185
rect 23478 4111 23534 4120
rect 23202 3496 23258 3505
rect 23202 3431 23258 3440
rect 21638 2544 21694 2553
rect 21638 2479 21694 2488
rect 17498 1728 17554 1737
rect 17498 1663 17554 1672
rect 16486 1592 16542 1601
rect 16486 1527 16542 1536
rect 23216 480 23244 3431
rect 23492 921 23520 4111
rect 23584 2009 23612 7239
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23676 3641 23704 7142
rect 23754 6896 23810 6905
rect 23754 6831 23756 6840
rect 23808 6831 23810 6840
rect 23756 6802 23808 6808
rect 23768 6458 23796 6802
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23662 3632 23718 3641
rect 23662 3567 23718 3576
rect 23570 2000 23626 2009
rect 23570 1935 23626 1944
rect 23478 912 23534 921
rect 23478 847 23534 856
rect 3146 368 3202 377
rect 3146 303 3202 312
rect 4618 0 4674 480
rect 13910 0 13966 480
rect 23202 0 23258 480
rect 23860 377 23888 7398
rect 23940 7404 23992 7410
rect 23940 7346 23992 7352
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 23938 6760 23994 6769
rect 23938 6695 23940 6704
rect 23992 6695 23994 6704
rect 23940 6666 23992 6672
rect 24136 4593 24164 7346
rect 24228 7177 24256 8327
rect 24320 7857 24348 8486
rect 24688 8294 24716 8978
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24674 7984 24730 7993
rect 24674 7919 24676 7928
rect 24728 7919 24730 7928
rect 24676 7890 24728 7896
rect 24306 7848 24362 7857
rect 24306 7783 24362 7792
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24688 7546 24716 7890
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24674 7440 24730 7449
rect 24674 7375 24730 7384
rect 24688 7342 24716 7375
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24214 7168 24270 7177
rect 24214 7103 24270 7112
rect 24780 6866 24808 9030
rect 25042 9007 25098 9016
rect 25056 8430 25084 9007
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 25332 7478 25360 16934
rect 25424 15473 25452 19366
rect 25516 18426 25544 21383
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25410 15464 25466 15473
rect 25410 15399 25466 15408
rect 25608 14618 25636 22918
rect 25700 19417 25728 23258
rect 25792 21350 25820 23695
rect 25884 21962 25912 27520
rect 26528 24426 26556 27520
rect 27080 24857 27108 27520
rect 27066 24848 27122 24857
rect 27066 24783 27122 24792
rect 26160 24398 26556 24426
rect 26160 22778 26188 24398
rect 27632 24041 27660 27520
rect 27618 24032 27674 24041
rect 27618 23967 27674 23976
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 25872 21956 25924 21962
rect 25872 21898 25924 21904
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25686 19408 25742 19417
rect 25686 19343 25742 19352
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25792 18426 25820 18702
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25686 17504 25742 17513
rect 25686 17439 25742 17448
rect 25596 14612 25648 14618
rect 25596 14554 25648 14560
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25516 12889 25544 13126
rect 25502 12880 25558 12889
rect 25502 12815 25558 12824
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25424 12447 25452 12582
rect 25410 12438 25466 12447
rect 25410 12373 25466 12382
rect 25596 12300 25648 12306
rect 25596 12242 25648 12248
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25502 12200 25558 12209
rect 25424 11762 25452 12174
rect 25502 12135 25558 12144
rect 25412 11756 25464 11762
rect 25412 11698 25464 11704
rect 25410 11112 25466 11121
rect 25410 11047 25466 11056
rect 25424 8634 25452 11047
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25516 8129 25544 12135
rect 25608 11286 25636 12242
rect 25700 11898 25728 17439
rect 25778 16280 25834 16289
rect 25778 16215 25834 16224
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25596 11280 25648 11286
rect 25594 11248 25596 11257
rect 25648 11248 25650 11257
rect 25594 11183 25650 11192
rect 25792 10810 25820 16215
rect 25884 13258 25912 20198
rect 26238 18728 26294 18737
rect 26238 18663 26294 18672
rect 26252 18426 26280 18663
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25884 10810 25912 13194
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25872 10804 25924 10810
rect 25872 10746 25924 10752
rect 25884 10606 25912 10746
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 25502 8120 25558 8129
rect 25976 8090 26004 17478
rect 26054 13968 26110 13977
rect 26054 13903 26110 13912
rect 26068 10742 26096 13903
rect 26056 10736 26108 10742
rect 26056 10678 26108 10684
rect 25502 8055 25558 8064
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 25320 7472 25372 7478
rect 25320 7414 25372 7420
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24766 5264 24822 5273
rect 24766 5199 24822 5208
rect 24122 4584 24178 4593
rect 24122 4519 24178 4528
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24780 3233 24808 5199
rect 24766 3224 24822 3233
rect 24766 3159 24822 3168
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23846 368 23902 377
rect 23846 303 23902 312
<< via2 >>
rect 4158 27648 4214 27704
rect 1858 26560 1914 26616
rect 1122 20304 1178 20360
rect 846 18944 902 19000
rect 1306 25336 1362 25392
rect 1766 25200 1822 25256
rect 1582 23296 1638 23352
rect 1950 23044 2006 23080
rect 1950 23024 1952 23044
rect 1952 23024 2004 23044
rect 2004 23024 2006 23044
rect 1490 20032 1546 20088
rect 1674 19896 1730 19952
rect 1582 17448 1638 17504
rect 1582 17176 1638 17232
rect 1582 15680 1638 15736
rect 2134 24656 2190 24712
rect 2502 22752 2558 22808
rect 2042 21548 2098 21584
rect 2042 21528 2044 21548
rect 2044 21528 2096 21548
rect 2096 21528 2098 21548
rect 2410 21800 2466 21856
rect 2778 24792 2834 24848
rect 2870 24248 2926 24304
rect 2778 23468 2780 23488
rect 2780 23468 2832 23488
rect 2832 23468 2834 23488
rect 2778 23432 2834 23468
rect 2686 22208 2742 22264
rect 2778 21392 2834 21448
rect 3054 25336 3110 25392
rect 3054 21936 3110 21992
rect 2410 20440 2466 20496
rect 2318 19488 2374 19544
rect 1582 15156 1638 15192
rect 1582 15136 1584 15156
rect 1584 15136 1636 15156
rect 1636 15136 1638 15156
rect 1582 14592 1638 14648
rect 1490 13912 1546 13968
rect 1950 18808 2006 18864
rect 2226 19236 2282 19272
rect 2226 19216 2228 19236
rect 2228 19216 2280 19236
rect 2280 19216 2282 19236
rect 1582 13368 1638 13424
rect 1766 12280 1822 12336
rect 2042 15972 2098 16008
rect 2042 15952 2044 15972
rect 2044 15952 2096 15972
rect 2096 15952 2098 15972
rect 2226 17856 2282 17912
rect 2410 16904 2466 16960
rect 2778 20576 2834 20632
rect 2226 16224 2282 16280
rect 2778 19624 2834 19680
rect 3606 27104 3662 27160
rect 3330 24556 3332 24576
rect 3332 24556 3384 24576
rect 3384 24556 3386 24576
rect 3330 24520 3386 24556
rect 3330 23704 3386 23760
rect 3238 21256 3294 21312
rect 3146 20440 3202 20496
rect 2962 17312 3018 17368
rect 2594 16088 2650 16144
rect 2410 14456 2466 14512
rect 2042 12708 2098 12744
rect 2042 12688 2044 12708
rect 2044 12688 2096 12708
rect 2096 12688 2098 12708
rect 2778 15816 2834 15872
rect 3882 26016 3938 26072
rect 3606 21936 3662 21992
rect 3974 25200 4030 25256
rect 3698 21392 3754 21448
rect 3146 19080 3202 19136
rect 3330 20324 3386 20360
rect 3330 20304 3332 20324
rect 3332 20304 3384 20324
rect 3384 20304 3386 20324
rect 3054 16088 3110 16144
rect 3882 21528 3938 21584
rect 23754 27648 23810 27704
rect 4158 23432 4214 23488
rect 4066 22344 4122 22400
rect 4526 23704 4582 23760
rect 4986 22652 4988 22672
rect 4988 22652 5040 22672
rect 5040 22652 5042 22672
rect 4986 22616 5042 22652
rect 5354 24384 5410 24440
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5998 24792 6054 24848
rect 6642 25880 6698 25936
rect 7010 24792 7066 24848
rect 7286 24812 7342 24848
rect 7286 24792 7288 24812
rect 7288 24792 7340 24812
rect 7340 24792 7342 24812
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5354 23568 5410 23624
rect 4342 21936 4398 21992
rect 4158 21528 4214 21584
rect 4066 21020 4068 21040
rect 4068 21020 4120 21040
rect 4120 21020 4122 21040
rect 4066 20984 4122 21020
rect 3606 19116 3608 19136
rect 3608 19116 3660 19136
rect 3660 19116 3662 19136
rect 3606 19080 3662 19116
rect 3606 18944 3662 19000
rect 3514 18672 3570 18728
rect 2962 14864 3018 14920
rect 2870 14728 2926 14784
rect 2686 12860 2688 12880
rect 2688 12860 2740 12880
rect 2740 12860 2742 12880
rect 2686 12824 2742 12860
rect 3054 13232 3110 13288
rect 3146 12824 3202 12880
rect 3146 12552 3202 12608
rect 2962 11736 3018 11792
rect 2410 10376 2466 10432
rect 3514 15680 3570 15736
rect 3514 14456 3570 14512
rect 3146 9424 3202 9480
rect 2226 9016 2282 9072
rect 3882 18536 3938 18592
rect 3882 17720 3938 17776
rect 4526 21972 4528 21992
rect 4528 21972 4580 21992
rect 4580 21972 4582 21992
rect 4526 21936 4582 21972
rect 4434 21800 4490 21856
rect 4434 21528 4490 21584
rect 4434 20576 4490 20632
rect 4526 19080 4582 19136
rect 3974 17040 4030 17096
rect 4066 16904 4122 16960
rect 3882 16652 3938 16688
rect 4250 16788 4306 16824
rect 4250 16768 4252 16788
rect 4252 16768 4304 16788
rect 4304 16768 4306 16788
rect 3882 16632 3884 16652
rect 3884 16632 3936 16652
rect 3936 16632 3938 16652
rect 4342 15428 4398 15464
rect 4342 15408 4344 15428
rect 4344 15408 4396 15428
rect 4396 15408 4398 15428
rect 4710 17332 4766 17368
rect 4710 17312 4712 17332
rect 4712 17312 4764 17332
rect 4764 17312 4766 17332
rect 5262 22752 5318 22808
rect 6090 23976 6146 24032
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 6458 23296 6514 23352
rect 6090 22344 6146 22400
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6090 21664 6146 21720
rect 5998 21392 6054 21448
rect 6642 24656 6698 24712
rect 7194 24112 7250 24168
rect 6918 22616 6974 22672
rect 7010 22480 7066 22536
rect 5998 21020 6000 21040
rect 6000 21020 6052 21040
rect 6052 21020 6054 21040
rect 5998 20984 6054 21020
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5170 19760 5226 19816
rect 5998 19896 6054 19952
rect 5446 19488 5502 19544
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5538 19352 5594 19408
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5814 18028 5816 18048
rect 5816 18028 5868 18048
rect 5868 18028 5870 18048
rect 5814 17992 5870 18028
rect 5354 17584 5410 17640
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 4526 14456 4582 14512
rect 4710 13912 4766 13968
rect 4986 16904 5042 16960
rect 4986 16496 5042 16552
rect 4710 12416 4766 12472
rect 4434 11328 4490 11384
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6734 21392 6790 21448
rect 6182 17992 6238 18048
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5538 15000 5594 15056
rect 5354 14356 5356 14376
rect 5356 14356 5408 14376
rect 5408 14356 5410 14376
rect 5354 14320 5410 14356
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5630 12824 5686 12880
rect 6366 16088 6422 16144
rect 6826 20712 6882 20768
rect 7010 20440 7066 20496
rect 6826 20032 6882 20088
rect 6550 16224 6606 16280
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 4710 11056 4766 11112
rect 6734 17876 6790 17912
rect 6734 17856 6736 17876
rect 6736 17856 6788 17876
rect 6788 17856 6790 17876
rect 7746 23432 7802 23488
rect 7470 22888 7526 22944
rect 7194 22752 7250 22808
rect 7286 21428 7288 21448
rect 7288 21428 7340 21448
rect 7340 21428 7342 21448
rect 7286 21392 7342 21428
rect 7010 17720 7066 17776
rect 7470 18400 7526 18456
rect 7194 17312 7250 17368
rect 7378 17720 7434 17776
rect 7010 15952 7066 16008
rect 7010 15544 7066 15600
rect 7102 13912 7158 13968
rect 8114 24404 8170 24440
rect 8114 24384 8116 24404
rect 8116 24384 8168 24404
rect 8168 24384 8170 24404
rect 8298 24248 8354 24304
rect 8114 23296 8170 23352
rect 8298 23160 8354 23216
rect 8666 23468 8668 23488
rect 8668 23468 8720 23488
rect 8720 23468 8722 23488
rect 8666 23432 8722 23468
rect 8666 23160 8722 23216
rect 8298 21936 8354 21992
rect 7930 21528 7986 21584
rect 7838 19252 7840 19272
rect 7840 19252 7892 19272
rect 7892 19252 7894 19272
rect 7838 19216 7894 19252
rect 7838 18964 7894 19000
rect 7838 18944 7840 18964
rect 7840 18944 7892 18964
rect 7892 18944 7894 18964
rect 7654 17584 7710 17640
rect 7746 17312 7802 17368
rect 7286 14184 7342 14240
rect 7470 15680 7526 15736
rect 7286 13232 7342 13288
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 4066 10648 4122 10704
rect 3882 10376 3938 10432
rect 3606 9424 3662 9480
rect 2962 6840 3018 6896
rect 2962 6024 3018 6080
rect 4066 9968 4122 10024
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 3974 9560 4030 9616
rect 4066 9288 4122 9344
rect 3974 8880 4030 8936
rect 7930 16632 7986 16688
rect 7838 16496 7894 16552
rect 7746 14340 7802 14376
rect 7746 14320 7748 14340
rect 7748 14320 7800 14340
rect 7800 14320 7802 14340
rect 7930 16224 7986 16280
rect 7838 12552 7894 12608
rect 8022 15544 8078 15600
rect 6918 9152 6974 9208
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 9402 25880 9458 25936
rect 8666 20868 8722 20904
rect 8666 20848 8668 20868
rect 8668 20848 8720 20868
rect 8720 20848 8722 20868
rect 8850 20848 8906 20904
rect 8298 19352 8354 19408
rect 8942 19352 8998 19408
rect 8758 18844 8760 18864
rect 8760 18844 8812 18864
rect 8812 18844 8814 18864
rect 8758 18808 8814 18844
rect 8574 18128 8630 18184
rect 8298 17992 8354 18048
rect 8206 16904 8262 16960
rect 8114 14728 8170 14784
rect 8850 16496 8906 16552
rect 8850 15816 8906 15872
rect 8758 15544 8814 15600
rect 8298 15444 8300 15464
rect 8300 15444 8352 15464
rect 8352 15444 8354 15464
rect 8298 15408 8354 15444
rect 8114 13388 8170 13424
rect 8114 13368 8116 13388
rect 8116 13368 8168 13388
rect 8168 13368 8170 13388
rect 8114 13198 8170 13254
rect 8850 15000 8906 15056
rect 8666 13504 8722 13560
rect 8390 11328 8446 11384
rect 9586 21936 9642 21992
rect 9770 21936 9826 21992
rect 9678 20032 9734 20088
rect 9034 15000 9090 15056
rect 9586 19216 9642 19272
rect 9402 18536 9458 18592
rect 9678 19080 9734 19136
rect 9402 17176 9458 17232
rect 9034 13096 9090 13152
rect 9126 12708 9182 12744
rect 9126 12688 9128 12708
rect 9128 12688 9180 12708
rect 9180 12688 9182 12708
rect 9678 17040 9734 17096
rect 9678 16940 9680 16960
rect 9680 16940 9732 16960
rect 9732 16940 9734 16960
rect 9678 16904 9734 16940
rect 9586 14220 9588 14240
rect 9588 14220 9640 14240
rect 9640 14220 9642 14240
rect 9586 14184 9642 14220
rect 9494 12688 9550 12744
rect 9402 11600 9458 11656
rect 9218 11192 9274 11248
rect 7562 8200 7618 8256
rect 8022 8200 8078 8256
rect 7562 7656 7618 7712
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 10046 24520 10102 24576
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10690 25472 10746 25528
rect 10690 24656 10746 24712
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10966 25220 11022 25256
rect 10966 25200 10968 25220
rect 10968 25200 11020 25220
rect 11020 25200 11022 25220
rect 11150 24792 11206 24848
rect 10874 24112 10930 24168
rect 10138 23704 10194 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 11426 24792 11482 24848
rect 11518 24556 11520 24576
rect 11520 24556 11572 24576
rect 11572 24556 11574 24576
rect 11518 24520 11574 24556
rect 11426 24248 11482 24304
rect 11518 23976 11574 24032
rect 10966 23432 11022 23488
rect 11150 23160 11206 23216
rect 11426 23160 11482 23216
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10598 22108 10600 22128
rect 10600 22108 10652 22128
rect 10652 22108 10654 22128
rect 10598 22072 10654 22108
rect 11334 22616 11390 22672
rect 11426 22480 11482 22536
rect 11794 23976 11850 24032
rect 11702 22888 11758 22944
rect 10506 21548 10562 21584
rect 10506 21528 10508 21548
rect 10508 21528 10560 21548
rect 10560 21528 10562 21548
rect 10046 21256 10102 21312
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 9862 18536 9918 18592
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18944 10194 19000
rect 9954 17720 10010 17776
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10138 15680 10194 15736
rect 9954 14184 10010 14240
rect 9862 9324 9864 9344
rect 9864 9324 9916 9344
rect 9916 9324 9918 9344
rect 9862 9288 9918 9324
rect 10598 14884 10654 14920
rect 10598 14864 10600 14884
rect 10600 14864 10652 14884
rect 10652 14864 10654 14884
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10138 14456 10194 14512
rect 10046 12416 10102 12472
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 11058 21664 11114 21720
rect 11058 21256 11114 21312
rect 11610 21256 11666 21312
rect 10966 21020 10968 21040
rect 10968 21020 11020 21040
rect 11020 21020 11022 21040
rect 10966 20984 11022 21020
rect 10874 20576 10930 20632
rect 10874 20340 10876 20360
rect 10876 20340 10928 20360
rect 10928 20340 10930 20360
rect 10874 20304 10930 20340
rect 10874 20168 10930 20224
rect 10782 16768 10838 16824
rect 11058 19352 11114 19408
rect 11518 20748 11520 20768
rect 11520 20748 11572 20768
rect 11572 20748 11574 20768
rect 11518 20712 11574 20748
rect 11610 19796 11612 19816
rect 11612 19796 11664 19816
rect 11664 19796 11666 19816
rect 11610 19760 11666 19796
rect 11150 19116 11152 19136
rect 11152 19116 11204 19136
rect 11204 19116 11206 19136
rect 11150 19080 11206 19116
rect 11242 18708 11244 18728
rect 11244 18708 11296 18728
rect 11296 18708 11298 18728
rect 11242 18672 11298 18708
rect 11426 17196 11482 17232
rect 11426 17176 11428 17196
rect 11428 17176 11480 17196
rect 11480 17176 11482 17196
rect 12070 23740 12072 23760
rect 12072 23740 12124 23760
rect 12124 23740 12126 23760
rect 12070 23704 12126 23740
rect 12070 22480 12126 22536
rect 12254 23840 12310 23896
rect 12438 22888 12494 22944
rect 11978 20440 12034 20496
rect 12438 22208 12494 22264
rect 12714 24656 12770 24712
rect 12714 22380 12716 22400
rect 12716 22380 12768 22400
rect 12768 22380 12770 22400
rect 12714 22344 12770 22380
rect 12622 21428 12624 21448
rect 12624 21428 12676 21448
rect 12676 21428 12678 21448
rect 12622 21392 12678 21428
rect 12070 19624 12126 19680
rect 12622 18672 12678 18728
rect 12622 18400 12678 18456
rect 12530 18264 12586 18320
rect 11702 16652 11758 16688
rect 10874 16224 10930 16280
rect 10782 15816 10838 15872
rect 10966 15700 11022 15736
rect 10966 15680 10968 15700
rect 10968 15680 11020 15700
rect 11020 15680 11022 15700
rect 11058 15408 11114 15464
rect 10782 15272 10838 15328
rect 11702 16632 11704 16652
rect 11704 16632 11756 16652
rect 11756 16632 11758 16652
rect 10782 13504 10838 13560
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10046 11056 10102 11112
rect 10138 10376 10194 10432
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10046 10104 10102 10160
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11426 12824 11482 12880
rect 11426 12164 11482 12200
rect 11426 12144 11428 12164
rect 11428 12144 11480 12164
rect 11480 12144 11482 12164
rect 11150 11736 11206 11792
rect 11702 12008 11758 12064
rect 11794 11620 11850 11656
rect 11794 11600 11796 11620
rect 11796 11600 11848 11620
rect 11848 11600 11850 11620
rect 11426 9696 11482 9752
rect 10782 7928 10838 7984
rect 9770 7384 9826 7440
rect 4066 7112 4122 7168
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 4066 5344 4122 5400
rect 3882 4800 3938 4856
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 4066 4528 4122 4584
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 3974 3984 4030 4040
rect 3330 3576 3386 3632
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 4066 3712 4122 3768
rect 3974 3168 4030 3224
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 4066 3032 4122 3088
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 3514 2624 3570 2680
rect 11702 2488 11758 2544
rect 4618 2352 4674 2408
rect 3514 1536 3570 1592
rect 3330 856 3386 912
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 11886 3576 11942 3632
rect 12990 23296 13046 23352
rect 12898 22752 12954 22808
rect 12806 15700 12862 15736
rect 12806 15680 12808 15700
rect 12808 15680 12860 15700
rect 12860 15680 12862 15700
rect 12898 15000 12954 15056
rect 12162 14320 12218 14376
rect 12346 14340 12402 14376
rect 12346 14320 12348 14340
rect 12348 14320 12400 14340
rect 12400 14320 12402 14340
rect 13174 20848 13230 20904
rect 13082 17312 13138 17368
rect 14922 25744 14978 25800
rect 13450 23432 13506 23488
rect 13542 22616 13598 22672
rect 13358 21528 13414 21584
rect 13910 24792 13966 24848
rect 13726 24656 13782 24712
rect 13910 24384 13966 24440
rect 13726 24148 13728 24168
rect 13728 24148 13780 24168
rect 13780 24148 13782 24168
rect 13726 24112 13782 24148
rect 14002 23976 14058 24032
rect 14370 24792 14426 24848
rect 14094 23024 14150 23080
rect 14278 22480 14334 22536
rect 13818 20984 13874 21040
rect 13634 20848 13690 20904
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 13450 20712 13506 20768
rect 14094 20712 14150 20768
rect 13358 19216 13414 19272
rect 13266 15408 13322 15464
rect 13358 15308 13360 15328
rect 13360 15308 13412 15328
rect 13412 15308 13414 15328
rect 13358 15272 13414 15308
rect 13174 14592 13230 14648
rect 13726 18808 13782 18864
rect 13818 18572 13820 18592
rect 13820 18572 13872 18592
rect 13872 18572 13874 18592
rect 13818 18536 13874 18572
rect 13542 16904 13598 16960
rect 13910 16632 13966 16688
rect 13542 15952 13598 16008
rect 12070 11192 12126 11248
rect 12530 12688 12586 12744
rect 13082 13232 13138 13288
rect 12346 9152 12402 9208
rect 11978 3440 12034 3496
rect 11978 2388 11980 2408
rect 11980 2388 12032 2408
rect 12032 2388 12034 2408
rect 11978 2352 12034 2388
rect 13082 12688 13138 12744
rect 12898 11056 12954 11112
rect 13542 13640 13598 13696
rect 13450 13368 13506 13424
rect 13266 13232 13322 13288
rect 13266 12824 13322 12880
rect 13174 10240 13230 10296
rect 13726 15680 13782 15736
rect 14370 17312 14426 17368
rect 14554 23860 14610 23896
rect 14554 23840 14556 23860
rect 14556 23840 14608 23860
rect 14608 23840 14610 23860
rect 14554 23568 14610 23624
rect 14554 22888 14610 22944
rect 14646 20576 14702 20632
rect 14186 16224 14242 16280
rect 14186 14184 14242 14240
rect 13910 13096 13966 13152
rect 14002 12824 14058 12880
rect 13818 11192 13874 11248
rect 13634 10512 13690 10568
rect 13634 10376 13690 10432
rect 13634 9560 13690 9616
rect 14094 11872 14150 11928
rect 12806 7284 12808 7304
rect 12808 7284 12860 7304
rect 12860 7284 12862 7304
rect 12806 7248 12862 7284
rect 14186 11328 14242 11384
rect 14186 9968 14242 10024
rect 14370 15852 14372 15872
rect 14372 15852 14424 15872
rect 14424 15852 14426 15872
rect 14370 15816 14426 15852
rect 14370 15544 14426 15600
rect 14554 12416 14610 12472
rect 14554 12280 14610 12336
rect 14462 12008 14518 12064
rect 14462 10104 14518 10160
rect 14462 9696 14518 9752
rect 14278 9560 14334 9616
rect 14186 7656 14242 7712
rect 14094 6840 14150 6896
rect 12714 6704 12770 6760
rect 14554 7112 14610 7168
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14830 23296 14886 23352
rect 14922 23024 14978 23080
rect 15106 23060 15108 23080
rect 15108 23060 15160 23080
rect 15160 23060 15162 23080
rect 15106 23024 15162 23060
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15198 22652 15200 22672
rect 15200 22652 15252 22672
rect 15252 22652 15254 22672
rect 15198 22616 15254 22652
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15382 24656 15438 24712
rect 15566 23976 15622 24032
rect 15566 22208 15622 22264
rect 15290 21528 15346 21584
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14830 20032 14886 20088
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15014 19080 15070 19136
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15106 17620 15108 17640
rect 15108 17620 15160 17640
rect 15160 17620 15162 17640
rect 15106 17584 15162 17620
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14830 15816 14886 15872
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15474 15952 15530 16008
rect 15474 15680 15530 15736
rect 15382 14184 15438 14240
rect 15382 13640 15438 13696
rect 15474 13504 15530 13560
rect 15934 24656 15990 24712
rect 15842 24248 15898 24304
rect 15750 23840 15806 23896
rect 15842 21392 15898 21448
rect 17038 25472 17094 25528
rect 17590 25880 17646 25936
rect 17222 25336 17278 25392
rect 16670 24792 16726 24848
rect 16578 24112 16634 24168
rect 16762 24112 16818 24168
rect 16394 22888 16450 22944
rect 17774 24656 17830 24712
rect 17038 23976 17094 24032
rect 17314 23160 17370 23216
rect 16762 23024 16818 23080
rect 17498 23044 17554 23080
rect 17498 23024 17500 23044
rect 17500 23024 17552 23044
rect 17552 23024 17554 23044
rect 16486 22752 16542 22808
rect 16394 21256 16450 21312
rect 15750 16904 15806 16960
rect 15750 15272 15806 15328
rect 16026 15952 16082 16008
rect 15934 15136 15990 15192
rect 15750 13388 15806 13424
rect 15750 13368 15752 13388
rect 15752 13368 15804 13388
rect 15804 13368 15806 13388
rect 15658 11736 15714 11792
rect 15566 11464 15622 11520
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15474 9832 15530 9888
rect 15658 9560 15714 9616
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15382 8336 15438 8392
rect 15106 8200 15162 8256
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14646 6704 14702 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15750 9424 15806 9480
rect 16302 16360 16358 16416
rect 18050 22380 18052 22400
rect 18052 22380 18104 22400
rect 18104 22380 18106 22400
rect 18050 22344 18106 22380
rect 17590 21972 17592 21992
rect 17592 21972 17644 21992
rect 17644 21972 17646 21992
rect 16762 17584 16818 17640
rect 16302 13132 16304 13152
rect 16304 13132 16356 13152
rect 16356 13132 16358 13152
rect 16302 13096 16358 13132
rect 17590 21936 17646 21972
rect 17406 20576 17462 20632
rect 17498 20440 17554 20496
rect 16854 15272 16910 15328
rect 16210 12144 16266 12200
rect 16118 11736 16174 11792
rect 17038 12688 17094 12744
rect 17222 19216 17278 19272
rect 17406 18672 17462 18728
rect 17222 17584 17278 17640
rect 17222 15408 17278 15464
rect 17130 10648 17186 10704
rect 17406 15544 17462 15600
rect 18234 24384 18290 24440
rect 18142 20848 18198 20904
rect 18418 23296 18474 23352
rect 19246 24792 19302 24848
rect 18878 24556 18880 24576
rect 18880 24556 18932 24576
rect 18932 24556 18934 24576
rect 18878 24520 18934 24556
rect 19338 24656 19394 24712
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19522 24248 19578 24304
rect 19430 23432 19486 23488
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 20258 22924 20260 22944
rect 20260 22924 20312 22944
rect 20312 22924 20314 22944
rect 20258 22888 20314 22924
rect 18786 22480 18842 22536
rect 19982 22480 20038 22536
rect 18326 18148 18382 18184
rect 18326 18128 18328 18148
rect 18328 18128 18380 18148
rect 18380 18128 18382 18148
rect 18326 17720 18382 17776
rect 18050 13096 18106 13152
rect 17682 12688 17738 12744
rect 17314 9968 17370 10024
rect 16670 9444 16726 9480
rect 16670 9424 16672 9444
rect 16672 9424 16724 9444
rect 16724 9424 16726 9444
rect 16118 8916 16120 8936
rect 16120 8916 16172 8936
rect 16172 8916 16174 8936
rect 15842 7792 15898 7848
rect 16118 8880 16174 8916
rect 16762 8200 16818 8256
rect 16486 6704 16542 6760
rect 14370 5888 14426 5944
rect 16394 5908 16450 5944
rect 16394 5888 16396 5908
rect 16396 5888 16448 5908
rect 16448 5888 16450 5908
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 11794 1536 11850 1592
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 17038 9288 17094 9344
rect 17038 9016 17094 9072
rect 17406 6840 17462 6896
rect 16854 5208 16910 5264
rect 17958 11772 17960 11792
rect 17960 11772 18012 11792
rect 18012 11772 18014 11792
rect 17958 11736 18014 11772
rect 17866 11464 17922 11520
rect 17682 10648 17738 10704
rect 17958 11348 18014 11384
rect 17958 11328 17960 11348
rect 17960 11328 18012 11348
rect 18012 11328 18014 11348
rect 18878 22072 18934 22128
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19706 21956 19762 21992
rect 19706 21936 19708 21956
rect 19708 21936 19760 21956
rect 19760 21936 19762 21956
rect 19246 21800 19302 21856
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 18510 18128 18566 18184
rect 18694 17176 18750 17232
rect 18694 16632 18750 16688
rect 18510 14864 18566 14920
rect 18510 12688 18566 12744
rect 18142 10920 18198 10976
rect 18878 11872 18934 11928
rect 17866 9560 17922 9616
rect 18602 9696 18658 9752
rect 18510 8900 18566 8936
rect 18510 8880 18512 8900
rect 18512 8880 18564 8900
rect 18564 8880 18566 8900
rect 17682 8064 17738 8120
rect 18142 5072 18198 5128
rect 19522 20440 19578 20496
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19246 17040 19302 17096
rect 19154 16788 19210 16824
rect 19154 16768 19156 16788
rect 19156 16768 19208 16788
rect 19208 16768 19210 16788
rect 20534 19760 20590 19816
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19338 15816 19394 15872
rect 19246 14612 19302 14648
rect 19246 14592 19248 14612
rect 19248 14592 19300 14612
rect 19300 14592 19302 14612
rect 19246 14456 19302 14512
rect 19154 13232 19210 13288
rect 18970 10376 19026 10432
rect 19246 12688 19302 12744
rect 19246 11872 19302 11928
rect 19154 9832 19210 9888
rect 19338 11600 19394 11656
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20074 19080 20130 19136
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19982 15136 20038 15192
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20166 14728 20222 14784
rect 21362 25336 21418 25392
rect 21270 24792 21326 24848
rect 20718 24248 20774 24304
rect 20718 23568 20774 23624
rect 20902 21548 20958 21584
rect 20902 21528 20904 21548
rect 20904 21528 20956 21548
rect 20956 21528 20958 21548
rect 21086 20304 21142 20360
rect 22742 24792 22798 24848
rect 21914 24248 21970 24304
rect 22374 24656 22430 24712
rect 22650 24692 22652 24712
rect 22652 24692 22704 24712
rect 22704 24692 22706 24712
rect 22650 24656 22706 24692
rect 21454 22072 21510 22128
rect 21546 21956 21602 21992
rect 21546 21936 21548 21956
rect 21548 21936 21600 21956
rect 21600 21936 21602 21956
rect 20810 18128 20866 18184
rect 20718 15408 20774 15464
rect 20074 11328 20130 11384
rect 20074 10920 20130 10976
rect 19982 10512 20038 10568
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19982 9832 20038 9888
rect 19522 9560 19578 9616
rect 19430 9288 19486 9344
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19430 8608 19486 8664
rect 19706 8472 19762 8528
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19338 7112 19394 7168
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 18786 6296 18842 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20074 6704 20130 6760
rect 20258 9696 20314 9752
rect 20442 11464 20498 11520
rect 20718 14320 20774 14376
rect 20718 12552 20774 12608
rect 20626 12144 20682 12200
rect 20534 8880 20590 8936
rect 20902 8744 20958 8800
rect 20534 8372 20536 8392
rect 20536 8372 20588 8392
rect 20588 8372 20590 8392
rect 20534 8336 20590 8372
rect 20902 8336 20958 8392
rect 21178 18128 21234 18184
rect 21362 18828 21418 18864
rect 21362 18808 21364 18828
rect 21364 18808 21416 18828
rect 21416 18808 21418 18828
rect 21914 18808 21970 18864
rect 22374 18284 22430 18320
rect 22374 18264 22376 18284
rect 22376 18264 22428 18284
rect 22428 18264 22430 18284
rect 22282 17584 22338 17640
rect 22190 16360 22246 16416
rect 21270 14068 21326 14104
rect 21270 14048 21272 14068
rect 21272 14048 21324 14068
rect 21324 14048 21326 14068
rect 21454 14592 21510 14648
rect 21914 13776 21970 13832
rect 21270 11056 21326 11112
rect 21638 9424 21694 9480
rect 21086 7520 21142 7576
rect 20166 4664 20222 4720
rect 19982 4120 20038 4176
rect 17498 3984 17554 4040
rect 18510 3984 18566 4040
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 17498 3576 17554 3632
rect 17406 3032 17462 3088
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22006 9444 22062 9480
rect 22006 9424 22008 9444
rect 22008 9424 22060 9444
rect 22060 9424 22062 9444
rect 22006 8880 22062 8936
rect 22374 16088 22430 16144
rect 22282 14456 22338 14512
rect 23570 25744 23626 25800
rect 24674 26560 24730 26616
rect 24398 26016 24454 26072
rect 23018 24112 23074 24168
rect 22926 23840 22982 23896
rect 23018 23024 23074 23080
rect 22926 20868 22982 20904
rect 22926 20848 22928 20868
rect 22928 20848 22980 20868
rect 22980 20848 22982 20868
rect 22926 19896 22982 19952
rect 23386 18808 23442 18864
rect 23478 17992 23534 18048
rect 22282 11736 22338 11792
rect 22190 8064 22246 8120
rect 22466 11636 22468 11656
rect 22468 11636 22520 11656
rect 22520 11636 22522 11656
rect 22466 11600 22522 11636
rect 22650 15000 22706 15056
rect 22742 12860 22744 12880
rect 22744 12860 22796 12880
rect 22796 12860 22798 12880
rect 22742 12824 22798 12860
rect 22558 9016 22614 9072
rect 23294 16904 23350 16960
rect 23754 23704 23810 23760
rect 23754 23024 23810 23080
rect 23662 21936 23718 21992
rect 24490 25356 24546 25392
rect 24490 25336 24492 25356
rect 24492 25336 24544 25356
rect 24544 25336 24546 25356
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 25336 24822 25392
rect 25318 27104 25374 27160
rect 25134 24792 25190 24848
rect 24030 23432 24086 23488
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24950 23704 25006 23760
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25042 22616 25098 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 23754 20576 23810 20632
rect 23662 18708 23664 18728
rect 23664 18708 23716 18728
rect 23716 18708 23718 18728
rect 23662 18672 23718 18708
rect 23478 15272 23534 15328
rect 23478 14184 23534 14240
rect 23110 13232 23166 13288
rect 22558 8336 22614 8392
rect 22374 6024 22430 6080
rect 23294 12688 23350 12744
rect 23754 15680 23810 15736
rect 23478 12416 23534 12472
rect 23478 11328 23534 11384
rect 23478 8200 23534 8256
rect 23294 6840 23350 6896
rect 23662 12552 23718 12608
rect 23662 11600 23718 11656
rect 23662 8880 23718 8936
rect 23662 8608 23718 8664
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24858 20440 24914 20496
rect 24674 19624 24730 19680
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24306 19352 24362 19408
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24122 16088 24178 16144
rect 24398 16632 24454 16688
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 25410 24792 25466 24848
rect 25226 23432 25282 23488
rect 25410 23976 25466 24032
rect 25778 23704 25834 23760
rect 25226 22516 25228 22536
rect 25228 22516 25280 22536
rect 25280 22516 25282 22536
rect 25226 22480 25282 22516
rect 25502 22480 25558 22536
rect 25134 21936 25190 21992
rect 25410 21936 25466 21992
rect 25318 21428 25320 21448
rect 25320 21428 25372 21448
rect 25372 21428 25374 21448
rect 25318 21392 25374 21428
rect 25502 21392 25558 21448
rect 24766 18536 24822 18592
rect 25226 19216 25282 19272
rect 24122 13812 24124 13832
rect 24124 13812 24176 13832
rect 24176 13812 24178 13832
rect 24122 13776 24178 13812
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25042 16940 25044 16960
rect 25044 16940 25096 16960
rect 25096 16940 25098 16960
rect 25042 16904 25098 16940
rect 25134 16768 25190 16824
rect 25226 14864 25282 14920
rect 24030 11872 24086 11928
rect 23846 9868 23848 9888
rect 23848 9868 23900 9888
rect 23900 9868 23902 9888
rect 23846 9832 23902 9868
rect 24674 13676 24676 13696
rect 24676 13676 24728 13696
rect 24728 13676 24730 13696
rect 24674 13640 24730 13676
rect 24766 13368 24822 13424
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24490 12416 24546 12472
rect 24674 12436 24730 12472
rect 24674 12416 24676 12436
rect 24676 12416 24728 12436
rect 24728 12416 24730 12436
rect 24674 12280 24730 12336
rect 24398 12164 24454 12200
rect 24398 12144 24400 12164
rect 24400 12144 24452 12164
rect 24452 12144 24454 12164
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24306 11464 24362 11520
rect 24674 11328 24730 11384
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24306 10512 24362 10568
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24582 9152 24638 9208
rect 25042 12280 25098 12336
rect 25226 13232 25282 13288
rect 25226 12824 25282 12880
rect 24950 10648 25006 10704
rect 24950 9968 25006 10024
rect 25134 9868 25136 9888
rect 25136 9868 25188 9888
rect 25188 9868 25190 9888
rect 25134 9832 25190 9868
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24030 8336 24086 8392
rect 24214 8336 24270 8392
rect 23662 7520 23718 7576
rect 23938 8084 23994 8120
rect 23938 8064 23940 8084
rect 23940 8064 23992 8084
rect 23992 8064 23994 8084
rect 23570 7248 23626 7304
rect 23478 5072 23534 5128
rect 22466 4528 22522 4584
rect 23478 4120 23534 4176
rect 23202 3440 23258 3496
rect 21638 2488 21694 2544
rect 17498 1672 17554 1728
rect 16486 1536 16542 1592
rect 23754 6860 23810 6896
rect 23754 6840 23756 6860
rect 23756 6840 23808 6860
rect 23808 6840 23810 6860
rect 23662 3576 23718 3632
rect 23570 1944 23626 2000
rect 23478 856 23534 912
rect 3146 312 3202 368
rect 23938 6724 23994 6760
rect 23938 6704 23940 6724
rect 23940 6704 23992 6724
rect 23992 6704 23994 6724
rect 24674 7948 24730 7984
rect 24674 7928 24676 7948
rect 24676 7928 24728 7948
rect 24728 7928 24730 7948
rect 24306 7792 24362 7848
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24674 7384 24730 7440
rect 24214 7112 24270 7168
rect 25042 9016 25098 9072
rect 25410 15408 25466 15464
rect 27066 24792 27122 24848
rect 27618 23976 27674 24032
rect 25686 19352 25742 19408
rect 25686 17448 25742 17504
rect 25502 12824 25558 12880
rect 25410 12382 25466 12438
rect 25502 12144 25558 12200
rect 25410 11056 25466 11112
rect 25778 16224 25834 16280
rect 25594 11228 25596 11248
rect 25596 11228 25648 11248
rect 25648 11228 25650 11248
rect 25594 11192 25650 11228
rect 26238 18672 26294 18728
rect 25502 8064 25558 8120
rect 26054 13912 26110 13968
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24766 5208 24822 5264
rect 24122 4528 24178 4584
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24766 3168 24822 3224
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23846 312 23902 368
<< metal3 >>
rect 0 27706 480 27736
rect 4153 27706 4219 27709
rect 0 27704 4219 27706
rect 0 27648 4158 27704
rect 4214 27648 4219 27704
rect 0 27646 4219 27648
rect 0 27616 480 27646
rect 4153 27643 4219 27646
rect 23749 27706 23815 27709
rect 27520 27706 28000 27736
rect 23749 27704 28000 27706
rect 23749 27648 23754 27704
rect 23810 27648 28000 27704
rect 23749 27646 28000 27648
rect 23749 27643 23815 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 3601 27162 3667 27165
rect 0 27160 3667 27162
rect 0 27104 3606 27160
rect 3662 27104 3667 27160
rect 0 27102 3667 27104
rect 0 27072 480 27102
rect 3601 27099 3667 27102
rect 25313 27162 25379 27165
rect 27520 27162 28000 27192
rect 25313 27160 28000 27162
rect 25313 27104 25318 27160
rect 25374 27104 28000 27160
rect 25313 27102 28000 27104
rect 25313 27099 25379 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 1853 26618 1919 26621
rect 0 26616 1919 26618
rect 0 26560 1858 26616
rect 1914 26560 1919 26616
rect 0 26558 1919 26560
rect 0 26528 480 26558
rect 1853 26555 1919 26558
rect 24669 26618 24735 26621
rect 27520 26618 28000 26648
rect 24669 26616 28000 26618
rect 24669 26560 24674 26616
rect 24730 26560 28000 26616
rect 24669 26558 28000 26560
rect 24669 26555 24735 26558
rect 27520 26528 28000 26558
rect 0 26074 480 26104
rect 3877 26074 3943 26077
rect 0 26072 3943 26074
rect 0 26016 3882 26072
rect 3938 26016 3943 26072
rect 0 26014 3943 26016
rect 0 25984 480 26014
rect 3877 26011 3943 26014
rect 24393 26074 24459 26077
rect 27520 26074 28000 26104
rect 24393 26072 28000 26074
rect 24393 26016 24398 26072
rect 24454 26016 28000 26072
rect 24393 26014 28000 26016
rect 24393 26011 24459 26014
rect 27520 25984 28000 26014
rect 6637 25938 6703 25941
rect 9397 25938 9463 25941
rect 17585 25938 17651 25941
rect 6637 25936 17651 25938
rect 6637 25880 6642 25936
rect 6698 25880 9402 25936
rect 9458 25880 17590 25936
rect 17646 25880 17651 25936
rect 6637 25878 17651 25880
rect 6637 25875 6703 25878
rect 9397 25875 9463 25878
rect 17585 25875 17651 25878
rect 14917 25802 14983 25805
rect 23565 25802 23631 25805
rect 14917 25800 23631 25802
rect 14917 25744 14922 25800
rect 14978 25744 23570 25800
rect 23626 25744 23631 25800
rect 14917 25742 23631 25744
rect 14917 25739 14983 25742
rect 23565 25739 23631 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 10685 25530 10751 25533
rect 17033 25530 17099 25533
rect 10685 25528 17099 25530
rect 10685 25472 10690 25528
rect 10746 25472 17038 25528
rect 17094 25472 17099 25528
rect 10685 25470 17099 25472
rect 10685 25467 10751 25470
rect 17033 25467 17099 25470
rect 0 25394 480 25424
rect 1301 25394 1367 25397
rect 0 25392 1367 25394
rect 0 25336 1306 25392
rect 1362 25336 1367 25392
rect 0 25334 1367 25336
rect 0 25304 480 25334
rect 1301 25331 1367 25334
rect 3049 25394 3115 25397
rect 9622 25394 9628 25396
rect 3049 25392 9628 25394
rect 3049 25336 3054 25392
rect 3110 25336 9628 25392
rect 3049 25334 9628 25336
rect 3049 25331 3115 25334
rect 9622 25332 9628 25334
rect 9692 25394 9698 25396
rect 17217 25394 17283 25397
rect 9692 25392 17283 25394
rect 9692 25336 17222 25392
rect 17278 25336 17283 25392
rect 9692 25334 17283 25336
rect 9692 25332 9698 25334
rect 17217 25331 17283 25334
rect 21357 25394 21423 25397
rect 24485 25394 24551 25397
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 21357 25392 28000 25394
rect 21357 25336 21362 25392
rect 21418 25336 24490 25392
rect 24546 25336 24766 25392
rect 24822 25336 28000 25392
rect 21357 25334 28000 25336
rect 21357 25331 21423 25334
rect 24485 25331 24551 25334
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 1761 25258 1827 25261
rect 3969 25258 4035 25261
rect 1761 25256 4035 25258
rect 1761 25200 1766 25256
rect 1822 25200 3974 25256
rect 4030 25200 4035 25256
rect 1761 25198 4035 25200
rect 1761 25195 1827 25198
rect 3969 25195 4035 25198
rect 10961 25258 11027 25261
rect 23790 25258 23796 25260
rect 10961 25256 23796 25258
rect 10961 25200 10966 25256
rect 11022 25200 23796 25256
rect 10961 25198 23796 25200
rect 10961 25195 11027 25198
rect 23790 25196 23796 25198
rect 23860 25196 23866 25260
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 2773 24850 2839 24853
rect 0 24848 2839 24850
rect 0 24792 2778 24848
rect 2834 24792 2839 24848
rect 0 24790 2839 24792
rect 0 24760 480 24790
rect 2773 24787 2839 24790
rect 5993 24850 6059 24853
rect 7005 24850 7071 24853
rect 5993 24848 7071 24850
rect 5993 24792 5998 24848
rect 6054 24792 7010 24848
rect 7066 24792 7071 24848
rect 5993 24790 7071 24792
rect 5993 24787 6059 24790
rect 7005 24787 7071 24790
rect 7281 24850 7347 24853
rect 11145 24850 11211 24853
rect 7281 24848 11211 24850
rect 7281 24792 7286 24848
rect 7342 24792 11150 24848
rect 11206 24792 11211 24848
rect 7281 24790 11211 24792
rect 7281 24787 7347 24790
rect 11145 24787 11211 24790
rect 11421 24850 11487 24853
rect 13905 24850 13971 24853
rect 11421 24848 13971 24850
rect 11421 24792 11426 24848
rect 11482 24792 13910 24848
rect 13966 24792 13971 24848
rect 11421 24790 13971 24792
rect 11421 24787 11487 24790
rect 13905 24787 13971 24790
rect 14365 24850 14431 24853
rect 16665 24850 16731 24853
rect 14365 24848 16731 24850
rect 14365 24792 14370 24848
rect 14426 24792 16670 24848
rect 16726 24792 16731 24848
rect 14365 24790 16731 24792
rect 14365 24787 14431 24790
rect 16665 24787 16731 24790
rect 19241 24850 19307 24853
rect 21265 24850 21331 24853
rect 19241 24848 21331 24850
rect 19241 24792 19246 24848
rect 19302 24792 21270 24848
rect 21326 24792 21331 24848
rect 19241 24790 21331 24792
rect 19241 24787 19307 24790
rect 21265 24787 21331 24790
rect 22737 24850 22803 24853
rect 25129 24850 25195 24853
rect 22737 24848 25195 24850
rect 22737 24792 22742 24848
rect 22798 24792 25134 24848
rect 25190 24792 25195 24848
rect 22737 24790 25195 24792
rect 22737 24787 22803 24790
rect 25129 24787 25195 24790
rect 25405 24850 25471 24853
rect 27061 24850 27127 24853
rect 27520 24850 28000 24880
rect 25405 24848 27127 24850
rect 25405 24792 25410 24848
rect 25466 24792 27066 24848
rect 27122 24792 27127 24848
rect 25405 24790 27127 24792
rect 25405 24787 25471 24790
rect 27061 24787 27127 24790
rect 27294 24790 28000 24850
rect 2129 24714 2195 24717
rect 6637 24714 6703 24717
rect 2129 24712 6703 24714
rect 2129 24656 2134 24712
rect 2190 24656 6642 24712
rect 6698 24656 6703 24712
rect 2129 24654 6703 24656
rect 2129 24651 2195 24654
rect 6637 24651 6703 24654
rect 10685 24714 10751 24717
rect 12709 24714 12775 24717
rect 10685 24712 12775 24714
rect 10685 24656 10690 24712
rect 10746 24656 12714 24712
rect 12770 24656 12775 24712
rect 10685 24654 12775 24656
rect 10685 24651 10751 24654
rect 12709 24651 12775 24654
rect 13721 24714 13787 24717
rect 15377 24714 15443 24717
rect 13721 24712 15443 24714
rect 13721 24656 13726 24712
rect 13782 24656 15382 24712
rect 15438 24656 15443 24712
rect 13721 24654 15443 24656
rect 13721 24651 13787 24654
rect 15377 24651 15443 24654
rect 15929 24714 15995 24717
rect 17769 24714 17835 24717
rect 15929 24712 17835 24714
rect 15929 24656 15934 24712
rect 15990 24656 17774 24712
rect 17830 24656 17835 24712
rect 15929 24654 17835 24656
rect 15929 24651 15995 24654
rect 17769 24651 17835 24654
rect 19333 24714 19399 24717
rect 22369 24714 22435 24717
rect 19333 24712 22435 24714
rect 19333 24656 19338 24712
rect 19394 24656 22374 24712
rect 22430 24656 22435 24712
rect 19333 24654 22435 24656
rect 19333 24651 19399 24654
rect 22369 24651 22435 24654
rect 22645 24714 22711 24717
rect 27294 24714 27354 24790
rect 27520 24760 28000 24790
rect 22645 24712 27354 24714
rect 22645 24656 22650 24712
rect 22706 24656 27354 24712
rect 22645 24654 27354 24656
rect 22645 24651 22711 24654
rect 3325 24578 3391 24581
rect 10041 24578 10107 24581
rect 3325 24576 10107 24578
rect 3325 24520 3330 24576
rect 3386 24520 10046 24576
rect 10102 24520 10107 24576
rect 3325 24518 10107 24520
rect 3325 24515 3391 24518
rect 10041 24515 10107 24518
rect 11513 24578 11579 24581
rect 18873 24578 18939 24581
rect 11513 24576 18939 24578
rect 11513 24520 11518 24576
rect 11574 24520 18878 24576
rect 18934 24520 18939 24576
rect 11513 24518 18939 24520
rect 11513 24515 11579 24518
rect 18873 24515 18939 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 5349 24442 5415 24445
rect 8109 24442 8175 24445
rect 5349 24440 8175 24442
rect 5349 24384 5354 24440
rect 5410 24384 8114 24440
rect 8170 24384 8175 24440
rect 5349 24382 8175 24384
rect 5349 24379 5415 24382
rect 8109 24379 8175 24382
rect 13905 24442 13971 24445
rect 18229 24442 18295 24445
rect 13905 24440 18295 24442
rect 13905 24384 13910 24440
rect 13966 24384 18234 24440
rect 18290 24384 18295 24440
rect 13905 24382 18295 24384
rect 13905 24379 13971 24382
rect 18229 24379 18295 24382
rect 0 24306 480 24336
rect 2865 24306 2931 24309
rect 0 24304 2931 24306
rect 0 24248 2870 24304
rect 2926 24248 2931 24304
rect 0 24246 2931 24248
rect 0 24216 480 24246
rect 2865 24243 2931 24246
rect 8293 24306 8359 24309
rect 11421 24306 11487 24309
rect 8293 24304 11487 24306
rect 8293 24248 8298 24304
rect 8354 24248 11426 24304
rect 11482 24248 11487 24304
rect 8293 24246 11487 24248
rect 8293 24243 8359 24246
rect 11421 24243 11487 24246
rect 15837 24306 15903 24309
rect 19517 24306 19583 24309
rect 15837 24304 19583 24306
rect 15837 24248 15842 24304
rect 15898 24248 19522 24304
rect 19578 24248 19583 24304
rect 15837 24246 19583 24248
rect 15837 24243 15903 24246
rect 19517 24243 19583 24246
rect 20713 24306 20779 24309
rect 21909 24306 21975 24309
rect 27520 24306 28000 24336
rect 20713 24304 28000 24306
rect 20713 24248 20718 24304
rect 20774 24248 21914 24304
rect 21970 24248 28000 24304
rect 20713 24246 28000 24248
rect 20713 24243 20779 24246
rect 21909 24243 21975 24246
rect 27520 24216 28000 24246
rect 7189 24170 7255 24173
rect 10869 24170 10935 24173
rect 7189 24168 10935 24170
rect 7189 24112 7194 24168
rect 7250 24112 10874 24168
rect 10930 24112 10935 24168
rect 7189 24110 10935 24112
rect 7189 24107 7255 24110
rect 10869 24107 10935 24110
rect 13721 24170 13787 24173
rect 16573 24170 16639 24173
rect 13721 24168 16639 24170
rect 13721 24112 13726 24168
rect 13782 24112 16578 24168
rect 16634 24112 16639 24168
rect 13721 24110 16639 24112
rect 13721 24107 13787 24110
rect 16573 24107 16639 24110
rect 16757 24170 16823 24173
rect 23013 24170 23079 24173
rect 16757 24168 23079 24170
rect 16757 24112 16762 24168
rect 16818 24112 23018 24168
rect 23074 24112 23079 24168
rect 16757 24110 23079 24112
rect 16757 24107 16823 24110
rect 23013 24107 23079 24110
rect 6085 24034 6151 24037
rect 11513 24034 11579 24037
rect 6085 24032 11579 24034
rect 6085 23976 6090 24032
rect 6146 23976 11518 24032
rect 11574 23976 11579 24032
rect 6085 23974 11579 23976
rect 6085 23971 6151 23974
rect 11513 23971 11579 23974
rect 11789 24034 11855 24037
rect 13997 24034 14063 24037
rect 11789 24032 14063 24034
rect 11789 23976 11794 24032
rect 11850 23976 14002 24032
rect 14058 23976 14063 24032
rect 11789 23974 14063 23976
rect 11789 23971 11855 23974
rect 13997 23971 14063 23974
rect 15561 24034 15627 24037
rect 17033 24034 17099 24037
rect 15561 24032 17099 24034
rect 15561 23976 15566 24032
rect 15622 23976 17038 24032
rect 17094 23976 17099 24032
rect 15561 23974 17099 23976
rect 15561 23971 15627 23974
rect 17033 23971 17099 23974
rect 25405 24034 25471 24037
rect 27613 24034 27679 24037
rect 25405 24032 27679 24034
rect 25405 23976 25410 24032
rect 25466 23976 27618 24032
rect 27674 23976 27679 24032
rect 25405 23974 27679 23976
rect 25405 23971 25471 23974
rect 27613 23971 27679 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 12249 23898 12315 23901
rect 14549 23898 14615 23901
rect 12249 23896 14615 23898
rect 12249 23840 12254 23896
rect 12310 23840 14554 23896
rect 14610 23840 14615 23896
rect 12249 23838 14615 23840
rect 12249 23835 12315 23838
rect 14549 23835 14615 23838
rect 15745 23898 15811 23901
rect 22921 23898 22987 23901
rect 15745 23896 22987 23898
rect 15745 23840 15750 23896
rect 15806 23840 22926 23896
rect 22982 23840 22987 23896
rect 15745 23838 22987 23840
rect 15745 23835 15811 23838
rect 22921 23835 22987 23838
rect 0 23762 480 23792
rect 3325 23762 3391 23765
rect 0 23760 3391 23762
rect 0 23704 3330 23760
rect 3386 23704 3391 23760
rect 0 23702 3391 23704
rect 0 23672 480 23702
rect 3325 23699 3391 23702
rect 4521 23762 4587 23765
rect 10133 23762 10199 23765
rect 12065 23762 12131 23765
rect 4521 23760 12131 23762
rect 4521 23704 4526 23760
rect 4582 23704 10138 23760
rect 10194 23704 12070 23760
rect 12126 23704 12131 23760
rect 4521 23702 12131 23704
rect 4521 23699 4587 23702
rect 10133 23699 10199 23702
rect 12065 23699 12131 23702
rect 23749 23762 23815 23765
rect 24945 23762 25011 23765
rect 23749 23760 25011 23762
rect 23749 23704 23754 23760
rect 23810 23704 24950 23760
rect 25006 23704 25011 23760
rect 23749 23702 25011 23704
rect 23749 23699 23815 23702
rect 24945 23699 25011 23702
rect 25773 23762 25839 23765
rect 27520 23762 28000 23792
rect 25773 23760 28000 23762
rect 25773 23704 25778 23760
rect 25834 23704 28000 23760
rect 25773 23702 28000 23704
rect 25773 23699 25839 23702
rect 27520 23672 28000 23702
rect 5349 23626 5415 23629
rect 14549 23626 14615 23629
rect 20713 23626 20779 23629
rect 2776 23624 5415 23626
rect 2776 23568 5354 23624
rect 5410 23568 5415 23624
rect 2776 23566 5415 23568
rect 2776 23493 2836 23566
rect 5349 23563 5415 23566
rect 9998 23566 10748 23626
rect 2773 23488 2839 23493
rect 2773 23432 2778 23488
rect 2834 23432 2839 23488
rect 2773 23427 2839 23432
rect 4153 23490 4219 23493
rect 7741 23490 7807 23493
rect 8661 23490 8727 23493
rect 4153 23488 8727 23490
rect 4153 23432 4158 23488
rect 4214 23432 7746 23488
rect 7802 23432 8666 23488
rect 8722 23432 8727 23488
rect 4153 23430 8727 23432
rect 4153 23427 4219 23430
rect 7741 23427 7807 23430
rect 8661 23427 8727 23430
rect 1577 23354 1643 23357
rect 6453 23354 6519 23357
rect 1577 23352 6519 23354
rect 1577 23296 1582 23352
rect 1638 23296 6458 23352
rect 6514 23296 6519 23352
rect 1577 23294 6519 23296
rect 1577 23291 1643 23294
rect 6453 23291 6519 23294
rect 8109 23354 8175 23357
rect 9998 23354 10058 23566
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 8109 23352 10058 23354
rect 8109 23296 8114 23352
rect 8170 23296 10058 23352
rect 8109 23294 10058 23296
rect 10688 23354 10748 23566
rect 14549 23624 20779 23626
rect 14549 23568 14554 23624
rect 14610 23568 20718 23624
rect 20774 23568 20779 23624
rect 14549 23566 20779 23568
rect 14549 23563 14615 23566
rect 20713 23563 20779 23566
rect 10961 23490 11027 23493
rect 13445 23490 13511 23493
rect 19425 23490 19491 23493
rect 10961 23488 19491 23490
rect 10961 23432 10966 23488
rect 11022 23432 13450 23488
rect 13506 23432 19430 23488
rect 19486 23432 19491 23488
rect 10961 23430 19491 23432
rect 10961 23427 11027 23430
rect 13445 23427 13511 23430
rect 19425 23427 19491 23430
rect 24025 23490 24091 23493
rect 25221 23490 25287 23493
rect 24025 23488 25287 23490
rect 24025 23432 24030 23488
rect 24086 23432 25226 23488
rect 25282 23432 25287 23488
rect 24025 23430 25287 23432
rect 24025 23427 24091 23430
rect 25221 23427 25287 23430
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 12985 23354 13051 23357
rect 10688 23352 13051 23354
rect 10688 23296 12990 23352
rect 13046 23296 13051 23352
rect 10688 23294 13051 23296
rect 8109 23291 8175 23294
rect 12985 23291 13051 23294
rect 14825 23354 14891 23357
rect 18413 23354 18479 23357
rect 14825 23352 18479 23354
rect 14825 23296 14830 23352
rect 14886 23296 18418 23352
rect 18474 23296 18479 23352
rect 14825 23294 18479 23296
rect 14825 23291 14891 23294
rect 18413 23291 18479 23294
rect 0 23218 480 23248
rect 8293 23218 8359 23221
rect 0 23216 8359 23218
rect 0 23160 8298 23216
rect 8354 23160 8359 23216
rect 0 23158 8359 23160
rect 0 23128 480 23158
rect 8293 23155 8359 23158
rect 8661 23218 8727 23221
rect 11145 23218 11211 23221
rect 8661 23216 11211 23218
rect 8661 23160 8666 23216
rect 8722 23160 11150 23216
rect 11206 23160 11211 23216
rect 8661 23158 11211 23160
rect 8661 23155 8727 23158
rect 11145 23155 11211 23158
rect 11421 23218 11487 23221
rect 17309 23218 17375 23221
rect 27520 23218 28000 23248
rect 11421 23216 17375 23218
rect 11421 23160 11426 23216
rect 11482 23160 17314 23216
rect 17370 23160 17375 23216
rect 11421 23158 17375 23160
rect 11421 23155 11487 23158
rect 17309 23155 17375 23158
rect 23798 23158 28000 23218
rect 23798 23085 23858 23158
rect 27520 23128 28000 23158
rect 1945 23082 2011 23085
rect 14089 23082 14155 23085
rect 14917 23082 14983 23085
rect 1945 23080 14983 23082
rect 1945 23024 1950 23080
rect 2006 23024 14094 23080
rect 14150 23024 14922 23080
rect 14978 23024 14983 23080
rect 1945 23022 14983 23024
rect 1945 23019 2011 23022
rect 14089 23019 14155 23022
rect 14917 23019 14983 23022
rect 15101 23082 15167 23085
rect 16757 23082 16823 23085
rect 15101 23080 16823 23082
rect 15101 23024 15106 23080
rect 15162 23024 16762 23080
rect 16818 23024 16823 23080
rect 15101 23022 16823 23024
rect 15101 23019 15167 23022
rect 16757 23019 16823 23022
rect 17493 23082 17559 23085
rect 23013 23082 23079 23085
rect 17493 23080 23079 23082
rect 17493 23024 17498 23080
rect 17554 23024 23018 23080
rect 23074 23024 23079 23080
rect 17493 23022 23079 23024
rect 17493 23019 17559 23022
rect 23013 23019 23079 23022
rect 23749 23080 23858 23085
rect 23749 23024 23754 23080
rect 23810 23024 23858 23080
rect 23749 23022 23858 23024
rect 23749 23019 23815 23022
rect 7465 22946 7531 22949
rect 11697 22946 11763 22949
rect 7465 22944 11763 22946
rect 7465 22888 7470 22944
rect 7526 22888 11702 22944
rect 11758 22888 11763 22944
rect 7465 22886 11763 22888
rect 7465 22883 7531 22886
rect 11697 22883 11763 22886
rect 12433 22946 12499 22949
rect 14549 22946 14615 22949
rect 12433 22944 14615 22946
rect 12433 22888 12438 22944
rect 12494 22888 14554 22944
rect 14610 22888 14615 22944
rect 12433 22886 14615 22888
rect 12433 22883 12499 22886
rect 14549 22883 14615 22886
rect 16389 22946 16455 22949
rect 20253 22946 20319 22949
rect 16389 22944 20319 22946
rect 16389 22888 16394 22944
rect 16450 22888 20258 22944
rect 20314 22888 20319 22944
rect 16389 22886 20319 22888
rect 16389 22883 16455 22886
rect 20253 22883 20319 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2497 22810 2563 22813
rect 5257 22810 5323 22813
rect 2497 22808 5323 22810
rect 2497 22752 2502 22808
rect 2558 22752 5262 22808
rect 5318 22752 5323 22808
rect 2497 22750 5323 22752
rect 2497 22747 2563 22750
rect 5257 22747 5323 22750
rect 7189 22810 7255 22813
rect 12893 22810 12959 22813
rect 7189 22808 12959 22810
rect 7189 22752 7194 22808
rect 7250 22752 12898 22808
rect 12954 22752 12959 22808
rect 7189 22750 12959 22752
rect 7189 22747 7255 22750
rect 12893 22747 12959 22750
rect 16481 22810 16547 22813
rect 16481 22808 23674 22810
rect 16481 22752 16486 22808
rect 16542 22752 23674 22808
rect 16481 22750 23674 22752
rect 16481 22747 16547 22750
rect 4981 22674 5047 22677
rect 6913 22674 6979 22677
rect 4981 22672 6979 22674
rect 4981 22616 4986 22672
rect 5042 22616 6918 22672
rect 6974 22616 6979 22672
rect 4981 22614 6979 22616
rect 4981 22611 5047 22614
rect 6913 22611 6979 22614
rect 11329 22674 11395 22677
rect 13537 22674 13603 22677
rect 15193 22674 15259 22677
rect 11329 22672 15259 22674
rect 11329 22616 11334 22672
rect 11390 22616 13542 22672
rect 13598 22616 15198 22672
rect 15254 22616 15259 22672
rect 11329 22614 15259 22616
rect 23614 22674 23674 22750
rect 25037 22674 25103 22677
rect 23614 22672 25103 22674
rect 23614 22616 25042 22672
rect 25098 22616 25103 22672
rect 23614 22614 25103 22616
rect 11329 22611 11395 22614
rect 13537 22611 13603 22614
rect 15193 22611 15259 22614
rect 25037 22611 25103 22614
rect 0 22538 480 22568
rect 7005 22538 7071 22541
rect 11421 22538 11487 22541
rect 0 22536 7071 22538
rect 0 22480 7010 22536
rect 7066 22480 7071 22536
rect 0 22478 7071 22480
rect 0 22448 480 22478
rect 7005 22475 7071 22478
rect 7606 22536 11487 22538
rect 7606 22480 11426 22536
rect 11482 22480 11487 22536
rect 7606 22478 11487 22480
rect 4061 22402 4127 22405
rect 6085 22402 6151 22405
rect 4061 22400 6151 22402
rect 4061 22344 4066 22400
rect 4122 22344 6090 22400
rect 6146 22344 6151 22400
rect 4061 22342 6151 22344
rect 4061 22339 4127 22342
rect 6085 22339 6151 22342
rect 2681 22266 2747 22269
rect 7606 22266 7666 22478
rect 11421 22475 11487 22478
rect 12065 22538 12131 22541
rect 14273 22538 14339 22541
rect 18781 22538 18847 22541
rect 12065 22536 12634 22538
rect 12065 22480 12070 22536
rect 12126 22480 12634 22536
rect 12065 22478 12634 22480
rect 12065 22475 12131 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 12433 22266 12499 22269
rect 2681 22264 7666 22266
rect 2681 22208 2686 22264
rect 2742 22208 7666 22264
rect 2681 22206 7666 22208
rect 11056 22264 12499 22266
rect 11056 22208 12438 22264
rect 12494 22208 12499 22264
rect 11056 22206 12499 22208
rect 12574 22266 12634 22478
rect 14273 22536 18847 22538
rect 14273 22480 14278 22536
rect 14334 22480 18786 22536
rect 18842 22480 18847 22536
rect 14273 22478 18847 22480
rect 14273 22475 14339 22478
rect 18781 22475 18847 22478
rect 19977 22538 20043 22541
rect 25221 22538 25287 22541
rect 19977 22536 25287 22538
rect 19977 22480 19982 22536
rect 20038 22480 25226 22536
rect 25282 22480 25287 22536
rect 19977 22478 25287 22480
rect 19977 22475 20043 22478
rect 25221 22475 25287 22478
rect 25497 22538 25563 22541
rect 27520 22538 28000 22568
rect 25497 22536 28000 22538
rect 25497 22480 25502 22536
rect 25558 22480 28000 22536
rect 25497 22478 28000 22480
rect 25497 22475 25563 22478
rect 27520 22448 28000 22478
rect 12709 22402 12775 22405
rect 18045 22402 18111 22405
rect 12709 22400 18111 22402
rect 12709 22344 12714 22400
rect 12770 22344 18050 22400
rect 18106 22344 18111 22400
rect 12709 22342 18111 22344
rect 12709 22339 12775 22342
rect 18045 22339 18111 22342
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 15561 22266 15627 22269
rect 12574 22264 15627 22266
rect 12574 22208 15566 22264
rect 15622 22208 15627 22264
rect 12574 22206 15627 22208
rect 2681 22203 2747 22206
rect 10593 22130 10659 22133
rect 11056 22130 11116 22206
rect 12433 22203 12499 22206
rect 15561 22203 15627 22206
rect 10593 22128 11116 22130
rect 10593 22072 10598 22128
rect 10654 22072 11116 22128
rect 10593 22070 11116 22072
rect 18873 22130 18939 22133
rect 21449 22130 21515 22133
rect 18873 22128 21515 22130
rect 18873 22072 18878 22128
rect 18934 22072 21454 22128
rect 21510 22072 21515 22128
rect 18873 22070 21515 22072
rect 10593 22067 10659 22070
rect 18873 22067 18939 22070
rect 21449 22067 21515 22070
rect 0 21994 480 22024
rect 3049 21994 3115 21997
rect 0 21992 3115 21994
rect 0 21936 3054 21992
rect 3110 21936 3115 21992
rect 0 21934 3115 21936
rect 0 21904 480 21934
rect 3049 21931 3115 21934
rect 3601 21994 3667 21997
rect 4337 21994 4403 21997
rect 3601 21992 4403 21994
rect 3601 21936 3606 21992
rect 3662 21936 4342 21992
rect 4398 21936 4403 21992
rect 3601 21934 4403 21936
rect 3601 21931 3667 21934
rect 4337 21931 4403 21934
rect 4521 21994 4587 21997
rect 8293 21994 8359 21997
rect 4521 21992 8359 21994
rect 4521 21936 4526 21992
rect 4582 21936 8298 21992
rect 8354 21936 8359 21992
rect 4521 21934 8359 21936
rect 4521 21931 4587 21934
rect 8293 21931 8359 21934
rect 9581 21994 9647 21997
rect 9765 21994 9831 21997
rect 9581 21992 9831 21994
rect 9581 21936 9586 21992
rect 9642 21936 9770 21992
rect 9826 21936 9831 21992
rect 9581 21934 9831 21936
rect 9581 21931 9647 21934
rect 9765 21931 9831 21934
rect 17585 21994 17651 21997
rect 19701 21994 19767 21997
rect 17585 21992 19767 21994
rect 17585 21936 17590 21992
rect 17646 21936 19706 21992
rect 19762 21936 19767 21992
rect 17585 21934 19767 21936
rect 17585 21931 17651 21934
rect 19701 21931 19767 21934
rect 21541 21994 21607 21997
rect 23657 21994 23723 21997
rect 25129 21994 25195 21997
rect 21541 21992 23723 21994
rect 21541 21936 21546 21992
rect 21602 21936 23662 21992
rect 23718 21936 23723 21992
rect 21541 21934 23723 21936
rect 21541 21931 21607 21934
rect 23657 21931 23723 21934
rect 23798 21992 25195 21994
rect 23798 21936 25134 21992
rect 25190 21936 25195 21992
rect 23798 21934 25195 21936
rect 2405 21858 2471 21861
rect 4429 21858 4495 21861
rect 2405 21856 4495 21858
rect 2405 21800 2410 21856
rect 2466 21800 4434 21856
rect 4490 21800 4495 21856
rect 2405 21798 4495 21800
rect 2405 21795 2471 21798
rect 4429 21795 4495 21798
rect 19241 21858 19307 21861
rect 23798 21858 23858 21934
rect 25129 21931 25195 21934
rect 25405 21994 25471 21997
rect 27520 21994 28000 22024
rect 25405 21992 28000 21994
rect 25405 21936 25410 21992
rect 25466 21936 28000 21992
rect 25405 21934 28000 21936
rect 25405 21931 25471 21934
rect 27520 21904 28000 21934
rect 19241 21856 23858 21858
rect 19241 21800 19246 21856
rect 19302 21800 23858 21856
rect 19241 21798 23858 21800
rect 19241 21795 19307 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 6085 21722 6151 21725
rect 11053 21722 11119 21725
rect 6085 21720 11119 21722
rect 6085 21664 6090 21720
rect 6146 21664 11058 21720
rect 11114 21664 11119 21720
rect 6085 21662 11119 21664
rect 6085 21659 6151 21662
rect 11053 21659 11119 21662
rect 2037 21586 2103 21589
rect 3877 21586 3943 21589
rect 4153 21586 4219 21589
rect 2037 21584 4219 21586
rect 2037 21528 2042 21584
rect 2098 21528 3882 21584
rect 3938 21528 4158 21584
rect 4214 21528 4219 21584
rect 2037 21526 4219 21528
rect 2037 21523 2103 21526
rect 3877 21523 3943 21526
rect 4153 21523 4219 21526
rect 4429 21586 4495 21589
rect 7925 21586 7991 21589
rect 4429 21584 7991 21586
rect 4429 21528 4434 21584
rect 4490 21528 7930 21584
rect 7986 21528 7991 21584
rect 4429 21526 7991 21528
rect 4429 21523 4495 21526
rect 7925 21523 7991 21526
rect 10501 21586 10567 21589
rect 13353 21586 13419 21589
rect 15285 21586 15351 21589
rect 20897 21586 20963 21589
rect 10501 21584 20963 21586
rect 10501 21528 10506 21584
rect 10562 21528 13358 21584
rect 13414 21528 15290 21584
rect 15346 21528 20902 21584
rect 20958 21528 20963 21584
rect 10501 21526 20963 21528
rect 10501 21523 10567 21526
rect 13353 21523 13419 21526
rect 15285 21523 15351 21526
rect 20897 21523 20963 21526
rect 0 21450 480 21480
rect 2773 21450 2839 21453
rect 0 21448 2839 21450
rect 0 21392 2778 21448
rect 2834 21392 2839 21448
rect 0 21390 2839 21392
rect 0 21360 480 21390
rect 2773 21387 2839 21390
rect 3693 21450 3759 21453
rect 5993 21450 6059 21453
rect 3693 21448 6059 21450
rect 3693 21392 3698 21448
rect 3754 21392 5998 21448
rect 6054 21392 6059 21448
rect 3693 21390 6059 21392
rect 3693 21387 3759 21390
rect 5993 21387 6059 21390
rect 6729 21450 6795 21453
rect 7281 21450 7347 21453
rect 12617 21450 12683 21453
rect 6729 21448 12683 21450
rect 6729 21392 6734 21448
rect 6790 21392 7286 21448
rect 7342 21392 12622 21448
rect 12678 21392 12683 21448
rect 6729 21390 12683 21392
rect 6729 21387 6795 21390
rect 7281 21387 7347 21390
rect 12617 21387 12683 21390
rect 15837 21450 15903 21453
rect 25313 21450 25379 21453
rect 15837 21448 25379 21450
rect 15837 21392 15842 21448
rect 15898 21392 25318 21448
rect 25374 21392 25379 21448
rect 15837 21390 25379 21392
rect 15837 21387 15903 21390
rect 25313 21387 25379 21390
rect 25497 21450 25563 21453
rect 27520 21450 28000 21480
rect 25497 21448 28000 21450
rect 25497 21392 25502 21448
rect 25558 21392 28000 21448
rect 25497 21390 28000 21392
rect 25497 21387 25563 21390
rect 27520 21360 28000 21390
rect 3233 21314 3299 21317
rect 10041 21314 10107 21317
rect 3233 21312 10107 21314
rect 3233 21256 3238 21312
rect 3294 21256 10046 21312
rect 10102 21256 10107 21312
rect 3233 21254 10107 21256
rect 3233 21251 3299 21254
rect 10041 21251 10107 21254
rect 11053 21314 11119 21317
rect 11605 21314 11671 21317
rect 16389 21314 16455 21317
rect 11053 21312 16455 21314
rect 11053 21256 11058 21312
rect 11114 21256 11610 21312
rect 11666 21256 16394 21312
rect 16450 21256 16455 21312
rect 11053 21254 16455 21256
rect 11053 21251 11119 21254
rect 11605 21251 11671 21254
rect 16389 21251 16455 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 4061 21042 4127 21045
rect 5993 21042 6059 21045
rect 4061 21040 6059 21042
rect 4061 20984 4066 21040
rect 4122 20984 5998 21040
rect 6054 20984 6059 21040
rect 4061 20982 6059 20984
rect 4061 20979 4127 20982
rect 5993 20979 6059 20982
rect 10961 21042 11027 21045
rect 13813 21042 13879 21045
rect 10961 21040 13879 21042
rect 10961 20984 10966 21040
rect 11022 20984 13818 21040
rect 13874 20984 13879 21040
rect 10961 20982 13879 20984
rect 10961 20979 11027 20982
rect 13813 20979 13879 20982
rect 0 20906 480 20936
rect 8661 20906 8727 20909
rect 0 20904 8727 20906
rect 0 20848 8666 20904
rect 8722 20848 8727 20904
rect 0 20846 8727 20848
rect 0 20816 480 20846
rect 8661 20843 8727 20846
rect 8845 20906 8911 20909
rect 13169 20906 13235 20909
rect 8845 20904 13235 20906
rect 8845 20848 8850 20904
rect 8906 20848 13174 20904
rect 13230 20848 13235 20904
rect 8845 20846 13235 20848
rect 8845 20843 8911 20846
rect 13169 20843 13235 20846
rect 13629 20906 13695 20909
rect 18137 20906 18203 20909
rect 13629 20904 18203 20906
rect 13629 20848 13634 20904
rect 13690 20848 18142 20904
rect 18198 20848 18203 20904
rect 13629 20846 18203 20848
rect 13629 20843 13695 20846
rect 18137 20843 18203 20846
rect 22921 20906 22987 20909
rect 27520 20906 28000 20936
rect 22921 20904 28000 20906
rect 22921 20848 22926 20904
rect 22982 20848 28000 20904
rect 22921 20846 28000 20848
rect 22921 20843 22987 20846
rect 27520 20816 28000 20846
rect 6821 20770 6887 20773
rect 11513 20770 11579 20773
rect 6821 20768 11579 20770
rect 6821 20712 6826 20768
rect 6882 20712 11518 20768
rect 11574 20712 11579 20768
rect 6821 20710 11579 20712
rect 6821 20707 6887 20710
rect 11513 20707 11579 20710
rect 13445 20770 13511 20773
rect 14089 20770 14155 20773
rect 13445 20768 14155 20770
rect 13445 20712 13450 20768
rect 13506 20712 14094 20768
rect 14150 20712 14155 20768
rect 13445 20710 14155 20712
rect 13445 20707 13511 20710
rect 14089 20707 14155 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 2773 20634 2839 20637
rect 4429 20634 4495 20637
rect 2773 20632 4495 20634
rect 2773 20576 2778 20632
rect 2834 20576 4434 20632
rect 4490 20576 4495 20632
rect 2773 20574 4495 20576
rect 2773 20571 2839 20574
rect 4429 20571 4495 20574
rect 10869 20634 10935 20637
rect 14641 20634 14707 20637
rect 10869 20632 14707 20634
rect 10869 20576 10874 20632
rect 10930 20576 14646 20632
rect 14702 20576 14707 20632
rect 10869 20574 14707 20576
rect 10869 20571 10935 20574
rect 14641 20571 14707 20574
rect 17401 20634 17467 20637
rect 23749 20634 23815 20637
rect 17401 20632 23815 20634
rect 17401 20576 17406 20632
rect 17462 20576 23754 20632
rect 23810 20576 23815 20632
rect 17401 20574 23815 20576
rect 17401 20571 17467 20574
rect 23749 20571 23815 20574
rect 2405 20498 2471 20501
rect 3141 20498 3207 20501
rect 7005 20498 7071 20501
rect 2405 20496 2928 20498
rect 2405 20440 2410 20496
rect 2466 20440 2928 20496
rect 2405 20438 2928 20440
rect 2405 20435 2471 20438
rect 0 20362 480 20392
rect 1117 20362 1183 20365
rect 0 20360 1183 20362
rect 0 20304 1122 20360
rect 1178 20304 1183 20360
rect 0 20302 1183 20304
rect 2868 20362 2928 20438
rect 3141 20496 7071 20498
rect 3141 20440 3146 20496
rect 3202 20440 7010 20496
rect 7066 20440 7071 20496
rect 3141 20438 7071 20440
rect 3141 20435 3207 20438
rect 7005 20435 7071 20438
rect 11973 20498 12039 20501
rect 17493 20498 17559 20501
rect 11973 20496 17559 20498
rect 11973 20440 11978 20496
rect 12034 20440 17498 20496
rect 17554 20440 17559 20496
rect 11973 20438 17559 20440
rect 11973 20435 12039 20438
rect 17493 20435 17559 20438
rect 19517 20498 19583 20501
rect 24853 20498 24919 20501
rect 19517 20496 24919 20498
rect 19517 20440 19522 20496
rect 19578 20440 24858 20496
rect 24914 20440 24919 20496
rect 19517 20438 24919 20440
rect 19517 20435 19583 20438
rect 24853 20435 24919 20438
rect 3325 20362 3391 20365
rect 10869 20362 10935 20365
rect 19374 20362 19380 20364
rect 2868 20360 10935 20362
rect 2868 20304 3330 20360
rect 3386 20304 10874 20360
rect 10930 20304 10935 20360
rect 2868 20302 10935 20304
rect 0 20272 480 20302
rect 1117 20299 1183 20302
rect 3325 20299 3391 20302
rect 10869 20299 10935 20302
rect 11056 20302 19380 20362
rect 10869 20226 10935 20229
rect 11056 20226 11116 20302
rect 19374 20300 19380 20302
rect 19444 20300 19450 20364
rect 21081 20362 21147 20365
rect 27520 20362 28000 20392
rect 21081 20360 28000 20362
rect 21081 20304 21086 20360
rect 21142 20304 28000 20360
rect 21081 20302 28000 20304
rect 21081 20299 21147 20302
rect 27520 20272 28000 20302
rect 10869 20224 11116 20226
rect 10869 20168 10874 20224
rect 10930 20168 11116 20224
rect 10869 20166 11116 20168
rect 10869 20163 10935 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1485 20090 1551 20093
rect 6821 20090 6887 20093
rect 9673 20092 9739 20093
rect 1485 20088 6887 20090
rect 1485 20032 1490 20088
rect 1546 20032 6826 20088
rect 6882 20032 6887 20088
rect 1485 20030 6887 20032
rect 1485 20027 1551 20030
rect 6821 20027 6887 20030
rect 9622 20028 9628 20092
rect 9692 20090 9739 20092
rect 14825 20090 14891 20093
rect 9692 20088 9784 20090
rect 9734 20032 9784 20088
rect 9692 20030 9784 20032
rect 14825 20088 15946 20090
rect 14825 20032 14830 20088
rect 14886 20032 15946 20088
rect 14825 20030 15946 20032
rect 9692 20028 9739 20030
rect 9673 20027 9739 20028
rect 14825 20027 14891 20030
rect 1669 19954 1735 19957
rect 5993 19954 6059 19957
rect 1669 19952 6059 19954
rect 1669 19896 1674 19952
rect 1730 19896 5998 19952
rect 6054 19896 6059 19952
rect 1669 19894 6059 19896
rect 15886 19954 15946 20030
rect 22921 19954 22987 19957
rect 15886 19952 22987 19954
rect 15886 19896 22926 19952
rect 22982 19896 22987 19952
rect 15886 19894 22987 19896
rect 1669 19891 1735 19894
rect 5993 19891 6059 19894
rect 22921 19891 22987 19894
rect 5165 19818 5231 19821
rect 11605 19818 11671 19821
rect 5165 19816 11671 19818
rect 5165 19760 5170 19816
rect 5226 19760 11610 19816
rect 11666 19760 11671 19816
rect 5165 19758 11671 19760
rect 5165 19755 5231 19758
rect 11605 19755 11671 19758
rect 19374 19756 19380 19820
rect 19444 19818 19450 19820
rect 20529 19818 20595 19821
rect 19444 19816 20595 19818
rect 19444 19760 20534 19816
rect 20590 19760 20595 19816
rect 19444 19758 20595 19760
rect 19444 19756 19450 19758
rect 20529 19755 20595 19758
rect 0 19682 480 19712
rect 2773 19682 2839 19685
rect 0 19680 2839 19682
rect 0 19624 2778 19680
rect 2834 19624 2839 19680
rect 0 19622 2839 19624
rect 0 19592 480 19622
rect 2773 19619 2839 19622
rect 9990 19620 9996 19684
rect 10060 19682 10066 19684
rect 12065 19682 12131 19685
rect 10060 19680 12131 19682
rect 10060 19624 12070 19680
rect 12126 19624 12131 19680
rect 10060 19622 12131 19624
rect 10060 19620 10066 19622
rect 12065 19619 12131 19622
rect 24669 19682 24735 19685
rect 27520 19682 28000 19712
rect 24669 19680 28000 19682
rect 24669 19624 24674 19680
rect 24730 19624 28000 19680
rect 24669 19622 28000 19624
rect 24669 19619 24735 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19622
rect 24277 19551 24597 19552
rect 2313 19546 2379 19549
rect 5441 19546 5507 19549
rect 2313 19544 5507 19546
rect 2313 19488 2318 19544
rect 2374 19488 5446 19544
rect 5502 19488 5507 19544
rect 2313 19486 5507 19488
rect 2313 19483 2379 19486
rect 5441 19483 5507 19486
rect 5533 19410 5599 19413
rect 8293 19410 8359 19413
rect 5533 19408 8359 19410
rect 5533 19352 5538 19408
rect 5594 19352 8298 19408
rect 8354 19352 8359 19408
rect 5533 19350 8359 19352
rect 5533 19347 5599 19350
rect 8293 19347 8359 19350
rect 8937 19410 9003 19413
rect 11053 19410 11119 19413
rect 8937 19408 11119 19410
rect 8937 19352 8942 19408
rect 8998 19352 11058 19408
rect 11114 19352 11119 19408
rect 8937 19350 11119 19352
rect 8937 19347 9003 19350
rect 11053 19347 11119 19350
rect 24301 19410 24367 19413
rect 25681 19410 25747 19413
rect 24301 19408 25747 19410
rect 24301 19352 24306 19408
rect 24362 19352 25686 19408
rect 25742 19352 25747 19408
rect 24301 19350 25747 19352
rect 24301 19347 24367 19350
rect 25681 19347 25747 19350
rect 2221 19274 2287 19277
rect 7833 19274 7899 19277
rect 2221 19272 7899 19274
rect 2221 19216 2226 19272
rect 2282 19216 7838 19272
rect 7894 19216 7899 19272
rect 2221 19214 7899 19216
rect 2221 19211 2287 19214
rect 7833 19211 7899 19214
rect 9581 19274 9647 19277
rect 13353 19274 13419 19277
rect 9581 19272 13419 19274
rect 9581 19216 9586 19272
rect 9642 19216 13358 19272
rect 13414 19216 13419 19272
rect 9581 19214 13419 19216
rect 9581 19211 9647 19214
rect 13353 19211 13419 19214
rect 17217 19274 17283 19277
rect 25221 19274 25287 19277
rect 17217 19272 25287 19274
rect 17217 19216 17222 19272
rect 17278 19216 25226 19272
rect 25282 19216 25287 19272
rect 17217 19214 25287 19216
rect 17217 19211 17283 19214
rect 25221 19211 25287 19214
rect 0 19138 480 19168
rect 3141 19138 3207 19141
rect 0 19136 3207 19138
rect 0 19080 3146 19136
rect 3202 19080 3207 19136
rect 0 19078 3207 19080
rect 0 19048 480 19078
rect 3141 19075 3207 19078
rect 3601 19138 3667 19141
rect 4521 19138 4587 19141
rect 9673 19138 9739 19141
rect 3601 19136 9739 19138
rect 3601 19080 3606 19136
rect 3662 19080 4526 19136
rect 4582 19080 9678 19136
rect 9734 19080 9739 19136
rect 3601 19078 9739 19080
rect 3601 19075 3667 19078
rect 4521 19075 4587 19078
rect 9673 19075 9739 19078
rect 11145 19138 11211 19141
rect 15009 19138 15075 19141
rect 11145 19136 15075 19138
rect 11145 19080 11150 19136
rect 11206 19080 15014 19136
rect 15070 19080 15075 19136
rect 11145 19078 15075 19080
rect 11145 19075 11211 19078
rect 15009 19075 15075 19078
rect 20069 19138 20135 19141
rect 27520 19138 28000 19168
rect 20069 19136 28000 19138
rect 20069 19080 20074 19136
rect 20130 19080 28000 19136
rect 20069 19078 28000 19080
rect 20069 19075 20135 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 841 19002 907 19005
rect 3601 19002 3667 19005
rect 841 19000 3667 19002
rect 841 18944 846 19000
rect 902 18944 3606 19000
rect 3662 18944 3667 19000
rect 841 18942 3667 18944
rect 841 18939 907 18942
rect 3601 18939 3667 18942
rect 7833 19002 7899 19005
rect 10133 19002 10199 19005
rect 7833 19000 10199 19002
rect 7833 18944 7838 19000
rect 7894 18944 10138 19000
rect 10194 18944 10199 19000
rect 7833 18942 10199 18944
rect 7833 18939 7899 18942
rect 10133 18939 10199 18942
rect 1945 18866 2011 18869
rect 8753 18866 8819 18869
rect 1945 18864 8819 18866
rect 1945 18808 1950 18864
rect 2006 18808 8758 18864
rect 8814 18808 8819 18864
rect 1945 18806 8819 18808
rect 1945 18803 2011 18806
rect 8753 18803 8819 18806
rect 13721 18866 13787 18869
rect 21357 18866 21423 18869
rect 13721 18864 21423 18866
rect 13721 18808 13726 18864
rect 13782 18808 21362 18864
rect 21418 18808 21423 18864
rect 13721 18806 21423 18808
rect 13721 18803 13787 18806
rect 21357 18803 21423 18806
rect 21909 18866 21975 18869
rect 23381 18866 23447 18869
rect 21909 18864 23447 18866
rect 21909 18808 21914 18864
rect 21970 18808 23386 18864
rect 23442 18808 23447 18864
rect 21909 18806 23447 18808
rect 21909 18803 21975 18806
rect 23381 18803 23447 18806
rect 3509 18730 3575 18733
rect 11237 18730 11303 18733
rect 3509 18728 11303 18730
rect 3509 18672 3514 18728
rect 3570 18672 11242 18728
rect 11298 18672 11303 18728
rect 3509 18670 11303 18672
rect 3509 18667 3575 18670
rect 11237 18667 11303 18670
rect 12617 18730 12683 18733
rect 17401 18730 17467 18733
rect 12617 18728 17467 18730
rect 12617 18672 12622 18728
rect 12678 18672 17406 18728
rect 17462 18672 17467 18728
rect 12617 18670 17467 18672
rect 12617 18667 12683 18670
rect 17401 18667 17467 18670
rect 23657 18730 23723 18733
rect 26233 18730 26299 18733
rect 23657 18728 26299 18730
rect 23657 18672 23662 18728
rect 23718 18672 26238 18728
rect 26294 18672 26299 18728
rect 23657 18670 26299 18672
rect 23657 18667 23723 18670
rect 26233 18667 26299 18670
rect 0 18594 480 18624
rect 3877 18594 3943 18597
rect 0 18592 3943 18594
rect 0 18536 3882 18592
rect 3938 18536 3943 18592
rect 0 18534 3943 18536
rect 0 18504 480 18534
rect 3877 18531 3943 18534
rect 9397 18594 9463 18597
rect 9857 18594 9923 18597
rect 13813 18594 13879 18597
rect 9397 18592 13879 18594
rect 9397 18536 9402 18592
rect 9458 18536 9862 18592
rect 9918 18536 13818 18592
rect 13874 18536 13879 18592
rect 9397 18534 13879 18536
rect 9397 18531 9463 18534
rect 9857 18531 9923 18534
rect 13813 18531 13879 18534
rect 24761 18594 24827 18597
rect 27520 18594 28000 18624
rect 24761 18592 28000 18594
rect 24761 18536 24766 18592
rect 24822 18536 28000 18592
rect 24761 18534 28000 18536
rect 24761 18531 24827 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 27520 18504 28000 18534
rect 24277 18463 24597 18464
rect 7465 18458 7531 18461
rect 12617 18458 12683 18461
rect 7465 18456 12683 18458
rect 7465 18400 7470 18456
rect 7526 18400 12622 18456
rect 12678 18400 12683 18456
rect 7465 18398 12683 18400
rect 7465 18395 7531 18398
rect 12617 18395 12683 18398
rect 12525 18322 12591 18325
rect 22369 18322 22435 18325
rect 12525 18320 22435 18322
rect 12525 18264 12530 18320
rect 12586 18264 22374 18320
rect 22430 18264 22435 18320
rect 12525 18262 22435 18264
rect 12525 18259 12591 18262
rect 22369 18259 22435 18262
rect 8569 18186 8635 18189
rect 18321 18186 18387 18189
rect 8569 18184 18387 18186
rect 8569 18128 8574 18184
rect 8630 18128 18326 18184
rect 18382 18128 18387 18184
rect 8569 18126 18387 18128
rect 8569 18123 8635 18126
rect 18321 18123 18387 18126
rect 18505 18186 18571 18189
rect 20805 18186 20871 18189
rect 21173 18186 21239 18189
rect 18505 18184 21239 18186
rect 18505 18128 18510 18184
rect 18566 18128 20810 18184
rect 20866 18128 21178 18184
rect 21234 18128 21239 18184
rect 18505 18126 21239 18128
rect 18505 18123 18571 18126
rect 20805 18123 20871 18126
rect 21173 18123 21239 18126
rect 0 18050 480 18080
rect 5809 18050 5875 18053
rect 0 18048 5875 18050
rect 0 17992 5814 18048
rect 5870 17992 5875 18048
rect 0 17990 5875 17992
rect 0 17960 480 17990
rect 5809 17987 5875 17990
rect 6177 18050 6243 18053
rect 8293 18050 8359 18053
rect 6177 18048 8359 18050
rect 6177 17992 6182 18048
rect 6238 17992 8298 18048
rect 8354 17992 8359 18048
rect 6177 17990 8359 17992
rect 6177 17987 6243 17990
rect 8293 17987 8359 17990
rect 23473 18050 23539 18053
rect 27520 18050 28000 18080
rect 23473 18048 28000 18050
rect 23473 17992 23478 18048
rect 23534 17992 28000 18048
rect 23473 17990 28000 17992
rect 23473 17987 23539 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 2221 17914 2287 17917
rect 6729 17914 6795 17917
rect 2221 17912 6795 17914
rect 2221 17856 2226 17912
rect 2282 17856 6734 17912
rect 6790 17856 6795 17912
rect 2221 17854 6795 17856
rect 2221 17851 2287 17854
rect 6729 17851 6795 17854
rect 3877 17778 3943 17781
rect 7005 17778 7071 17781
rect 3877 17776 7071 17778
rect 3877 17720 3882 17776
rect 3938 17720 7010 17776
rect 7066 17720 7071 17776
rect 3877 17718 7071 17720
rect 3877 17715 3943 17718
rect 7005 17715 7071 17718
rect 7373 17778 7439 17781
rect 9949 17778 10015 17781
rect 18321 17778 18387 17781
rect 7373 17776 18387 17778
rect 7373 17720 7378 17776
rect 7434 17720 9954 17776
rect 10010 17720 18326 17776
rect 18382 17720 18387 17776
rect 7373 17718 18387 17720
rect 7373 17715 7439 17718
rect 9949 17715 10015 17718
rect 18321 17715 18387 17718
rect 5349 17642 5415 17645
rect 7649 17642 7715 17645
rect 5349 17640 7715 17642
rect 5349 17584 5354 17640
rect 5410 17584 7654 17640
rect 7710 17584 7715 17640
rect 5349 17582 7715 17584
rect 5349 17579 5415 17582
rect 7649 17579 7715 17582
rect 15101 17642 15167 17645
rect 16757 17642 16823 17645
rect 15101 17640 16823 17642
rect 15101 17584 15106 17640
rect 15162 17584 16762 17640
rect 16818 17584 16823 17640
rect 15101 17582 16823 17584
rect 15101 17579 15167 17582
rect 16757 17579 16823 17582
rect 17217 17642 17283 17645
rect 22277 17642 22343 17645
rect 17217 17640 22343 17642
rect 17217 17584 17222 17640
rect 17278 17584 22282 17640
rect 22338 17584 22343 17640
rect 17217 17582 22343 17584
rect 17217 17579 17283 17582
rect 22277 17579 22343 17582
rect 0 17506 480 17536
rect 1577 17506 1643 17509
rect 0 17504 1643 17506
rect 0 17448 1582 17504
rect 1638 17448 1643 17504
rect 0 17446 1643 17448
rect 0 17416 480 17446
rect 1577 17443 1643 17446
rect 25681 17506 25747 17509
rect 27520 17506 28000 17536
rect 25681 17504 28000 17506
rect 25681 17448 25686 17504
rect 25742 17448 28000 17504
rect 25681 17446 28000 17448
rect 25681 17443 25747 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 2957 17370 3023 17373
rect 4705 17370 4771 17373
rect 2957 17368 4771 17370
rect 2957 17312 2962 17368
rect 3018 17312 4710 17368
rect 4766 17312 4771 17368
rect 2957 17310 4771 17312
rect 2957 17307 3023 17310
rect 4705 17307 4771 17310
rect 7189 17370 7255 17373
rect 7741 17370 7807 17373
rect 13077 17370 13143 17373
rect 7189 17368 13143 17370
rect 7189 17312 7194 17368
rect 7250 17312 7746 17368
rect 7802 17312 13082 17368
rect 13138 17312 13143 17368
rect 7189 17310 13143 17312
rect 7189 17307 7255 17310
rect 7741 17307 7807 17310
rect 13077 17307 13143 17310
rect 14222 17308 14228 17372
rect 14292 17370 14298 17372
rect 14365 17370 14431 17373
rect 14292 17368 14431 17370
rect 14292 17312 14370 17368
rect 14426 17312 14431 17368
rect 14292 17310 14431 17312
rect 14292 17308 14298 17310
rect 14365 17307 14431 17310
rect 1577 17234 1643 17237
rect 9397 17234 9463 17237
rect 1577 17232 9463 17234
rect 1577 17176 1582 17232
rect 1638 17176 9402 17232
rect 9458 17176 9463 17232
rect 1577 17174 9463 17176
rect 1577 17171 1643 17174
rect 9397 17171 9463 17174
rect 11421 17234 11487 17237
rect 18689 17234 18755 17237
rect 11421 17232 18755 17234
rect 11421 17176 11426 17232
rect 11482 17176 18694 17232
rect 18750 17176 18755 17232
rect 11421 17174 18755 17176
rect 11421 17171 11487 17174
rect 18689 17171 18755 17174
rect 3969 17098 4035 17101
rect 7966 17098 7972 17100
rect 3969 17096 7972 17098
rect 3969 17040 3974 17096
rect 4030 17040 7972 17096
rect 3969 17038 7972 17040
rect 3969 17035 4035 17038
rect 7966 17036 7972 17038
rect 8036 17036 8042 17100
rect 9673 17098 9739 17101
rect 19241 17098 19307 17101
rect 9673 17096 19307 17098
rect 9673 17040 9678 17096
rect 9734 17040 19246 17096
rect 19302 17040 19307 17096
rect 9673 17038 19307 17040
rect 9673 17035 9739 17038
rect 19241 17035 19307 17038
rect 2405 16962 2471 16965
rect 4061 16962 4127 16965
rect 2405 16960 4127 16962
rect 2405 16904 2410 16960
rect 2466 16904 4066 16960
rect 4122 16904 4127 16960
rect 2405 16902 4127 16904
rect 2405 16899 2471 16902
rect 4061 16899 4127 16902
rect 4981 16962 5047 16965
rect 8201 16962 8267 16965
rect 9673 16962 9739 16965
rect 4981 16960 9739 16962
rect 4981 16904 4986 16960
rect 5042 16904 8206 16960
rect 8262 16904 9678 16960
rect 9734 16904 9739 16960
rect 4981 16902 9739 16904
rect 4981 16899 5047 16902
rect 8201 16899 8267 16902
rect 9673 16899 9739 16902
rect 13537 16962 13603 16965
rect 15745 16962 15811 16965
rect 13537 16960 15811 16962
rect 13537 16904 13542 16960
rect 13598 16904 15750 16960
rect 15806 16904 15811 16960
rect 13537 16902 15811 16904
rect 13537 16899 13603 16902
rect 15745 16899 15811 16902
rect 23289 16962 23355 16965
rect 25037 16962 25103 16965
rect 23289 16960 25103 16962
rect 23289 16904 23294 16960
rect 23350 16904 25042 16960
rect 25098 16904 25103 16960
rect 23289 16902 25103 16904
rect 23289 16899 23355 16902
rect 25037 16899 25103 16902
rect 10277 16896 10597 16897
rect 0 16826 480 16856
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4245 16826 4311 16829
rect 0 16824 4311 16826
rect 0 16768 4250 16824
rect 4306 16768 4311 16824
rect 0 16766 4311 16768
rect 0 16736 480 16766
rect 4245 16763 4311 16766
rect 10777 16826 10843 16829
rect 19149 16826 19215 16829
rect 10777 16824 19215 16826
rect 10777 16768 10782 16824
rect 10838 16768 19154 16824
rect 19210 16768 19215 16824
rect 10777 16766 19215 16768
rect 10777 16763 10843 16766
rect 19149 16763 19215 16766
rect 25129 16826 25195 16829
rect 27520 16826 28000 16856
rect 25129 16824 28000 16826
rect 25129 16768 25134 16824
rect 25190 16768 28000 16824
rect 25129 16766 28000 16768
rect 25129 16763 25195 16766
rect 27520 16736 28000 16766
rect 3877 16690 3943 16693
rect 7925 16690 7991 16693
rect 3877 16688 7991 16690
rect 3877 16632 3882 16688
rect 3938 16632 7930 16688
rect 7986 16632 7991 16688
rect 3877 16630 7991 16632
rect 3877 16627 3943 16630
rect 7925 16627 7991 16630
rect 11697 16690 11763 16693
rect 13905 16690 13971 16693
rect 11697 16688 13971 16690
rect 11697 16632 11702 16688
rect 11758 16632 13910 16688
rect 13966 16632 13971 16688
rect 11697 16630 13971 16632
rect 11697 16627 11763 16630
rect 13905 16627 13971 16630
rect 18689 16690 18755 16693
rect 24393 16690 24459 16693
rect 18689 16688 24459 16690
rect 18689 16632 18694 16688
rect 18750 16632 24398 16688
rect 24454 16632 24459 16688
rect 18689 16630 24459 16632
rect 18689 16627 18755 16630
rect 24393 16627 24459 16630
rect 4981 16554 5047 16557
rect 7833 16554 7899 16557
rect 4981 16552 7899 16554
rect 4981 16496 4986 16552
rect 5042 16496 7838 16552
rect 7894 16496 7899 16552
rect 4981 16494 7899 16496
rect 4981 16491 5047 16494
rect 7833 16491 7899 16494
rect 8845 16554 8911 16557
rect 8845 16552 16314 16554
rect 8845 16496 8850 16552
rect 8906 16496 16314 16552
rect 8845 16494 16314 16496
rect 8845 16491 8911 16494
rect 16254 16421 16314 16494
rect 16254 16418 16363 16421
rect 22185 16418 22251 16421
rect 16254 16416 22251 16418
rect 16254 16360 16302 16416
rect 16358 16360 22190 16416
rect 22246 16360 22251 16416
rect 16254 16358 22251 16360
rect 16297 16355 16363 16358
rect 22185 16355 22251 16358
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 2221 16282 2287 16285
rect 6545 16282 6611 16285
rect 7925 16282 7991 16285
rect 0 16280 2287 16282
rect 0 16224 2226 16280
rect 2282 16224 2287 16280
rect 0 16222 2287 16224
rect 0 16192 480 16222
rect 2221 16219 2287 16222
rect 6088 16280 7991 16282
rect 6088 16224 6550 16280
rect 6606 16224 7930 16280
rect 7986 16224 7991 16280
rect 6088 16222 7991 16224
rect 2589 16146 2655 16149
rect 3049 16146 3115 16149
rect 6088 16146 6148 16222
rect 6545 16219 6611 16222
rect 7925 16219 7991 16222
rect 10869 16282 10935 16285
rect 14181 16282 14247 16285
rect 10869 16280 14247 16282
rect 10869 16224 10874 16280
rect 10930 16224 14186 16280
rect 14242 16224 14247 16280
rect 10869 16222 14247 16224
rect 10869 16219 10935 16222
rect 14181 16219 14247 16222
rect 25773 16282 25839 16285
rect 27520 16282 28000 16312
rect 25773 16280 28000 16282
rect 25773 16224 25778 16280
rect 25834 16224 28000 16280
rect 25773 16222 28000 16224
rect 25773 16219 25839 16222
rect 27520 16192 28000 16222
rect 2589 16144 6148 16146
rect 2589 16088 2594 16144
rect 2650 16088 3054 16144
rect 3110 16088 6148 16144
rect 2589 16086 6148 16088
rect 6361 16146 6427 16149
rect 22369 16146 22435 16149
rect 6361 16144 22435 16146
rect 6361 16088 6366 16144
rect 6422 16088 22374 16144
rect 22430 16088 22435 16144
rect 6361 16086 22435 16088
rect 2589 16083 2655 16086
rect 3049 16083 3115 16086
rect 6361 16083 6427 16086
rect 22369 16083 22435 16086
rect 24117 16144 24183 16149
rect 24117 16088 24122 16144
rect 24178 16088 24183 16144
rect 24117 16083 24183 16088
rect 2037 16010 2103 16013
rect 7005 16010 7071 16013
rect 2037 16008 7071 16010
rect 2037 15952 2042 16008
rect 2098 15952 7010 16008
rect 7066 15952 7071 16008
rect 2037 15950 7071 15952
rect 2037 15947 2103 15950
rect 7005 15947 7071 15950
rect 13537 16010 13603 16013
rect 15469 16010 15535 16013
rect 13537 16008 15535 16010
rect 13537 15952 13542 16008
rect 13598 15952 15474 16008
rect 15530 15952 15535 16008
rect 13537 15950 15535 15952
rect 13537 15947 13603 15950
rect 15469 15947 15535 15950
rect 16021 16010 16087 16013
rect 24120 16010 24180 16083
rect 16021 16008 24180 16010
rect 16021 15952 16026 16008
rect 16082 15952 24180 16008
rect 16021 15950 24180 15952
rect 16021 15947 16087 15950
rect 2773 15874 2839 15877
rect 8845 15874 8911 15877
rect 2773 15872 8911 15874
rect 2773 15816 2778 15872
rect 2834 15816 8850 15872
rect 8906 15816 8911 15872
rect 2773 15814 8911 15816
rect 2773 15811 2839 15814
rect 8845 15811 8911 15814
rect 10777 15874 10843 15877
rect 14365 15874 14431 15877
rect 10777 15872 14431 15874
rect 10777 15816 10782 15872
rect 10838 15816 14370 15872
rect 14426 15816 14431 15872
rect 10777 15814 14431 15816
rect 10777 15811 10843 15814
rect 14365 15811 14431 15814
rect 14825 15874 14891 15877
rect 19333 15874 19399 15877
rect 14825 15872 19399 15874
rect 14825 15816 14830 15872
rect 14886 15816 19338 15872
rect 19394 15816 19399 15872
rect 14825 15814 19399 15816
rect 14825 15811 14891 15814
rect 19333 15811 19399 15814
rect 10277 15808 10597 15809
rect 0 15738 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 1577 15738 1643 15741
rect 0 15736 1643 15738
rect 0 15680 1582 15736
rect 1638 15680 1643 15736
rect 0 15678 1643 15680
rect 0 15648 480 15678
rect 1577 15675 1643 15678
rect 3509 15738 3575 15741
rect 7465 15738 7531 15741
rect 3509 15736 7531 15738
rect 3509 15680 3514 15736
rect 3570 15680 7470 15736
rect 7526 15680 7531 15736
rect 3509 15678 7531 15680
rect 3509 15675 3575 15678
rect 7465 15675 7531 15678
rect 9990 15676 9996 15740
rect 10060 15738 10066 15740
rect 10133 15738 10199 15741
rect 10060 15736 10199 15738
rect 10060 15680 10138 15736
rect 10194 15680 10199 15736
rect 10060 15678 10199 15680
rect 10060 15676 10066 15678
rect 10133 15675 10199 15678
rect 10961 15738 11027 15741
rect 12801 15738 12867 15741
rect 10961 15736 12867 15738
rect 10961 15680 10966 15736
rect 11022 15680 12806 15736
rect 12862 15680 12867 15736
rect 10961 15678 12867 15680
rect 10961 15675 11027 15678
rect 12801 15675 12867 15678
rect 13721 15738 13787 15741
rect 15469 15738 15535 15741
rect 13721 15736 15535 15738
rect 13721 15680 13726 15736
rect 13782 15680 15474 15736
rect 15530 15680 15535 15736
rect 13721 15678 15535 15680
rect 13721 15675 13787 15678
rect 15469 15675 15535 15678
rect 23749 15738 23815 15741
rect 27520 15738 28000 15768
rect 23749 15736 28000 15738
rect 23749 15680 23754 15736
rect 23810 15680 28000 15736
rect 23749 15678 28000 15680
rect 23749 15675 23815 15678
rect 27520 15648 28000 15678
rect 7005 15602 7071 15605
rect 8017 15602 8083 15605
rect 7005 15600 8083 15602
rect 7005 15544 7010 15600
rect 7066 15544 8022 15600
rect 8078 15544 8083 15600
rect 7005 15542 8083 15544
rect 7005 15539 7071 15542
rect 8017 15539 8083 15542
rect 8753 15602 8819 15605
rect 14365 15602 14431 15605
rect 17401 15602 17467 15605
rect 8753 15600 14290 15602
rect 8753 15544 8758 15600
rect 8814 15544 14290 15600
rect 8753 15542 14290 15544
rect 8753 15539 8819 15542
rect 4337 15466 4403 15469
rect 8293 15466 8359 15469
rect 4337 15464 8359 15466
rect 4337 15408 4342 15464
rect 4398 15408 8298 15464
rect 8354 15408 8359 15464
rect 4337 15406 8359 15408
rect 4337 15403 4403 15406
rect 8293 15403 8359 15406
rect 11053 15466 11119 15469
rect 13261 15466 13327 15469
rect 11053 15464 13327 15466
rect 11053 15408 11058 15464
rect 11114 15408 13266 15464
rect 13322 15408 13327 15464
rect 11053 15406 13327 15408
rect 14230 15466 14290 15542
rect 14365 15600 17467 15602
rect 14365 15544 14370 15600
rect 14426 15544 17406 15600
rect 17462 15544 17467 15600
rect 14365 15542 17467 15544
rect 14365 15539 14431 15542
rect 17401 15539 17467 15542
rect 17217 15466 17283 15469
rect 14230 15464 17283 15466
rect 14230 15408 17222 15464
rect 17278 15408 17283 15464
rect 14230 15406 17283 15408
rect 11053 15403 11119 15406
rect 13261 15403 13327 15406
rect 17217 15403 17283 15406
rect 20713 15466 20779 15469
rect 25405 15466 25471 15469
rect 20713 15464 25471 15466
rect 20713 15408 20718 15464
rect 20774 15408 25410 15464
rect 25466 15408 25471 15464
rect 20713 15406 25471 15408
rect 20713 15403 20779 15406
rect 25405 15403 25471 15406
rect 10777 15330 10843 15333
rect 13353 15330 13419 15333
rect 10777 15328 13419 15330
rect 10777 15272 10782 15328
rect 10838 15272 13358 15328
rect 13414 15272 13419 15328
rect 10777 15270 13419 15272
rect 10777 15267 10843 15270
rect 13353 15267 13419 15270
rect 15745 15330 15811 15333
rect 16849 15330 16915 15333
rect 23473 15330 23539 15333
rect 15745 15328 23539 15330
rect 15745 15272 15750 15328
rect 15806 15272 16854 15328
rect 16910 15272 23478 15328
rect 23534 15272 23539 15328
rect 15745 15270 23539 15272
rect 15745 15267 15811 15270
rect 16849 15267 16915 15270
rect 23473 15267 23539 15270
rect 5610 15264 5930 15265
rect 0 15194 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 1577 15194 1643 15197
rect 0 15192 1643 15194
rect 0 15136 1582 15192
rect 1638 15136 1643 15192
rect 0 15134 1643 15136
rect 0 15104 480 15134
rect 1577 15131 1643 15134
rect 15929 15194 15995 15197
rect 19977 15194 20043 15197
rect 27520 15194 28000 15224
rect 15929 15192 20043 15194
rect 15929 15136 15934 15192
rect 15990 15136 19982 15192
rect 20038 15136 20043 15192
rect 15929 15134 20043 15136
rect 15929 15131 15995 15134
rect 19977 15131 20043 15134
rect 24672 15134 28000 15194
rect 5533 15058 5599 15061
rect 8845 15058 8911 15061
rect 5533 15056 8911 15058
rect 5533 15000 5538 15056
rect 5594 15000 8850 15056
rect 8906 15000 8911 15056
rect 5533 14998 8911 15000
rect 5533 14995 5599 14998
rect 8845 14995 8911 14998
rect 9029 15058 9095 15061
rect 12893 15058 12959 15061
rect 9029 15056 12959 15058
rect 9029 15000 9034 15056
rect 9090 15000 12898 15056
rect 12954 15000 12959 15056
rect 9029 14998 12959 15000
rect 9029 14995 9095 14998
rect 12893 14995 12959 14998
rect 22645 15058 22711 15061
rect 24672 15058 24732 15134
rect 27520 15104 28000 15134
rect 22645 15056 24732 15058
rect 22645 15000 22650 15056
rect 22706 15000 24732 15056
rect 22645 14998 24732 15000
rect 22645 14995 22711 14998
rect 2957 14922 3023 14925
rect 10593 14922 10659 14925
rect 2957 14920 10659 14922
rect 2957 14864 2962 14920
rect 3018 14864 10598 14920
rect 10654 14864 10659 14920
rect 2957 14862 10659 14864
rect 2957 14859 3023 14862
rect 10593 14859 10659 14862
rect 18505 14922 18571 14925
rect 25221 14922 25287 14925
rect 18505 14920 25287 14922
rect 18505 14864 18510 14920
rect 18566 14864 25226 14920
rect 25282 14864 25287 14920
rect 18505 14862 25287 14864
rect 18505 14859 18571 14862
rect 25221 14859 25287 14862
rect 2865 14786 2931 14789
rect 8109 14786 8175 14789
rect 2865 14784 8175 14786
rect 2865 14728 2870 14784
rect 2926 14728 8114 14784
rect 8170 14728 8175 14784
rect 2865 14726 8175 14728
rect 2865 14723 2931 14726
rect 8109 14723 8175 14726
rect 20161 14786 20227 14789
rect 23422 14786 23428 14788
rect 20161 14784 23428 14786
rect 20161 14728 20166 14784
rect 20222 14728 23428 14784
rect 20161 14726 23428 14728
rect 20161 14723 20227 14726
rect 23422 14724 23428 14726
rect 23492 14724 23498 14788
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1577 14650 1643 14653
rect 0 14648 1643 14650
rect 0 14592 1582 14648
rect 1638 14592 1643 14648
rect 0 14590 1643 14592
rect 0 14560 480 14590
rect 1577 14587 1643 14590
rect 13169 14650 13235 14653
rect 19241 14650 19307 14653
rect 13169 14648 19307 14650
rect 13169 14592 13174 14648
rect 13230 14592 19246 14648
rect 19302 14592 19307 14648
rect 13169 14590 19307 14592
rect 13169 14587 13235 14590
rect 19241 14587 19307 14590
rect 21449 14650 21515 14653
rect 27520 14650 28000 14680
rect 21449 14648 28000 14650
rect 21449 14592 21454 14648
rect 21510 14592 28000 14648
rect 21449 14590 28000 14592
rect 21449 14587 21515 14590
rect 27520 14560 28000 14590
rect 2405 14514 2471 14517
rect 3509 14514 3575 14517
rect 2405 14512 3575 14514
rect 2405 14456 2410 14512
rect 2466 14456 3514 14512
rect 3570 14456 3575 14512
rect 2405 14454 3575 14456
rect 2405 14451 2471 14454
rect 3509 14451 3575 14454
rect 4521 14514 4587 14517
rect 10133 14514 10199 14517
rect 4521 14512 10199 14514
rect 4521 14456 4526 14512
rect 4582 14456 10138 14512
rect 10194 14456 10199 14512
rect 4521 14454 10199 14456
rect 4521 14451 4587 14454
rect 10133 14451 10199 14454
rect 19241 14514 19307 14517
rect 22277 14514 22343 14517
rect 19241 14512 22343 14514
rect 19241 14456 19246 14512
rect 19302 14456 22282 14512
rect 22338 14456 22343 14512
rect 19241 14454 22343 14456
rect 19241 14451 19307 14454
rect 22277 14451 22343 14454
rect 5349 14378 5415 14381
rect 7741 14378 7807 14381
rect 5349 14376 7807 14378
rect 5349 14320 5354 14376
rect 5410 14320 7746 14376
rect 7802 14320 7807 14376
rect 5349 14318 7807 14320
rect 5349 14315 5415 14318
rect 7741 14315 7807 14318
rect 9622 14316 9628 14380
rect 9692 14378 9698 14380
rect 12157 14378 12223 14381
rect 9692 14376 12223 14378
rect 9692 14320 12162 14376
rect 12218 14320 12223 14376
rect 9692 14318 12223 14320
rect 9692 14316 9698 14318
rect 12157 14315 12223 14318
rect 12341 14378 12407 14381
rect 20713 14378 20779 14381
rect 12341 14376 20779 14378
rect 12341 14320 12346 14376
rect 12402 14320 20718 14376
rect 20774 14320 20779 14376
rect 12341 14318 20779 14320
rect 12341 14315 12407 14318
rect 20713 14315 20779 14318
rect 7281 14242 7347 14245
rect 9581 14242 9647 14245
rect 9949 14242 10015 14245
rect 14181 14242 14247 14245
rect 7281 14240 9460 14242
rect 7281 14184 7286 14240
rect 7342 14184 9460 14240
rect 7281 14182 9460 14184
rect 7281 14179 7347 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 9400 14106 9460 14182
rect 9581 14240 14247 14242
rect 9581 14184 9586 14240
rect 9642 14184 9954 14240
rect 10010 14184 14186 14240
rect 14242 14184 14247 14240
rect 9581 14182 14247 14184
rect 9581 14179 9647 14182
rect 9949 14179 10015 14182
rect 14181 14179 14247 14182
rect 15377 14242 15443 14245
rect 23473 14242 23539 14245
rect 15377 14240 23539 14242
rect 15377 14184 15382 14240
rect 15438 14184 23478 14240
rect 23534 14184 23539 14240
rect 15377 14182 23539 14184
rect 15377 14179 15443 14182
rect 23473 14179 23539 14182
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 9622 14106 9628 14108
rect 9400 14046 9628 14106
rect 9622 14044 9628 14046
rect 9692 14044 9698 14108
rect 21265 14106 21331 14109
rect 20118 14104 21331 14106
rect 20118 14048 21270 14104
rect 21326 14048 21331 14104
rect 20118 14046 21331 14048
rect 0 13970 480 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 0 13880 480 13910
rect 1485 13907 1551 13910
rect 4705 13970 4771 13973
rect 7097 13970 7163 13973
rect 4705 13968 7163 13970
rect 4705 13912 4710 13968
rect 4766 13912 7102 13968
rect 7158 13912 7163 13968
rect 4705 13910 7163 13912
rect 4705 13907 4771 13910
rect 7097 13907 7163 13910
rect 14222 13908 14228 13972
rect 14292 13970 14298 13972
rect 20118 13970 20178 14046
rect 21265 14043 21331 14046
rect 14292 13910 20178 13970
rect 26049 13970 26115 13973
rect 27520 13970 28000 14000
rect 26049 13968 28000 13970
rect 26049 13912 26054 13968
rect 26110 13912 28000 13968
rect 26049 13910 28000 13912
rect 14292 13908 14298 13910
rect 26049 13907 26115 13910
rect 27520 13880 28000 13910
rect 21909 13834 21975 13837
rect 24117 13834 24183 13837
rect 21909 13832 24183 13834
rect 21909 13776 21914 13832
rect 21970 13776 24122 13832
rect 24178 13776 24183 13832
rect 21909 13774 24183 13776
rect 21909 13771 21975 13774
rect 24117 13771 24183 13774
rect 8150 13636 8156 13700
rect 8220 13636 8226 13700
rect 13537 13698 13603 13701
rect 15377 13698 15443 13701
rect 24669 13700 24735 13701
rect 24669 13698 24716 13700
rect 13537 13696 15443 13698
rect 13537 13640 13542 13696
rect 13598 13640 15382 13696
rect 15438 13640 15443 13696
rect 13537 13638 15443 13640
rect 24624 13696 24716 13698
rect 24624 13640 24674 13696
rect 24624 13638 24716 13640
rect 8158 13562 8218 13636
rect 13537 13635 13603 13638
rect 15377 13635 15443 13638
rect 24669 13636 24716 13638
rect 24780 13636 24786 13700
rect 24669 13635 24735 13636
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 8661 13562 8727 13565
rect 8158 13560 8727 13562
rect 8158 13504 8666 13560
rect 8722 13504 8727 13560
rect 8158 13502 8727 13504
rect 8661 13499 8727 13502
rect 10777 13562 10843 13565
rect 15469 13562 15535 13565
rect 10777 13560 15535 13562
rect 10777 13504 10782 13560
rect 10838 13504 15474 13560
rect 15530 13504 15535 13560
rect 10777 13502 15535 13504
rect 10777 13499 10843 13502
rect 15469 13499 15535 13502
rect 0 13426 480 13456
rect 1577 13426 1643 13429
rect 0 13424 1643 13426
rect 0 13368 1582 13424
rect 1638 13368 1643 13424
rect 0 13366 1643 13368
rect 0 13336 480 13366
rect 1577 13363 1643 13366
rect 8109 13426 8175 13429
rect 13445 13426 13511 13429
rect 8109 13424 13511 13426
rect 8109 13368 8114 13424
rect 8170 13368 13450 13424
rect 13506 13368 13511 13424
rect 8109 13366 13511 13368
rect 8109 13363 8175 13366
rect 13445 13363 13511 13366
rect 15745 13426 15811 13429
rect 24761 13426 24827 13429
rect 27520 13426 28000 13456
rect 15745 13424 22938 13426
rect 15745 13368 15750 13424
rect 15806 13368 22938 13424
rect 15745 13366 22938 13368
rect 15745 13363 15811 13366
rect 3049 13290 3115 13293
rect 7281 13290 7347 13293
rect 13077 13290 13143 13293
rect 3049 13288 7347 13290
rect 3049 13232 3054 13288
rect 3110 13232 7286 13288
rect 7342 13232 7347 13288
rect 8112 13288 13143 13290
rect 8112 13259 13082 13288
rect 3049 13230 7347 13232
rect 3049 13227 3115 13230
rect 7281 13227 7347 13230
rect 8109 13254 13082 13259
rect 8109 13198 8114 13254
rect 8170 13232 13082 13254
rect 13138 13232 13143 13288
rect 8170 13230 13143 13232
rect 8170 13198 8175 13230
rect 13077 13227 13143 13230
rect 13261 13290 13327 13293
rect 19149 13290 19215 13293
rect 13261 13288 19215 13290
rect 13261 13232 13266 13288
rect 13322 13232 19154 13288
rect 19210 13232 19215 13288
rect 13261 13230 19215 13232
rect 13261 13227 13327 13230
rect 19149 13227 19215 13230
rect 8109 13193 8175 13198
rect 9029 13154 9095 13157
rect 13905 13154 13971 13157
rect 9029 13152 13971 13154
rect 9029 13096 9034 13152
rect 9090 13096 13910 13152
rect 13966 13096 13971 13152
rect 9029 13094 13971 13096
rect 9029 13091 9095 13094
rect 13905 13091 13971 13094
rect 16297 13154 16363 13157
rect 18045 13154 18111 13157
rect 16297 13152 18111 13154
rect 16297 13096 16302 13152
rect 16358 13096 18050 13152
rect 18106 13096 18111 13152
rect 16297 13094 18111 13096
rect 16297 13091 16363 13094
rect 18045 13091 18111 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 0 12882 480 12912
rect 2681 12882 2747 12885
rect 0 12880 2747 12882
rect 0 12824 2686 12880
rect 2742 12824 2747 12880
rect 0 12822 2747 12824
rect 0 12792 480 12822
rect 2681 12819 2747 12822
rect 3141 12882 3207 12885
rect 5625 12882 5691 12885
rect 3141 12880 5691 12882
rect 3141 12824 3146 12880
rect 3202 12824 5630 12880
rect 5686 12824 5691 12880
rect 3141 12822 5691 12824
rect 3141 12819 3207 12822
rect 5625 12819 5691 12822
rect 11421 12882 11487 12885
rect 13261 12882 13327 12885
rect 11421 12880 13327 12882
rect 11421 12824 11426 12880
rect 11482 12824 13266 12880
rect 13322 12824 13327 12880
rect 11421 12822 13327 12824
rect 11421 12819 11487 12822
rect 13261 12819 13327 12822
rect 13997 12882 14063 12885
rect 22737 12882 22803 12885
rect 13997 12880 22803 12882
rect 13997 12824 14002 12880
rect 14058 12824 22742 12880
rect 22798 12824 22803 12880
rect 13997 12822 22803 12824
rect 22878 12882 22938 13366
rect 24761 13424 28000 13426
rect 24761 13368 24766 13424
rect 24822 13368 28000 13424
rect 24761 13366 28000 13368
rect 24761 13363 24827 13366
rect 27520 13336 28000 13366
rect 23105 13290 23171 13293
rect 25221 13290 25287 13293
rect 23105 13288 25287 13290
rect 23105 13232 23110 13288
rect 23166 13232 25226 13288
rect 25282 13232 25287 13288
rect 23105 13230 25287 13232
rect 23105 13227 23171 13230
rect 25221 13227 25287 13230
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 25221 12882 25287 12885
rect 22878 12880 25287 12882
rect 22878 12824 25226 12880
rect 25282 12824 25287 12880
rect 22878 12822 25287 12824
rect 13997 12819 14063 12822
rect 22737 12819 22803 12822
rect 25221 12819 25287 12822
rect 25497 12882 25563 12885
rect 27520 12882 28000 12912
rect 25497 12880 28000 12882
rect 25497 12824 25502 12880
rect 25558 12824 28000 12880
rect 25497 12822 28000 12824
rect 25497 12819 25563 12822
rect 27520 12792 28000 12822
rect 2037 12746 2103 12749
rect 9121 12746 9187 12749
rect 2037 12744 9187 12746
rect 2037 12688 2042 12744
rect 2098 12688 9126 12744
rect 9182 12688 9187 12744
rect 2037 12686 9187 12688
rect 2037 12683 2103 12686
rect 9121 12683 9187 12686
rect 9489 12746 9555 12749
rect 12525 12746 12591 12749
rect 9489 12744 12591 12746
rect 9489 12688 9494 12744
rect 9550 12688 12530 12744
rect 12586 12688 12591 12744
rect 9489 12686 12591 12688
rect 9489 12683 9555 12686
rect 12525 12683 12591 12686
rect 13077 12746 13143 12749
rect 17033 12746 17099 12749
rect 17677 12746 17743 12749
rect 13077 12744 17743 12746
rect 13077 12688 13082 12744
rect 13138 12688 17038 12744
rect 17094 12688 17682 12744
rect 17738 12688 17743 12744
rect 13077 12686 17743 12688
rect 13077 12683 13143 12686
rect 17033 12683 17099 12686
rect 17677 12683 17743 12686
rect 18505 12746 18571 12749
rect 19241 12746 19307 12749
rect 23289 12746 23355 12749
rect 18505 12744 23355 12746
rect 18505 12688 18510 12744
rect 18566 12688 19246 12744
rect 19302 12688 23294 12744
rect 23350 12688 23355 12744
rect 18505 12686 23355 12688
rect 18505 12683 18571 12686
rect 19241 12683 19307 12686
rect 23289 12683 23355 12686
rect 3141 12610 3207 12613
rect 7833 12610 7899 12613
rect 3141 12608 7899 12610
rect 3141 12552 3146 12608
rect 3202 12552 7838 12608
rect 7894 12552 7899 12608
rect 3141 12550 7899 12552
rect 3141 12547 3207 12550
rect 7833 12547 7899 12550
rect 20713 12610 20779 12613
rect 23657 12610 23723 12613
rect 20713 12608 23723 12610
rect 20713 12552 20718 12608
rect 20774 12552 23662 12608
rect 23718 12552 23723 12608
rect 20713 12550 23723 12552
rect 20713 12547 20779 12550
rect 23657 12547 23723 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 4705 12474 4771 12477
rect 10041 12474 10107 12477
rect 4705 12472 10107 12474
rect 4705 12416 4710 12472
rect 4766 12416 10046 12472
rect 10102 12416 10107 12472
rect 4705 12414 10107 12416
rect 4705 12411 4771 12414
rect 10041 12411 10107 12414
rect 14549 12472 14615 12477
rect 14549 12416 14554 12472
rect 14610 12416 14615 12472
rect 14549 12411 14615 12416
rect 23473 12474 23539 12477
rect 24485 12474 24551 12477
rect 24669 12474 24735 12477
rect 23473 12472 23674 12474
rect 23473 12416 23478 12472
rect 23534 12416 23674 12472
rect 23473 12414 23674 12416
rect 23473 12411 23539 12414
rect 0 12338 480 12368
rect 14552 12341 14612 12411
rect 1761 12338 1827 12341
rect 0 12336 1827 12338
rect 0 12280 1766 12336
rect 1822 12280 1827 12336
rect 0 12278 1827 12280
rect 0 12248 480 12278
rect 1761 12275 1827 12278
rect 14549 12336 14615 12341
rect 14549 12280 14554 12336
rect 14610 12280 14615 12336
rect 14549 12275 14615 12280
rect 23614 12338 23674 12414
rect 24485 12472 24735 12474
rect 24485 12416 24490 12472
rect 24546 12416 24674 12472
rect 24730 12416 24735 12472
rect 24485 12414 24735 12416
rect 24485 12411 24551 12414
rect 24669 12411 24735 12414
rect 25405 12440 25471 12443
rect 25405 12438 25514 12440
rect 25405 12382 25410 12438
rect 25466 12382 25514 12438
rect 25405 12377 25514 12382
rect 24669 12338 24735 12341
rect 23614 12336 24735 12338
rect 23614 12280 24674 12336
rect 24730 12280 24735 12336
rect 23614 12278 24735 12280
rect 24669 12275 24735 12278
rect 25037 12338 25103 12341
rect 25454 12338 25514 12377
rect 27520 12338 28000 12368
rect 25037 12336 25330 12338
rect 25037 12280 25042 12336
rect 25098 12280 25330 12336
rect 25037 12278 25330 12280
rect 25454 12278 28000 12338
rect 25037 12275 25103 12278
rect 11421 12202 11487 12205
rect 16205 12202 16271 12205
rect 11421 12200 16271 12202
rect 11421 12144 11426 12200
rect 11482 12144 16210 12200
rect 16266 12144 16271 12200
rect 11421 12142 16271 12144
rect 11421 12139 11487 12142
rect 16205 12139 16271 12142
rect 20621 12202 20687 12205
rect 24393 12202 24459 12205
rect 20621 12200 24459 12202
rect 20621 12144 20626 12200
rect 20682 12144 24398 12200
rect 24454 12144 24459 12200
rect 20621 12142 24459 12144
rect 25270 12202 25330 12278
rect 27520 12248 28000 12278
rect 25497 12202 25563 12205
rect 25270 12200 25563 12202
rect 25270 12144 25502 12200
rect 25558 12144 25563 12200
rect 25270 12142 25563 12144
rect 20621 12139 20687 12142
rect 24393 12139 24459 12142
rect 25497 12139 25563 12142
rect 11697 12066 11763 12069
rect 14457 12066 14523 12069
rect 11697 12064 14523 12066
rect 11697 12008 11702 12064
rect 11758 12008 14462 12064
rect 14518 12008 14523 12064
rect 11697 12006 14523 12008
rect 11697 12003 11763 12006
rect 14457 12003 14523 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 14089 11930 14155 11933
rect 14222 11930 14228 11932
rect 14089 11928 14228 11930
rect 14089 11872 14094 11928
rect 14150 11872 14228 11928
rect 14089 11870 14228 11872
rect 14089 11867 14155 11870
rect 14222 11868 14228 11870
rect 14292 11868 14298 11932
rect 18873 11930 18939 11933
rect 19241 11930 19307 11933
rect 24025 11930 24091 11933
rect 18873 11928 24091 11930
rect 18873 11872 18878 11928
rect 18934 11872 19246 11928
rect 19302 11872 24030 11928
rect 24086 11872 24091 11928
rect 18873 11870 24091 11872
rect 18873 11867 18939 11870
rect 19241 11867 19307 11870
rect 24025 11867 24091 11870
rect 0 11794 480 11824
rect 2957 11794 3023 11797
rect 0 11792 3023 11794
rect 0 11736 2962 11792
rect 3018 11736 3023 11792
rect 0 11734 3023 11736
rect 0 11704 480 11734
rect 2957 11731 3023 11734
rect 11145 11794 11211 11797
rect 15653 11794 15719 11797
rect 11145 11792 15719 11794
rect 11145 11736 11150 11792
rect 11206 11736 15658 11792
rect 15714 11736 15719 11792
rect 11145 11734 15719 11736
rect 11145 11731 11211 11734
rect 15653 11731 15719 11734
rect 16113 11794 16179 11797
rect 17953 11794 18019 11797
rect 16113 11792 18019 11794
rect 16113 11736 16118 11792
rect 16174 11736 17958 11792
rect 18014 11736 18019 11792
rect 16113 11734 18019 11736
rect 16113 11731 16179 11734
rect 17953 11731 18019 11734
rect 22277 11794 22343 11797
rect 27520 11794 28000 11824
rect 22277 11792 28000 11794
rect 22277 11736 22282 11792
rect 22338 11736 28000 11792
rect 22277 11734 28000 11736
rect 22277 11731 22343 11734
rect 27520 11704 28000 11734
rect 9397 11658 9463 11661
rect 11789 11658 11855 11661
rect 9397 11656 11855 11658
rect 9397 11600 9402 11656
rect 9458 11600 11794 11656
rect 11850 11600 11855 11656
rect 9397 11598 11855 11600
rect 9397 11595 9463 11598
rect 11789 11595 11855 11598
rect 19333 11658 19399 11661
rect 22461 11658 22527 11661
rect 19333 11656 22527 11658
rect 19333 11600 19338 11656
rect 19394 11600 22466 11656
rect 22522 11600 22527 11656
rect 19333 11598 22527 11600
rect 19333 11595 19399 11598
rect 22461 11595 22527 11598
rect 23422 11596 23428 11660
rect 23492 11658 23498 11660
rect 23657 11658 23723 11661
rect 23492 11656 23723 11658
rect 23492 11600 23662 11656
rect 23718 11600 23723 11656
rect 23492 11598 23723 11600
rect 23492 11596 23498 11598
rect 23657 11595 23723 11598
rect 15561 11522 15627 11525
rect 17861 11522 17927 11525
rect 15561 11520 17927 11522
rect 15561 11464 15566 11520
rect 15622 11464 17866 11520
rect 17922 11464 17927 11520
rect 15561 11462 17927 11464
rect 15561 11459 15627 11462
rect 17861 11459 17927 11462
rect 20437 11522 20503 11525
rect 24301 11522 24367 11525
rect 20437 11520 24367 11522
rect 20437 11464 20442 11520
rect 20498 11464 24306 11520
rect 24362 11464 24367 11520
rect 20437 11462 24367 11464
rect 20437 11459 20503 11462
rect 24301 11459 24367 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 4429 11386 4495 11389
rect 8385 11386 8451 11389
rect 4429 11384 8451 11386
rect 4429 11328 4434 11384
rect 4490 11328 8390 11384
rect 8446 11328 8451 11384
rect 4429 11326 8451 11328
rect 4429 11323 4495 11326
rect 8385 11323 8451 11326
rect 14181 11386 14247 11389
rect 17953 11386 18019 11389
rect 14181 11384 18019 11386
rect 14181 11328 14186 11384
rect 14242 11328 17958 11384
rect 18014 11328 18019 11384
rect 14181 11326 18019 11328
rect 14181 11323 14247 11326
rect 17953 11323 18019 11326
rect 20069 11386 20135 11389
rect 23473 11386 23539 11389
rect 20069 11384 23539 11386
rect 20069 11328 20074 11384
rect 20130 11328 23478 11384
rect 23534 11328 23539 11384
rect 20069 11326 23539 11328
rect 20069 11323 20135 11326
rect 23473 11323 23539 11326
rect 24669 11386 24735 11389
rect 24669 11384 25882 11386
rect 24669 11328 24674 11384
rect 24730 11328 25882 11384
rect 24669 11326 25882 11328
rect 24669 11323 24735 11326
rect 9213 11250 9279 11253
rect 12065 11250 12131 11253
rect 9213 11248 12131 11250
rect 9213 11192 9218 11248
rect 9274 11192 12070 11248
rect 12126 11192 12131 11248
rect 9213 11190 12131 11192
rect 9213 11187 9279 11190
rect 12065 11187 12131 11190
rect 13813 11250 13879 11253
rect 25589 11250 25655 11253
rect 13813 11248 25655 11250
rect 13813 11192 13818 11248
rect 13874 11192 25594 11248
rect 25650 11192 25655 11248
rect 13813 11190 25655 11192
rect 13813 11187 13879 11190
rect 25589 11187 25655 11190
rect 0 11114 480 11144
rect 4705 11114 4771 11117
rect 0 11112 4771 11114
rect 0 11056 4710 11112
rect 4766 11056 4771 11112
rect 0 11054 4771 11056
rect 0 11024 480 11054
rect 4705 11051 4771 11054
rect 10041 11114 10107 11117
rect 12893 11114 12959 11117
rect 10041 11112 12959 11114
rect 10041 11056 10046 11112
rect 10102 11056 12898 11112
rect 12954 11056 12959 11112
rect 10041 11054 12959 11056
rect 10041 11051 10107 11054
rect 12893 11051 12959 11054
rect 21265 11114 21331 11117
rect 25405 11114 25471 11117
rect 21265 11112 25471 11114
rect 21265 11056 21270 11112
rect 21326 11056 25410 11112
rect 25466 11056 25471 11112
rect 21265 11054 25471 11056
rect 25822 11114 25882 11326
rect 27520 11114 28000 11144
rect 25822 11054 28000 11114
rect 21265 11051 21331 11054
rect 25405 11051 25471 11054
rect 27520 11024 28000 11054
rect 18137 10978 18203 10981
rect 20069 10978 20135 10981
rect 18137 10976 20135 10978
rect 18137 10920 18142 10976
rect 18198 10920 20074 10976
rect 20130 10920 20135 10976
rect 18137 10918 20135 10920
rect 18137 10915 18203 10918
rect 20069 10915 20135 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 4061 10706 4127 10709
rect 17125 10706 17191 10709
rect 4061 10704 17191 10706
rect 4061 10648 4066 10704
rect 4122 10648 17130 10704
rect 17186 10648 17191 10704
rect 4061 10646 17191 10648
rect 4061 10643 4127 10646
rect 17125 10643 17191 10646
rect 17677 10706 17743 10709
rect 24945 10706 25011 10709
rect 17677 10704 25011 10706
rect 17677 10648 17682 10704
rect 17738 10648 24950 10704
rect 25006 10648 25011 10704
rect 17677 10646 25011 10648
rect 17677 10643 17743 10646
rect 24945 10643 25011 10646
rect 0 10570 480 10600
rect 13629 10570 13695 10573
rect 0 10568 13695 10570
rect 0 10512 13634 10568
rect 13690 10512 13695 10568
rect 0 10510 13695 10512
rect 0 10480 480 10510
rect 13629 10507 13695 10510
rect 19977 10570 20043 10573
rect 24301 10570 24367 10573
rect 27520 10570 28000 10600
rect 19977 10568 24367 10570
rect 19977 10512 19982 10568
rect 20038 10512 24306 10568
rect 24362 10512 24367 10568
rect 19977 10510 24367 10512
rect 19977 10507 20043 10510
rect 24301 10507 24367 10510
rect 24902 10510 28000 10570
rect 2405 10434 2471 10437
rect 3877 10434 3943 10437
rect 10133 10434 10199 10437
rect 2405 10432 3802 10434
rect 2405 10376 2410 10432
rect 2466 10376 3802 10432
rect 2405 10374 3802 10376
rect 2405 10371 2471 10374
rect 3742 10162 3802 10374
rect 3877 10432 10199 10434
rect 3877 10376 3882 10432
rect 3938 10376 10138 10432
rect 10194 10376 10199 10432
rect 3877 10374 10199 10376
rect 3877 10371 3943 10374
rect 10133 10371 10199 10374
rect 13629 10434 13695 10437
rect 18965 10434 19031 10437
rect 13629 10432 19031 10434
rect 13629 10376 13634 10432
rect 13690 10376 18970 10432
rect 19026 10376 19031 10432
rect 13629 10374 19031 10376
rect 13629 10371 13695 10374
rect 18965 10371 19031 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 13169 10298 13235 10301
rect 13169 10296 14658 10298
rect 13169 10240 13174 10296
rect 13230 10240 14658 10296
rect 13169 10238 14658 10240
rect 13169 10235 13235 10238
rect 10041 10162 10107 10165
rect 14457 10162 14523 10165
rect 3742 10160 14523 10162
rect 3742 10104 10046 10160
rect 10102 10104 14462 10160
rect 14518 10104 14523 10160
rect 3742 10102 14523 10104
rect 14598 10162 14658 10238
rect 24902 10162 24962 10510
rect 27520 10480 28000 10510
rect 14598 10102 24962 10162
rect 10041 10099 10107 10102
rect 14457 10099 14523 10102
rect 0 10026 480 10056
rect 4061 10026 4127 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 480 9966
rect 4061 9963 4127 9966
rect 14181 10026 14247 10029
rect 17309 10026 17375 10029
rect 24945 10026 25011 10029
rect 27520 10026 28000 10056
rect 14181 10024 17375 10026
rect 14181 9968 14186 10024
rect 14242 9968 17314 10024
rect 17370 9968 17375 10024
rect 14181 9966 17375 9968
rect 14181 9963 14247 9966
rect 17309 9963 17375 9966
rect 24120 9966 24778 10026
rect 15469 9890 15535 9893
rect 19149 9890 19215 9893
rect 15469 9888 19215 9890
rect 15469 9832 15474 9888
rect 15530 9832 19154 9888
rect 19210 9832 19215 9888
rect 15469 9830 19215 9832
rect 15469 9827 15535 9830
rect 19149 9827 19215 9830
rect 19977 9890 20043 9893
rect 23841 9890 23907 9893
rect 19977 9888 23907 9890
rect 19977 9832 19982 9888
rect 20038 9832 23846 9888
rect 23902 9832 23907 9888
rect 19977 9830 23907 9832
rect 19977 9827 20043 9830
rect 23841 9827 23907 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 11421 9754 11487 9757
rect 14457 9754 14523 9757
rect 11421 9752 14523 9754
rect 11421 9696 11426 9752
rect 11482 9696 14462 9752
rect 14518 9696 14523 9752
rect 11421 9694 14523 9696
rect 11421 9691 11487 9694
rect 14457 9691 14523 9694
rect 18597 9754 18663 9757
rect 20253 9754 20319 9757
rect 24120 9754 24180 9966
rect 24718 9890 24778 9966
rect 24945 10024 28000 10026
rect 24945 9968 24950 10024
rect 25006 9968 28000 10024
rect 24945 9966 28000 9968
rect 24945 9963 25011 9966
rect 27520 9936 28000 9966
rect 25129 9890 25195 9893
rect 24718 9888 25195 9890
rect 24718 9832 25134 9888
rect 25190 9832 25195 9888
rect 24718 9830 25195 9832
rect 25129 9827 25195 9830
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 18597 9752 24180 9754
rect 18597 9696 18602 9752
rect 18658 9696 20258 9752
rect 20314 9696 24180 9752
rect 18597 9694 24180 9696
rect 18597 9691 18663 9694
rect 20253 9691 20319 9694
rect 3969 9618 4035 9621
rect 13629 9618 13695 9621
rect 3969 9616 13695 9618
rect 3969 9560 3974 9616
rect 4030 9560 13634 9616
rect 13690 9560 13695 9616
rect 3969 9558 13695 9560
rect 3969 9555 4035 9558
rect 13629 9555 13695 9558
rect 14273 9618 14339 9621
rect 15653 9618 15719 9621
rect 14273 9616 15719 9618
rect 14273 9560 14278 9616
rect 14334 9560 15658 9616
rect 15714 9560 15719 9616
rect 14273 9558 15719 9560
rect 14273 9555 14339 9558
rect 15653 9555 15719 9558
rect 17861 9618 17927 9621
rect 19517 9618 19583 9621
rect 17861 9616 19583 9618
rect 17861 9560 17866 9616
rect 17922 9560 19522 9616
rect 19578 9560 19583 9616
rect 17861 9558 19583 9560
rect 17861 9555 17927 9558
rect 19517 9555 19583 9558
rect 0 9482 480 9512
rect 3141 9482 3207 9485
rect 0 9480 3207 9482
rect 0 9424 3146 9480
rect 3202 9424 3207 9480
rect 0 9422 3207 9424
rect 0 9392 480 9422
rect 3141 9419 3207 9422
rect 3601 9482 3667 9485
rect 15745 9482 15811 9485
rect 3601 9480 15811 9482
rect 3601 9424 3606 9480
rect 3662 9424 15750 9480
rect 15806 9424 15811 9480
rect 3601 9422 15811 9424
rect 3601 9419 3667 9422
rect 15745 9419 15811 9422
rect 16665 9482 16731 9485
rect 21633 9482 21699 9485
rect 16665 9480 21699 9482
rect 16665 9424 16670 9480
rect 16726 9424 21638 9480
rect 21694 9424 21699 9480
rect 16665 9422 21699 9424
rect 16665 9419 16731 9422
rect 21633 9419 21699 9422
rect 22001 9482 22067 9485
rect 27520 9482 28000 9512
rect 22001 9480 28000 9482
rect 22001 9424 22006 9480
rect 22062 9424 28000 9480
rect 22001 9422 28000 9424
rect 22001 9419 22067 9422
rect 27520 9392 28000 9422
rect 4061 9346 4127 9349
rect 9857 9346 9923 9349
rect 4061 9344 9923 9346
rect 4061 9288 4066 9344
rect 4122 9288 9862 9344
rect 9918 9288 9923 9344
rect 4061 9286 9923 9288
rect 4061 9283 4127 9286
rect 9857 9283 9923 9286
rect 17033 9346 17099 9349
rect 19425 9346 19491 9349
rect 17033 9344 19491 9346
rect 17033 9288 17038 9344
rect 17094 9288 19430 9344
rect 19486 9288 19491 9344
rect 17033 9286 19491 9288
rect 17033 9283 17099 9286
rect 19425 9283 19491 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 6913 9210 6979 9213
rect 12341 9210 12407 9213
rect 24577 9210 24643 9213
rect 24710 9210 24716 9212
rect 6913 9208 8218 9210
rect 6913 9152 6918 9208
rect 6974 9152 8218 9208
rect 6913 9150 8218 9152
rect 6913 9147 6979 9150
rect 2221 9074 2287 9077
rect 8158 9074 8218 9150
rect 12341 9208 17234 9210
rect 12341 9152 12346 9208
rect 12402 9152 17234 9208
rect 12341 9150 17234 9152
rect 12341 9147 12407 9150
rect 17033 9074 17099 9077
rect 2221 9072 7666 9074
rect 2221 9016 2226 9072
rect 2282 9016 7666 9072
rect 2221 9014 7666 9016
rect 8158 9072 17099 9074
rect 8158 9016 17038 9072
rect 17094 9016 17099 9072
rect 8158 9014 17099 9016
rect 17174 9074 17234 9150
rect 22372 9208 24716 9210
rect 22372 9152 24582 9208
rect 24638 9152 24716 9208
rect 22372 9150 24716 9152
rect 22372 9074 22432 9150
rect 24577 9147 24643 9150
rect 24710 9148 24716 9150
rect 24780 9148 24786 9212
rect 17174 9014 22432 9074
rect 22553 9074 22619 9077
rect 25037 9074 25103 9077
rect 22553 9072 25103 9074
rect 22553 9016 22558 9072
rect 22614 9016 25042 9072
rect 25098 9016 25103 9072
rect 22553 9014 25103 9016
rect 2221 9011 2287 9014
rect 0 8938 480 8968
rect 3969 8938 4035 8941
rect 0 8936 4035 8938
rect 0 8880 3974 8936
rect 4030 8880 4035 8936
rect 0 8878 4035 8880
rect 7606 8938 7666 9014
rect 17033 9011 17099 9014
rect 22553 9011 22619 9014
rect 25037 9011 25103 9014
rect 16113 8938 16179 8941
rect 18505 8938 18571 8941
rect 7606 8878 15946 8938
rect 0 8848 480 8878
rect 3969 8875 4035 8878
rect 15886 8802 15946 8878
rect 16113 8936 18571 8938
rect 16113 8880 16118 8936
rect 16174 8880 18510 8936
rect 18566 8880 18571 8936
rect 16113 8878 18571 8880
rect 16113 8875 16179 8878
rect 18505 8875 18571 8878
rect 20529 8938 20595 8941
rect 22001 8938 22067 8941
rect 20529 8936 22067 8938
rect 20529 8880 20534 8936
rect 20590 8880 22006 8936
rect 22062 8880 22067 8936
rect 20529 8878 22067 8880
rect 20529 8875 20595 8878
rect 22001 8875 22067 8878
rect 23657 8938 23723 8941
rect 27520 8938 28000 8968
rect 23657 8936 28000 8938
rect 23657 8880 23662 8936
rect 23718 8880 28000 8936
rect 23657 8878 28000 8880
rect 23657 8875 23723 8878
rect 27520 8848 28000 8878
rect 20897 8802 20963 8805
rect 15886 8800 20963 8802
rect 15886 8744 20902 8800
rect 20958 8744 20963 8800
rect 15886 8742 20963 8744
rect 20897 8739 20963 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 19425 8666 19491 8669
rect 23657 8666 23723 8669
rect 19425 8664 23723 8666
rect 19425 8608 19430 8664
rect 19486 8608 23662 8664
rect 23718 8608 23723 8664
rect 19425 8606 23723 8608
rect 19425 8603 19491 8606
rect 23657 8603 23723 8606
rect 19701 8530 19767 8533
rect 19701 8528 24226 8530
rect 19701 8472 19706 8528
rect 19762 8472 24226 8528
rect 19701 8470 24226 8472
rect 19701 8467 19767 8470
rect 24166 8397 24226 8470
rect 15377 8394 15443 8397
rect 20529 8394 20595 8397
rect 9998 8334 10794 8394
rect 0 8258 480 8288
rect 7557 8258 7623 8261
rect 0 8256 7623 8258
rect 0 8200 7562 8256
rect 7618 8200 7623 8256
rect 0 8198 7623 8200
rect 0 8168 480 8198
rect 7557 8195 7623 8198
rect 8017 8258 8083 8261
rect 9998 8258 10058 8334
rect 8017 8256 10058 8258
rect 8017 8200 8022 8256
rect 8078 8200 10058 8256
rect 8017 8198 10058 8200
rect 10734 8258 10794 8334
rect 15377 8392 20595 8394
rect 15377 8336 15382 8392
rect 15438 8336 20534 8392
rect 20590 8336 20595 8392
rect 15377 8334 20595 8336
rect 15377 8331 15443 8334
rect 20529 8331 20595 8334
rect 20897 8394 20963 8397
rect 22553 8394 22619 8397
rect 24025 8394 24091 8397
rect 20897 8392 22386 8394
rect 20897 8336 20902 8392
rect 20958 8336 22386 8392
rect 20897 8334 22386 8336
rect 20897 8331 20963 8334
rect 15101 8258 15167 8261
rect 16757 8258 16823 8261
rect 10734 8198 15026 8258
rect 8017 8195 8083 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 14966 8122 15026 8198
rect 15101 8256 16823 8258
rect 15101 8200 15106 8256
rect 15162 8200 16762 8256
rect 16818 8200 16823 8256
rect 15101 8198 16823 8200
rect 22326 8258 22386 8334
rect 22553 8392 24091 8394
rect 22553 8336 22558 8392
rect 22614 8336 24030 8392
rect 24086 8336 24091 8392
rect 22553 8334 24091 8336
rect 24166 8392 24275 8397
rect 24166 8336 24214 8392
rect 24270 8336 24275 8392
rect 24166 8334 24275 8336
rect 22553 8331 22619 8334
rect 24025 8331 24091 8334
rect 24209 8331 24275 8334
rect 23473 8258 23539 8261
rect 27520 8258 28000 8288
rect 22326 8256 23539 8258
rect 22326 8200 23478 8256
rect 23534 8200 23539 8256
rect 22326 8198 23539 8200
rect 15101 8195 15167 8198
rect 16757 8195 16823 8198
rect 23473 8195 23539 8198
rect 23614 8198 28000 8258
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 17677 8122 17743 8125
rect 14966 8120 17743 8122
rect 14966 8064 17682 8120
rect 17738 8064 17743 8120
rect 14966 8062 17743 8064
rect 17677 8059 17743 8062
rect 22185 8122 22251 8125
rect 23614 8122 23674 8198
rect 27520 8168 28000 8198
rect 22185 8120 23674 8122
rect 22185 8064 22190 8120
rect 22246 8064 23674 8120
rect 22185 8062 23674 8064
rect 23933 8122 23999 8125
rect 25497 8122 25563 8125
rect 23933 8120 25563 8122
rect 23933 8064 23938 8120
rect 23994 8064 25502 8120
rect 25558 8064 25563 8120
rect 23933 8062 25563 8064
rect 22185 8059 22251 8062
rect 23933 8059 23999 8062
rect 25497 8059 25563 8062
rect 10777 7986 10843 7989
rect 24669 7986 24735 7989
rect 10777 7984 24735 7986
rect 10777 7928 10782 7984
rect 10838 7928 24674 7984
rect 24730 7928 24735 7984
rect 10777 7926 24735 7928
rect 10777 7923 10843 7926
rect 24669 7923 24735 7926
rect 15837 7850 15903 7853
rect 5398 7848 15903 7850
rect 5398 7792 15842 7848
rect 15898 7792 15903 7848
rect 5398 7790 15903 7792
rect 0 7714 480 7744
rect 5398 7714 5458 7790
rect 15837 7787 15903 7790
rect 24301 7850 24367 7853
rect 24301 7848 24732 7850
rect 24301 7792 24306 7848
rect 24362 7792 24732 7848
rect 24301 7790 24732 7792
rect 24301 7787 24367 7790
rect 0 7654 5458 7714
rect 7557 7714 7623 7717
rect 14181 7714 14247 7717
rect 7557 7712 14247 7714
rect 7557 7656 7562 7712
rect 7618 7656 14186 7712
rect 14242 7656 14247 7712
rect 7557 7654 14247 7656
rect 24672 7714 24732 7790
rect 27520 7714 28000 7744
rect 24672 7654 28000 7714
rect 0 7624 480 7654
rect 7557 7651 7623 7654
rect 14181 7651 14247 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 21081 7578 21147 7581
rect 23657 7578 23723 7581
rect 21081 7576 23723 7578
rect 21081 7520 21086 7576
rect 21142 7520 23662 7576
rect 23718 7520 23723 7576
rect 21081 7518 23723 7520
rect 21081 7515 21147 7518
rect 23657 7515 23723 7518
rect 9765 7442 9831 7445
rect 24669 7442 24735 7445
rect 9765 7440 24735 7442
rect 9765 7384 9770 7440
rect 9826 7384 24674 7440
rect 24730 7384 24735 7440
rect 9765 7382 24735 7384
rect 9765 7379 9831 7382
rect 24669 7379 24735 7382
rect 12801 7306 12867 7309
rect 23565 7306 23631 7309
rect 12801 7304 23631 7306
rect 12801 7248 12806 7304
rect 12862 7248 23570 7304
rect 23626 7248 23631 7304
rect 12801 7246 23631 7248
rect 12801 7243 12867 7246
rect 23565 7243 23631 7246
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 14549 7170 14615 7173
rect 19333 7170 19399 7173
rect 14549 7168 19399 7170
rect 14549 7112 14554 7168
rect 14610 7112 19338 7168
rect 19394 7112 19399 7168
rect 14549 7110 19399 7112
rect 14549 7107 14615 7110
rect 19333 7107 19399 7110
rect 24209 7170 24275 7173
rect 27520 7170 28000 7200
rect 24209 7168 28000 7170
rect 24209 7112 24214 7168
rect 24270 7112 28000 7168
rect 24209 7110 28000 7112
rect 24209 7107 24275 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 27520 7080 28000 7110
rect 19610 7039 19930 7040
rect 2957 6898 3023 6901
rect 14089 6898 14155 6901
rect 2957 6896 14155 6898
rect 2957 6840 2962 6896
rect 3018 6840 14094 6896
rect 14150 6840 14155 6896
rect 2957 6838 14155 6840
rect 2957 6835 3023 6838
rect 14089 6835 14155 6838
rect 17401 6898 17467 6901
rect 23289 6898 23355 6901
rect 23749 6900 23815 6901
rect 23749 6898 23796 6900
rect 17401 6896 23355 6898
rect 17401 6840 17406 6896
rect 17462 6840 23294 6896
rect 23350 6840 23355 6896
rect 17401 6838 23355 6840
rect 23704 6896 23796 6898
rect 23704 6840 23754 6896
rect 23704 6838 23796 6840
rect 17401 6835 17467 6838
rect 23289 6835 23355 6838
rect 23749 6836 23796 6838
rect 23860 6836 23866 6900
rect 23749 6835 23815 6836
rect 12709 6762 12775 6765
rect 5398 6760 12775 6762
rect 5398 6704 12714 6760
rect 12770 6704 12775 6760
rect 5398 6702 12775 6704
rect 0 6626 480 6656
rect 5398 6626 5458 6702
rect 12709 6699 12775 6702
rect 14641 6762 14707 6765
rect 16481 6762 16547 6765
rect 14641 6760 16547 6762
rect 14641 6704 14646 6760
rect 14702 6704 16486 6760
rect 16542 6704 16547 6760
rect 14641 6702 16547 6704
rect 14641 6699 14707 6702
rect 16481 6699 16547 6702
rect 20069 6762 20135 6765
rect 23933 6762 23999 6765
rect 20069 6760 23999 6762
rect 20069 6704 20074 6760
rect 20130 6704 23938 6760
rect 23994 6704 23999 6760
rect 20069 6702 23999 6704
rect 20069 6699 20135 6702
rect 23933 6699 23999 6702
rect 27520 6626 28000 6656
rect 0 6566 5458 6626
rect 24902 6566 28000 6626
rect 0 6536 480 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 18781 6354 18847 6357
rect 24902 6354 24962 6566
rect 27520 6536 28000 6566
rect 18781 6352 24962 6354
rect 18781 6296 18786 6352
rect 18842 6296 24962 6352
rect 18781 6294 24962 6296
rect 18781 6291 18847 6294
rect 0 6082 480 6112
rect 2957 6082 3023 6085
rect 0 6080 3023 6082
rect 0 6024 2962 6080
rect 3018 6024 3023 6080
rect 0 6022 3023 6024
rect 0 5992 480 6022
rect 2957 6019 3023 6022
rect 22369 6082 22435 6085
rect 27520 6082 28000 6112
rect 22369 6080 28000 6082
rect 22369 6024 22374 6080
rect 22430 6024 28000 6080
rect 22369 6022 28000 6024
rect 22369 6019 22435 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 14365 5946 14431 5949
rect 16389 5946 16455 5949
rect 14365 5944 16455 5946
rect 14365 5888 14370 5944
rect 14426 5888 16394 5944
rect 16450 5888 16455 5944
rect 14365 5886 16455 5888
rect 14365 5883 14431 5886
rect 16389 5883 16455 5886
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 4061 5402 4127 5405
rect 27520 5402 28000 5432
rect 0 5400 4127 5402
rect 0 5344 4066 5400
rect 4122 5344 4127 5400
rect 0 5342 4127 5344
rect 0 5312 480 5342
rect 4061 5339 4127 5342
rect 24902 5342 28000 5402
rect 16849 5266 16915 5269
rect 24761 5266 24827 5269
rect 16849 5264 24827 5266
rect 16849 5208 16854 5264
rect 16910 5208 24766 5264
rect 24822 5208 24827 5264
rect 16849 5206 24827 5208
rect 16849 5203 16915 5206
rect 24761 5203 24827 5206
rect 18137 5130 18203 5133
rect 23473 5130 23539 5133
rect 24902 5130 24962 5342
rect 27520 5312 28000 5342
rect 18137 5128 22064 5130
rect 18137 5072 18142 5128
rect 18198 5072 22064 5128
rect 18137 5070 22064 5072
rect 18137 5067 18203 5070
rect 22004 4994 22064 5070
rect 23473 5128 24962 5130
rect 23473 5072 23478 5128
rect 23534 5072 24962 5128
rect 23473 5070 24962 5072
rect 23473 5067 23539 5070
rect 22004 4934 22248 4994
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3877 4858 3943 4861
rect 0 4856 3943 4858
rect 0 4800 3882 4856
rect 3938 4800 3943 4856
rect 0 4798 3943 4800
rect 22188 4858 22248 4934
rect 27520 4858 28000 4888
rect 22188 4798 28000 4858
rect 0 4768 480 4798
rect 3877 4795 3943 4798
rect 27520 4768 28000 4798
rect 20161 4722 20227 4725
rect 3926 4720 20227 4722
rect 3926 4664 20166 4720
rect 20222 4664 20227 4720
rect 3926 4662 20227 4664
rect 0 4314 480 4344
rect 3926 4314 3986 4662
rect 20161 4659 20227 4662
rect 4061 4586 4127 4589
rect 22461 4586 22527 4589
rect 4061 4584 22527 4586
rect 4061 4528 4066 4584
rect 4122 4528 22466 4584
rect 22522 4528 22527 4584
rect 4061 4526 22527 4528
rect 4061 4523 4127 4526
rect 22461 4523 22527 4526
rect 24117 4586 24183 4589
rect 24117 4584 24732 4586
rect 24117 4528 24122 4584
rect 24178 4528 24732 4584
rect 24117 4526 24732 4528
rect 24117 4523 24183 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 0 4254 3986 4314
rect 24672 4314 24732 4526
rect 27520 4314 28000 4344
rect 24672 4254 28000 4314
rect 0 4224 480 4254
rect 27520 4224 28000 4254
rect 19977 4178 20043 4181
rect 23473 4178 23539 4181
rect 19977 4176 23539 4178
rect 19977 4120 19982 4176
rect 20038 4120 23478 4176
rect 23534 4120 23539 4176
rect 19977 4118 23539 4120
rect 19977 4115 20043 4118
rect 23473 4115 23539 4118
rect 3969 4042 4035 4045
rect 17493 4042 17559 4045
rect 3969 4040 17559 4042
rect 3969 3984 3974 4040
rect 4030 3984 17498 4040
rect 17554 3984 17559 4040
rect 3969 3982 17559 3984
rect 3969 3979 4035 3982
rect 17493 3979 17559 3982
rect 18505 4042 18571 4045
rect 18505 4040 22064 4042
rect 18505 3984 18510 4040
rect 18566 3984 22064 4040
rect 18505 3982 22064 3984
rect 18505 3979 18571 3982
rect 22004 3906 22064 3982
rect 22004 3846 22248 3906
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 4061 3770 4127 3773
rect 0 3768 4127 3770
rect 0 3712 4066 3768
rect 4122 3712 4127 3768
rect 0 3710 4127 3712
rect 22188 3770 22248 3846
rect 27520 3770 28000 3800
rect 22188 3710 28000 3770
rect 0 3680 480 3710
rect 4061 3707 4127 3710
rect 27520 3680 28000 3710
rect 3325 3634 3391 3637
rect 11881 3634 11947 3637
rect 3325 3632 11947 3634
rect 3325 3576 3330 3632
rect 3386 3576 11886 3632
rect 11942 3576 11947 3632
rect 3325 3574 11947 3576
rect 3325 3571 3391 3574
rect 11881 3571 11947 3574
rect 17493 3634 17559 3637
rect 23657 3634 23723 3637
rect 17493 3632 23723 3634
rect 17493 3576 17498 3632
rect 17554 3576 23662 3632
rect 23718 3576 23723 3632
rect 17493 3574 23723 3576
rect 17493 3571 17559 3574
rect 23657 3571 23723 3574
rect 11973 3498 12039 3501
rect 23197 3498 23263 3501
rect 11973 3496 23263 3498
rect 11973 3440 11978 3496
rect 12034 3440 23202 3496
rect 23258 3440 23263 3496
rect 11973 3438 23263 3440
rect 11973 3435 12039 3438
rect 23197 3435 23263 3438
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 3969 3226 4035 3229
rect 0 3224 4035 3226
rect 0 3168 3974 3224
rect 4030 3168 4035 3224
rect 0 3166 4035 3168
rect 0 3136 480 3166
rect 3969 3163 4035 3166
rect 24761 3226 24827 3229
rect 27520 3226 28000 3256
rect 24761 3224 28000 3226
rect 24761 3168 24766 3224
rect 24822 3168 28000 3224
rect 24761 3166 28000 3168
rect 24761 3163 24827 3166
rect 27520 3136 28000 3166
rect 4061 3090 4127 3093
rect 17401 3090 17467 3093
rect 4061 3088 17467 3090
rect 4061 3032 4066 3088
rect 4122 3032 17406 3088
rect 17462 3032 17467 3088
rect 4061 3030 17467 3032
rect 4061 3027 4127 3030
rect 17401 3027 17467 3030
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 3509 2682 3575 2685
rect 3190 2680 3575 2682
rect 3190 2624 3514 2680
rect 3570 2624 3575 2680
rect 3190 2622 3575 2624
rect 0 2546 480 2576
rect 3190 2546 3250 2622
rect 3509 2619 3575 2622
rect 11697 2546 11763 2549
rect 0 2486 3250 2546
rect 3374 2544 11763 2546
rect 3374 2488 11702 2544
rect 11758 2488 11763 2544
rect 3374 2486 11763 2488
rect 0 2456 480 2486
rect 0 2002 480 2032
rect 3374 2002 3434 2486
rect 11697 2483 11763 2486
rect 21633 2546 21699 2549
rect 27520 2546 28000 2576
rect 21633 2544 28000 2546
rect 21633 2488 21638 2544
rect 21694 2488 28000 2544
rect 21633 2486 28000 2488
rect 21633 2483 21699 2486
rect 27520 2456 28000 2486
rect 4613 2410 4679 2413
rect 11973 2410 12039 2413
rect 4613 2408 12039 2410
rect 4613 2352 4618 2408
rect 4674 2352 11978 2408
rect 12034 2352 12039 2408
rect 4613 2350 12039 2352
rect 4613 2347 4679 2350
rect 11973 2347 12039 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 0 1942 3434 2002
rect 23565 2002 23631 2005
rect 27520 2002 28000 2032
rect 23565 2000 28000 2002
rect 23565 1944 23570 2000
rect 23626 1944 28000 2000
rect 23565 1942 28000 1944
rect 0 1912 480 1942
rect 23565 1939 23631 1942
rect 27520 1912 28000 1942
rect 17493 1730 17559 1733
rect 3374 1728 17559 1730
rect 3374 1672 17498 1728
rect 17554 1672 17559 1728
rect 3374 1670 17559 1672
rect 0 1458 480 1488
rect 3374 1458 3434 1670
rect 17493 1667 17559 1670
rect 3509 1594 3575 1597
rect 11789 1594 11855 1597
rect 3509 1592 11855 1594
rect 3509 1536 3514 1592
rect 3570 1536 11794 1592
rect 11850 1536 11855 1592
rect 3509 1534 11855 1536
rect 3509 1531 3575 1534
rect 11789 1531 11855 1534
rect 16481 1594 16547 1597
rect 16481 1592 27538 1594
rect 16481 1536 16486 1592
rect 16542 1536 27538 1592
rect 16481 1534 27538 1536
rect 16481 1531 16547 1534
rect 0 1398 3434 1458
rect 27478 1488 27538 1534
rect 27478 1398 28000 1488
rect 0 1368 480 1398
rect 27520 1368 28000 1398
rect 0 914 480 944
rect 3325 914 3391 917
rect 0 912 3391 914
rect 0 856 3330 912
rect 3386 856 3391 912
rect 0 854 3391 856
rect 0 824 480 854
rect 3325 851 3391 854
rect 23473 914 23539 917
rect 27520 914 28000 944
rect 23473 912 28000 914
rect 23473 856 23478 912
rect 23534 856 28000 912
rect 23473 854 28000 856
rect 23473 851 23539 854
rect 27520 824 28000 854
rect 0 370 480 400
rect 3141 370 3207 373
rect 0 368 3207 370
rect 0 312 3146 368
rect 3202 312 3207 368
rect 0 310 3207 312
rect 0 280 480 310
rect 3141 307 3207 310
rect 23841 370 23907 373
rect 27520 370 28000 400
rect 23841 368 28000 370
rect 23841 312 23846 368
rect 23902 312 28000 368
rect 23841 310 28000 312
rect 23841 307 23907 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 9628 25332 9692 25396
rect 23796 25196 23860 25260
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 19380 20300 19444 20364
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 9628 20088 9692 20092
rect 9628 20032 9678 20088
rect 9678 20032 9692 20088
rect 9628 20028 9692 20032
rect 19380 19756 19444 19820
rect 9996 19620 10060 19684
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 14228 17308 14292 17372
rect 7972 17036 8036 17100
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 9996 15676 10060 15740
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 23428 14724 23492 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 9628 14316 9692 14380
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 9628 14044 9692 14108
rect 14228 13908 14292 13972
rect 8156 13636 8220 13700
rect 24716 13696 24780 13700
rect 24716 13640 24730 13696
rect 24730 13640 24780 13696
rect 24716 13636 24780 13640
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 14228 11868 14292 11932
rect 23428 11596 23492 11660
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 24716 9148 24780 9212
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 23796 6896 23860 6900
rect 23796 6840 23810 6896
rect 23810 6840 23860 6896
rect 23796 6836 23860 6840
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 9627 25396 9693 25397
rect 9627 25332 9628 25396
rect 9692 25332 9693 25396
rect 9627 25331 9693 25332
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 9630 20093 9690 25331
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9627 20092 9693 20093
rect 9627 20028 9628 20092
rect 9692 20028 9693 20092
rect 9627 20027 9693 20028
rect 9995 19684 10061 19685
rect 9995 19620 9996 19684
rect 10060 19620 10061 19684
rect 9995 19619 10061 19620
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 7971 17100 8037 17101
rect 7971 17036 7972 17100
rect 8036 17036 8037 17100
rect 7971 17035 8037 17036
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 7974 13290 8034 17035
rect 9998 15741 10058 19619
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 23795 25260 23861 25261
rect 23795 25196 23796 25260
rect 23860 25196 23861 25260
rect 23795 25195 23861 25196
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19379 20364 19445 20365
rect 19379 20300 19380 20364
rect 19444 20300 19445 20364
rect 19379 20299 19445 20300
rect 19382 19821 19442 20299
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19379 19820 19445 19821
rect 19379 19756 19380 19820
rect 19444 19756 19445 19820
rect 19379 19755 19445 19756
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14227 17372 14293 17373
rect 14227 17308 14228 17372
rect 14292 17308 14293 17372
rect 14227 17307 14293 17308
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 9995 15740 10061 15741
rect 9995 15676 9996 15740
rect 10060 15676 10061 15740
rect 9995 15675 10061 15676
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 9627 14380 9693 14381
rect 9627 14316 9628 14380
rect 9692 14316 9693 14380
rect 9627 14315 9693 14316
rect 9630 14109 9690 14315
rect 9627 14108 9693 14109
rect 9627 14044 9628 14108
rect 9692 14044 9693 14108
rect 9627 14043 9693 14044
rect 8155 13700 8221 13701
rect 8155 13636 8156 13700
rect 8220 13636 8221 13700
rect 8155 13635 8221 13636
rect 8158 13290 8218 13635
rect 7974 13230 8218 13290
rect 10277 13632 10597 14656
rect 14230 13973 14290 17307
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14227 13972 14293 13973
rect 14227 13908 14228 13972
rect 14292 13908 14293 13972
rect 14227 13907 14293 13908
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 14230 11933 14290 13907
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14227 11932 14293 11933
rect 14227 11868 14228 11932
rect 14292 11868 14293 11932
rect 14227 11867 14293 11868
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 23427 14788 23493 14789
rect 23427 14724 23428 14788
rect 23492 14724 23493 14788
rect 23427 14723 23493 14724
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 23430 11661 23490 14723
rect 23427 11660 23493 11661
rect 23427 11596 23428 11660
rect 23492 11596 23493 11660
rect 23427 11595 23493 11596
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 23798 6901 23858 25195
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24715 13700 24781 13701
rect 24715 13636 24716 13700
rect 24780 13636 24781 13700
rect 24715 13635 24781 13636
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24718 9213 24778 13635
rect 24715 9212 24781 9213
rect 24715 9148 24716 9212
rect 24780 9148 24781 9212
rect 24715 9147 24781 9148
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 23795 6900 23861 6901
rect 23795 6836 23796 6900
rect 23860 6836 23861 6900
rect 23795 6835 23861 6836
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604666999
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604666999
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604666999
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604666999
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604666999
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604666999
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604666999
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604666999
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604666999
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604666999
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604666999
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604666999
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1604666999
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604666999
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604666999
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604666999
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604666999
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604666999
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604666999
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604666999
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604666999
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604666999
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604666999
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604666999
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604666999
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604666999
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604666999
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604666999
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604666999
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604666999
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604666999
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604666999
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604666999
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604666999
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604666999
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604666999
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604666999
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604666999
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604666999
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604666999
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604666999
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604666999
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604666999
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604666999
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604666999
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604666999
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604666999
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604666999
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604666999
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604666999
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604666999
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604666999
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604666999
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604666999
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604666999
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604666999
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604666999
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604666999
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604666999
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604666999
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604666999
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604666999
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604666999
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604666999
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604666999
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604666999
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604666999
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604666999
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604666999
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604666999
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604666999
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604666999
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604666999
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604666999
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604666999
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604666999
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604666999
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604666999
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604666999
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604666999
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604666999
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604666999
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604666999
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604666999
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_163
timestamp 1604666999
transform 1 0 16100 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_159
timestamp 1604666999
transform 1 0 15732 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_168
timestamp 1604666999
transform 1 0 16560 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604666999
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_172
timestamp 1604666999
transform 1 0 16928 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_175
timestamp 1604666999
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_187
timestamp 1604666999
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604666999
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604666999
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_199
timestamp 1604666999
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1604666999
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604666999
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604666999
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604666999
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604666999
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604666999
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1604666999
transform 1 0 24012 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604666999
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1604666999
transform 1 0 25116 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_273
timestamp 1604666999
transform 1 0 26220 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604666999
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604666999
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604666999
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604666999
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604666999
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604666999
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1604666999
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604666999
transform 1 0 17020 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_164
timestamp 1604666999
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_168
timestamp 1604666999
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_172
timestamp 1604666999
transform 1 0 16928 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1604666999
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_186
timestamp 1604666999
transform 1 0 18216 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_196
timestamp 1604666999
transform 1 0 19136 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_200
timestamp 1604666999
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1604666999
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1604666999
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604666999
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604666999
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _033_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 24748 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 23736 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_239
timestamp 1604666999
transform 1 0 23092 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_245
timestamp 1604666999
transform 1 0 23644 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_249
timestamp 1604666999
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_260
timestamp 1604666999
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1604666999
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604666999
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604666999
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604666999
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604666999
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604666999
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604666999
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_110
timestamp 1604666999
transform 1 0 11224 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1604666999
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1604666999
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_127
timestamp 1604666999
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_133
timestamp 1604666999
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_136
timestamp 1604666999
transform 1 0 13616 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604666999
transform 1 0 15088 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_148
timestamp 1604666999
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_155
timestamp 1604666999
transform 1 0 15364 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_159
timestamp 1604666999
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1604666999
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604666999
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604666999
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1604666999
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1604666999
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604666999
transform 1 0 21160 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_210
timestamp 1604666999
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_214
timestamp 1604666999
transform 1 0 20792 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604666999
transform 1 0 22540 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_221
timestamp 1604666999
transform 1 0 21436 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604666999
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 24656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 24104 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_240
timestamp 1604666999
transform 1 0 23184 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_248
timestamp 1604666999
transform 1 0 23920 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_252
timestamp 1604666999
transform 1 0 24288 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_259
timestamp 1604666999
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_263
timestamp 1604666999
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_267
timestamp 1604666999
transform 1 0 25668 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_275
timestamp 1604666999
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604666999
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604666999
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604666999
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604666999
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 13432 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1604666999
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1604666999
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1604666999
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1604666999
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_147
timestamp 1604666999
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16468 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_159
timestamp 1604666999
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 1604666999
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18952 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_186
timestamp 1604666999
transform 1 0 18216 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1604666999
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_207
timestamp 1604666999
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_211
timestamp 1604666999
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604666999
transform 1 0 21528 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22632 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 21988 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_221
timestamp 1604666999
transform 1 0 21436 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_225
timestamp 1604666999
transform 1 0 21804 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_229
timestamp 1604666999
transform 1 0 22172 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_233
timestamp 1604666999
transform 1 0 22540 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_237
timestamp 1604666999
transform 1 0 22908 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23644 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 24656 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_248
timestamp 1604666999
transform 1 0 23920 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_259
timestamp 1604666999
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1604666999
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604666999
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604666999
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604666999
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604666999
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604666999
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604666999
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_98
timestamp 1604666999
transform 1 0 10120 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_106
timestamp 1604666999
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_111
timestamp 1604666999
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1604666999
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1604666999
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12880 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_137
timestamp 1604666999
transform 1 0 13708 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_141
timestamp 1604666999
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_154
timestamp 1604666999
transform 1 0 15272 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1604666999
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_163
timestamp 1604666999
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604666999
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_187
timestamp 1604666999
transform 1 0 18308 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604666999
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1604666999
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_191
timestamp 1604666999
transform 1 0 18676 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1604666999
transform 1 0 19320 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_207
timestamp 1604666999
transform 1 0 20148 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1604666999
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1604666999
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21252 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_228
timestamp 1604666999
transform 1 0 22080 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_234
timestamp 1604666999
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_238
timestamp 1604666999
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604666999
transform 1 0 24012 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604666999
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1604666999
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_252
timestamp 1604666999
transform 1 0 24288 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_257
timestamp 1604666999
transform 1 0 24748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25024 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_263
timestamp 1604666999
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_267
timestamp 1604666999
transform 1 0 25668 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_275
timestamp 1604666999
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604666999
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604666999
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604666999
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604666999
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604666999
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1604666999
transform 1 0 10212 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 11868 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13432 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_126
timestamp 1604666999
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_130
timestamp 1604666999
transform 1 0 13064 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15548 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1604666999
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_147
timestamp 1604666999
transform 1 0 14628 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 17112 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1604666999
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp 1604666999
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_193
timestamp 1604666999
transform 1 0 18860 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1604666999
transform 1 0 19228 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19780 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_200
timestamp 1604666999
transform 1 0 19504 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_206
timestamp 1604666999
transform 1 0 20056 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 22448 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1604666999
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1604666999
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_241
timestamp 1604666999
transform 1 0 23276 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1604666999
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_259
timestamp 1604666999
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1604666999
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604666999
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604666999
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604666999
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604666999
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604666999
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604666999
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604666999
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_86
timestamp 1604666999
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1604666999
transform 1 0 8464 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_99
timestamp 1604666999
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1604666999
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1604666999
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10028 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_106
timestamp 1604666999
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 10580 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1604666999
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1604666999
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604666999
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604666999
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1604666999
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_127
timestamp 1604666999
transform 1 0 12788 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604666999
transform 1 0 12512 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 1604666999
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12144 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13708 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_14_147
timestamp 1604666999
transform 1 0 14628 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_139
timestamp 1604666999
transform 1 0 13892 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604666999
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1604666999
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_158
timestamp 1604666999
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16008 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604666999
transform 1 0 16192 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1604666999
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_173
timestamp 1604666999
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1604666999
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_185
timestamp 1604666999
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1604666999
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_184
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_189
timestamp 1604666999
transform 1 0 18492 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18308 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_205
timestamp 1604666999
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_201
timestamp 1604666999
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1604666999
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_210
timestamp 1604666999
transform 1 0 20424 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_206
timestamp 1604666999
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1604666999
transform 1 0 21160 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604666999
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_216
timestamp 1604666999
transform 1 0 20976 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_225
timestamp 1604666999
transform 1 0 21804 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1604666999
transform 1 0 21528 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_219
timestamp 1604666999
transform 1 0 21252 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21620 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_236
timestamp 1604666999
transform 1 0 22816 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_232
timestamp 1604666999
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21896 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_245
timestamp 1604666999
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1604666999
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_249
timestamp 1604666999
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604666999
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604666999
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604666999
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_259
timestamp 1604666999
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1604666999
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604666999
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_275
timestamp 1604666999
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604666999
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_263
timestamp 1604666999
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604666999
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604666999
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604666999
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604666999
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_70
timestamp 1604666999
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_73
timestamp 1604666999
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_77
timestamp 1604666999
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1604666999
transform 1 0 8556 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_85
timestamp 1604666999
transform 1 0 8924 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_97
timestamp 1604666999
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_34.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_101
timestamp 1604666999
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604666999
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604666999
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1604666999
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1604666999
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1604666999
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1604666999
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1604666999
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_174
timestamp 1604666999
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18216 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604666999
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1604666999
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 21068 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19872 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_199
timestamp 1604666999
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_203
timestamp 1604666999
transform 1 0 19780 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_207
timestamp 1604666999
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_213
timestamp 1604666999
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604666999
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604666999
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_254
timestamp 1604666999
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604666999
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604666999
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_258
timestamp 1604666999
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1604666999
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_270
timestamp 1604666999
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604666999
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604666999
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_44
timestamp 1604666999
transform 1 0 5152 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_48
timestamp 1604666999
transform 1 0 5520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1604666999
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_55
timestamp 1604666999
transform 1 0 6164 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604666999
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_63
timestamp 1604666999
transform 1 0 6900 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_68
timestamp 1604666999
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1604666999
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_84
timestamp 1604666999
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604666999
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_96
timestamp 1604666999
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_36.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1604666999
transform 1 0 10304 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_104
timestamp 1604666999
transform 1 0 10672 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_116
timestamp 1604666999
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 12512 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1604666999
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1604666999
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_137
timestamp 1604666999
transform 1 0 13708 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604666999
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1604666999
transform 1 0 14076 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_145
timestamp 1604666999
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_173
timestamp 1604666999
transform 1 0 17020 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_178
timestamp 1604666999
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 18308 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_182
timestamp 1604666999
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 1604666999
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604666999
transform 1 0 21068 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604666999
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1604666999
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 22080 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604666999
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_220
timestamp 1604666999
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1604666999
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_1_
timestamp 1604666999
transform 1 0 24564 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_247
timestamp 1604666999
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_251
timestamp 1604666999
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_264
timestamp 1604666999
transform 1 0 25392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_268
timestamp 1604666999
transform 1 0 25760 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604666999
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604666999
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_6
timestamp 1604666999
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_10
timestamp 1604666999
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_14
timestamp 1604666999
transform 1 0 2392 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_19
timestamp 1604666999
transform 1 0 2852 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_31
timestamp 1604666999
transform 1 0 3956 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1604666999
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1604666999
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_47
timestamp 1604666999
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1604666999
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_55
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604666999
transform 1 0 7636 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_67
timestamp 1604666999
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_34.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1604666999
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1604666999
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1604666999
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_36.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604666999
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604666999
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604666999
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13248 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_128
timestamp 1604666999
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_151
timestamp 1604666999
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_156
timestamp 1604666999
transform 1 0 15456 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15732 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_168
timestamp 1604666999
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_172
timestamp 1604666999
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_176
timestamp 1604666999
transform 1 0 17296 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1604666999
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1604666999
transform 1 0 19228 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19872 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_201
timestamp 1604666999
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604666999
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604666999
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_223
timestamp 1604666999
transform 1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1604666999
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604666999
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604666999
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_254
timestamp 1604666999
transform 1 0 24472 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604666999
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604666999
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_260
timestamp 1604666999
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_266
timestamp 1604666999
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_270
timestamp 1604666999
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_274
timestamp 1604666999
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604666999
transform 1 0 1564 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604666999
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604666999
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_9
timestamp 1604666999
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_13
timestamp 1604666999
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1604666999
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1604666999
transform 1 0 3312 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1604666999
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_38
timestamp 1604666999
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_42
timestamp 1604666999
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_46
timestamp 1604666999
transform 1 0 5336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_58
timestamp 1604666999
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1604666999
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1604666999
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1604666999
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_30.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_83
timestamp 1604666999
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1604666999
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604666999
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11500 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_102
timestamp 1604666999
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1604666999
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1604666999
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_132
timestamp 1604666999
transform 1 0 13248 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1604666999
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604666999
transform 1 0 14168 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1604666999
transform 1 0 14076 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_145
timestamp 1604666999
transform 1 0 14444 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_173
timestamp 1604666999
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_177
timestamp 1604666999
transform 1 0 17388 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18308 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 1604666999
transform 1 0 17940 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_186
timestamp 1604666999
transform 1 0 18216 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1604666999
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1604666999
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604666999
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 22356 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_223
timestamp 1604666999
transform 1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_228
timestamp 1604666999
transform 1 0 22080 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1604666999
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_254
timestamp 1604666999
transform 1 0 24472 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604666999
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1604666999
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1604666999
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1604666999
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604666999
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1604666999
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1604666999
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604666999
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp 1604666999
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1604666999
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604666999
transform 1 0 2484 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604666999
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1604666999
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1604666999
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1604666999
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604666999
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 3588 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604666999
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_30
timestamp 1604666999
transform 1 0 3864 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1604666999
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1604666999
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1604666999
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604666999
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604666999
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604666999
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1604666999
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_62
timestamp 1604666999
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_70
timestamp 1604666999
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1604666999
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_71
timestamp 1604666999
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_88
timestamp 1604666999
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_84
timestamp 1604666999
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_85
timestamp 1604666999
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604666999
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9292 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1604666999
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1604666999
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9936 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604666999
transform 1 0 10948 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp 1604666999
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_106
timestamp 1604666999
transform 1 0 10856 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_110
timestamp 1604666999
transform 1 0 11224 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_115
timestamp 1604666999
transform 1 0 11684 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_119
timestamp 1604666999
transform 1 0 12052 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_122
timestamp 1604666999
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1604666999
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604666999
transform 1 0 12512 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1604666999
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_34.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_20_146
timestamp 1604666999
transform 1 0 14536 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_142
timestamp 1604666999
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1604666999
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1604666999
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1604666999
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1604666999
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15088 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_166
timestamp 1604666999
transform 1 0 16376 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1604666999
transform 1 0 16008 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_168
timestamp 1604666999
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_165
timestamp 1604666999
transform 1 0 16284 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_161
timestamp 1604666999
transform 1 0 15916 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604666999
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604666999
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16928 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16744 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604666999
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1604666999
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1604666999
transform 1 0 18492 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1604666999
transform 1 0 18860 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18676 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1604666999
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1604666999
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1604666999
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604666999
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_218
timestamp 1604666999
transform 1 0 21160 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_214
timestamp 1604666999
transform 1 0 20792 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1604666999
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21252 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21896 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21712 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 1604666999
transform 1 0 21436 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_235
timestamp 1604666999
transform 1 0 22724 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_238
timestamp 1604666999
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_242
timestamp 1604666999
transform 1 0 23368 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604666999
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23184 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 23552 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 23736 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_255
timestamp 1604666999
transform 1 0 24564 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_254
timestamp 1604666999
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_266
timestamp 1604666999
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1604666999
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604666999
transform 1 0 25208 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604666999
transform 1 0 25300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1604666999
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_274
timestamp 1604666999
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_270
timestamp 1604666999
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604666999
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604666999
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604666999
transform 1 0 2484 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1604666999
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1604666999
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1604666999
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604666999
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1604666999
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1604666999
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604666999
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604666999
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1604666999
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_30.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_65
timestamp 1604666999
transform 1 0 7084 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604666999
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9568 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1604666999
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1604666999
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_111
timestamp 1604666999
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1604666999
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1604666999
transform 1 0 12052 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13432 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_126
timestamp 1604666999
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_130
timestamp 1604666999
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_153
timestamp 1604666999
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1604666999
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15916 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_170
timestamp 1604666999
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_174
timestamp 1604666999
transform 1 0 17112 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18584 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_180
timestamp 1604666999
transform 1 0 17664 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1604666999
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1604666999
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604666999
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1604666999
transform 1 0 21436 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_230
timestamp 1604666999
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_234
timestamp 1604666999
transform 1 0 22632 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604666999
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_254
timestamp 1604666999
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604666999
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604666999
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_258
timestamp 1604666999
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_266
timestamp 1604666999
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_270
timestamp 1604666999
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_274
timestamp 1604666999
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1604666999
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1604666999
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604666999
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604666999
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1604666999
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 6348 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604666999
transform 1 0 4784 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_49
timestamp 1604666999
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_53
timestamp 1604666999
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1604666999
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1604666999
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604666999
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1604666999
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1604666999
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12144 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_123
timestamp 1604666999
transform 1 0 12420 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1604666999
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1604666999
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1604666999
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_158
timestamp 1604666999
transform 1 0 15640 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16192 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_163
timestamp 1604666999
transform 1 0 16100 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18676 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1604666999
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_187
timestamp 1604666999
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_200
timestamp 1604666999
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_204
timestamp 1604666999
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1604666999
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1604666999
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22908 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_234
timestamp 1604666999
transform 1 0 22632 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 23828 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 23276 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_239
timestamp 1604666999
transform 1 0 23092 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_243
timestamp 1604666999
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_256
timestamp 1604666999
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25392 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_260
timestamp 1604666999
transform 1 0 25024 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267
timestamp 1604666999
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2668 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_7
timestamp 1604666999
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_12
timestamp 1604666999
transform 1 0 2208 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_26
timestamp 1604666999
transform 1 0 3496 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_30
timestamp 1604666999
transform 1 0 3864 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1604666999
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_37
timestamp 1604666999
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_41
timestamp 1604666999
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604666999
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604666999
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 7728 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_66
timestamp 1604666999
transform 1 0 7176 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1604666999
transform 1 0 9476 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1604666999
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_28.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604666999
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604666999
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604666999
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1604666999
transform 1 0 12696 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1604666999
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14628 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_141
timestamp 1604666999
transform 1 0 14076 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1604666999
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_170
timestamp 1604666999
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_174
timestamp 1604666999
transform 1 0 17112 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604666999
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1604666999
transform 1 0 18860 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19596 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_199
timestamp 1604666999
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604666999
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604666999
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_220
timestamp 1604666999
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_224
timestamp 1604666999
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_228
timestamp 1604666999
transform 1 0 22080 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604666999
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 23828 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604666999
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_256
timestamp 1604666999
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604666999
transform 1 0 25392 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604666999
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_260
timestamp 1604666999
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1604666999
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_272
timestamp 1604666999
transform 1 0 26128 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604666999
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2024 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604666999
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_7
timestamp 1604666999
transform 1 0 1748 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1604666999
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604666999
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5888 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_44
timestamp 1604666999
transform 1 0 5152 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_49
timestamp 1604666999
transform 1 0 5612 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_71
timestamp 1604666999
transform 1 0 7636 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_76
timestamp 1604666999
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9844 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_80
timestamp 1604666999
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604666999
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604666999
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11408 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_104
timestamp 1604666999
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_108
timestamp 1604666999
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_131
timestamp 1604666999
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1604666999
transform 1 0 13524 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 13892 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 15456 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_142
timestamp 1604666999
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1604666999
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1604666999
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16468 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_159
timestamp 1604666999
transform 1 0 15732 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604666999
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1604666999
transform 1 0 18216 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_190
timestamp 1604666999
transform 1 0 18584 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1604666999
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604666999
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604666999
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 21528 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_24_219
timestamp 1604666999
transform 1 0 21252 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 24012 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23460 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_241
timestamp 1604666999
transform 1 0 23276 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_245
timestamp 1604666999
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1604666999
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1604666999
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604666999
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2576 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604666999
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1604666999
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp 1604666999
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_35
timestamp 1604666999
transform 1 0 4324 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1604666999
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604666999
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604666999
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9844 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1604666999
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1604666999
transform 1 0 8924 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1604666999
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604666999
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604666999
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_28.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604666999
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1604666999
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_149
timestamp 1604666999
transform 1 0 14812 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_155
timestamp 1604666999
transform 1 0 15364 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_158
timestamp 1604666999
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1604666999
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1604666999
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604666999
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604666999
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1604666999
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_197
timestamp 1604666999
transform 1 0 19228 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604666999
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_201
timestamp 1604666999
transform 1 0 19596 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_213
timestamp 1604666999
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1604666999
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604666999
transform 1 0 21436 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1604666999
transform 1 0 22264 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604666999
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604666999
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_264
timestamp 1604666999
transform 1 0 25392 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604666999
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1604666999
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_6
timestamp 1604666999
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_10
timestamp 1604666999
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 2024 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604666999
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1604666999
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1604666999
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1604666999
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_36
timestamp 1604666999
transform 1 0 4416 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1604666999
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_40
timestamp 1604666999
transform 1 0 4784 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_58
timestamp 1604666999
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_54
timestamp 1604666999
transform 1 0 6072 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1604666999
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5428 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_66
timestamp 1604666999
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1604666999
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604666999
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_74
timestamp 1604666999
transform 1 0 7912 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_70
timestamp 1604666999
transform 1 0 7544 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1604666999
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 7728 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7912 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8004 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1604666999
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_83
timestamp 1604666999
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_98
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_94
timestamp 1604666999
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9844 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_102
timestamp 1604666999
transform 1 0 10488 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_108
timestamp 1604666999
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_104
timestamp 1604666999
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604666999
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604666999
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_28.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11408 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_126
timestamp 1604666999
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_134
timestamp 1604666999
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_130
timestamp 1604666999
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_131
timestamp 1604666999
transform 1 0 13156 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13708 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_142
timestamp 1604666999
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604666999
transform 1 0 13892 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1604666999
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_150
timestamp 1604666999
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_156
timestamp 1604666999
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1604666999
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_164
timestamp 1604666999
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_160
timestamp 1604666999
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_161
timestamp 1604666999
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1604666999
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16284 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604666999
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1604666999
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_184
timestamp 1604666999
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18768 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18584 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_26_205
timestamp 1604666999
transform 1 0 19964 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_201
timestamp 1604666999
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 1604666999
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1604666999
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604666999
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21068 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 23000 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604666999
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1604666999
transform 1 0 22080 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_234
timestamp 1604666999
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1604666999
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_257
timestamp 1604666999
transform 1 0 24748 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604666999
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604666999
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_269
timestamp 1604666999
transform 1 0 25852 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1604666999
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_268
timestamp 1604666999
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604666999
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1472 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604666999
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_36
timestamp 1604666999
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 4784 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1604666999
transform 1 0 6532 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604666999
transform 1 0 7268 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1604666999
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1604666999
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_80
timestamp 1604666999
transform 1 0 8464 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604666999
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604666999
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11408 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_102
timestamp 1604666999
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_107
timestamp 1604666999
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_131
timestamp 1604666999
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_135
timestamp 1604666999
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604666999
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15364 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_139
timestamp 1604666999
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604666999
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1604666999
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_154
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16928 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_164
timestamp 1604666999
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1604666999
transform 1 0 16560 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 1604666999
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_195
timestamp 1604666999
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604666999
transform 1 0 19688 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_199
timestamp 1604666999
transform 1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604666999
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604666999
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_234
timestamp 1604666999
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_238
timestamp 1604666999
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 23368 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 24748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_251
timestamp 1604666999
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_255
timestamp 1604666999
transform 1 0 24564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604666999
transform 1 0 24932 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604666999
transform 1 0 25484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_263
timestamp 1604666999
transform 1 0 25300 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_267
timestamp 1604666999
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1604666999
transform 1 0 1472 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 1604666999
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_17
timestamp 1604666999
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 3128 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604666999
transform 1 0 5612 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604666999
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1604666999
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_45
timestamp 1604666999
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604666999
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604666999
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7820 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_65
timestamp 1604666999
transform 1 0 7084 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_70
timestamp 1604666999
transform 1 0 7544 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9384 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_82
timestamp 1604666999
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1604666999
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1604666999
transform 1 0 11132 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1604666999
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_136
timestamp 1604666999
transform 1 0 13616 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 14260 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_140
timestamp 1604666999
transform 1 0 13984 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604666999
transform 1 0 16928 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1604666999
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1604666999
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_170
timestamp 1604666999
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1604666999
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604666999
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604666999
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1604666999
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604666999
transform 1 0 20056 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_201
timestamp 1604666999
transform 1 0 19596 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1604666999
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21896 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1604666999
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_225
timestamp 1604666999
transform 1 0 21804 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_235
timestamp 1604666999
transform 1 0 22724 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 24748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604666999
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_254
timestamp 1604666999
transform 1 0 24472 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604666999
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 26128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_259
timestamp 1604666999
transform 1 0 24932 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_266
timestamp 1604666999
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_270
timestamp 1604666999
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_274
timestamp 1604666999
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1604666999
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_16
timestamp 1604666999
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604666999
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1604666999
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604666999
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604666999
transform 1 0 5796 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1604666999
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_45
timestamp 1604666999
transform 1 0 5244 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_60
timestamp 1604666999
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1604666999
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1604666999
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9844 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_81
timestamp 1604666999
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1604666999
transform 1 0 8924 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_89
timestamp 1604666999
transform 1 0 9292 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11408 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp 1604666999
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 1604666999
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_131
timestamp 1604666999
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1604666999
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_139
timestamp 1604666999
transform 1 0 13892 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604666999
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_145
timestamp 1604666999
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1604666999
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_158
timestamp 1604666999
transform 1 0 15640 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 15916 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 17480 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1604666999
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_174
timestamp 1604666999
transform 1 0 17112 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19044 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_187
timestamp 1604666999
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_191
timestamp 1604666999
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_204
timestamp 1604666999
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1604666999
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 21620 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 22632 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23000 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_219
timestamp 1604666999
transform 1 0 21252 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_232
timestamp 1604666999
transform 1 0 22448 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_236
timestamp 1604666999
transform 1 0 22816 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604666999
transform 1 0 24748 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604666999
transform 1 0 23184 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 24196 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 24564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_249
timestamp 1604666999
transform 1 0 24012 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1604666999
transform 1 0 24380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 25760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_266
timestamp 1604666999
transform 1 0 25576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_270
timestamp 1604666999
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604666999
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1840 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1604666999
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1604666999
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1604666999
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1604666999
transform 1 0 3036 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1604666999
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1604666999
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604666999
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604666999
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604666999
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604666999
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_75
timestamp 1604666999
transform 1 0 8004 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_80
timestamp 1604666999
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_84
timestamp 1604666999
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1604666999
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1604666999
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604666999
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604666999
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12972 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1604666999
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14536 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_142
timestamp 1604666999
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604666999
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_165
timestamp 1604666999
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1604666999
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1604666999
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_177
timestamp 1604666999
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20884 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604666999
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1604666999
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1604666999
transform 1 0 20148 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1604666999
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_234
timestamp 1604666999
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1604666999
transform 1 0 23000 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_264
timestamp 1604666999
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_268
timestamp 1604666999
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_272
timestamp 1604666999
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_276
timestamp 1604666999
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1604666999
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_6
timestamp 1604666999
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1604666999
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1604666999
transform 1 0 3220 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1604666999
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5796 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_41
timestamp 1604666999
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1604666999
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_50
timestamp 1604666999
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604666999
transform 1 0 8280 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1604666999
transform 1 0 7544 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_74
timestamp 1604666999
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1604666999
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_86
timestamp 1604666999
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1604666999
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12052 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11592 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_112
timestamp 1604666999
transform 1 0 11408 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_116
timestamp 1604666999
transform 1 0 11776 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604666999
transform 1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1604666999
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1604666999
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_132
timestamp 1604666999
transform 1 0 13248 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1604666999
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604666999
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604666999
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604666999
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1604666999
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_167
timestamp 1604666999
transform 1 0 16468 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_172
timestamp 1604666999
transform 1 0 16928 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18308 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1604666999
transform 1 0 17572 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1604666999
transform 1 0 17940 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_186
timestamp 1604666999
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604666999
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1604666999
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_210
timestamp 1604666999
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21988 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21804 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_219
timestamp 1604666999
transform 1 0 21252 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_223
timestamp 1604666999
transform 1 0 21620 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 24472 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 23920 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_246
timestamp 1604666999
transform 1 0 23736 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1604666999
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 25484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_263
timestamp 1604666999
transform 1 0 25300 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1604666999
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_6
timestamp 1604666999
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604666999
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604666999
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_10
timestamp 1604666999
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604666999
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604666999
transform 1 0 2852 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604666999
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1604666999
transform 1 0 3680 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_34
timestamp 1604666999
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4416 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_45
timestamp 1604666999
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_51
timestamp 1604666999
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1604666999
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604666999
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_55
timestamp 1604666999
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_59
timestamp 1604666999
transform 1 0 6532 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604666999
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6348 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6716 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6900 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_76
timestamp 1604666999
transform 1 0 8096 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_72
timestamp 1604666999
transform 1 0 7728 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1604666999
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1604666999
transform 1 0 7636 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 7912 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604666999
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_84
timestamp 1604666999
transform 1 0 8832 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_97
timestamp 1604666999
transform 1 0 10028 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1604666999
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 10212 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 8556 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_34_101
timestamp 1604666999
transform 1 0 10396 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_104
timestamp 1604666999
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_100
timestamp 1604666999
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10488 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604666999
transform 1 0 11040 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_115
timestamp 1604666999
transform 1 0 11684 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_111
timestamp 1604666999
transform 1 0 11316 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1604666999
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_111
timestamp 1604666999
transform 1 0 11316 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1604666999
transform 1 0 12052 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604666999
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 13248 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1604666999
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_128
timestamp 1604666999
transform 1 0 12880 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1604666999
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604666999
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_146
timestamp 1604666999
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_142
timestamp 1604666999
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604666999
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604666999
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_150
timestamp 1604666999
transform 1 0 14904 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604666999
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604666999
transform 1 0 15640 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15364 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16744 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_174
timestamp 1604666999
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_178
timestamp 1604666999
transform 1 0 17480 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_162
timestamp 1604666999
transform 1 0 16008 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_168
timestamp 1604666999
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1604666999
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1604666999
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17664 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_193
timestamp 1604666999
transform 1 0 18860 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1604666999
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1604666999
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18676 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19044 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_206
timestamp 1604666999
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1604666999
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_210
timestamp 1604666999
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_212
timestamp 1604666999
transform 1 0 20608 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_209
timestamp 1604666999
transform 1 0 20332 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20424 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20976 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604666999
transform 1 0 22724 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604666999
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_235
timestamp 1604666999
transform 1 0 22724 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1604666999
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_228
timestamp 1604666999
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_232
timestamp 1604666999
transform 1 0 22448 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_244
timestamp 1604666999
transform 1 0 23552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_239
timestamp 1604666999
transform 1 0 23092 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_239
timestamp 1604666999
transform 1 0 23092 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 23368 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604666999
transform 1 0 23828 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_256
timestamp 1604666999
transform 1 0 24656 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604666999
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_260
timestamp 1604666999
transform 1 0 25024 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_266
timestamp 1604666999
transform 1 0 25576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 1604666999
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604666999
transform 1 0 25208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 24840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604666999
transform 1 0 25208 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604666999
transform 1 0 25392 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_267
timestamp 1604666999
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_270
timestamp 1604666999
transform 1 0 25944 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604666999
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604666999
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604666999
transform 1 0 1564 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_14
timestamp 1604666999
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_18
timestamp 1604666999
transform 1 0 2760 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 3312 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_43
timestamp 1604666999
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_47
timestamp 1604666999
transform 1 0 5428 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_53
timestamp 1604666999
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1604666999
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_71
timestamp 1604666999
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_75
timestamp 1604666999
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_79
timestamp 1604666999
transform 1 0 8372 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_84
timestamp 1604666999
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_97
timestamp 1604666999
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_101
timestamp 1604666999
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604666999
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13248 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12604 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_123
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_127
timestamp 1604666999
transform 1 0 12788 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_151
timestamp 1604666999
transform 1 0 14996 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_155
timestamp 1604666999
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_158
timestamp 1604666999
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_162
timestamp 1604666999
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1604666999
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18952 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18768 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604666999
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_184
timestamp 1604666999
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_189
timestamp 1604666999
transform 1 0 18492 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_213
timestamp 1604666999
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_217
timestamp 1604666999
transform 1 0 21068 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21436 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 22448 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1604666999
transform 1 0 22264 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_234
timestamp 1604666999
transform 1 0 22632 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 23736 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 24748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604666999
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_245
timestamp 1604666999
transform 1 0 23644 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_255
timestamp 1604666999
transform 1 0 24564 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604666999
transform 1 0 25300 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604666999
transform 1 0 25852 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_259
timestamp 1604666999
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_267
timestamp 1604666999
transform 1 0 25668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_271
timestamp 1604666999
transform 1 0 26036 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604666999
transform 1 0 1564 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_14
timestamp 1604666999
transform 1 0 2392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_18
timestamp 1604666999
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3312 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 2944 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3680 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_22
timestamp 1604666999
transform 1 0 3128 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1604666999
transform 1 0 3496 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_30
timestamp 1604666999
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6164 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5060 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5428 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_41
timestamp 1604666999
transform 1 0 4876 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_45
timestamp 1604666999
transform 1 0 5244 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_49
timestamp 1604666999
transform 1 0 5612 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1604666999
transform 1 0 5980 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8096 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_74
timestamp 1604666999
transform 1 0 7912 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_78
timestamp 1604666999
transform 1 0 8280 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9844 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8464 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_82
timestamp 1604666999
transform 1 0 8648 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604666999
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11408 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 11224 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_104
timestamp 1604666999
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_108
timestamp 1604666999
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_131
timestamp 1604666999
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1604666999
transform 1 0 13524 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13892 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604666999
transform 1 0 14076 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1604666999
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604666999
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1604666999
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1604666999
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604666999
transform 1 0 15640 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1604666999
transform 1 0 16744 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 16560 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_162
timestamp 1604666999
transform 1 0 16008 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_166
timestamp 1604666999
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18308 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18124 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17756 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_179
timestamp 1604666999
transform 1 0 17572 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_183
timestamp 1604666999
transform 1 0 17940 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604666999
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_206
timestamp 1604666999
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_210
timestamp 1604666999
transform 1 0 20424 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_215
timestamp 1604666999
transform 1 0 20884 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604666999
transform 1 0 21804 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 21436 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_223
timestamp 1604666999
transform 1 0 21620 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_234
timestamp 1604666999
transform 1 0 22632 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604666999
transform 1 0 23368 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 24380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 24748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 23184 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_251
timestamp 1604666999
transform 1 0 24196 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_255
timestamp 1604666999
transform 1 0 24564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604666999
transform 1 0 24932 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604666999
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604666999
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 1748 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1604666999
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604666999
transform 1 0 3312 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 3128 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_20
timestamp 1604666999
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_33
timestamp 1604666999
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_37
timestamp 1604666999
transform 1 0 4508 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4876 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5888 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_50
timestamp 1604666999
transform 1 0 5704 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_54
timestamp 1604666999
transform 1 0 6072 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_58
timestamp 1604666999
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8004 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 7452 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_66
timestamp 1604666999
transform 1 0 7176 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1604666999
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 9936 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_94
timestamp 1604666999
transform 1 0 9752 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_98
timestamp 1604666999
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10488 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11500 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11868 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_111
timestamp 1604666999
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_115
timestamp 1604666999
transform 1 0 11684 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_119
timestamp 1604666999
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12880 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 12604 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_127
timestamp 1604666999
transform 1 0 12788 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_131
timestamp 1604666999
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_135
timestamp 1604666999
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 13892 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_158
timestamp 1604666999
transform 1 0 15640 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_162
timestamp 1604666999
transform 1 0 16008 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_165
timestamp 1604666999
transform 1 0 16284 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604666999
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604666999
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_193
timestamp 1604666999
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1604666999
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 19596 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604666999
transform 1 0 22448 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 21528 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 21896 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604666999
transform 1 0 22264 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_220
timestamp 1604666999
transform 1 0 21344 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_224
timestamp 1604666999
transform 1 0 21712 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_228
timestamp 1604666999
transform 1 0 22080 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1604666999
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604666999
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_254
timestamp 1604666999
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604666999
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604666999
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_258
timestamp 1604666999
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_266
timestamp 1604666999
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_270
timestamp 1604666999
transform 1 0 25944 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604666999
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1604666999
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_6
timestamp 1604666999
transform 1 0 1656 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_10
timestamp 1604666999
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 4600 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1604666999
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1604666999
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_36
timestamp 1604666999
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4876 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_38_40
timestamp 1604666999
transform 1 0 4784 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_60
timestamp 1604666999
transform 1 0 6624 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_64
timestamp 1604666999
transform 1 0 6992 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_68
timestamp 1604666999
transform 1 0 7360 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_71
timestamp 1604666999
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_84
timestamp 1604666999
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604666999
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11500 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_102
timestamp 1604666999
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_106
timestamp 1604666999
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_110
timestamp 1604666999
transform 1 0 11224 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_132
timestamp 1604666999
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1604666999
transform 1 0 13616 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_140
timestamp 1604666999
transform 1 0 13984 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604666999
transform 1 0 14076 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1604666999
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604666999
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1604666999
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_158
timestamp 1604666999
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_154
timestamp 1604666999
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 15456 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16100 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_162
timestamp 1604666999
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18308 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19044 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_182
timestamp 1604666999
transform 1 0 17848 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_186
timestamp 1604666999
transform 1 0 18216 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_189
timestamp 1604666999
transform 1 0 18492 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_193
timestamp 1604666999
transform 1 0 18860 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_206
timestamp 1604666999
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1604666999
transform 1 0 20424 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_215
timestamp 1604666999
transform 1 0 20884 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 21528 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 21344 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_219
timestamp 1604666999
transform 1 0 21252 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604666999
transform 1 0 24012 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 23460 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 23828 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_241
timestamp 1604666999
transform 1 0 23276 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_245
timestamp 1604666999
transform 1 0 23644 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604666999
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 25024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604666999
transform 1 0 25392 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_258
timestamp 1604666999
transform 1 0 24840 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_262
timestamp 1604666999
transform 1 0 25208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_266
timestamp 1604666999
transform 1 0 25576 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604666999
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604666999
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_6
timestamp 1604666999
transform 1 0 1656 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_6
timestamp 1604666999
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 1840 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_10
timestamp 1604666999
transform 1 0 2024 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_10
timestamp 1604666999
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 2208 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2392 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1604666999
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_23
timestamp 1604666999
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_27
timestamp 1604666999
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_23
timestamp 1604666999
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 3772 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1604666999
transform 1 0 4140 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 3956 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_46
timestamp 1604666999
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_42
timestamp 1604666999
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_58
timestamp 1604666999
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1604666999
transform 1 0 6072 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_50
timestamp 1604666999
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6256 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5888 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5704 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_69
timestamp 1604666999
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_66
timestamp 1604666999
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604666999
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_73
timestamp 1604666999
transform 1 0 7820 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_74
timestamp 1604666999
transform 1 0 7912 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1604666999
transform 1 0 7544 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7636 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8004 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604666999
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604666999
transform 1 0 8188 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604666999
transform 1 0 8188 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_89
timestamp 1604666999
transform 1 0 9292 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1604666999
transform 1 0 8924 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_81
timestamp 1604666999
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_86
timestamp 1604666999
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9108 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8740 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_96
timestamp 1604666999
transform 1 0 9936 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_90
timestamp 1604666999
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10120 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 9752 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10672 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11684 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1604666999
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_117
timestamp 1604666999
transform 1 0 11868 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_100
timestamp 1604666999
transform 1 0 10304 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1604666999
transform 1 0 11500 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_117
timestamp 1604666999
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_127
timestamp 1604666999
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_123
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12604 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12236 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1604666999
transform 1 0 13432 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_130
timestamp 1604666999
transform 1 0 13064 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13248 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12972 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_145
timestamp 1604666999
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_140
timestamp 1604666999
transform 1 0 13984 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_148
timestamp 1604666999
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604666999
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604666999
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_158
timestamp 1604666999
transform 1 0 15640 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1604666999
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1604666999
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_152
timestamp 1604666999
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 15456 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604666999
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15456 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 17296 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15732 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17112 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_175
timestamp 1604666999
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_168
timestamp 1604666999
transform 1 0 16560 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_185
timestamp 1604666999
transform 1 0 18124 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_184
timestamp 1604666999
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604666999
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604666999
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18308 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_40_193
timestamp 1604666999
transform 1 0 18860 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_189
timestamp 1604666999
transform 1 0 18492 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_196
timestamp 1604666999
transform 1 0 19136 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604666999
transform 1 0 18952 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19320 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604666999
transform 1 0 19136 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_207
timestamp 1604666999
transform 1 0 20148 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_204
timestamp 1604666999
transform 1 0 19872 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_200
timestamp 1604666999
transform 1 0 19504 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_207
timestamp 1604666999
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1604666999
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604666999
transform 1 0 19964 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19872 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_215
timestamp 1604666999
transform 1 0 20884 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_212
timestamp 1604666999
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_211
timestamp 1604666999
transform 1 0 20516 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 21160 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604666999
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 20884 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21712 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21528 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 22724 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_234
timestamp 1604666999
transform 1 0 22632 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_220
timestamp 1604666999
transform 1 0 21344 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_233
timestamp 1604666999
transform 1 0 22540 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_237
timestamp 1604666999
transform 1 0 22908 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1604666999
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_239
timestamp 1604666999
transform 1 0 23092 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 23276 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604666999
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1604666999
transform 1 0 23276 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_254
timestamp 1604666999
transform 1 0 24472 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1604666999
transform 1 0 24104 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1604666999
transform 1 0 24472 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 24288 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604666999
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_266
timestamp 1604666999
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_260
timestamp 1604666999
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1604666999
transform 1 0 24840 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604666999
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604666999
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_276
timestamp 1604666999
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_270
timestamp 1604666999
transform 1 0 25944 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604666999
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 1564 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 2576 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_14
timestamp 1604666999
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_18
timestamp 1604666999
transform 1 0 2760 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 3128 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 2944 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604666999
transform 1 0 5612 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604666999
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 5244 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_41
timestamp 1604666999
transform 1 0 4876 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_47
timestamp 1604666999
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604666999
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604666999
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_71
timestamp 1604666999
transform 1 0 7636 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_75
timestamp 1604666999
transform 1 0 8004 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_78
timestamp 1604666999
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8464 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1604666999
transform 1 0 10212 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 11316 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_105
timestamp 1604666999
transform 1 0 10764 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_109
timestamp 1604666999
transform 1 0 11132 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604666999
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604666999
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604666999
transform 1 0 12972 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_138
timestamp 1604666999
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604666999
transform 1 0 14996 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_142
timestamp 1604666999
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_146
timestamp 1604666999
transform 1 0 14536 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604666999
transform 1 0 16560 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 16008 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17112 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604666999
transform 1 0 17480 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_160
timestamp 1604666999
transform 1 0 15824 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_164
timestamp 1604666999
transform 1 0 16192 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_172
timestamp 1604666999
transform 1 0 16928 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_176
timestamp 1604666999
transform 1 0 17296 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604666999
transform 1 0 19044 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604666999
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604666999
transform 1 0 18492 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604666999
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1604666999
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_187
timestamp 1604666999
transform 1 0 18308 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_191
timestamp 1604666999
transform 1 0 18676 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20424 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 20240 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 19872 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_199
timestamp 1604666999
transform 1 0 19412 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_203
timestamp 1604666999
transform 1 0 19780 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_206
timestamp 1604666999
transform 1 0 20056 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21988 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 21436 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_219
timestamp 1604666999
transform 1 0 21252 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_223
timestamp 1604666999
transform 1 0 21620 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_236
timestamp 1604666999
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1604666999
transform 1 0 23644 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604666999
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_240
timestamp 1604666999
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_254
timestamp 1604666999
transform 1 0 24472 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604666999
transform 1 0 25208 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 25024 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25760 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_258
timestamp 1604666999
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_266
timestamp 1604666999
transform 1 0 25576 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_270
timestamp 1604666999
transform 1 0 25944 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_276
timestamp 1604666999
transform 1 0 26496 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 1840 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_6
timestamp 1604666999
transform 1 0 1656 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_10
timestamp 1604666999
transform 1 0 2024 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 4600 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_23
timestamp 1604666999
transform 1 0 3220 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1604666999
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_36
timestamp 1604666999
transform 1 0 4416 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5244 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5060 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604666999
transform 1 0 6256 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_40
timestamp 1604666999
transform 1 0 4784 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_54
timestamp 1604666999
transform 1 0 6072 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_58
timestamp 1604666999
transform 1 0 6440 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8096 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 7084 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7544 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 7912 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_63
timestamp 1604666999
transform 1 0 6900 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_68
timestamp 1604666999
transform 1 0 7360 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_72
timestamp 1604666999
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9936 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1604666999
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_89
timestamp 1604666999
transform 1 0 9292 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_94
timestamp 1604666999
transform 1 0 9752 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_99
timestamp 1604666999
transform 1 0 10212 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10948 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 10396 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_103
timestamp 1604666999
transform 1 0 10580 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_116
timestamp 1604666999
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12604 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604666999
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_120
timestamp 1604666999
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_134
timestamp 1604666999
transform 1 0 13432 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604666999
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15456 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604666999
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_142
timestamp 1604666999
transform 1 0 14168 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1604666999
transform 1 0 14628 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_153
timestamp 1604666999
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604666999
transform 1 0 17112 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604666999
transform 1 0 16560 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_165
timestamp 1604666999
transform 1 0 16284 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_170
timestamp 1604666999
transform 1 0 16744 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_178
timestamp 1604666999
transform 1 0 17480 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604666999
transform 1 0 18400 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604666999
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_187
timestamp 1604666999
transform 1 0 18308 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_192
timestamp 1604666999
transform 1 0 18768 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604666999
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604666999
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_204
timestamp 1604666999
transform 1 0 19872 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1604666999
transform 1 0 20332 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_218
timestamp 1604666999
transform 1 0 21160 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604666999
transform 1 0 22816 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604666999
transform 1 0 21712 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604666999
transform 1 0 22264 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 22632 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604666999
transform 1 0 21528 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_228
timestamp 1604666999
transform 1 0 22080 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_232
timestamp 1604666999
transform 1 0 22448 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604666999
transform 1 0 24012 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604666999
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 23644 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_240
timestamp 1604666999
transform 1 0 23184 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_244
timestamp 1604666999
transform 1 0 23552 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_247
timestamp 1604666999
transform 1 0 23828 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25576 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604666999
transform 1 0 25208 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_258
timestamp 1604666999
transform 1 0 24840 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_264
timestamp 1604666999
transform 1 0 25392 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_269
timestamp 1604666999
transform 1 0 25852 0 -1 25568
box -38 -48 774 592
<< labels >>
rlabel metal2 s 13910 0 13966 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 23202 0 23258 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21904 480 22024 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 27520 824 28000 944 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 27520 4224 28000 4344 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 4894 27520 4950 28000 6 chany_top_in[0]
port 82 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[10]
port 83 nsew default input
rlabel metal2 s 11334 27520 11390 28000 6 chany_top_in[11]
port 84 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[12]
port 85 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 86 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 87 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 88 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 89 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 90 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 91 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_in[19]
port 92 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[1]
port 93 nsew default input
rlabel metal2 s 6090 27520 6146 28000 6 chany_top_in[2]
port 94 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[3]
port 95 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[4]
port 96 nsew default input
rlabel metal2 s 7838 27520 7894 28000 6 chany_top_in[5]
port 97 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[6]
port 98 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[7]
port 99 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[8]
port 100 nsew default input
rlabel metal2 s 10138 27520 10194 28000 6 chany_top_in[9]
port 101 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[0]
port 102 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[10]
port 103 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[11]
port 104 nsew default tristate
rlabel metal2 s 23570 27520 23626 28000 6 chany_top_out[12]
port 105 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[13]
port 106 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[14]
port 107 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[15]
port 108 nsew default tristate
rlabel metal2 s 25870 27520 25926 28000 6 chany_top_out[16]
port 109 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[17]
port 110 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[18]
port 111 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 chany_top_out[19]
port 112 nsew default tristate
rlabel metal2 s 17130 27520 17186 28000 6 chany_top_out[1]
port 113 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 114 nsew default tristate
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_out[3]
port 115 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_top_out[4]
port 116 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[5]
port 117 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[6]
port 118 nsew default tristate
rlabel metal2 s 20626 27520 20682 28000 6 chany_top_out[7]
port 119 nsew default tristate
rlabel metal2 s 21270 27520 21326 28000 6 chany_top_out[8]
port 120 nsew default tristate
rlabel metal2 s 21822 27520 21878 28000 6 chany_top_out[9]
port 121 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 122 nsew default input
rlabel metal3 s 0 23672 480 23792 6 left_top_grid_pin_42_
port 123 nsew default input
rlabel metal3 s 0 24216 480 24336 6 left_top_grid_pin_43_
port 124 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 125 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 126 nsew default input
rlabel metal3 s 0 25984 480 26104 6 left_top_grid_pin_46_
port 127 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 128 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 129 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 130 nsew default input
rlabel metal2 s 4618 0 4674 480 6 prog_clk
port 131 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_1_
port 132 nsew default input
rlabel metal3 s 27520 23672 28000 23792 6 right_top_grid_pin_42_
port 133 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 right_top_grid_pin_43_
port 134 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 135 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 136 nsew default input
rlabel metal3 s 27520 25984 28000 26104 6 right_top_grid_pin_46_
port 137 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 138 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 139 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 140 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 141 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 142 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 143 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 top_left_grid_pin_37_
port 144 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 top_left_grid_pin_38_
port 145 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 146 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 top_left_grid_pin_40_
port 147 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 top_left_grid_pin_41_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
