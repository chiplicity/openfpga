magic
tech sky130A
magscale 1 2
timestamp 1606150568
<< locali >>
rect 84997 202199 85031 208965
rect 84537 192407 84571 201961
rect 122533 182819 122567 192305
rect 74693 134199 74727 134369
rect 116185 134131 116219 134301
rect 128547 134233 128639 134267
rect 125753 134131 125787 134233
rect 128605 134199 128639 134233
rect 64205 99927 64239 100029
rect 65125 99927 65159 100301
rect 72761 100199 72795 100369
rect 74693 99927 74727 100301
rect 74785 99927 74819 100097
rect 80305 99927 80339 100165
rect 99533 99995 99567 100097
rect 106525 99995 106559 100233
rect 116093 100131 116127 100233
rect 26209 96799 26243 96969
rect 74693 51375 74727 51545
rect 87205 51171 87239 51273
rect 96773 51171 96807 51409
rect 116185 51239 116219 51409
rect 125753 51307 125787 51409
rect 128547 51273 128605 51307
rect 74049 18055 74083 18429
rect 65217 17647 65251 17749
<< viali >>
rect 84997 208965 85031 208999
rect 84997 202165 85031 202199
rect 84537 201961 84571 201995
rect 84537 192373 84571 192407
rect 122533 192305 122567 192339
rect 122533 182785 122567 182819
rect 91713 141441 91747 141475
rect 78097 134709 78131 134743
rect 74693 134369 74727 134403
rect 74693 134165 74727 134199
rect 116185 134301 116219 134335
rect 116185 134097 116219 134131
rect 125753 134233 125787 134267
rect 128513 134233 128547 134267
rect 128605 134165 128639 134199
rect 125753 134097 125787 134131
rect 91437 133621 91471 133655
rect 85181 106829 85215 106863
rect 91069 104653 91103 104687
rect 72761 100369 72795 100403
rect 65125 100301 65159 100335
rect 64205 100029 64239 100063
rect 64205 99893 64239 99927
rect 72761 100165 72795 100199
rect 74693 100301 74727 100335
rect 65125 99893 65159 99927
rect 106525 100233 106559 100267
rect 80305 100165 80339 100199
rect 74693 99893 74727 99927
rect 74785 100097 74819 100131
rect 74785 99893 74819 99927
rect 99533 100097 99567 100131
rect 99533 99961 99567 99995
rect 116093 100233 116127 100267
rect 116093 100097 116127 100131
rect 106525 99961 106559 99995
rect 80305 99893 80339 99927
rect 26209 96969 26243 97003
rect 26209 96765 26243 96799
rect 74693 51545 74727 51579
rect 74693 51341 74727 51375
rect 96773 51409 96807 51443
rect 87205 51273 87239 51307
rect 87205 51137 87239 51171
rect 116185 51409 116219 51443
rect 125753 51409 125787 51443
rect 125753 51273 125787 51307
rect 128513 51273 128547 51307
rect 128605 51273 128639 51307
rect 116185 51205 116219 51239
rect 96773 51137 96807 51171
rect 74049 18429 74083 18463
rect 74049 18021 74083 18055
rect 65217 17749 65251 17783
rect 65217 17613 65251 17647
<< metal1 >>
rect 80198 216504 80204 216556
rect 80256 216544 80262 216556
rect 89766 216544 89772 216556
rect 80256 216516 89772 216544
rect 80256 216504 80262 216516
rect 89766 216504 89772 216516
rect 89824 216504 89830 216556
rect 83142 216436 83148 216488
rect 83200 216476 83206 216488
rect 153798 216476 153804 216488
rect 83200 216448 153804 216476
rect 83200 216436 83206 216448
rect 153798 216436 153804 216448
rect 153856 216436 153862 216488
rect 155546 216436 155552 216488
rect 155604 216476 155610 216488
rect 185814 216476 185820 216488
rect 155604 216448 185820 216476
rect 155604 216436 155610 216448
rect 185814 216436 185820 216448
rect 185872 216436 185878 216488
rect 22698 213104 22704 213156
rect 22756 213144 22762 213156
rect 56738 213144 56744 213156
rect 22756 213116 56744 213144
rect 22756 213104 22762 213116
rect 56738 213104 56744 213116
rect 56796 213104 56802 213156
rect 66490 213104 66496 213156
rect 66548 213144 66554 213156
rect 115066 213144 115072 213156
rect 66548 213116 115072 213144
rect 66548 213104 66554 213116
rect 115066 213104 115072 213116
rect 115124 213104 115130 213156
rect 56186 211676 56192 211728
rect 56244 211716 56250 211728
rect 56738 211716 56744 211728
rect 56244 211688 56744 211716
rect 56244 211676 56250 211688
rect 56738 211676 56744 211688
rect 56796 211716 56802 211728
rect 96482 211716 96488 211728
rect 56796 211688 96488 211716
rect 56796 211676 56802 211688
rect 96482 211676 96488 211688
rect 96540 211716 96546 211728
rect 128866 211716 128872 211728
rect 96540 211688 128872 211716
rect 96540 211676 96546 211688
rect 128866 211676 128872 211688
rect 128924 211676 128930 211728
rect 25826 210996 25832 211048
rect 25884 211036 25890 211048
rect 76518 211036 76524 211048
rect 25884 211008 76524 211036
rect 25884 210996 25890 211008
rect 76518 210996 76524 211008
rect 76576 210996 76582 211048
rect 121782 210996 121788 211048
rect 121840 211036 121846 211048
rect 151590 211036 151596 211048
rect 121840 211008 151596 211036
rect 121840 210996 121846 211008
rect 151590 210996 151596 211008
rect 151648 210996 151654 211048
rect 57658 210928 57664 210980
rect 57716 210968 57722 210980
rect 148278 210968 148284 210980
rect 57716 210940 148284 210968
rect 57716 210928 57722 210940
rect 148278 210928 148284 210940
rect 148336 210928 148342 210980
rect 28126 210588 28132 210640
rect 28184 210588 28190 210640
rect 105958 210588 105964 210640
rect 106016 210588 106022 210640
rect 28144 210356 28172 210588
rect 47262 210384 47268 210436
rect 47320 210424 47326 210436
rect 59866 210424 59872 210436
rect 47320 210396 59872 210424
rect 47320 210384 47326 210396
rect 59866 210384 59872 210396
rect 59924 210384 59930 210436
rect 69802 210356 69808 210368
rect 28144 210328 69808 210356
rect 69802 210316 69808 210328
rect 69860 210316 69866 210368
rect 105976 210356 106004 210588
rect 128866 210384 128872 210436
rect 128924 210424 128930 210436
rect 192070 210424 192076 210436
rect 128924 210396 192076 210424
rect 128924 210384 128930 210396
rect 192070 210384 192076 210396
rect 192128 210384 192134 210436
rect 141470 210356 141476 210368
rect 105976 210328 141476 210356
rect 141470 210316 141476 210328
rect 141528 210316 141534 210368
rect 156834 210316 156840 210368
rect 156892 210356 156898 210368
rect 160330 210356 160336 210368
rect 156892 210328 160336 210356
rect 156892 210316 156898 210328
rect 160330 210316 160336 210328
rect 160388 210316 160394 210368
rect 13314 209568 13320 209620
rect 13372 209608 13378 209620
rect 191702 209608 191708 209620
rect 13372 209580 191708 209608
rect 13372 209568 13378 209580
rect 191702 209568 191708 209580
rect 191760 209568 191766 209620
rect 84985 208999 85043 209005
rect 84985 208965 84997 208999
rect 85031 208996 85043 208999
rect 88570 208996 88576 209008
rect 85031 208968 88576 208996
rect 85031 208965 85043 208968
rect 84985 208959 85043 208965
rect 88570 208956 88576 208968
rect 88628 208956 88634 209008
rect 159042 207188 159048 207240
rect 159100 207228 159106 207240
rect 160514 207228 160520 207240
rect 159100 207200 160520 207228
rect 159100 207188 159106 207200
rect 160514 207188 160520 207200
rect 160572 207188 160578 207240
rect 159042 206780 159048 206832
rect 159100 206820 159106 206832
rect 160606 206820 160612 206832
rect 159100 206792 160612 206820
rect 159100 206780 159106 206792
rect 160606 206780 160612 206792
rect 160664 206780 160670 206832
rect 122150 205352 122156 205404
rect 122208 205392 122214 205404
rect 124358 205392 124364 205404
rect 122208 205364 124364 205392
rect 122208 205352 122214 205364
rect 124358 205352 124364 205364
rect 124416 205352 124422 205404
rect 49286 204672 49292 204724
rect 49344 204712 49350 204724
rect 50482 204712 50488 204724
rect 49344 204684 50488 204712
rect 49344 204672 49350 204684
rect 50482 204672 50488 204684
rect 50540 204672 50546 204724
rect 159042 203380 159048 203432
rect 159100 203420 159106 203432
rect 160514 203420 160520 203432
rect 159100 203392 160520 203420
rect 159100 203380 159106 203392
rect 160514 203380 160520 203392
rect 160572 203380 160578 203432
rect 84982 202196 84988 202208
rect 84943 202168 84988 202196
rect 84982 202156 84988 202168
rect 85040 202156 85046 202208
rect 120862 202020 120868 202072
rect 120920 202060 120926 202072
rect 122426 202060 122432 202072
rect 120920 202032 122432 202060
rect 120920 202020 120926 202032
rect 122426 202020 122432 202032
rect 122484 202020 122490 202072
rect 84525 201995 84583 202001
rect 84525 201961 84537 201995
rect 84571 201992 84583 201995
rect 84982 201992 84988 202004
rect 84571 201964 84988 201992
rect 84571 201961 84583 201964
rect 84525 201955 84583 201961
rect 84982 201952 84988 201964
rect 85040 201952 85046 202004
rect 158950 201884 158956 201936
rect 159008 201924 159014 201936
rect 160606 201924 160612 201936
rect 159008 201896 160612 201924
rect 159008 201884 159014 201896
rect 160606 201884 160612 201896
rect 160664 201884 160670 201936
rect 87190 201272 87196 201324
rect 87248 201312 87254 201324
rect 88938 201312 88944 201324
rect 87248 201284 88944 201312
rect 87248 201272 87254 201284
rect 88938 201272 88944 201284
rect 88996 201272 89002 201324
rect 87190 199300 87196 199352
rect 87248 199340 87254 199352
rect 88938 199340 88944 199352
rect 87248 199312 88944 199340
rect 87248 199300 87254 199312
rect 88938 199300 88944 199312
rect 88996 199300 89002 199352
rect 158950 198688 158956 198740
rect 159008 198728 159014 198740
rect 160514 198728 160520 198740
rect 159008 198700 160520 198728
rect 159008 198688 159014 198700
rect 160514 198688 160520 198700
rect 160572 198688 160578 198740
rect 87190 197532 87196 197584
rect 87248 197572 87254 197584
rect 88938 197572 88944 197584
rect 87248 197544 88944 197572
rect 87248 197532 87254 197544
rect 88938 197532 88944 197544
rect 88996 197532 89002 197584
rect 121782 196512 121788 196564
rect 121840 196552 121846 196564
rect 124174 196552 124180 196564
rect 121840 196524 124180 196552
rect 121840 196512 121846 196524
rect 124174 196512 124180 196524
rect 124232 196512 124238 196564
rect 158950 195356 158956 195408
rect 159008 195396 159014 195408
rect 160514 195396 160520 195408
rect 159008 195368 160520 195396
rect 159008 195356 159014 195368
rect 160514 195356 160520 195368
rect 160572 195356 160578 195408
rect 122242 194132 122248 194184
rect 122300 194172 122306 194184
rect 123346 194172 123352 194184
rect 122300 194144 123352 194172
rect 122300 194132 122306 194144
rect 123346 194132 123352 194144
rect 123404 194132 123410 194184
rect 50298 192364 50304 192416
rect 50356 192404 50362 192416
rect 50482 192404 50488 192416
rect 50356 192376 50488 192404
rect 50356 192364 50362 192376
rect 50482 192364 50488 192376
rect 50540 192364 50546 192416
rect 84522 192404 84528 192416
rect 84483 192376 84528 192404
rect 84522 192364 84528 192376
rect 84580 192364 84586 192416
rect 122518 192336 122524 192348
rect 122479 192308 122524 192336
rect 122518 192296 122524 192308
rect 122576 192296 122582 192348
rect 87190 192092 87196 192144
rect 87248 192132 87254 192144
rect 88846 192132 88852 192144
rect 87248 192104 88852 192132
rect 87248 192092 87254 192104
rect 88846 192092 88852 192104
rect 88904 192092 88910 192144
rect 122150 191480 122156 191532
rect 122208 191520 122214 191532
rect 123346 191520 123352 191532
rect 122208 191492 123352 191520
rect 122208 191480 122214 191492
rect 123346 191480 123352 191492
rect 123404 191480 123410 191532
rect 194738 191004 194744 191056
rect 194796 191044 194802 191056
rect 196854 191044 196860 191056
rect 194796 191016 196860 191044
rect 194796 191004 194802 191016
rect 196854 191004 196860 191016
rect 196912 191004 196918 191056
rect 158950 190868 158956 190920
rect 159008 190908 159014 190920
rect 160606 190908 160612 190920
rect 159008 190880 160612 190908
rect 159008 190868 159014 190880
rect 160606 190868 160612 190880
rect 160664 190868 160670 190920
rect 121966 188760 121972 188812
rect 122024 188800 122030 188812
rect 123346 188800 123352 188812
rect 122024 188772 123352 188800
rect 122024 188760 122030 188772
rect 123346 188760 123352 188772
rect 123404 188760 123410 188812
rect 87190 188216 87196 188268
rect 87248 188256 87254 188268
rect 88662 188256 88668 188268
rect 87248 188228 88668 188256
rect 87248 188216 87254 188228
rect 88662 188216 88668 188228
rect 88720 188216 88726 188268
rect 87098 186856 87104 186908
rect 87156 186896 87162 186908
rect 88570 186896 88576 186908
rect 87156 186868 88576 186896
rect 87156 186856 87162 186868
rect 88570 186856 88576 186868
rect 88628 186856 88634 186908
rect 122886 185972 122892 186024
rect 122944 186012 122950 186024
rect 126474 186012 126480 186024
rect 122944 185984 126480 186012
rect 122944 185972 122950 185984
rect 126474 185972 126480 185984
rect 126532 185972 126538 186024
rect 87006 185904 87012 185956
rect 87064 185944 87070 185956
rect 88570 185944 88576 185956
rect 87064 185916 88576 185944
rect 87064 185904 87070 185916
rect 88570 185904 88576 185916
rect 88628 185904 88634 185956
rect 122978 185700 122984 185752
rect 123036 185740 123042 185752
rect 126566 185740 126572 185752
rect 123036 185712 126572 185740
rect 123036 185700 123042 185712
rect 126566 185700 126572 185712
rect 126624 185700 126630 185752
rect 85718 185632 85724 185684
rect 85776 185672 85782 185684
rect 88570 185672 88576 185684
rect 85776 185644 88576 185672
rect 85776 185632 85782 185644
rect 88570 185632 88576 185644
rect 88628 185632 88634 185684
rect 157478 185564 157484 185616
rect 157536 185604 157542 185616
rect 160606 185604 160612 185616
rect 157536 185576 160612 185604
rect 157536 185564 157542 185576
rect 160606 185564 160612 185576
rect 160664 185564 160670 185616
rect 49930 185496 49936 185548
rect 49988 185536 49994 185548
rect 52046 185536 52052 185548
rect 49988 185508 52052 185536
rect 49988 185496 49994 185508
rect 52046 185496 52052 185508
rect 52104 185496 52110 185548
rect 158858 185496 158864 185548
rect 158916 185536 158922 185548
rect 160514 185536 160520 185548
rect 158916 185508 160520 185536
rect 158916 185496 158922 185508
rect 160514 185496 160520 185508
rect 160572 185496 160578 185548
rect 84522 185292 84528 185344
rect 84580 185292 84586 185344
rect 84246 185224 84252 185276
rect 84304 185264 84310 185276
rect 84540 185264 84568 185292
rect 84304 185236 84568 185264
rect 84304 185224 84310 185236
rect 122886 184204 122892 184256
rect 122944 184244 122950 184256
rect 124450 184244 124456 184256
rect 122944 184216 124456 184244
rect 122944 184204 122950 184216
rect 124450 184204 124456 184216
rect 124508 184204 124514 184256
rect 86454 184136 86460 184188
rect 86512 184176 86518 184188
rect 88662 184176 88668 184188
rect 86512 184148 88668 184176
rect 86512 184136 86518 184148
rect 88662 184136 88668 184148
rect 88720 184136 88726 184188
rect 122334 184136 122340 184188
rect 122392 184176 122398 184188
rect 125462 184176 125468 184188
rect 122392 184148 125468 184176
rect 122392 184136 122398 184148
rect 125462 184136 125468 184148
rect 125520 184136 125526 184188
rect 85166 184068 85172 184120
rect 85224 184108 85230 184120
rect 88570 184108 88576 184120
rect 85224 184080 88576 184108
rect 85224 184068 85230 184080
rect 88570 184068 88576 184080
rect 88628 184068 88634 184120
rect 122978 184068 122984 184120
rect 123036 184108 123042 184120
rect 124542 184108 124548 184120
rect 123036 184080 124548 184108
rect 123036 184068 123042 184080
rect 124542 184068 124548 184080
rect 124600 184068 124606 184120
rect 158214 184068 158220 184120
rect 158272 184108 158278 184120
rect 160330 184108 160336 184120
rect 158272 184080 160336 184108
rect 158272 184068 158278 184080
rect 160330 184068 160336 184080
rect 160388 184068 160394 184120
rect 122521 182819 122579 182825
rect 122521 182785 122533 182819
rect 122567 182816 122579 182819
rect 122610 182816 122616 182828
rect 122567 182788 122616 182816
rect 122567 182785 122579 182788
rect 122521 182779 122579 182785
rect 122610 182776 122616 182788
rect 122668 182776 122674 182828
rect 55376 182720 55496 182748
rect 50390 182572 50396 182624
rect 50448 182612 50454 182624
rect 55376 182612 55404 182720
rect 55468 182692 55496 182720
rect 86546 182708 86552 182760
rect 86604 182748 86610 182760
rect 88570 182748 88576 182760
rect 86604 182720 88576 182748
rect 86604 182708 86610 182720
rect 88570 182708 88576 182720
rect 88628 182708 88634 182760
rect 158306 182708 158312 182760
rect 158364 182748 158370 182760
rect 160330 182748 160336 182760
rect 158364 182720 160336 182748
rect 158364 182708 158370 182720
rect 160330 182708 160336 182720
rect 160388 182708 160394 182760
rect 55450 182640 55456 182692
rect 55508 182640 55514 182692
rect 122610 182640 122616 182692
rect 122668 182680 122674 182692
rect 127578 182680 127584 182692
rect 122668 182652 127584 182680
rect 122668 182640 122674 182652
rect 127578 182640 127584 182652
rect 127636 182640 127642 182692
rect 50448 182584 55404 182612
rect 50448 182572 50454 182584
rect 67134 182436 67140 182488
rect 67192 182476 67198 182488
rect 69802 182476 69808 182488
rect 67192 182448 69808 182476
rect 67192 182436 67198 182448
rect 69802 182436 69808 182448
rect 69860 182436 69866 182488
rect 70446 182436 70452 182488
rect 70504 182476 70510 182488
rect 74034 182476 74040 182488
rect 70504 182448 74040 182476
rect 70504 182436 70510 182448
rect 74034 182436 74040 182448
rect 74092 182436 74098 182488
rect 143678 182436 143684 182488
rect 143736 182476 143742 182488
rect 147542 182476 147548 182488
rect 143736 182448 147548 182476
rect 143736 182436 143742 182448
rect 147542 182436 147548 182448
rect 147600 182436 147606 182488
rect 66030 182368 66036 182420
rect 66088 182408 66094 182420
rect 68330 182408 68336 182420
rect 66088 182380 68336 182408
rect 66088 182368 66094 182380
rect 68330 182368 68336 182380
rect 68388 182368 68394 182420
rect 69342 182368 69348 182420
rect 69400 182408 69406 182420
rect 72654 182408 72660 182420
rect 69400 182380 72660 182408
rect 69400 182368 69406 182380
rect 72654 182368 72660 182380
rect 72712 182368 72718 182420
rect 137238 182368 137244 182420
rect 137296 182408 137302 182420
rect 138986 182408 138992 182420
rect 137296 182380 138992 182408
rect 137296 182368 137302 182380
rect 138986 182368 138992 182380
rect 139044 182368 139050 182420
rect 139446 182368 139452 182420
rect 139504 182408 139510 182420
rect 141838 182408 141844 182420
rect 139504 182380 141844 182408
rect 139504 182368 139510 182380
rect 141838 182368 141844 182380
rect 141896 182368 141902 182420
rect 142758 182368 142764 182420
rect 142816 182408 142822 182420
rect 146070 182408 146076 182420
rect 142816 182380 146076 182408
rect 142816 182368 142822 182380
rect 146070 182368 146076 182380
rect 146128 182368 146134 182420
rect 68238 182300 68244 182352
rect 68296 182340 68302 182352
rect 71182 182340 71188 182352
rect 68296 182312 71188 182340
rect 68296 182300 68302 182312
rect 71182 182300 71188 182312
rect 71240 182300 71246 182352
rect 144874 182300 144880 182352
rect 144932 182340 144938 182352
rect 148922 182340 148928 182352
rect 144932 182312 148928 182340
rect 144932 182300 144938 182312
rect 148922 182300 148928 182312
rect 148980 182300 148986 182352
rect 146070 182232 146076 182284
rect 146128 182272 146134 182284
rect 150394 182272 150400 182284
rect 146128 182244 150400 182272
rect 146128 182232 146134 182244
rect 150394 182232 150400 182244
rect 150452 182232 150458 182284
rect 134938 182164 134944 182216
rect 134996 182204 135002 182216
rect 136134 182204 136140 182216
rect 134996 182176 136140 182204
rect 134996 182164 135002 182176
rect 136134 182164 136140 182176
rect 136192 182164 136198 182216
rect 73758 182028 73764 182080
rect 73816 182068 73822 182080
rect 78358 182068 78364 182080
rect 73816 182040 78364 182068
rect 73816 182028 73822 182040
rect 78358 182028 78364 182040
rect 78416 182028 78422 182080
rect 136134 182028 136140 182080
rect 136192 182068 136198 182080
rect 137514 182068 137520 182080
rect 136192 182040 137520 182068
rect 136192 182028 136198 182040
rect 137514 182028 137520 182040
rect 137572 182028 137578 182080
rect 138158 181960 138164 182012
rect 138216 182000 138222 182012
rect 140366 182000 140372 182012
rect 138216 181972 140372 182000
rect 138216 181960 138222 181972
rect 140366 181960 140372 181972
rect 140424 181960 140430 182012
rect 61522 181892 61528 181944
rect 61580 181932 61586 181944
rect 62626 181932 62632 181944
rect 61580 181904 62632 181932
rect 61580 181892 61586 181904
rect 62626 181892 62632 181904
rect 62684 181892 62690 181944
rect 147174 181824 147180 181876
rect 147232 181864 147238 181876
rect 151774 181864 151780 181876
rect 147232 181836 151780 181864
rect 147232 181824 147238 181836
rect 151774 181824 151780 181836
rect 151832 181824 151838 181876
rect 62626 181756 62632 181808
rect 62684 181796 62690 181808
rect 64098 181796 64104 181808
rect 62684 181768 64104 181796
rect 62684 181756 62690 181768
rect 64098 181756 64104 181768
rect 64156 181756 64162 181808
rect 74862 181756 74868 181808
rect 74920 181796 74926 181808
rect 79738 181796 79744 181808
rect 74920 181768 79744 181796
rect 74920 181756 74926 181768
rect 79738 181756 79744 181768
rect 79796 181756 79802 181808
rect 64926 181416 64932 181468
rect 64984 181456 64990 181468
rect 66950 181456 66956 181468
rect 64984 181428 66956 181456
rect 64984 181416 64990 181428
rect 66950 181416 66956 181428
rect 67008 181416 67014 181468
rect 72654 181416 72660 181468
rect 72712 181456 72718 181468
rect 76886 181456 76892 181468
rect 72712 181428 76892 181456
rect 72712 181416 72718 181428
rect 76886 181416 76892 181428
rect 76944 181416 76950 181468
rect 140550 181416 140556 181468
rect 140608 181456 140614 181468
rect 143218 181456 143224 181468
rect 140608 181428 143224 181456
rect 140608 181416 140614 181428
rect 143218 181416 143224 181428
rect 143276 181416 143282 181468
rect 148278 181416 148284 181468
rect 148336 181456 148342 181468
rect 153246 181456 153252 181468
rect 148336 181428 153252 181456
rect 148336 181416 148342 181428
rect 153246 181416 153252 181428
rect 153304 181416 153310 181468
rect 63822 181348 63828 181400
rect 63880 181388 63886 181400
rect 65478 181388 65484 181400
rect 63880 181360 65484 181388
rect 63880 181348 63886 181360
rect 65478 181348 65484 181360
rect 65536 181348 65542 181400
rect 71550 181348 71556 181400
rect 71608 181388 71614 181400
rect 75506 181388 75512 181400
rect 71608 181360 75512 181388
rect 71608 181348 71614 181360
rect 75506 181348 75512 181360
rect 75564 181348 75570 181400
rect 141654 181348 141660 181400
rect 141712 181388 141718 181400
rect 144690 181388 144696 181400
rect 141712 181360 144696 181388
rect 141712 181348 141718 181360
rect 144690 181348 144696 181360
rect 144748 181348 144754 181400
rect 175694 181348 175700 181400
rect 175752 181388 175758 181400
rect 176430 181388 176436 181400
rect 175752 181360 176436 181388
rect 175752 181348 175758 181360
rect 176430 181348 176436 181360
rect 176488 181348 176494 181400
rect 20858 181280 20864 181332
rect 20916 181320 20922 181332
rect 26102 181320 26108 181332
rect 20916 181292 26108 181320
rect 20916 181280 20922 181292
rect 26102 181280 26108 181292
rect 26160 181280 26166 181332
rect 29966 181280 29972 181332
rect 30024 181320 30030 181332
rect 31346 181320 31352 181332
rect 30024 181292 31352 181320
rect 30024 181280 30030 181292
rect 31346 181280 31352 181292
rect 31404 181280 31410 181332
rect 31898 181280 31904 181332
rect 31956 181320 31962 181332
rect 32818 181320 32824 181332
rect 31956 181292 32824 181320
rect 31956 181280 31962 181292
rect 32818 181280 32824 181292
rect 32876 181280 32882 181332
rect 33186 181280 33192 181332
rect 33244 181320 33250 181332
rect 33646 181320 33652 181332
rect 33244 181292 33652 181320
rect 33244 181280 33250 181292
rect 33646 181280 33652 181292
rect 33704 181280 33710 181332
rect 36866 181280 36872 181332
rect 36924 181320 36930 181332
rect 37694 181320 37700 181332
rect 36924 181292 37700 181320
rect 36924 181280 36930 181292
rect 37694 181280 37700 181292
rect 37752 181280 37758 181332
rect 38890 181280 38896 181332
rect 38948 181320 38954 181332
rect 41006 181320 41012 181332
rect 38948 181292 41012 181320
rect 38948 181280 38954 181292
rect 41006 181280 41012 181292
rect 41064 181280 41070 181332
rect 106694 181280 106700 181332
rect 106752 181320 106758 181332
rect 107982 181320 107988 181332
rect 106752 181292 107988 181320
rect 106752 181280 106758 181292
rect 107982 181280 107988 181292
rect 108040 181280 108046 181332
rect 108350 181280 108356 181332
rect 108408 181320 108414 181332
rect 109822 181320 109828 181332
rect 108408 181292 109828 181320
rect 108408 181280 108414 181292
rect 109822 181280 109828 181292
rect 109880 181280 109886 181332
rect 130430 181280 130436 181332
rect 130488 181320 130494 181332
rect 190966 181320 190972 181332
rect 130488 181292 190972 181320
rect 130488 181280 130494 181292
rect 190966 181280 190972 181292
rect 191024 181280 191030 181332
rect 27758 181212 27764 181264
rect 27816 181252 27822 181264
rect 30426 181252 30432 181264
rect 27816 181224 30432 181252
rect 27816 181212 27822 181224
rect 30426 181212 30432 181224
rect 30484 181212 30490 181264
rect 37418 181212 37424 181264
rect 37476 181252 37482 181264
rect 38430 181252 38436 181264
rect 37476 181224 38436 181252
rect 37476 181212 37482 181224
rect 38430 181212 38436 181224
rect 38488 181212 38494 181264
rect 107154 181212 107160 181264
rect 107212 181252 107218 181264
rect 108166 181252 108172 181264
rect 107212 181224 108172 181252
rect 107212 181212 107218 181224
rect 108166 181212 108172 181224
rect 108224 181212 108230 181264
rect 168978 181212 168984 181264
rect 169036 181252 169042 181264
rect 170450 181252 170456 181264
rect 169036 181224 170456 181252
rect 169036 181212 169042 181224
rect 170450 181212 170456 181224
rect 170508 181212 170514 181264
rect 176430 181212 176436 181264
rect 176488 181252 176494 181264
rect 177258 181252 177264 181264
rect 176488 181224 177264 181252
rect 176488 181212 176494 181224
rect 177258 181212 177264 181224
rect 177316 181212 177322 181264
rect 177534 181212 177540 181264
rect 177592 181252 177598 181264
rect 178270 181252 178276 181264
rect 177592 181224 178276 181252
rect 177592 181212 177598 181224
rect 178270 181212 178276 181224
rect 178328 181212 178334 181264
rect 179098 181212 179104 181264
rect 179156 181252 179162 181264
rect 180478 181252 180484 181264
rect 179156 181224 180484 181252
rect 179156 181212 179162 181224
rect 180478 181212 180484 181224
rect 180536 181212 180542 181264
rect 182870 181212 182876 181264
rect 182928 181252 182934 181264
rect 185998 181252 186004 181264
rect 182928 181224 186004 181252
rect 182928 181212 182934 181224
rect 185998 181212 186004 181224
rect 186056 181212 186062 181264
rect 37694 181144 37700 181196
rect 37752 181184 37758 181196
rect 39074 181184 39080 181196
rect 37752 181156 39080 181184
rect 37752 181144 37758 181156
rect 39074 181144 39080 181156
rect 39132 181144 39138 181196
rect 40454 181144 40460 181196
rect 40512 181184 40518 181196
rect 43582 181184 43588 181196
rect 40512 181156 43588 181184
rect 40512 181144 40518 181156
rect 43582 181144 43588 181156
rect 43640 181144 43646 181196
rect 106234 181144 106240 181196
rect 106292 181184 106298 181196
rect 107062 181184 107068 181196
rect 106292 181156 107068 181184
rect 106292 181144 106298 181156
rect 107062 181144 107068 181156
rect 107120 181144 107126 181196
rect 107522 181144 107528 181196
rect 107580 181184 107586 181196
rect 108718 181184 108724 181196
rect 107580 181156 108724 181184
rect 107580 181144 107586 181156
rect 108718 181144 108724 181156
rect 108776 181144 108782 181196
rect 109086 181144 109092 181196
rect 109144 181184 109150 181196
rect 110926 181184 110932 181196
rect 109144 181156 110932 181184
rect 109144 181144 109150 181156
rect 110926 181144 110932 181156
rect 110984 181144 110990 181196
rect 168426 181144 168432 181196
rect 168484 181184 168490 181196
rect 170082 181184 170088 181196
rect 168484 181156 170088 181184
rect 168484 181144 168490 181156
rect 170082 181144 170088 181156
rect 170140 181144 170146 181196
rect 176798 181144 176804 181196
rect 176856 181184 176862 181196
rect 177810 181184 177816 181196
rect 176856 181156 177816 181184
rect 176856 181144 176862 181156
rect 177810 181144 177816 181156
rect 177868 181144 177874 181196
rect 178086 181144 178092 181196
rect 178144 181184 178150 181196
rect 179374 181184 179380 181196
rect 178144 181156 179380 181184
rect 178144 181144 178150 181156
rect 179374 181144 179380 181156
rect 179432 181144 179438 181196
rect 182410 181144 182416 181196
rect 182468 181184 182474 181196
rect 185446 181184 185452 181196
rect 182468 181156 185452 181184
rect 182468 181144 182474 181156
rect 185446 181144 185452 181156
rect 185504 181144 185510 181196
rect 38430 181076 38436 181128
rect 38488 181116 38494 181128
rect 40362 181116 40368 181128
rect 38488 181088 40368 181116
rect 38488 181076 38494 181088
rect 40362 181076 40368 181088
rect 40420 181076 40426 181128
rect 177626 181076 177632 181128
rect 177684 181116 177690 181128
rect 178822 181116 178828 181128
rect 177684 181088 178828 181116
rect 177684 181076 177690 181088
rect 178822 181076 178828 181088
rect 178880 181076 178886 181128
rect 181214 181076 181220 181128
rect 181272 181116 181278 181128
rect 183790 181116 183796 181128
rect 181272 181088 183796 181116
rect 181272 181076 181278 181088
rect 183790 181076 183796 181088
rect 183848 181076 183854 181128
rect 28586 181008 28592 181060
rect 28644 181048 28650 181060
rect 30886 181048 30892 181060
rect 28644 181020 30892 181048
rect 28644 181008 28650 181020
rect 30886 181008 30892 181020
rect 30944 181008 30950 181060
rect 40086 181008 40092 181060
rect 40144 181048 40150 181060
rect 43030 181048 43036 181060
rect 40144 181020 43036 181048
rect 40144 181008 40150 181020
rect 43030 181008 43036 181020
rect 43088 181008 43094 181060
rect 108718 181008 108724 181060
rect 108776 181048 108782 181060
rect 110742 181048 110748 181060
rect 108776 181020 110748 181048
rect 108776 181008 108782 181020
rect 110742 181008 110748 181020
rect 110800 181008 110806 181060
rect 183606 181008 183612 181060
rect 183664 181048 183670 181060
rect 187102 181048 187108 181060
rect 183664 181020 187108 181048
rect 183664 181008 183670 181020
rect 187102 181008 187108 181020
rect 187160 181008 187166 181060
rect 163182 180940 163188 180992
rect 163240 180980 163246 180992
rect 167874 180980 167880 180992
rect 163240 180952 167880 180980
rect 163240 180940 163246 180952
rect 167874 180940 167880 180952
rect 167932 180940 167938 180992
rect 180846 180940 180852 180992
rect 180904 180980 180910 180992
rect 183238 180980 183244 180992
rect 180904 180952 183244 180980
rect 180904 180940 180910 180952
rect 183238 180940 183244 180952
rect 183296 180940 183302 180992
rect 27298 180872 27304 180924
rect 27356 180912 27362 180924
rect 30058 180912 30064 180924
rect 27356 180884 30064 180912
rect 27356 180872 27362 180884
rect 30058 180872 30064 180884
rect 30116 180872 30122 180924
rect 39626 180872 39632 180924
rect 39684 180912 39690 180924
rect 42294 180912 42300 180924
rect 39684 180884 42300 180912
rect 39684 180872 39690 180884
rect 42294 180872 42300 180884
rect 42352 180872 42358 180924
rect 99334 180872 99340 180924
rect 99392 180912 99398 180924
rect 99794 180912 99800 180924
rect 99392 180884 99800 180912
rect 99392 180872 99398 180884
rect 99794 180872 99800 180884
rect 99852 180872 99858 180924
rect 181674 180872 181680 180924
rect 181732 180912 181738 180924
rect 184342 180912 184348 180924
rect 181732 180884 184348 180912
rect 181732 180872 181738 180884
rect 184342 180872 184348 180884
rect 184400 180872 184406 180924
rect 183238 180804 183244 180856
rect 183296 180844 183302 180856
rect 186550 180844 186556 180856
rect 183296 180816 186556 180844
rect 183296 180804 183302 180816
rect 186550 180804 186556 180816
rect 186608 180804 186614 180856
rect 105958 180736 105964 180788
rect 106016 180776 106022 180788
rect 106510 180776 106516 180788
rect 106016 180748 106516 180776
rect 106016 180736 106022 180748
rect 106510 180736 106516 180748
rect 106568 180736 106574 180788
rect 182042 180736 182048 180788
rect 182100 180776 182106 180788
rect 184894 180776 184900 180788
rect 182100 180748 184900 180776
rect 182100 180736 182106 180748
rect 184894 180736 184900 180748
rect 184952 180736 184958 180788
rect 39258 180600 39264 180652
rect 39316 180640 39322 180652
rect 41742 180640 41748 180652
rect 39316 180612 41748 180640
rect 39316 180600 39322 180612
rect 41742 180600 41748 180612
rect 41800 180600 41806 180652
rect 168518 180600 168524 180652
rect 168576 180640 168582 180652
rect 190414 180640 190420 180652
rect 168576 180612 190420 180640
rect 168576 180600 168582 180612
rect 190414 180600 190420 180612
rect 190472 180600 190478 180652
rect 26378 180532 26384 180584
rect 26436 180572 26442 180584
rect 27850 180572 27856 180584
rect 26436 180544 27856 180572
rect 26436 180532 26442 180544
rect 27850 180532 27856 180544
rect 27908 180532 27914 180584
rect 178454 180532 178460 180584
rect 178512 180572 178518 180584
rect 179926 180572 179932 180584
rect 178512 180544 179932 180572
rect 178512 180532 178518 180544
rect 179926 180532 179932 180544
rect 179984 180532 179990 180584
rect 30518 180464 30524 180516
rect 30576 180504 30582 180516
rect 32082 180504 32088 180516
rect 30576 180476 32088 180504
rect 30576 180464 30582 180476
rect 32082 180464 32088 180476
rect 32140 180464 32146 180516
rect 24722 180396 24728 180448
rect 24780 180436 24786 180448
rect 26562 180436 26568 180448
rect 24780 180408 26568 180436
rect 24780 180396 24786 180408
rect 26562 180396 26568 180408
rect 26620 180396 26626 180448
rect 25366 180328 25372 180380
rect 25424 180368 25430 180380
rect 28862 180368 28868 180380
rect 25424 180340 28868 180368
rect 25424 180328 25430 180340
rect 28862 180328 28868 180340
rect 28920 180328 28926 180380
rect 31254 180328 31260 180380
rect 31312 180368 31318 180380
rect 32450 180368 32456 180380
rect 31312 180340 32456 180368
rect 31312 180328 31318 180340
rect 32450 180328 32456 180340
rect 32508 180328 32514 180380
rect 22790 180260 22796 180312
rect 22848 180300 22854 180312
rect 26378 180300 26384 180312
rect 22848 180272 26384 180300
rect 22848 180260 22854 180272
rect 26378 180260 26384 180272
rect 26436 180260 26442 180312
rect 92158 180260 92164 180312
rect 92216 180300 92222 180312
rect 94366 180300 94372 180312
rect 92216 180272 94372 180300
rect 92216 180260 92222 180272
rect 94366 180260 94372 180272
rect 94424 180260 94430 180312
rect 110558 180260 110564 180312
rect 110616 180300 110622 180312
rect 113502 180300 113508 180312
rect 110616 180272 113508 180300
rect 110616 180260 110622 180272
rect 113502 180260 113508 180272
rect 113560 180260 113566 180312
rect 23434 180192 23440 180244
rect 23492 180232 23498 180244
rect 25366 180232 25372 180244
rect 23492 180204 25372 180232
rect 23492 180192 23498 180204
rect 25366 180192 25372 180204
rect 25424 180192 25430 180244
rect 26010 180192 26016 180244
rect 26068 180232 26074 180244
rect 27942 180232 27948 180244
rect 26068 180204 27948 180232
rect 26068 180192 26074 180204
rect 27942 180192 27948 180204
rect 28000 180192 28006 180244
rect 29138 180192 29144 180244
rect 29196 180232 29202 180244
rect 31254 180232 31260 180244
rect 29196 180204 31260 180232
rect 29196 180192 29202 180204
rect 31254 180192 31260 180204
rect 31312 180192 31318 180244
rect 92434 180192 92440 180244
rect 92492 180232 92498 180244
rect 93262 180232 93268 180244
rect 92492 180204 93268 180232
rect 92492 180192 92498 180204
rect 93262 180192 93268 180204
rect 93320 180192 93326 180244
rect 98874 180192 98880 180244
rect 98932 180232 98938 180244
rect 99610 180232 99616 180244
rect 98932 180204 99616 180232
rect 98932 180192 98938 180204
rect 99610 180192 99616 180204
rect 99668 180192 99674 180244
rect 107798 180192 107804 180244
rect 107856 180232 107862 180244
rect 109362 180232 109368 180244
rect 107856 180204 109368 180232
rect 107856 180192 107862 180204
rect 109362 180192 109368 180204
rect 109420 180192 109426 180244
rect 111110 180192 111116 180244
rect 111168 180232 111174 180244
rect 113686 180232 113692 180244
rect 111168 180204 113692 180232
rect 111168 180192 111174 180204
rect 113686 180192 113692 180204
rect 113744 180192 113750 180244
rect 24078 180124 24084 180176
rect 24136 180164 24142 180176
rect 27758 180164 27764 180176
rect 24136 180136 27764 180164
rect 24136 180124 24142 180136
rect 27758 180124 27764 180136
rect 27816 180124 27822 180176
rect 92710 180164 92716 180176
rect 91992 180136 92716 180164
rect 21502 180056 21508 180108
rect 21560 180096 21566 180108
rect 26470 180096 26476 180108
rect 21560 180068 26476 180096
rect 21560 180056 21566 180068
rect 26470 180056 26476 180068
rect 26528 180056 26534 180108
rect 38062 180056 38068 180108
rect 38120 180096 38126 180108
rect 39718 180096 39724 180108
rect 38120 180068 39724 180096
rect 38120 180056 38126 180068
rect 39718 180056 39724 180068
rect 39776 180056 39782 180108
rect 91992 180040 92020 180136
rect 92710 180124 92716 180136
rect 92768 180124 92774 180176
rect 111570 180124 111576 180176
rect 111628 180164 111634 180176
rect 114238 180164 114244 180176
rect 111628 180136 114244 180164
rect 111628 180124 111634 180136
rect 114238 180124 114244 180136
rect 114296 180124 114302 180176
rect 169530 180124 169536 180176
rect 169588 180164 169594 180176
rect 170818 180164 170824 180176
rect 169588 180136 170824 180164
rect 169588 180124 169594 180136
rect 170818 180124 170824 180136
rect 170876 180124 170882 180176
rect 179282 180124 179288 180176
rect 179340 180164 179346 180176
rect 181030 180164 181036 180176
rect 179340 180136 181036 180164
rect 179340 180124 179346 180136
rect 181030 180124 181036 180136
rect 181088 180124 181094 180176
rect 92342 180056 92348 180108
rect 92400 180096 92406 180108
rect 94918 180096 94924 180108
rect 92400 180068 94924 180096
rect 92400 180056 92406 180068
rect 94918 180056 94924 180068
rect 94976 180056 94982 180108
rect 97770 180056 97776 180108
rect 97828 180096 97834 180108
rect 98690 180096 98696 180108
rect 97828 180068 98696 180096
rect 97828 180056 97834 180068
rect 98690 180056 98696 180068
rect 98748 180056 98754 180108
rect 110282 180056 110288 180108
rect 110340 180096 110346 180108
rect 112582 180096 112588 180108
rect 110340 180068 112588 180096
rect 110340 180056 110346 180068
rect 112582 180056 112588 180068
rect 112640 180056 112646 180108
rect 180754 180056 180760 180108
rect 180812 180096 180818 180108
rect 182686 180096 182692 180108
rect 180812 180068 182692 180096
rect 180812 180056 180818 180068
rect 182686 180056 182692 180068
rect 182744 180056 182750 180108
rect 184066 180056 184072 180108
rect 184124 180096 184130 180108
rect 187654 180096 187660 180108
rect 184124 180068 187660 180096
rect 184124 180056 184130 180068
rect 187654 180056 187660 180068
rect 187712 180056 187718 180108
rect 22146 179988 22152 180040
rect 22204 180028 22210 180040
rect 26838 180028 26844 180040
rect 22204 180000 26844 180028
rect 22204 179988 22210 180000
rect 26838 179988 26844 180000
rect 26896 179988 26902 180040
rect 91974 179988 91980 180040
rect 92032 179988 92038 180040
rect 92066 179988 92072 180040
rect 92124 180028 92130 180040
rect 92434 180028 92440 180040
rect 92124 180000 92440 180028
rect 92124 179988 92130 180000
rect 92434 179988 92440 180000
rect 92492 179988 92498 180040
rect 92618 179988 92624 180040
rect 92676 180028 92682 180040
rect 95470 180028 95476 180040
rect 92676 180000 95476 180028
rect 92676 179988 92682 180000
rect 95470 179988 95476 180000
rect 95528 179988 95534 180040
rect 97218 179988 97224 180040
rect 97276 180028 97282 180040
rect 98230 180028 98236 180040
rect 97276 180000 98236 180028
rect 97276 179988 97282 180000
rect 98230 179988 98236 180000
rect 98288 179988 98294 180040
rect 109914 179988 109920 180040
rect 109972 180028 109978 180040
rect 112030 180028 112036 180040
rect 109972 180000 112036 180028
rect 109972 179988 109978 180000
rect 112030 179988 112036 180000
rect 112088 179988 112094 180040
rect 112214 179988 112220 180040
rect 112272 180028 112278 180040
rect 115342 180028 115348 180040
rect 112272 180000 115348 180028
rect 112272 179988 112278 180000
rect 115342 179988 115348 180000
rect 115400 179988 115406 180040
rect 170634 179988 170640 180040
rect 170692 180028 170698 180040
rect 171646 180028 171652 180040
rect 170692 180000 171652 180028
rect 170692 179988 170698 180000
rect 171646 179988 171652 180000
rect 171704 179988 171710 180040
rect 179650 179988 179656 180040
rect 179708 180028 179714 180040
rect 181582 180028 181588 180040
rect 179708 180000 181588 180028
rect 179708 179988 179714 180000
rect 181582 179988 181588 180000
rect 181640 179988 181646 180040
rect 36222 179960 36228 179972
rect 36056 179932 36228 179960
rect 36056 179904 36084 179932
rect 36222 179920 36228 179932
rect 36280 179920 36286 179972
rect 92250 179920 92256 179972
rect 92308 179960 92314 179972
rect 94090 179960 94096 179972
rect 92308 179932 94096 179960
rect 92308 179920 92314 179932
rect 94090 179920 94096 179932
rect 94148 179920 94154 179972
rect 96666 179920 96672 179972
rect 96724 179960 96730 179972
rect 97770 179960 97776 179972
rect 96724 179932 97776 179960
rect 96724 179920 96730 179932
rect 97770 179920 97776 179932
rect 97828 179920 97834 179972
rect 98138 179920 98144 179972
rect 98196 179960 98202 179972
rect 98966 179960 98972 179972
rect 98196 179932 98972 179960
rect 98196 179920 98202 179932
rect 98966 179920 98972 179932
rect 99024 179920 99030 179972
rect 100714 179920 100720 179972
rect 100772 179960 100778 179972
rect 100990 179960 100996 179972
rect 100772 179932 100996 179960
rect 100772 179920 100778 179932
rect 100990 179920 100996 179932
rect 101048 179920 101054 179972
rect 105038 179920 105044 179972
rect 105096 179960 105102 179972
rect 105498 179960 105504 179972
rect 105096 179932 105504 179960
rect 105096 179920 105102 179932
rect 105498 179920 105504 179932
rect 105556 179920 105562 179972
rect 109546 179920 109552 179972
rect 109604 179960 109610 179972
rect 111478 179960 111484 179972
rect 109604 179932 111484 179960
rect 109604 179920 109610 179932
rect 111478 179920 111484 179932
rect 111536 179920 111542 179972
rect 111938 179920 111944 179972
rect 111996 179960 112002 179972
rect 114790 179960 114796 179972
rect 111996 179932 114796 179960
rect 111996 179920 112002 179932
rect 114790 179920 114796 179932
rect 114848 179920 114854 179972
rect 171186 179920 171192 179972
rect 171244 179960 171250 179972
rect 172014 179960 172020 179972
rect 171244 179932 172020 179960
rect 171244 179920 171250 179932
rect 172014 179920 172020 179932
rect 172072 179920 172078 179972
rect 180018 179920 180024 179972
rect 180076 179960 180082 179972
rect 182134 179960 182140 179972
rect 180076 179932 182140 179960
rect 180076 179920 180082 179932
rect 182134 179920 182140 179932
rect 182192 179920 182198 179972
rect 36038 179852 36044 179904
rect 36096 179852 36102 179904
rect 163090 179852 163096 179904
rect 163148 179892 163154 179904
rect 163274 179892 163280 179904
rect 163148 179864 163280 179892
rect 163148 179852 163154 179864
rect 163274 179852 163280 179864
rect 163332 179852 163338 179904
rect 113042 178492 113048 178544
rect 113100 178532 113106 178544
rect 116446 178532 116452 178544
rect 113100 178504 116452 178532
rect 113100 178492 113106 178504
rect 116446 178492 116452 178504
rect 116504 178492 116510 178544
rect 126566 178492 126572 178544
rect 126624 178532 126630 178544
rect 127670 178532 127676 178544
rect 126624 178504 127676 178532
rect 126624 178492 126630 178504
rect 127670 178492 127676 178504
rect 127728 178492 127734 178544
rect 25366 178424 25372 178476
rect 25424 178464 25430 178476
rect 27666 178464 27672 178476
rect 25424 178436 27672 178464
rect 25424 178424 25430 178436
rect 27666 178424 27672 178436
rect 27724 178424 27730 178476
rect 81578 178424 81584 178476
rect 81636 178464 81642 178476
rect 85166 178464 85172 178476
rect 81636 178436 85172 178464
rect 81636 178424 81642 178436
rect 85166 178424 85172 178436
rect 85224 178424 85230 178476
rect 113502 178424 113508 178476
rect 113560 178464 113566 178476
rect 116998 178464 117004 178476
rect 113560 178436 117004 178464
rect 113560 178424 113566 178436
rect 116998 178424 117004 178436
rect 117056 178424 117062 178476
rect 112674 178356 112680 178408
rect 112732 178396 112738 178408
rect 116262 178396 116268 178408
rect 112732 178368 116268 178396
rect 112732 178356 112738 178368
rect 116262 178356 116268 178368
rect 116320 178356 116326 178408
rect 124450 178356 124456 178408
rect 124508 178396 124514 178408
rect 126658 178396 126664 178408
rect 124508 178368 126664 178396
rect 124508 178356 124514 178368
rect 126658 178356 126664 178368
rect 126716 178356 126722 178408
rect 52046 178288 52052 178340
rect 52104 178328 52110 178340
rect 56002 178328 56008 178340
rect 52104 178300 56008 178328
rect 52104 178288 52110 178300
rect 56002 178288 56008 178300
rect 56060 178288 56066 178340
rect 26378 178152 26384 178204
rect 26436 178192 26442 178204
rect 27298 178192 27304 178204
rect 26436 178164 27304 178192
rect 26436 178152 26442 178164
rect 27298 178152 27304 178164
rect 27356 178152 27362 178204
rect 83786 178152 83792 178204
rect 83844 178192 83850 178204
rect 86454 178192 86460 178204
rect 83844 178164 86460 178192
rect 83844 178152 83850 178164
rect 86454 178152 86460 178164
rect 86512 178152 86518 178204
rect 80474 178016 80480 178068
rect 80532 178056 80538 178068
rect 87834 178056 87840 178068
rect 80532 178028 87840 178056
rect 80532 178016 80538 178028
rect 87834 178016 87840 178028
rect 87892 178016 87898 178068
rect 113962 178016 113968 178068
rect 114020 178056 114026 178068
rect 117550 178056 117556 178068
rect 114020 178028 117556 178056
rect 114020 178016 114026 178028
rect 117550 178016 117556 178028
rect 117608 178016 117614 178068
rect 153890 178016 153896 178068
rect 153948 178056 153954 178068
rect 161066 178056 161072 178068
rect 153948 178028 161072 178056
rect 153948 178016 153954 178028
rect 161066 178016 161072 178028
rect 161124 178016 161130 178068
rect 82682 177948 82688 178000
rect 82740 177988 82746 178000
rect 89214 177988 89220 178000
rect 82740 177960 89220 177988
rect 82740 177948 82746 177960
rect 89214 177948 89220 177960
rect 89272 177948 89278 178000
rect 151682 177948 151688 178000
rect 151740 177988 151746 178000
rect 158306 177988 158312 178000
rect 151740 177960 158312 177988
rect 151740 177948 151746 177960
rect 158306 177948 158312 177960
rect 158364 177948 158370 178000
rect 122426 177880 122432 177932
rect 122484 177920 122490 177932
rect 129970 177920 129976 177932
rect 122484 177892 129976 177920
rect 122484 177880 122490 177892
rect 129970 177880 129976 177892
rect 130028 177880 130034 177932
rect 50666 177812 50672 177864
rect 50724 177852 50730 177864
rect 58210 177852 58216 177864
rect 50724 177824 58216 177852
rect 50724 177812 50730 177824
rect 58210 177812 58216 177824
rect 58268 177812 58274 177864
rect 58302 177812 58308 177864
rect 58360 177852 58366 177864
rect 88202 177852 88208 177864
rect 58360 177824 88208 177852
rect 58360 177812 58366 177824
rect 88202 177812 88208 177824
rect 88260 177812 88266 177864
rect 128590 177812 128596 177864
rect 128648 177852 128654 177864
rect 161066 177852 161072 177864
rect 128648 177824 161072 177852
rect 128648 177812 128654 177824
rect 161066 177812 161072 177824
rect 161124 177812 161130 177864
rect 41650 177744 41656 177796
rect 41708 177784 41714 177796
rect 45790 177784 45796 177796
rect 41708 177756 45796 177784
rect 41708 177744 41714 177756
rect 45790 177744 45796 177756
rect 45848 177744 45854 177796
rect 154626 177744 154632 177796
rect 154684 177784 154690 177796
rect 161250 177784 161256 177796
rect 154684 177756 161256 177784
rect 154684 177744 154690 177756
rect 161250 177744 161256 177756
rect 161308 177744 161314 177796
rect 27850 177676 27856 177728
rect 27908 177716 27914 177728
rect 29690 177716 29696 177728
rect 27908 177688 29696 177716
rect 27908 177676 27914 177688
rect 29690 177676 29696 177688
rect 29748 177676 29754 177728
rect 50114 177676 50120 177728
rect 50172 177716 50178 177728
rect 53794 177716 53800 177728
rect 50172 177688 53800 177716
rect 50172 177676 50178 177688
rect 53794 177676 53800 177688
rect 53852 177676 53858 177728
rect 126474 177676 126480 177728
rect 126532 177716 126538 177728
rect 128774 177716 128780 177728
rect 126532 177688 128780 177716
rect 126532 177676 126538 177688
rect 128774 177676 128780 177688
rect 128832 177676 128838 177728
rect 159410 177676 159416 177728
rect 159468 177716 159474 177728
rect 160974 177716 160980 177728
rect 159468 177688 160980 177716
rect 159468 177676 159474 177688
rect 160974 177676 160980 177688
rect 161032 177676 161038 177728
rect 185262 177676 185268 177728
rect 185320 177716 185326 177728
rect 189310 177716 189316 177728
rect 185320 177688 189316 177716
rect 185320 177676 185326 177688
rect 189310 177676 189316 177688
rect 189368 177676 189374 177728
rect 27942 177608 27948 177660
rect 28000 177648 28006 177660
rect 29230 177648 29236 177660
rect 28000 177620 29236 177648
rect 28000 177608 28006 177620
rect 29230 177608 29236 177620
rect 29288 177608 29294 177660
rect 33370 177608 33376 177660
rect 33428 177648 33434 177660
rect 34106 177648 34112 177660
rect 33428 177620 34112 177648
rect 33428 177608 33434 177620
rect 34106 177608 34112 177620
rect 34164 177608 34170 177660
rect 41282 177608 41288 177660
rect 41340 177648 41346 177660
rect 44870 177648 44876 177660
rect 41340 177620 44876 177648
rect 41340 177608 41346 177620
rect 44870 177608 44876 177620
rect 44928 177608 44934 177660
rect 50022 177608 50028 177660
rect 50080 177648 50086 177660
rect 52690 177648 52696 177660
rect 50080 177620 52696 177648
rect 50080 177608 50086 177620
rect 52690 177608 52696 177620
rect 52748 177608 52754 177660
rect 75966 177608 75972 177660
rect 76024 177648 76030 177660
rect 80290 177648 80296 177660
rect 76024 177620 80296 177648
rect 76024 177608 76030 177620
rect 80290 177608 80296 177620
rect 80348 177608 80354 177660
rect 84890 177608 84896 177660
rect 84948 177648 84954 177660
rect 85718 177648 85724 177660
rect 84948 177620 85724 177648
rect 84948 177608 84954 177620
rect 85718 177608 85724 177620
rect 85776 177608 85782 177660
rect 99702 177608 99708 177660
rect 99760 177648 99766 177660
rect 100162 177648 100168 177660
rect 99760 177620 100168 177648
rect 99760 177608 99766 177620
rect 100162 177608 100168 177620
rect 100220 177608 100226 177660
rect 100254 177608 100260 177660
rect 100312 177648 100318 177660
rect 100714 177648 100720 177660
rect 100312 177620 100720 177648
rect 100312 177608 100318 177620
rect 100714 177608 100720 177620
rect 100772 177608 100778 177660
rect 104210 177608 104216 177660
rect 104268 177648 104274 177660
rect 104670 177648 104676 177660
rect 104268 177620 104676 177648
rect 104268 177608 104274 177620
rect 104670 177608 104676 177620
rect 104728 177608 104734 177660
rect 156098 177608 156104 177660
rect 156156 177648 156162 177660
rect 158214 177648 158220 177660
rect 156156 177620 158220 177648
rect 156156 177608 156162 177620
rect 158214 177608 158220 177620
rect 158272 177608 158278 177660
rect 158306 177608 158312 177660
rect 158364 177648 158370 177660
rect 158858 177648 158864 177660
rect 158364 177620 158864 177648
rect 158364 177608 158370 177620
rect 158858 177608 158864 177620
rect 158916 177608 158922 177660
rect 169990 177608 169996 177660
rect 170048 177648 170054 177660
rect 171278 177648 171284 177660
rect 170048 177620 171284 177648
rect 170048 177608 170054 177620
rect 171278 177608 171284 177620
rect 171336 177608 171342 177660
rect 172842 177608 172848 177660
rect 172900 177648 172906 177660
rect 173210 177648 173216 177660
rect 172900 177620 173216 177648
rect 172900 177608 172906 177620
rect 173210 177608 173216 177620
rect 173268 177608 173274 177660
rect 175602 177608 175608 177660
rect 175660 177648 175666 177660
rect 176154 177648 176160 177660
rect 175660 177620 176160 177648
rect 175660 177608 175666 177620
rect 176154 177608 176160 177620
rect 176212 177608 176218 177660
rect 184434 177608 184440 177660
rect 184492 177648 184498 177660
rect 188206 177648 188212 177660
rect 184492 177620 188212 177648
rect 184492 177608 184498 177620
rect 188206 177608 188212 177620
rect 188264 177608 188270 177660
rect 152786 177540 152792 177592
rect 152844 177580 152850 177592
rect 159594 177580 159600 177592
rect 152844 177552 159600 177580
rect 152844 177540 152850 177552
rect 159594 177540 159600 177552
rect 159652 177540 159658 177592
rect 185630 177540 185636 177592
rect 185688 177580 185694 177592
rect 189862 177580 189868 177592
rect 185688 177552 189868 177580
rect 185688 177540 185694 177552
rect 189862 177540 189868 177552
rect 189920 177540 189926 177592
rect 50206 177472 50212 177524
rect 50264 177512 50270 177524
rect 54898 177512 54904 177524
rect 50264 177484 54904 177512
rect 50264 177472 50270 177484
rect 54898 177472 54904 177484
rect 54956 177472 54962 177524
rect 85994 177472 86000 177524
rect 86052 177512 86058 177524
rect 87006 177512 87012 177524
rect 86052 177484 87012 177512
rect 86052 177472 86058 177484
rect 87006 177472 87012 177484
rect 87064 177472 87070 177524
rect 105498 177472 105504 177524
rect 105556 177512 105562 177524
rect 106142 177512 106148 177524
rect 105556 177484 106148 177512
rect 105556 177472 105562 177484
rect 106142 177472 106148 177484
rect 106200 177472 106206 177524
rect 26562 177404 26568 177456
rect 26620 177444 26626 177456
rect 28494 177444 28500 177456
rect 26620 177416 28500 177444
rect 26620 177404 26626 177416
rect 28494 177404 28500 177416
rect 28552 177404 28558 177456
rect 79370 177404 79376 177456
rect 79428 177444 79434 177456
rect 86546 177444 86552 177456
rect 79428 177416 86552 177444
rect 79428 177404 79434 177416
rect 86546 177404 86552 177416
rect 86604 177404 86610 177456
rect 184802 177404 184808 177456
rect 184860 177444 184866 177456
rect 188758 177444 188764 177456
rect 184860 177416 188764 177444
rect 184860 177404 184866 177416
rect 188758 177404 188764 177416
rect 188816 177404 188822 177456
rect 40822 177336 40828 177388
rect 40880 177376 40886 177388
rect 44410 177376 44416 177388
rect 40880 177348 44416 177376
rect 40880 177336 40886 177348
rect 44410 177336 44416 177348
rect 44468 177336 44474 177388
rect 51954 177336 51960 177388
rect 52012 177376 52018 177388
rect 57106 177376 57112 177388
rect 52012 177348 57112 177376
rect 52012 177336 52018 177348
rect 57106 177336 57112 177348
rect 57164 177336 57170 177388
rect 31990 177268 31996 177320
rect 32048 177308 32054 177320
rect 33278 177308 33284 177320
rect 32048 177280 33284 177308
rect 32048 177268 32054 177280
rect 33278 177268 33284 177280
rect 33336 177268 33342 177320
rect 171738 177200 171744 177252
rect 171796 177240 171802 177252
rect 172474 177240 172480 177252
rect 171796 177212 172480 177240
rect 171796 177200 171802 177212
rect 172474 177200 172480 177212
rect 172532 177200 172538 177252
rect 164378 174004 164384 174056
rect 164436 174044 164442 174056
rect 167138 174044 167144 174056
rect 164436 174016 167144 174044
rect 164436 174004 164442 174016
rect 167138 174004 167144 174016
rect 167196 174004 167202 174056
rect 188022 172984 188028 173036
rect 188080 173024 188086 173036
rect 196946 173024 196952 173036
rect 188080 172996 196952 173024
rect 188080 172984 188086 172996
rect 196946 172984 196952 172996
rect 197004 172984 197010 173036
rect 164286 172780 164292 172832
rect 164344 172820 164350 172832
rect 166770 172820 166776 172832
rect 164344 172792 166776 172820
rect 164344 172780 164350 172792
rect 166770 172780 166776 172792
rect 166828 172780 166834 172832
rect 92618 171692 92624 171744
rect 92676 171732 92682 171744
rect 95010 171732 95016 171744
rect 92676 171704 95016 171732
rect 92676 171692 92682 171704
rect 95010 171692 95016 171704
rect 95068 171692 95074 171744
rect 164010 171556 164016 171608
rect 164068 171596 164074 171608
rect 166218 171596 166224 171608
rect 164068 171568 166224 171596
rect 164068 171556 164074 171568
rect 166218 171556 166224 171568
rect 166276 171556 166282 171608
rect 163366 170332 163372 170384
rect 163424 170372 163430 170384
rect 165666 170372 165672 170384
rect 163424 170344 165672 170372
rect 163424 170332 163430 170344
rect 165666 170332 165672 170344
rect 165724 170332 165730 170384
rect 163182 169108 163188 169160
rect 163240 169148 163246 169160
rect 165114 169148 165120 169160
rect 163240 169120 165120 169148
rect 163240 169108 163246 169120
rect 165114 169108 165120 169120
rect 165172 169108 165178 169160
rect 91698 168904 91704 168956
rect 91756 168944 91762 168956
rect 94826 168944 94832 168956
rect 91756 168916 94832 168944
rect 91756 168904 91762 168916
rect 94826 168904 94832 168916
rect 94884 168904 94890 168956
rect 114054 168904 114060 168956
rect 114112 168944 114118 168956
rect 118930 168944 118936 168956
rect 114112 168916 118936 168944
rect 114112 168904 114118 168916
rect 118930 168904 118936 168916
rect 118988 168904 118994 168956
rect 13314 167544 13320 167596
rect 13372 167584 13378 167596
rect 22238 167584 22244 167596
rect 13372 167556 22244 167584
rect 13372 167544 13378 167556
rect 22238 167544 22244 167556
rect 22296 167544 22302 167596
rect 163182 165912 163188 165964
rect 163240 165952 163246 165964
rect 167506 165952 167512 165964
rect 163240 165924 167512 165952
rect 163240 165912 163246 165924
rect 167506 165912 167512 165924
rect 167564 165912 167570 165964
rect 91974 165844 91980 165896
rect 92032 165884 92038 165896
rect 94550 165884 94556 165896
rect 92032 165856 94556 165884
rect 92032 165844 92038 165856
rect 94550 165844 94556 165856
rect 94608 165844 94614 165896
rect 116538 164756 116544 164808
rect 116596 164796 116602 164808
rect 119574 164796 119580 164808
rect 116596 164768 119580 164796
rect 116596 164756 116602 164768
rect 119574 164756 119580 164768
rect 119632 164756 119638 164808
rect 188022 164756 188028 164808
rect 188080 164796 188086 164808
rect 197590 164796 197596 164808
rect 188080 164768 197596 164796
rect 188080 164756 188086 164768
rect 197590 164756 197596 164768
rect 197648 164756 197654 164808
rect 164286 164348 164292 164400
rect 164344 164388 164350 164400
rect 167322 164388 167328 164400
rect 164344 164360 167328 164388
rect 164344 164348 164350 164360
rect 167322 164348 167328 164360
rect 167380 164348 167386 164400
rect 164286 163124 164292 163176
rect 164344 163164 164350 163176
rect 167230 163164 167236 163176
rect 164344 163136 167236 163164
rect 164344 163124 164350 163136
rect 167230 163124 167236 163136
rect 167288 163124 167294 163176
rect 164470 162104 164476 162156
rect 164528 162144 164534 162156
rect 168426 162144 168432 162156
rect 164528 162116 168432 162144
rect 164528 162104 164534 162116
rect 168426 162104 168432 162116
rect 168484 162104 168490 162156
rect 92618 161900 92624 161952
rect 92676 161940 92682 161952
rect 95378 161940 95384 161952
rect 92676 161912 95384 161940
rect 92676 161900 92682 161912
rect 95378 161900 95384 161912
rect 95436 161900 95442 161952
rect 164286 161900 164292 161952
rect 164344 161940 164350 161952
rect 167966 161940 167972 161952
rect 164344 161912 167972 161940
rect 164344 161900 164350 161912
rect 167966 161900 167972 161912
rect 168024 161900 168030 161952
rect 91974 161152 91980 161204
rect 92032 161192 92038 161204
rect 94182 161192 94188 161204
rect 92032 161164 94188 161192
rect 92032 161152 92038 161164
rect 94182 161152 94188 161164
rect 94240 161152 94246 161204
rect 168518 160648 168524 160660
rect 164488 160620 168524 160648
rect 91974 160540 91980 160592
rect 92032 160580 92038 160592
rect 94090 160580 94096 160592
rect 92032 160552 94096 160580
rect 92032 160540 92038 160552
rect 94090 160540 94096 160552
rect 94148 160540 94154 160592
rect 164286 160540 164292 160592
rect 164344 160580 164350 160592
rect 164488 160580 164516 160620
rect 168518 160608 168524 160620
rect 168576 160608 168582 160660
rect 164344 160552 164516 160580
rect 164344 160540 164350 160552
rect 91974 159180 91980 159232
rect 92032 159220 92038 159232
rect 93998 159220 94004 159232
rect 92032 159192 94004 159220
rect 92032 159180 92038 159192
rect 93998 159180 94004 159192
rect 94056 159180 94062 159232
rect 164286 158228 164292 158280
rect 164344 158268 164350 158280
rect 168518 158268 168524 158280
rect 164344 158240 168524 158268
rect 164344 158228 164350 158240
rect 168518 158228 168524 158240
rect 168576 158228 168582 158280
rect 91790 157208 91796 157260
rect 91848 157248 91854 157260
rect 93998 157248 94004 157260
rect 91848 157220 94004 157248
rect 91848 157208 91854 157220
rect 93998 157208 94004 157220
rect 94056 157208 94062 157260
rect 164286 156936 164292 156988
rect 164344 156976 164350 156988
rect 168518 156976 168524 156988
rect 164344 156948 168524 156976
rect 164344 156936 164350 156948
rect 168518 156936 168524 156948
rect 168576 156936 168582 156988
rect 45054 156392 45060 156444
rect 45112 156432 45118 156444
rect 47814 156432 47820 156444
rect 45112 156404 47820 156432
rect 45112 156392 45118 156404
rect 47814 156392 47820 156404
rect 47872 156392 47878 156444
rect 164378 155304 164384 155356
rect 164436 155344 164442 155356
rect 167138 155344 167144 155356
rect 164436 155316 167144 155344
rect 164436 155304 164442 155316
rect 167138 155304 167144 155316
rect 167196 155304 167202 155356
rect 13406 155100 13412 155152
rect 13464 155140 13470 155152
rect 22330 155140 22336 155152
rect 13464 155112 22336 155140
rect 13464 155100 13470 155112
rect 22330 155100 22336 155112
rect 22388 155100 22394 155152
rect 163366 154488 163372 154540
rect 163424 154528 163430 154540
rect 167138 154528 167144 154540
rect 163424 154500 167144 154528
rect 163424 154488 163430 154500
rect 167138 154488 167144 154500
rect 167196 154488 167202 154540
rect 91422 154080 91428 154132
rect 91480 154120 91486 154132
rect 94734 154120 94740 154132
rect 91480 154092 94740 154120
rect 91480 154080 91486 154092
rect 94734 154080 94740 154092
rect 94792 154080 94798 154132
rect 91790 152516 91796 152568
rect 91848 152556 91854 152568
rect 95378 152556 95384 152568
rect 91848 152528 95384 152556
rect 91848 152516 91854 152528
rect 95378 152516 95384 152528
rect 95436 152516 95442 152568
rect 164378 152380 164384 152432
rect 164436 152420 164442 152432
rect 167230 152420 167236 152432
rect 164436 152392 167236 152420
rect 164436 152380 164442 152392
rect 167230 152380 167236 152392
rect 167288 152380 167294 152432
rect 91698 151564 91704 151616
rect 91756 151604 91762 151616
rect 94182 151604 94188 151616
rect 91756 151576 94188 151604
rect 91756 151564 91762 151576
rect 94182 151564 94188 151576
rect 94240 151564 94246 151616
rect 164378 151496 164384 151548
rect 164436 151536 164442 151548
rect 167322 151536 167328 151548
rect 164436 151508 167328 151536
rect 164436 151496 164442 151508
rect 167322 151496 167328 151508
rect 167380 151496 167386 151548
rect 164378 149728 164384 149780
rect 164436 149768 164442 149780
rect 167138 149768 167144 149780
rect 164436 149740 167144 149768
rect 164436 149728 164442 149740
rect 167138 149728 167144 149740
rect 167196 149728 167202 149780
rect 91422 149592 91428 149644
rect 91480 149632 91486 149644
rect 93998 149632 94004 149644
rect 91480 149604 94004 149632
rect 91480 149592 91486 149604
rect 93998 149592 94004 149604
rect 94056 149592 94062 149644
rect 163918 149592 163924 149644
rect 163976 149632 163982 149644
rect 167230 149632 167236 149644
rect 163976 149604 167236 149632
rect 163976 149592 163982 149604
rect 167230 149592 167236 149604
rect 167288 149592 167294 149644
rect 164378 148504 164384 148556
rect 164436 148544 164442 148556
rect 167046 148544 167052 148556
rect 164436 148516 167052 148544
rect 164436 148504 164442 148516
rect 167046 148504 167052 148516
rect 167104 148504 167110 148556
rect 13314 146804 13320 146856
rect 13372 146844 13378 146856
rect 22330 146844 22336 146856
rect 13372 146816 22336 146844
rect 13372 146804 13378 146816
rect 22330 146804 22336 146816
rect 22388 146804 22394 146856
rect 91422 146804 91428 146856
rect 91480 146844 91486 146856
rect 93538 146844 93544 146856
rect 91480 146816 93544 146844
rect 91480 146804 91486 146816
rect 93538 146804 93544 146816
rect 93596 146804 93602 146856
rect 164378 146804 164384 146856
rect 164436 146844 164442 146856
rect 167874 146844 167880 146856
rect 164436 146816 167880 146844
rect 164436 146804 164442 146816
rect 167874 146804 167880 146816
rect 167932 146804 167938 146856
rect 164378 145444 164384 145496
rect 164436 145484 164442 145496
rect 167966 145484 167972 145496
rect 164436 145456 167972 145484
rect 164436 145444 164442 145456
rect 167966 145444 167972 145456
rect 168024 145444 168030 145496
rect 91330 143540 91336 143592
rect 91388 143580 91394 143592
rect 94366 143580 94372 143592
rect 91388 143552 94372 143580
rect 91388 143540 91394 143552
rect 94366 143540 94372 143552
rect 94424 143540 94430 143592
rect 91790 142724 91796 142776
rect 91848 142764 91854 142776
rect 95654 142764 95660 142776
rect 91848 142736 95660 142764
rect 91848 142724 91854 142736
rect 95654 142724 95660 142736
rect 95712 142724 95718 142776
rect 91698 142656 91704 142708
rect 91756 142696 91762 142708
rect 95378 142696 95384 142708
rect 91756 142668 95384 142696
rect 91756 142656 91762 142668
rect 95378 142656 95384 142668
rect 95436 142656 95442 142708
rect 116814 142588 116820 142640
rect 116872 142628 116878 142640
rect 118930 142628 118936 142640
rect 116872 142600 118936 142628
rect 116872 142588 116878 142600
rect 118930 142588 118936 142600
rect 118988 142588 118994 142640
rect 164378 141568 164384 141620
rect 164436 141608 164442 141620
rect 167046 141608 167052 141620
rect 164436 141580 167052 141608
rect 164436 141568 164442 141580
rect 167046 141568 167052 141580
rect 167104 141568 167110 141620
rect 91698 141472 91704 141484
rect 91659 141444 91704 141472
rect 91698 141432 91704 141444
rect 91756 141432 91762 141484
rect 91790 141296 91796 141348
rect 91848 141336 91854 141348
rect 95010 141336 95016 141348
rect 91848 141308 95016 141336
rect 91848 141296 91854 141308
rect 95010 141296 95016 141308
rect 95068 141296 95074 141348
rect 92526 140004 92532 140056
rect 92584 140044 92590 140056
rect 93446 140044 93452 140056
rect 92584 140016 93452 140044
rect 92584 140004 92590 140016
rect 93446 140004 93452 140016
rect 93504 140004 93510 140056
rect 164286 140004 164292 140056
rect 164344 140044 164350 140056
rect 166402 140044 166408 140056
rect 164344 140016 166408 140044
rect 164344 140004 164350 140016
rect 166402 140004 166408 140016
rect 166460 140004 166466 140056
rect 92618 139936 92624 139988
rect 92676 139976 92682 139988
rect 93906 139976 93912 139988
rect 92676 139948 93912 139976
rect 92676 139936 92682 139948
rect 93906 139936 93912 139948
rect 93964 139936 93970 139988
rect 164378 139936 164384 139988
rect 164436 139976 164442 139988
rect 165850 139976 165856 139988
rect 164436 139948 165856 139976
rect 164436 139936 164442 139948
rect 165850 139936 165856 139948
rect 165908 139936 165914 139988
rect 188022 139188 188028 139240
rect 188080 139228 188086 139240
rect 192070 139228 192076 139240
rect 188080 139200 192076 139228
rect 188080 139188 188086 139200
rect 192070 139188 192076 139200
rect 192128 139228 192134 139240
rect 193450 139228 193456 139240
rect 192128 139200 193456 139228
rect 192128 139188 192134 139200
rect 193450 139188 193456 139200
rect 193508 139188 193514 139240
rect 48458 134700 48464 134752
rect 48516 134740 48522 134752
rect 78085 134743 78143 134749
rect 78085 134740 78097 134743
rect 48516 134712 78097 134740
rect 48516 134700 48522 134712
rect 78085 134709 78097 134712
rect 78131 134709 78143 134743
rect 78085 134703 78143 134709
rect 74681 134403 74739 134409
rect 74681 134369 74693 134403
rect 74727 134400 74739 134403
rect 82130 134400 82136 134412
rect 74727 134372 82136 134400
rect 74727 134369 74739 134372
rect 74681 134363 74739 134369
rect 82130 134360 82136 134372
rect 82188 134360 82194 134412
rect 84338 134360 84344 134412
rect 84396 134400 84402 134412
rect 145150 134400 145156 134412
rect 84396 134372 145156 134400
rect 84396 134360 84402 134372
rect 145150 134360 145156 134372
rect 145208 134360 145214 134412
rect 116173 134335 116231 134341
rect 116173 134332 116185 134335
rect 89968 134304 116185 134332
rect 23618 134224 23624 134276
rect 23676 134264 23682 134276
rect 27666 134264 27672 134276
rect 23676 134236 27672 134264
rect 23676 134224 23682 134236
rect 27666 134224 27672 134236
rect 27724 134224 27730 134276
rect 73206 134224 73212 134276
rect 73264 134264 73270 134276
rect 83602 134264 83608 134276
rect 73264 134236 83608 134264
rect 73264 134224 73270 134236
rect 83602 134224 83608 134236
rect 83660 134264 83666 134276
rect 84338 134264 84344 134276
rect 83660 134236 84344 134264
rect 83660 134224 83666 134236
rect 84338 134224 84344 134236
rect 84396 134224 84402 134276
rect 66582 134156 66588 134208
rect 66640 134196 66646 134208
rect 74681 134199 74739 134205
rect 74681 134196 74693 134199
rect 66640 134168 74693 134196
rect 66640 134156 66646 134168
rect 74681 134165 74693 134168
rect 74727 134165 74739 134199
rect 89968 134196 89996 134304
rect 116173 134301 116185 134304
rect 116219 134301 116231 134335
rect 116173 134295 116231 134301
rect 125741 134267 125799 134273
rect 125741 134233 125753 134267
rect 125787 134264 125799 134267
rect 128501 134267 128559 134273
rect 128501 134264 128513 134267
rect 125787 134236 128513 134264
rect 125787 134233 125799 134236
rect 125741 134227 125799 134233
rect 128501 134233 128513 134236
rect 128547 134233 128559 134267
rect 128501 134227 128559 134233
rect 74681 134159 74739 134165
rect 89784 134168 89996 134196
rect 128593 134199 128651 134205
rect 82130 134088 82136 134140
rect 82188 134128 82194 134140
rect 89784 134128 89812 134168
rect 128593 134165 128605 134199
rect 128639 134196 128651 134199
rect 138250 134196 138256 134208
rect 128639 134168 138256 134196
rect 128639 134165 128651 134168
rect 128593 134159 128651 134165
rect 138250 134156 138256 134168
rect 138308 134156 138314 134208
rect 82188 134100 89812 134128
rect 116173 134131 116231 134137
rect 82188 134088 82194 134100
rect 116173 134097 116185 134131
rect 116219 134128 116231 134131
rect 125741 134131 125799 134137
rect 125741 134128 125753 134131
rect 116219 134100 125753 134128
rect 116219 134097 116231 134100
rect 116173 134091 116231 134097
rect 125741 134097 125753 134100
rect 125787 134097 125799 134131
rect 125741 134091 125799 134097
rect 182410 134020 182416 134072
rect 182468 134060 182474 134072
rect 186366 134060 186372 134072
rect 182468 134032 186372 134060
rect 182468 134020 182474 134032
rect 186366 134020 186372 134032
rect 186424 134020 186430 134072
rect 27022 133952 27028 134004
rect 27080 133992 27086 134004
rect 29690 133992 29696 134004
rect 27080 133964 29696 133992
rect 27080 133952 27086 133964
rect 29690 133952 29696 133964
rect 29748 133952 29754 134004
rect 38430 133952 38436 134004
rect 38488 133992 38494 134004
rect 41558 133992 41564 134004
rect 38488 133964 41564 133992
rect 38488 133952 38494 133964
rect 41558 133952 41564 133964
rect 41616 133952 41622 134004
rect 114054 133992 114060 134004
rect 104412 133964 114060 133992
rect 26286 133884 26292 133936
rect 26344 133924 26350 133936
rect 29230 133924 29236 133936
rect 26344 133896 29236 133924
rect 26344 133884 26350 133896
rect 29230 133884 29236 133896
rect 29288 133884 29294 133936
rect 37694 133884 37700 133936
rect 37752 133924 37758 133936
rect 40638 133924 40644 133936
rect 37752 133896 40644 133924
rect 37752 133884 37758 133896
rect 40638 133884 40644 133896
rect 40696 133884 40702 133936
rect 28310 133816 28316 133868
rect 28368 133856 28374 133868
rect 30426 133856 30432 133868
rect 28368 133828 30432 133856
rect 28368 133816 28374 133828
rect 30426 133816 30432 133828
rect 30484 133816 30490 133868
rect 31070 133816 31076 133868
rect 31128 133856 31134 133868
rect 32082 133856 32088 133868
rect 31128 133828 32088 133856
rect 31128 133816 31134 133828
rect 32082 133816 32088 133828
rect 32140 133816 32146 133868
rect 37234 133816 37240 133868
rect 37292 133856 37298 133868
rect 39994 133856 40000 133868
rect 37292 133828 40000 133856
rect 37292 133816 37298 133828
rect 39994 133816 40000 133828
rect 40052 133816 40058 133868
rect 40822 133816 40828 133868
rect 40880 133856 40886 133868
rect 43582 133856 43588 133868
rect 40880 133828 43588 133856
rect 40880 133816 40886 133828
rect 43582 133816 43588 133828
rect 43640 133816 43646 133868
rect 29690 133748 29696 133800
rect 29748 133788 29754 133800
rect 31254 133788 31260 133800
rect 29748 133760 31260 133788
rect 29748 133748 29754 133760
rect 31254 133748 31260 133760
rect 31312 133748 31318 133800
rect 34842 133748 34848 133800
rect 34900 133788 34906 133800
rect 35854 133788 35860 133800
rect 34900 133760 35860 133788
rect 34900 133748 34906 133760
rect 35854 133748 35860 133760
rect 35912 133748 35918 133800
rect 36498 133748 36504 133800
rect 36556 133788 36562 133800
rect 38614 133788 38620 133800
rect 36556 133760 38620 133788
rect 36556 133748 36562 133760
rect 38614 133748 38620 133760
rect 38672 133748 38678 133800
rect 41282 133748 41288 133800
rect 41340 133788 41346 133800
rect 44318 133788 44324 133800
rect 41340 133760 44324 133788
rect 41340 133748 41346 133760
rect 44318 133748 44324 133760
rect 44376 133748 44382 133800
rect 27666 133680 27672 133732
rect 27724 133720 27730 133732
rect 30058 133720 30064 133732
rect 27724 133692 30064 133720
rect 27724 133680 27730 133692
rect 30058 133680 30064 133692
rect 30116 133680 30122 133732
rect 40454 133680 40460 133732
rect 40512 133720 40518 133732
rect 43030 133720 43036 133732
rect 40512 133692 43036 133720
rect 40512 133680 40518 133692
rect 43030 133680 43036 133692
rect 43088 133680 43094 133732
rect 62350 133680 62356 133732
rect 62408 133720 62414 133732
rect 86546 133720 86552 133732
rect 62408 133692 86552 133720
rect 62408 133680 62414 133692
rect 86546 133680 86552 133692
rect 86604 133680 86610 133732
rect 38062 133612 38068 133664
rect 38120 133652 38126 133664
rect 41006 133652 41012 133664
rect 38120 133624 41012 133652
rect 38120 133612 38126 133624
rect 41006 133612 41012 133624
rect 41064 133612 41070 133664
rect 91425 133655 91483 133661
rect 91425 133621 91437 133655
rect 91471 133652 91483 133655
rect 104412 133652 104440 133964
rect 114054 133952 114060 133964
rect 114112 133952 114118 134004
rect 182870 133952 182876 134004
rect 182928 133992 182934 134004
rect 186458 133992 186464 134004
rect 182928 133964 186464 133992
rect 182928 133952 182934 133964
rect 186458 133952 186464 133964
rect 186516 133952 186522 134004
rect 107522 133884 107528 133936
rect 107580 133924 107586 133936
rect 110190 133924 110196 133936
rect 107580 133896 110196 133924
rect 107580 133884 107586 133896
rect 110190 133884 110196 133896
rect 110248 133884 110254 133936
rect 169254 133884 169260 133936
rect 169312 133924 169318 133936
rect 170450 133924 170456 133936
rect 169312 133896 170456 133924
rect 169312 133884 169318 133896
rect 170450 133884 170456 133896
rect 170508 133884 170514 133936
rect 178454 133884 178460 133936
rect 178512 133924 178518 133936
rect 180662 133924 180668 133936
rect 178512 133896 180668 133924
rect 178512 133884 178518 133896
rect 180662 133884 180668 133896
rect 180720 133884 180726 133936
rect 181214 133884 181220 133936
rect 181272 133924 181278 133936
rect 184710 133924 184716 133936
rect 181272 133896 184716 133924
rect 181272 133884 181278 133896
rect 184710 133884 184716 133896
rect 184768 133884 184774 133936
rect 169898 133816 169904 133868
rect 169956 133856 169962 133868
rect 170818 133856 170824 133868
rect 169956 133828 170824 133856
rect 169956 133816 169962 133828
rect 170818 133816 170824 133828
rect 170876 133816 170882 133868
rect 175602 133816 175608 133868
rect 175660 133856 175666 133868
rect 176706 133856 176712 133868
rect 175660 133828 176712 133856
rect 175660 133816 175666 133828
rect 176706 133816 176712 133828
rect 176764 133816 176770 133868
rect 177258 133816 177264 133868
rect 177316 133856 177322 133868
rect 179006 133856 179012 133868
rect 177316 133828 179012 133856
rect 177316 133816 177322 133828
rect 179006 133816 179012 133828
rect 179064 133816 179070 133868
rect 184434 133816 184440 133868
rect 184492 133856 184498 133868
rect 186826 133856 186832 133868
rect 184492 133828 186832 133856
rect 184492 133816 184498 133828
rect 186826 133816 186832 133828
rect 186884 133816 186890 133868
rect 108994 133748 109000 133800
rect 109052 133788 109058 133800
rect 110834 133788 110840 133800
rect 109052 133760 110840 133788
rect 109052 133748 109058 133760
rect 110834 133748 110840 133760
rect 110892 133748 110898 133800
rect 113962 133748 113968 133800
rect 114020 133788 114026 133800
rect 119482 133788 119488 133800
rect 114020 133760 119488 133788
rect 114020 133748 114026 133760
rect 119482 133748 119488 133760
rect 119540 133748 119546 133800
rect 168702 133748 168708 133800
rect 168760 133788 168766 133800
rect 170082 133788 170088 133800
rect 168760 133760 170088 133788
rect 168760 133748 168766 133760
rect 170082 133748 170088 133760
rect 170140 133748 170146 133800
rect 170450 133748 170456 133800
rect 170508 133788 170514 133800
rect 171278 133788 171284 133800
rect 170508 133760 171284 133788
rect 170508 133748 170514 133760
rect 171278 133748 171284 133760
rect 171336 133748 171342 133800
rect 175234 133748 175240 133800
rect 175292 133788 175298 133800
rect 176154 133788 176160 133800
rect 175292 133760 176160 133788
rect 175292 133748 175298 133760
rect 176154 133748 176160 133760
rect 176212 133748 176218 133800
rect 176430 133748 176436 133800
rect 176488 133788 176494 133800
rect 177810 133788 177816 133800
rect 176488 133760 177816 133788
rect 176488 133748 176494 133760
rect 177810 133748 177816 133760
rect 177868 133748 177874 133800
rect 183606 133748 183612 133800
rect 183664 133788 183670 133800
rect 185538 133788 185544 133800
rect 183664 133760 185544 133788
rect 183664 133748 183670 133760
rect 185538 133748 185544 133760
rect 185596 133748 185602 133800
rect 110282 133680 110288 133732
rect 110340 133720 110346 133732
rect 113226 133720 113232 133732
rect 110340 133692 113232 133720
rect 110340 133680 110346 133692
rect 113226 133680 113232 133692
rect 113284 133680 113290 133732
rect 113318 133680 113324 133732
rect 113376 133720 113382 133732
rect 118930 133720 118936 133732
rect 113376 133692 118936 133720
rect 113376 133680 113382 133692
rect 118930 133680 118936 133692
rect 118988 133680 118994 133732
rect 174866 133680 174872 133732
rect 174924 133720 174930 133732
rect 175602 133720 175608 133732
rect 174924 133692 175608 133720
rect 174924 133680 174930 133692
rect 175602 133680 175608 133692
rect 175660 133680 175666 133732
rect 176798 133680 176804 133732
rect 176856 133720 176862 133732
rect 178454 133720 178460 133732
rect 176856 133692 178460 133720
rect 176856 133680 176862 133692
rect 178454 133680 178460 133692
rect 178512 133680 178518 133732
rect 184066 133680 184072 133732
rect 184124 133720 184130 133732
rect 186642 133720 186648 133732
rect 184124 133692 186648 133720
rect 184124 133680 184130 133692
rect 186642 133680 186648 133692
rect 186700 133680 186706 133732
rect 91471 133624 104440 133652
rect 91471 133621 91483 133624
rect 91425 133615 91483 133621
rect 108350 133612 108356 133664
rect 108408 133652 108414 133664
rect 111386 133652 111392 133664
rect 108408 133624 111392 133652
rect 108408 133612 108414 133624
rect 111386 133612 111392 133624
rect 111444 133612 111450 133664
rect 181674 133612 181680 133664
rect 181732 133652 181738 133664
rect 185078 133652 185084 133664
rect 181732 133624 185084 133652
rect 181732 133612 181738 133624
rect 185078 133612 185084 133624
rect 185136 133612 185142 133664
rect 39258 133544 39264 133596
rect 39316 133584 39322 133596
rect 42938 133584 42944 133596
rect 39316 133556 42944 133584
rect 39316 133544 39322 133556
rect 42938 133544 42944 133556
rect 42996 133544 43002 133596
rect 109914 133544 109920 133596
rect 109972 133584 109978 133596
rect 113318 133584 113324 133596
rect 109972 133556 113324 133584
rect 109972 133544 109978 133556
rect 113318 133544 113324 133556
rect 113376 133544 113382 133596
rect 149658 133544 149664 133596
rect 149716 133584 149722 133596
rect 151590 133584 151596 133596
rect 149716 133556 151596 133584
rect 149716 133544 149722 133556
rect 151590 133544 151596 133556
rect 151648 133544 151654 133596
rect 184802 133544 184808 133596
rect 184860 133584 184866 133596
rect 187286 133584 187292 133596
rect 184860 133556 187292 133584
rect 184860 133544 184866 133556
rect 187286 133544 187292 133556
rect 187344 133544 187350 133596
rect 39626 133476 39632 133528
rect 39684 133516 39690 133528
rect 41834 133516 41840 133528
rect 39684 133488 41840 133516
rect 39684 133476 39690 133488
rect 41834 133476 41840 133488
rect 41892 133476 41898 133528
rect 108718 133476 108724 133528
rect 108776 133516 108782 133528
rect 111938 133516 111944 133528
rect 108776 133488 111944 133516
rect 108776 133476 108782 133488
rect 111938 133476 111944 133488
rect 111996 133476 112002 133528
rect 177626 133476 177632 133528
rect 177684 133516 177690 133528
rect 179558 133516 179564 133528
rect 177684 133488 179564 133516
rect 177684 133476 177690 133488
rect 179558 133476 179564 133488
rect 179616 133476 179622 133528
rect 180846 133476 180852 133528
rect 180904 133516 180910 133528
rect 182502 133516 182508 133528
rect 180904 133488 182508 133516
rect 180904 133476 180910 133488
rect 182502 133476 182508 133488
rect 182560 133476 182566 133528
rect 29046 133408 29052 133460
rect 29104 133448 29110 133460
rect 30886 133448 30892 133460
rect 29104 133420 30892 133448
rect 29104 133408 29110 133420
rect 30886 133408 30892 133420
rect 30944 133408 30950 133460
rect 34474 133408 34480 133460
rect 34532 133448 34538 133460
rect 35210 133448 35216 133460
rect 34532 133420 35216 133448
rect 34532 133408 34538 133420
rect 35210 133408 35216 133420
rect 35268 133408 35274 133460
rect 36866 133408 36872 133460
rect 36924 133448 36930 133460
rect 39258 133448 39264 133460
rect 36924 133420 39264 133448
rect 36924 133408 36930 133420
rect 39258 133408 39264 133420
rect 39316 133408 39322 133460
rect 40086 133408 40092 133460
rect 40144 133448 40150 133460
rect 42294 133448 42300 133460
rect 40144 133420 42300 133448
rect 40144 133408 40150 133420
rect 42294 133408 42300 133420
rect 42352 133408 42358 133460
rect 107154 133408 107160 133460
rect 107212 133448 107218 133460
rect 109638 133448 109644 133460
rect 107212 133420 109644 133448
rect 107212 133408 107218 133420
rect 109638 133408 109644 133420
rect 109696 133408 109702 133460
rect 183238 133408 183244 133460
rect 183296 133448 183302 133460
rect 185722 133448 185728 133460
rect 183296 133420 185728 133448
rect 183296 133408 183302 133420
rect 185722 133408 185728 133420
rect 185780 133408 185786 133460
rect 24998 133340 25004 133392
rect 25056 133380 25062 133392
rect 26102 133380 26108 133392
rect 25056 133352 26108 133380
rect 25056 133340 25062 133352
rect 26102 133340 26108 133352
rect 26160 133340 26166 133392
rect 38890 133340 38896 133392
rect 38948 133380 38954 133392
rect 42662 133380 42668 133392
rect 38948 133352 42668 133380
rect 38948 133340 38954 133352
rect 42662 133340 42668 133352
rect 42720 133340 42726 133392
rect 107798 133340 107804 133392
rect 107856 133380 107862 133392
rect 110558 133380 110564 133392
rect 107856 133352 110564 133380
rect 107856 133340 107862 133352
rect 110558 133340 110564 133352
rect 110616 133340 110622 133392
rect 111478 133340 111484 133392
rect 111536 133380 111542 133392
rect 114422 133380 114428 133392
rect 111536 133352 114428 133380
rect 111536 133340 111542 133352
rect 114422 133340 114428 133352
rect 114480 133340 114486 133392
rect 180018 133340 180024 133392
rect 180076 133380 180082 133392
rect 182962 133380 182968 133392
rect 180076 133352 182968 133380
rect 180076 133340 180082 133352
rect 182962 133340 182968 133352
rect 183020 133340 183026 133392
rect 30426 133272 30432 133324
rect 30484 133312 30490 133324
rect 31622 133312 31628 133324
rect 30484 133284 31628 133312
rect 30484 133272 30490 133284
rect 31622 133272 31628 133284
rect 31680 133272 31686 133324
rect 106694 133272 106700 133324
rect 106752 133312 106758 133324
rect 108994 133312 109000 133324
rect 106752 133284 109000 133312
rect 106752 133272 106758 133284
rect 108994 133272 109000 133284
rect 109052 133272 109058 133324
rect 111110 133272 111116 133324
rect 111168 133312 111174 133324
rect 113410 133312 113416 133324
rect 111168 133284 113416 133312
rect 111168 133272 111174 133284
rect 113410 133272 113416 133284
rect 113468 133272 113474 133324
rect 176062 133272 176068 133324
rect 176120 133312 176126 133324
rect 177258 133312 177264 133324
rect 176120 133284 177264 133312
rect 176120 133272 176126 133284
rect 177258 133272 177264 133284
rect 177316 133272 177322 133324
rect 178086 133272 178092 133324
rect 178144 133312 178150 133324
rect 180110 133312 180116 133324
rect 178144 133284 180116 133312
rect 178144 133272 178150 133284
rect 180110 133272 180116 133284
rect 180168 133272 180174 133324
rect 182042 133272 182048 133324
rect 182100 133312 182106 133324
rect 184802 133312 184808 133324
rect 182100 133284 184808 133312
rect 182100 133272 182106 133284
rect 184802 133272 184808 133284
rect 184860 133272 184866 133324
rect 24906 133204 24912 133256
rect 24964 133244 24970 133256
rect 28494 133244 28500 133256
rect 24964 133216 28500 133244
rect 24964 133204 24970 133216
rect 28494 133204 28500 133216
rect 28552 133204 28558 133256
rect 105498 133204 105504 133256
rect 105556 133244 105562 133256
rect 107246 133244 107252 133256
rect 105556 133216 107252 133244
rect 105556 133204 105562 133216
rect 107246 133204 107252 133216
rect 107304 133204 107310 133256
rect 111846 133204 111852 133256
rect 111904 133244 111910 133256
rect 114698 133244 114704 133256
rect 111904 133216 114704 133244
rect 111904 133204 111910 133216
rect 114698 133204 114704 133216
rect 114756 133204 114762 133256
rect 179282 133204 179288 133256
rect 179340 133244 179346 133256
rect 181858 133244 181864 133256
rect 179340 133216 181864 133244
rect 179340 133204 179346 133216
rect 181858 133204 181864 133216
rect 181916 133204 181922 133256
rect 185262 133204 185268 133256
rect 185320 133244 185326 133256
rect 190414 133244 190420 133256
rect 185320 133216 190420 133244
rect 185320 133204 185326 133216
rect 190414 133204 190420 133216
rect 190472 133204 190478 133256
rect 24262 133136 24268 133188
rect 24320 133176 24326 133188
rect 28034 133176 28040 133188
rect 24320 133148 28040 133176
rect 24320 133136 24326 133148
rect 28034 133136 28040 133148
rect 28092 133136 28098 133188
rect 35670 133136 35676 133188
rect 35728 133176 35734 133188
rect 37234 133176 37240 133188
rect 35728 133148 37240 133176
rect 35728 133136 35734 133148
rect 37234 133136 37240 133148
rect 37292 133136 37298 133188
rect 103566 133136 103572 133188
rect 103624 133176 103630 133188
rect 104946 133176 104952 133188
rect 103624 133148 104952 133176
rect 103624 133136 103630 133148
rect 104946 133136 104952 133148
rect 105004 133136 105010 133188
rect 105038 133136 105044 133188
rect 105096 133176 105102 133188
rect 106694 133176 106700 133188
rect 105096 133148 106700 133176
rect 105096 133136 105102 133148
rect 106694 133136 106700 133148
rect 106752 133136 106758 133188
rect 110466 133136 110472 133188
rect 110524 133176 110530 133188
rect 112582 133176 112588 133188
rect 110524 133148 112588 133176
rect 110524 133136 110530 133148
rect 112582 133136 112588 133148
rect 112640 133136 112646 133188
rect 112674 133136 112680 133188
rect 112732 133176 112738 133188
rect 116078 133176 116084 133188
rect 112732 133148 116084 133176
rect 112732 133136 112738 133148
rect 116078 133136 116084 133148
rect 116136 133136 116142 133188
rect 178822 133136 178828 133188
rect 178880 133176 178886 133188
rect 181306 133176 181312 133188
rect 178880 133148 181312 133176
rect 178880 133136 178886 133148
rect 181306 133136 181312 133148
rect 181364 133136 181370 133188
rect 25642 133068 25648 133120
rect 25700 133108 25706 133120
rect 28862 133108 28868 133120
rect 25700 133080 28868 133108
rect 25700 133068 25706 133080
rect 28862 133068 28868 133080
rect 28920 133068 28926 133120
rect 35302 133068 35308 133120
rect 35360 133108 35366 133120
rect 36498 133108 36504 133120
rect 35360 133080 36504 133108
rect 35360 133068 35366 133080
rect 36498 133068 36504 133080
rect 36556 133068 36562 133120
rect 41650 133068 41656 133120
rect 41708 133108 41714 133120
rect 47446 133108 47452 133120
rect 41708 133080 47452 133108
rect 41708 133068 41714 133080
rect 47446 133068 47452 133080
rect 47504 133068 47510 133120
rect 96758 133068 96764 133120
rect 96816 133108 96822 133120
rect 97770 133108 97776 133120
rect 96816 133080 97776 133108
rect 96816 133068 96822 133080
rect 97770 133068 97776 133080
rect 97828 133068 97834 133120
rect 97954 133068 97960 133120
rect 98012 133108 98018 133120
rect 98598 133108 98604 133120
rect 98012 133080 98604 133108
rect 98012 133068 98018 133080
rect 98598 133068 98604 133080
rect 98656 133068 98662 133120
rect 103474 133068 103480 133120
rect 103532 133108 103538 133120
rect 104394 133108 104400 133120
rect 103532 133080 104400 133108
rect 103532 133068 103538 133080
rect 104394 133068 104400 133080
rect 104452 133068 104458 133120
rect 104670 133068 104676 133120
rect 104728 133108 104734 133120
rect 106142 133108 106148 133120
rect 104728 133080 106148 133108
rect 104728 133068 104734 133080
rect 106142 133068 106148 133080
rect 106200 133068 106206 133120
rect 106326 133068 106332 133120
rect 106384 133108 106390 133120
rect 108442 133108 108448 133120
rect 106384 133080 108448 133108
rect 106384 133068 106390 133080
rect 108442 133068 108448 133080
rect 108500 133068 108506 133120
rect 112306 133068 112312 133120
rect 112364 133108 112370 133120
rect 114790 133108 114796 133120
rect 112364 133080 114796 133108
rect 112364 133068 112370 133080
rect 114790 133068 114796 133080
rect 114848 133068 114854 133120
rect 180478 133068 180484 133120
rect 180536 133108 180542 133120
rect 183514 133108 183520 133120
rect 180536 133080 183520 133108
rect 180536 133068 180542 133080
rect 183514 133068 183520 133080
rect 183572 133068 183578 133120
rect 22882 133000 22888 133052
rect 22940 133040 22946 133052
rect 27298 133040 27304 133052
rect 22940 133012 27304 133040
rect 22940 133000 22946 133012
rect 27298 133000 27304 133012
rect 27356 133000 27362 133052
rect 36038 133000 36044 133052
rect 36096 133040 36102 133052
rect 37878 133040 37884 133052
rect 36096 133012 37884 133040
rect 36096 133000 36102 133012
rect 37878 133000 37884 133012
rect 37936 133000 37942 133052
rect 97402 133000 97408 133052
rect 97460 133040 97466 133052
rect 98230 133040 98236 133052
rect 97460 133012 98236 133040
rect 97460 133000 97466 133012
rect 98230 133000 98236 133012
rect 98288 133000 98294 133052
rect 103106 133000 103112 133052
rect 103164 133040 103170 133052
rect 103750 133040 103756 133052
rect 103164 133012 103756 133040
rect 103164 133000 103170 133012
rect 103750 133000 103756 133012
rect 103808 133000 103814 133052
rect 104302 133000 104308 133052
rect 104360 133040 104366 133052
rect 105498 133040 105504 133052
rect 104360 133012 105504 133040
rect 104360 133000 104366 133012
rect 105498 133000 105504 133012
rect 105556 133000 105562 133052
rect 105958 133000 105964 133052
rect 106016 133040 106022 133052
rect 107890 133040 107896 133052
rect 106016 133012 107896 133040
rect 106016 133000 106022 133012
rect 107890 133000 107896 133012
rect 107948 133000 107954 133052
rect 109546 133000 109552 133052
rect 109604 133040 109610 133052
rect 112766 133040 112772 133052
rect 109604 133012 112772 133040
rect 109604 133000 109610 133012
rect 112766 133000 112772 133012
rect 112824 133000 112830 133052
rect 113134 133000 113140 133052
rect 113192 133040 113198 133052
rect 115710 133040 115716 133052
rect 113192 133012 115716 133040
rect 113192 133000 113198 133012
rect 115710 133000 115716 133012
rect 115768 133000 115774 133052
rect 179650 133000 179656 133052
rect 179708 133040 179714 133052
rect 182410 133040 182416 133052
rect 179708 133012 182416 133040
rect 179708 133000 179714 133012
rect 182410 133000 182416 133012
rect 182468 133000 182474 133052
rect 185630 133000 185636 133052
rect 185688 133040 185694 133052
rect 190966 133040 190972 133052
rect 185688 133012 190972 133040
rect 185688 133000 185694 133012
rect 190966 133000 190972 133012
rect 191024 133000 191030 133052
rect 92066 131572 92072 131624
rect 92124 131612 92130 131624
rect 92710 131612 92716 131624
rect 92124 131584 92716 131612
rect 92124 131572 92130 131584
rect 92710 131572 92716 131584
rect 92768 131572 92774 131624
rect 93446 131572 93452 131624
rect 93504 131612 93510 131624
rect 94458 131612 94464 131624
rect 93504 131584 94464 131612
rect 93504 131572 93510 131584
rect 94458 131572 94464 131584
rect 94516 131572 94522 131624
rect 110834 131572 110840 131624
rect 110892 131612 110898 131624
rect 112490 131612 112496 131624
rect 110892 131584 112496 131612
rect 110892 131572 110898 131584
rect 112490 131572 112496 131584
rect 112548 131572 112554 131624
rect 116078 131572 116084 131624
rect 116136 131612 116142 131624
rect 117734 131612 117740 131624
rect 116136 131584 117740 131612
rect 116136 131572 116142 131584
rect 117734 131572 117740 131584
rect 117792 131572 117798 131624
rect 114422 131504 114428 131556
rect 114480 131544 114486 131556
rect 115986 131544 115992 131556
rect 114480 131516 115992 131544
rect 114480 131504 114486 131516
rect 115986 131504 115992 131516
rect 116044 131504 116050 131556
rect 21502 131368 21508 131420
rect 21560 131408 21566 131420
rect 26470 131408 26476 131420
rect 21560 131380 26476 131408
rect 21560 131368 21566 131380
rect 26470 131368 26476 131380
rect 26528 131368 26534 131420
rect 43582 131368 43588 131420
rect 43640 131408 43646 131420
rect 46066 131408 46072 131420
rect 43640 131380 46072 131408
rect 43640 131368 43646 131380
rect 46066 131368 46072 131380
rect 46124 131368 46130 131420
rect 114698 131368 114704 131420
rect 114756 131408 114762 131420
rect 116630 131408 116636 131420
rect 114756 131380 116636 131408
rect 114756 131368 114762 131380
rect 116630 131368 116636 131380
rect 116688 131368 116694 131420
rect 22238 131232 22244 131284
rect 22296 131272 22302 131284
rect 26838 131272 26844 131284
rect 22296 131244 26844 131272
rect 22296 131232 22302 131244
rect 26838 131232 26844 131244
rect 26896 131232 26902 131284
rect 113226 131232 113232 131284
rect 113284 131272 113290 131284
rect 114238 131272 114244 131284
rect 113284 131244 114244 131272
rect 113284 131232 113290 131244
rect 114238 131232 114244 131244
rect 114296 131232 114302 131284
rect 114790 131232 114796 131284
rect 114848 131272 114854 131284
rect 117182 131272 117188 131284
rect 114848 131244 117188 131272
rect 114848 131232 114854 131244
rect 117182 131232 117188 131244
rect 117240 131232 117246 131284
rect 44318 131096 44324 131148
rect 44376 131136 44382 131148
rect 46802 131136 46808 131148
rect 44376 131108 46808 131136
rect 44376 131096 44382 131108
rect 46802 131096 46808 131108
rect 46860 131096 46866 131148
rect 91974 131096 91980 131148
rect 92032 131136 92038 131148
rect 96206 131136 96212 131148
rect 92032 131108 96212 131136
rect 92032 131096 92038 131108
rect 96206 131096 96212 131108
rect 96264 131096 96270 131148
rect 113410 131096 113416 131148
rect 113468 131136 113474 131148
rect 115434 131136 115440 131148
rect 113468 131108 115440 131136
rect 113468 131096 113474 131108
rect 115434 131096 115440 131108
rect 115492 131096 115498 131148
rect 115710 130960 115716 131012
rect 115768 131000 115774 131012
rect 118378 131000 118384 131012
rect 115768 130972 118384 131000
rect 115768 130960 115774 130972
rect 118378 130960 118384 130972
rect 118436 130960 118442 131012
rect 20214 130892 20220 130944
rect 20272 130932 20278 130944
rect 44410 130932 44416 130944
rect 20272 130904 44416 130932
rect 20272 130892 20278 130904
rect 44410 130892 44416 130904
rect 44468 130892 44474 130944
rect 168518 130892 168524 130944
rect 168576 130932 168582 130944
rect 191518 130932 191524 130944
rect 168576 130904 191524 130932
rect 168576 130892 168582 130904
rect 191518 130892 191524 130904
rect 191576 130892 191582 130944
rect 112582 130688 112588 130740
rect 112640 130728 112646 130740
rect 114882 130728 114888 130740
rect 112640 130700 114888 130728
rect 112640 130688 112646 130700
rect 114882 130688 114888 130700
rect 114940 130688 114946 130740
rect 185630 130552 185636 130604
rect 185688 130592 185694 130604
rect 188114 130592 188120 130604
rect 185688 130564 188120 130592
rect 185688 130552 185694 130564
rect 188114 130552 188120 130564
rect 188172 130552 188178 130604
rect 185722 130484 185728 130536
rect 185780 130524 185786 130536
rect 187562 130524 187568 130536
rect 185780 130496 187568 130524
rect 185780 130484 185786 130496
rect 187562 130484 187568 130496
rect 187620 130484 187626 130536
rect 43030 130416 43036 130468
rect 43088 130456 43094 130468
rect 45422 130456 45428 130468
rect 43088 130428 45428 130456
rect 43088 130416 43094 130428
rect 45422 130416 45428 130428
rect 45480 130416 45486 130468
rect 163734 130416 163740 130468
rect 163792 130456 163798 130468
rect 168150 130456 168156 130468
rect 163792 130428 168156 130456
rect 163792 130416 163798 130428
rect 168150 130416 168156 130428
rect 168208 130416 168214 130468
rect 186826 130416 186832 130468
rect 186884 130456 186890 130468
rect 189218 130456 189224 130468
rect 186884 130428 189224 130456
rect 186884 130416 186890 130428
rect 189218 130416 189224 130428
rect 189276 130416 189282 130468
rect 42294 130348 42300 130400
rect 42352 130388 42358 130400
rect 44686 130388 44692 130400
rect 42352 130360 44692 130388
rect 42352 130348 42358 130360
rect 44686 130348 44692 130360
rect 44744 130348 44750 130400
rect 163826 130348 163832 130400
rect 163884 130388 163890 130400
rect 167598 130388 167604 130400
rect 163884 130360 167604 130388
rect 163884 130348 163890 130360
rect 167598 130348 167604 130360
rect 167656 130348 167662 130400
rect 186642 130348 186648 130400
rect 186700 130388 186706 130400
rect 188666 130388 188672 130400
rect 186700 130360 188672 130388
rect 186700 130348 186706 130360
rect 188666 130348 188672 130360
rect 188724 130348 188730 130400
rect 20858 130280 20864 130332
rect 20916 130320 20922 130332
rect 24998 130320 25004 130332
rect 20916 130292 25004 130320
rect 20916 130280 20922 130292
rect 24998 130280 25004 130292
rect 25056 130280 25062 130332
rect 41834 130280 41840 130332
rect 41892 130320 41898 130332
rect 44042 130320 44048 130332
rect 41892 130292 44048 130320
rect 41892 130280 41898 130292
rect 44042 130280 44048 130292
rect 44100 130280 44106 130332
rect 163918 130280 163924 130332
rect 163976 130320 163982 130332
rect 165298 130320 165304 130332
rect 163976 130292 165304 130320
rect 163976 130280 163982 130292
rect 165298 130280 165304 130292
rect 165356 130280 165362 130332
rect 182502 130280 182508 130332
rect 182560 130320 182566 130332
rect 184158 130320 184164 130332
rect 182560 130292 184164 130320
rect 182560 130280 182566 130292
rect 184158 130280 184164 130292
rect 184216 130280 184222 130332
rect 184802 130280 184808 130332
rect 184860 130320 184866 130332
rect 185814 130320 185820 130332
rect 184860 130292 185820 130320
rect 184860 130280 184866 130292
rect 185814 130280 185820 130292
rect 185872 130280 185878 130332
rect 187286 130280 187292 130332
rect 187344 130320 187350 130332
rect 189862 130320 189868 130332
rect 187344 130292 189868 130320
rect 187344 130280 187350 130292
rect 189862 130280 189868 130292
rect 189920 130280 189926 130332
rect 121690 126880 121696 126932
rect 121748 126920 121754 126932
rect 123990 126920 123996 126932
rect 121748 126892 123996 126920
rect 121748 126880 121754 126892
rect 123990 126880 123996 126892
rect 124048 126880 124054 126932
rect 121782 126200 121788 126252
rect 121840 126240 121846 126252
rect 124358 126240 124364 126252
rect 121840 126212 124364 126240
rect 121840 126200 121846 126212
rect 124358 126200 124364 126212
rect 124416 126200 124422 126252
rect 121690 126132 121696 126184
rect 121748 126172 121754 126184
rect 123898 126172 123904 126184
rect 121748 126144 123904 126172
rect 121748 126132 121754 126144
rect 123898 126132 123904 126144
rect 123956 126132 123962 126184
rect 121690 125112 121696 125164
rect 121748 125152 121754 125164
rect 123714 125152 123720 125164
rect 121748 125124 123720 125152
rect 121748 125112 121754 125124
rect 123714 125112 123720 125124
rect 123772 125112 123778 125164
rect 87742 124568 87748 124620
rect 87800 124608 87806 124620
rect 88754 124608 88760 124620
rect 87800 124580 88760 124608
rect 87800 124568 87806 124580
rect 88754 124568 88760 124580
rect 88812 124568 88818 124620
rect 121690 123480 121696 123532
rect 121748 123520 121754 123532
rect 123530 123520 123536 123532
rect 121748 123492 123536 123520
rect 121748 123480 121754 123492
rect 123530 123480 123536 123492
rect 123588 123480 123594 123532
rect 121690 122120 121696 122172
rect 121748 122160 121754 122172
rect 123438 122160 123444 122172
rect 121748 122132 123444 122160
rect 121748 122120 121754 122132
rect 123438 122120 123444 122132
rect 123496 122120 123502 122172
rect 121690 121984 121696 122036
rect 121748 122024 121754 122036
rect 123346 122024 123352 122036
rect 121748 121996 123352 122024
rect 121748 121984 121754 121996
rect 123346 121984 123352 121996
rect 123404 121984 123410 122036
rect 121690 120896 121696 120948
rect 121748 120936 121754 120948
rect 124358 120936 124364 120948
rect 121748 120908 124364 120936
rect 121748 120896 121754 120908
rect 124358 120896 124364 120908
rect 124416 120896 124422 120948
rect 121690 119332 121696 119384
rect 121748 119372 121754 119384
rect 124266 119372 124272 119384
rect 121748 119344 124272 119372
rect 121748 119332 121754 119344
rect 124266 119332 124272 119344
rect 124324 119332 124330 119384
rect 51126 119264 51132 119316
rect 51184 119304 51190 119316
rect 51586 119304 51592 119316
rect 51184 119276 51592 119304
rect 51184 119264 51190 119276
rect 51586 119264 51592 119276
rect 51644 119264 51650 119316
rect 121690 118176 121696 118228
rect 121748 118216 121754 118228
rect 124358 118216 124364 118228
rect 121748 118188 124364 118216
rect 121748 118176 121754 118188
rect 124358 118176 124364 118188
rect 124416 118176 124422 118228
rect 123070 116544 123076 116596
rect 123128 116584 123134 116596
rect 124266 116584 124272 116596
rect 123128 116556 124272 116584
rect 123128 116544 123134 116556
rect 124266 116544 124272 116556
rect 124324 116544 124330 116596
rect 50574 116476 50580 116528
rect 50632 116516 50638 116528
rect 51586 116516 51592 116528
rect 50632 116488 51592 116516
rect 50632 116476 50638 116488
rect 51586 116476 51592 116488
rect 51644 116476 51650 116528
rect 121690 115660 121696 115712
rect 121748 115700 121754 115712
rect 124358 115700 124364 115712
rect 121748 115672 124364 115700
rect 121748 115660 121754 115672
rect 124358 115660 124364 115672
rect 124416 115660 124422 115712
rect 121690 115388 121696 115440
rect 121748 115428 121754 115440
rect 123990 115428 123996 115440
rect 121748 115400 123996 115428
rect 121748 115388 121754 115400
rect 123990 115388 123996 115400
rect 124048 115388 124054 115440
rect 121690 115116 121696 115168
rect 121748 115156 121754 115168
rect 124266 115156 124272 115168
rect 121748 115128 124272 115156
rect 121748 115116 121754 115128
rect 124266 115116 124272 115128
rect 124324 115116 124330 115168
rect 159042 115116 159048 115168
rect 159100 115156 159106 115168
rect 160606 115156 160612 115168
rect 159100 115128 160612 115156
rect 159100 115116 159106 115128
rect 160606 115116 160612 115128
rect 160664 115116 160670 115168
rect 121690 113960 121696 114012
rect 121748 114000 121754 114012
rect 123438 114000 123444 114012
rect 121748 113972 123444 114000
rect 121748 113960 121754 113972
rect 123438 113960 123444 113972
rect 123496 113960 123502 114012
rect 121690 112328 121696 112380
rect 121748 112368 121754 112380
rect 123346 112368 123352 112380
rect 121748 112340 123352 112368
rect 121748 112328 121754 112340
rect 123346 112328 123352 112340
rect 123404 112328 123410 112380
rect 51218 111240 51224 111292
rect 51276 111280 51282 111292
rect 51586 111280 51592 111292
rect 51276 111252 51592 111280
rect 51276 111240 51282 111252
rect 51586 111240 51592 111252
rect 51644 111240 51650 111292
rect 51218 111104 51224 111156
rect 51276 111144 51282 111156
rect 51678 111144 51684 111156
rect 51276 111116 51684 111144
rect 51276 111104 51282 111116
rect 51678 111104 51684 111116
rect 51736 111104 51742 111156
rect 121690 110968 121696 111020
rect 121748 111008 121754 111020
rect 124266 111008 124272 111020
rect 121748 110980 124272 111008
rect 121748 110968 121754 110980
rect 124266 110968 124272 110980
rect 124324 110968 124330 111020
rect 121690 109744 121696 109796
rect 121748 109784 121754 109796
rect 124358 109784 124364 109796
rect 121748 109756 124364 109784
rect 121748 109744 121754 109756
rect 124358 109744 124364 109756
rect 124416 109744 124422 109796
rect 121690 108724 121696 108776
rect 121748 108764 121754 108776
rect 123438 108764 123444 108776
rect 121748 108736 123444 108764
rect 121748 108724 121754 108736
rect 123438 108724 123444 108736
rect 123496 108724 123502 108776
rect 51218 108520 51224 108572
rect 51276 108560 51282 108572
rect 51586 108560 51592 108572
rect 51276 108532 51592 108560
rect 51276 108520 51282 108532
rect 51586 108520 51592 108532
rect 51644 108520 51650 108572
rect 85166 106860 85172 106872
rect 85127 106832 85172 106860
rect 85166 106820 85172 106832
rect 85224 106820 85230 106872
rect 121690 106820 121696 106872
rect 121748 106860 121754 106872
rect 124266 106860 124272 106872
rect 121748 106832 124272 106860
rect 121748 106820 121754 106832
rect 124266 106820 124272 106832
rect 124324 106820 124330 106872
rect 121690 105868 121696 105920
rect 121748 105908 121754 105920
rect 124358 105908 124364 105920
rect 121748 105880 124364 105908
rect 121748 105868 121754 105880
rect 124358 105868 124364 105880
rect 124416 105868 124422 105920
rect 121690 105596 121696 105648
rect 121748 105636 121754 105648
rect 124174 105636 124180 105648
rect 121748 105608 124180 105636
rect 121748 105596 121754 105608
rect 124174 105596 124180 105608
rect 124232 105596 124238 105648
rect 91054 104684 91060 104696
rect 91015 104656 91060 104684
rect 91054 104644 91060 104656
rect 91112 104644 91118 104696
rect 85902 104100 85908 104152
rect 85960 104140 85966 104152
rect 88662 104140 88668 104152
rect 85960 104112 88668 104140
rect 85960 104100 85966 104112
rect 88662 104100 88668 104112
rect 88720 104100 88726 104152
rect 121782 104100 121788 104152
rect 121840 104140 121846 104152
rect 126934 104140 126940 104152
rect 121840 104112 126940 104140
rect 121840 104100 121846 104112
rect 126934 104100 126940 104112
rect 126992 104100 126998 104152
rect 85810 104032 85816 104084
rect 85868 104072 85874 104084
rect 88570 104072 88576 104084
rect 85868 104044 88576 104072
rect 85868 104032 85874 104044
rect 88570 104032 88576 104044
rect 88628 104032 88634 104084
rect 121690 104032 121696 104084
rect 121748 104072 121754 104084
rect 127026 104072 127032 104084
rect 121748 104044 127032 104072
rect 121748 104032 121754 104044
rect 127026 104032 127032 104044
rect 127084 104032 127090 104084
rect 157570 104032 157576 104084
rect 157628 104072 157634 104084
rect 160330 104072 160336 104084
rect 157628 104044 160336 104072
rect 157628 104032 157634 104044
rect 160330 104032 160336 104044
rect 160388 104032 160394 104084
rect 50758 103012 50764 103064
rect 50816 103052 50822 103064
rect 54070 103052 54076 103064
rect 50816 103024 54076 103052
rect 50816 103012 50822 103024
rect 54070 103012 54076 103024
rect 54128 103012 54134 103064
rect 121690 102808 121696 102860
rect 121748 102848 121754 102860
rect 124542 102848 124548 102860
rect 121748 102820 124548 102848
rect 121748 102808 121754 102820
rect 124542 102808 124548 102820
rect 124600 102808 124606 102860
rect 51218 102740 51224 102792
rect 51276 102780 51282 102792
rect 55358 102780 55364 102792
rect 51276 102752 55364 102780
rect 51276 102740 51282 102752
rect 55358 102740 55364 102752
rect 55416 102740 55422 102792
rect 121782 102740 121788 102792
rect 121840 102780 121846 102792
rect 125922 102780 125928 102792
rect 121840 102752 125928 102780
rect 121840 102740 121846 102752
rect 125922 102740 125928 102752
rect 125980 102740 125986 102792
rect 127118 102740 127124 102792
rect 127176 102740 127182 102792
rect 121874 102672 121880 102724
rect 121932 102712 121938 102724
rect 127136 102712 127164 102740
rect 121932 102684 127164 102712
rect 121932 102672 121938 102684
rect 81578 101380 81584 101432
rect 81636 101420 81642 101432
rect 88662 101420 88668 101432
rect 81636 101392 88668 101420
rect 81636 101380 81642 101392
rect 88662 101380 88668 101392
rect 88720 101380 88726 101432
rect 152786 101380 152792 101432
rect 152844 101420 152850 101432
rect 160422 101420 160428 101432
rect 152844 101392 160428 101420
rect 152844 101380 152850 101392
rect 160422 101380 160428 101392
rect 160480 101380 160486 101432
rect 51218 101312 51224 101364
rect 51276 101352 51282 101364
rect 52598 101352 52604 101364
rect 51276 101324 52604 101352
rect 51276 101312 51282 101324
rect 52598 101312 52604 101324
rect 52656 101312 52662 101364
rect 80474 101312 80480 101364
rect 80532 101352 80538 101364
rect 88570 101352 88576 101364
rect 80532 101324 88576 101352
rect 80532 101312 80538 101324
rect 88570 101312 88576 101324
rect 88628 101312 88634 101364
rect 153890 101312 153896 101364
rect 153948 101352 153954 101364
rect 160330 101352 160336 101364
rect 153948 101324 160336 101352
rect 153948 101312 153954 101324
rect 160330 101312 160336 101324
rect 160388 101312 160394 101364
rect 18006 101244 18012 101296
rect 18064 101284 18070 101296
rect 58394 101284 58400 101296
rect 18064 101256 58400 101284
rect 18064 101244 18070 101256
rect 58394 101244 58400 101256
rect 58452 101244 58458 101296
rect 128958 101244 128964 101296
rect 129016 101284 129022 101296
rect 193542 101284 193548 101296
rect 129016 101256 193548 101284
rect 129016 101244 129022 101256
rect 193542 101244 193548 101256
rect 193600 101244 193606 101296
rect 116354 101040 116360 101092
rect 116412 101080 116418 101092
rect 127578 101080 127584 101092
rect 116412 101052 127584 101080
rect 116412 101040 116418 101052
rect 127578 101040 127584 101052
rect 127636 101040 127642 101092
rect 73758 100768 73764 100820
rect 73816 100808 73822 100820
rect 78358 100808 78364 100820
rect 73816 100780 78364 100808
rect 73816 100768 73822 100780
rect 78358 100768 78364 100780
rect 78416 100768 78422 100820
rect 127578 100564 127584 100616
rect 127636 100604 127642 100616
rect 190598 100604 190604 100616
rect 127636 100576 190604 100604
rect 127636 100564 127642 100576
rect 190598 100564 190604 100576
rect 190656 100604 190662 100616
rect 193450 100604 193456 100616
rect 190656 100576 193456 100604
rect 190656 100564 190662 100576
rect 193450 100564 193456 100576
rect 193508 100564 193514 100616
rect 71550 100360 71556 100412
rect 71608 100400 71614 100412
rect 72749 100403 72807 100409
rect 72749 100400 72761 100403
rect 71608 100372 72761 100400
rect 71608 100360 71614 100372
rect 72749 100369 72761 100372
rect 72795 100369 72807 100403
rect 72749 100363 72807 100369
rect 65113 100335 65171 100341
rect 65113 100301 65125 100335
rect 65159 100332 65171 100335
rect 74681 100335 74739 100341
rect 74681 100332 74693 100335
rect 65159 100304 74693 100332
rect 65159 100301 65171 100304
rect 65113 100295 65171 100301
rect 74681 100301 74693 100304
rect 74727 100301 74739 100335
rect 74681 100295 74739 100301
rect 106513 100267 106571 100273
rect 106513 100233 106525 100267
rect 106559 100264 106571 100267
rect 116081 100267 116139 100273
rect 116081 100264 116093 100267
rect 106559 100236 116093 100264
rect 106559 100233 106571 100236
rect 106513 100227 106571 100233
rect 116081 100233 116093 100236
rect 116127 100233 116139 100267
rect 116081 100227 116139 100233
rect 69342 100156 69348 100208
rect 69400 100196 69406 100208
rect 72654 100196 72660 100208
rect 69400 100168 72660 100196
rect 69400 100156 69406 100168
rect 72654 100156 72660 100168
rect 72712 100156 72718 100208
rect 72749 100199 72807 100205
rect 72749 100165 72761 100199
rect 72795 100196 72807 100199
rect 75506 100196 75512 100208
rect 72795 100168 75512 100196
rect 72795 100165 72807 100168
rect 72749 100159 72807 100165
rect 75506 100156 75512 100168
rect 75564 100156 75570 100208
rect 80293 100199 80351 100205
rect 80293 100196 80305 100199
rect 75616 100168 80305 100196
rect 64926 100088 64932 100140
rect 64984 100128 64990 100140
rect 66950 100128 66956 100140
rect 64984 100100 66956 100128
rect 64984 100088 64990 100100
rect 66950 100088 66956 100100
rect 67008 100088 67014 100140
rect 68238 100088 68244 100140
rect 68296 100128 68302 100140
rect 71182 100128 71188 100140
rect 68296 100100 71188 100128
rect 68296 100088 68302 100100
rect 71182 100088 71188 100100
rect 71240 100088 71246 100140
rect 74773 100131 74831 100137
rect 74773 100097 74785 100131
rect 74819 100128 74831 100131
rect 75616 100128 75644 100168
rect 80293 100165 80305 100168
rect 80339 100165 80351 100199
rect 80293 100159 80351 100165
rect 145978 100156 145984 100208
rect 146036 100196 146042 100208
rect 150394 100196 150400 100208
rect 146036 100168 150400 100196
rect 146036 100156 146042 100168
rect 150394 100156 150400 100168
rect 150452 100156 150458 100208
rect 74819 100100 75644 100128
rect 74819 100097 74831 100100
rect 74773 100091 74831 100097
rect 75966 100088 75972 100140
rect 76024 100128 76030 100140
rect 81210 100128 81216 100140
rect 76024 100100 81216 100128
rect 76024 100088 76030 100100
rect 81210 100088 81216 100100
rect 81268 100088 81274 100140
rect 95930 100088 95936 100140
rect 95988 100128 95994 100140
rect 99521 100131 99579 100137
rect 99521 100128 99533 100131
rect 95988 100100 99533 100128
rect 95988 100088 95994 100100
rect 99521 100097 99533 100100
rect 99567 100097 99579 100131
rect 99521 100091 99579 100097
rect 116081 100131 116139 100137
rect 116081 100097 116093 100131
rect 116127 100128 116139 100131
rect 116354 100128 116360 100140
rect 116127 100100 116360 100128
rect 116127 100097 116139 100100
rect 116081 100091 116139 100097
rect 116354 100088 116360 100100
rect 116412 100088 116418 100140
rect 144966 100088 144972 100140
rect 145024 100128 145030 100140
rect 148922 100128 148928 100140
rect 145024 100100 148928 100128
rect 145024 100088 145030 100100
rect 148922 100088 148928 100100
rect 148980 100088 148986 100140
rect 56738 100020 56744 100072
rect 56796 100060 56802 100072
rect 64193 100063 64251 100069
rect 64193 100060 64205 100063
rect 56796 100032 64205 100060
rect 56796 100020 56802 100032
rect 64193 100029 64205 100032
rect 64239 100029 64251 100063
rect 64193 100023 64251 100029
rect 67134 100020 67140 100072
rect 67192 100060 67198 100072
rect 69802 100060 69808 100072
rect 67192 100032 69808 100060
rect 67192 100020 67198 100032
rect 69802 100020 69808 100032
rect 69860 100020 69866 100072
rect 70446 100020 70452 100072
rect 70504 100060 70510 100072
rect 74034 100060 74040 100072
rect 70504 100032 74040 100060
rect 70504 100020 70510 100032
rect 74034 100020 74040 100032
rect 74092 100020 74098 100072
rect 74862 100020 74868 100072
rect 74920 100060 74926 100072
rect 79738 100060 79744 100072
rect 74920 100032 79744 100060
rect 74920 100020 74926 100032
rect 79738 100020 79744 100032
rect 79796 100020 79802 100072
rect 141654 100020 141660 100072
rect 141712 100060 141718 100072
rect 144690 100060 144696 100072
rect 141712 100032 144696 100060
rect 141712 100020 141718 100032
rect 144690 100020 144696 100032
rect 144748 100020 144754 100072
rect 148278 100020 148284 100072
rect 148336 100060 148342 100072
rect 153246 100060 153252 100072
rect 148336 100032 153252 100060
rect 148336 100020 148342 100032
rect 153246 100020 153252 100032
rect 153304 100020 153310 100072
rect 63822 99952 63828 100004
rect 63880 99992 63886 100004
rect 65478 99992 65484 100004
rect 63880 99964 65484 99992
rect 63880 99952 63886 99964
rect 65478 99952 65484 99964
rect 65536 99952 65542 100004
rect 66030 99952 66036 100004
rect 66088 99992 66094 100004
rect 68330 99992 68336 100004
rect 66088 99964 68336 99992
rect 66088 99952 66094 99964
rect 68330 99952 68336 99964
rect 68388 99952 68394 100004
rect 72654 99952 72660 100004
rect 72712 99992 72718 100004
rect 76886 99992 76892 100004
rect 72712 99964 76892 99992
rect 72712 99952 72718 99964
rect 76886 99952 76892 99964
rect 76944 99952 76950 100004
rect 99521 99995 99579 100001
rect 99521 99961 99533 99995
rect 99567 99992 99579 99995
rect 106513 99995 106571 100001
rect 106513 99992 106525 99995
rect 99567 99964 106525 99992
rect 99567 99961 99579 99964
rect 99521 99955 99579 99961
rect 106513 99961 106525 99964
rect 106559 99961 106571 99995
rect 106513 99955 106571 99961
rect 136042 99952 136048 100004
rect 136100 99992 136106 100004
rect 137514 99992 137520 100004
rect 136100 99964 137520 99992
rect 136100 99952 136106 99964
rect 137514 99952 137520 99964
rect 137572 99952 137578 100004
rect 138158 99952 138164 100004
rect 138216 99992 138222 100004
rect 140366 99992 140372 100004
rect 138216 99964 140372 99992
rect 138216 99952 138222 99964
rect 140366 99952 140372 99964
rect 140424 99952 140430 100004
rect 140550 99952 140556 100004
rect 140608 99992 140614 100004
rect 143218 99992 143224 100004
rect 140608 99964 143224 99992
rect 140608 99952 140614 99964
rect 143218 99952 143224 99964
rect 143276 99952 143282 100004
rect 143678 99952 143684 100004
rect 143736 99992 143742 100004
rect 147542 99992 147548 100004
rect 143736 99964 147548 99992
rect 143736 99952 143742 99964
rect 147542 99952 147548 99964
rect 147600 99952 147606 100004
rect 59314 99884 59320 99936
rect 59372 99924 59378 99936
rect 59774 99924 59780 99936
rect 59372 99896 59780 99924
rect 59372 99884 59378 99896
rect 59774 99884 59780 99896
rect 59832 99884 59838 99936
rect 60418 99884 60424 99936
rect 60476 99924 60482 99936
rect 61246 99924 61252 99936
rect 60476 99896 61252 99924
rect 60476 99884 60482 99896
rect 61246 99884 61252 99896
rect 61304 99884 61310 99936
rect 61522 99884 61528 99936
rect 61580 99924 61586 99936
rect 62626 99924 62632 99936
rect 61580 99896 62632 99924
rect 61580 99884 61586 99896
rect 62626 99884 62632 99896
rect 62684 99884 62690 99936
rect 62994 99884 63000 99936
rect 63052 99924 63058 99936
rect 64098 99924 64104 99936
rect 63052 99896 64104 99924
rect 63052 99884 63058 99896
rect 64098 99884 64104 99896
rect 64156 99884 64162 99936
rect 64193 99927 64251 99933
rect 64193 99893 64205 99927
rect 64239 99924 64251 99927
rect 65113 99927 65171 99933
rect 65113 99924 65125 99927
rect 64239 99896 65125 99924
rect 64239 99893 64251 99896
rect 64193 99887 64251 99893
rect 65113 99893 65125 99896
rect 65159 99893 65171 99927
rect 65113 99887 65171 99893
rect 74681 99927 74739 99933
rect 74681 99893 74693 99927
rect 74727 99924 74739 99927
rect 74773 99927 74831 99933
rect 74773 99924 74785 99927
rect 74727 99896 74785 99924
rect 74727 99893 74739 99896
rect 74681 99887 74739 99893
rect 74773 99893 74785 99896
rect 74819 99893 74831 99927
rect 74773 99887 74831 99893
rect 80293 99927 80351 99933
rect 80293 99893 80305 99927
rect 80339 99924 80351 99927
rect 95930 99924 95936 99936
rect 80339 99896 95936 99924
rect 80339 99893 80351 99896
rect 80293 99887 80351 99893
rect 95930 99884 95936 99896
rect 95988 99884 95994 99936
rect 97034 99884 97040 99936
rect 97092 99924 97098 99936
rect 130430 99924 130436 99936
rect 97092 99896 130436 99924
rect 97092 99884 97098 99896
rect 130430 99884 130436 99896
rect 130488 99884 130494 99936
rect 131258 99884 131264 99936
rect 131316 99924 131322 99936
rect 131810 99924 131816 99936
rect 131316 99896 131816 99924
rect 131316 99884 131322 99896
rect 131810 99884 131816 99896
rect 131868 99884 131874 99936
rect 132546 99884 132552 99936
rect 132604 99924 132610 99936
rect 133282 99924 133288 99936
rect 132604 99896 133288 99924
rect 132604 99884 132610 99896
rect 133282 99884 133288 99896
rect 133340 99884 133346 99936
rect 133834 99884 133840 99936
rect 133892 99924 133898 99936
rect 134662 99924 134668 99936
rect 133892 99896 134668 99924
rect 133892 99884 133898 99896
rect 134662 99884 134668 99896
rect 134720 99884 134726 99936
rect 134938 99884 134944 99936
rect 134996 99924 135002 99936
rect 136134 99924 136140 99936
rect 134996 99896 136140 99924
rect 134996 99884 135002 99896
rect 136134 99884 136140 99896
rect 136192 99884 136198 99936
rect 137238 99884 137244 99936
rect 137296 99924 137302 99936
rect 138986 99924 138992 99936
rect 137296 99896 138992 99924
rect 137296 99884 137302 99896
rect 138986 99884 138992 99896
rect 139044 99884 139050 99936
rect 139446 99884 139452 99936
rect 139504 99924 139510 99936
rect 141838 99924 141844 99936
rect 139504 99896 141844 99924
rect 139504 99884 139510 99896
rect 141838 99884 141844 99896
rect 141896 99884 141902 99936
rect 142758 99884 142764 99936
rect 142816 99924 142822 99936
rect 146070 99924 146076 99936
rect 142816 99896 146076 99924
rect 142816 99884 142822 99896
rect 146070 99884 146076 99896
rect 146128 99884 146134 99936
rect 147174 99884 147180 99936
rect 147232 99924 147238 99936
rect 151774 99924 151780 99936
rect 147232 99896 151780 99924
rect 147232 99884 147238 99896
rect 151774 99884 151780 99896
rect 151832 99884 151838 99936
rect 154626 99884 154632 99936
rect 154684 99924 154690 99936
rect 160974 99924 160980 99936
rect 154684 99896 160980 99924
rect 154684 99884 154690 99896
rect 160974 99884 160980 99896
rect 161032 99884 161038 99936
rect 56922 98456 56928 98508
rect 56980 98496 56986 98508
rect 97126 98496 97132 98508
rect 56980 98468 97132 98496
rect 56980 98456 56986 98468
rect 97126 98456 97132 98468
rect 97184 98456 97190 98508
rect 93354 98252 93360 98304
rect 93412 98292 93418 98304
rect 94366 98292 94372 98304
rect 93412 98264 94372 98292
rect 93412 98252 93418 98264
rect 94366 98252 94372 98264
rect 94424 98252 94430 98304
rect 92158 98116 92164 98168
rect 92216 98156 92222 98168
rect 94090 98156 94096 98168
rect 92216 98128 94096 98156
rect 92216 98116 92222 98128
rect 94090 98116 94096 98128
rect 94148 98116 94154 98168
rect 171002 98116 171008 98168
rect 171060 98156 171066 98168
rect 171646 98156 171652 98168
rect 171060 98128 171652 98156
rect 171060 98116 171066 98128
rect 171646 98116 171652 98128
rect 171704 98116 171710 98168
rect 182226 98116 182232 98168
rect 182284 98156 182290 98168
rect 183514 98156 183520 98168
rect 182284 98128 183520 98156
rect 182284 98116 182290 98128
rect 183514 98116 183520 98128
rect 183572 98116 183578 98168
rect 92342 98048 92348 98100
rect 92400 98088 92406 98100
rect 94918 98088 94924 98100
rect 92400 98060 94924 98088
rect 92400 98048 92406 98060
rect 94918 98048 94924 98060
rect 94976 98048 94982 98100
rect 21778 97776 21784 97828
rect 21836 97816 21842 97828
rect 23618 97816 23624 97828
rect 21836 97788 23624 97816
rect 21836 97776 21842 97788
rect 23618 97776 23624 97788
rect 23676 97776 23682 97828
rect 168518 97776 168524 97828
rect 168576 97816 168582 97828
rect 191518 97816 191524 97828
rect 168576 97788 191524 97816
rect 168576 97776 168582 97788
rect 191518 97776 191524 97788
rect 191576 97776 191582 97828
rect 179742 97640 179748 97692
rect 179800 97680 179806 97692
rect 181858 97680 181864 97692
rect 179800 97652 181864 97680
rect 179800 97640 179806 97652
rect 181858 97640 181864 97652
rect 181916 97640 181922 97692
rect 181582 97504 181588 97556
rect 181640 97544 181646 97556
rect 182410 97544 182416 97556
rect 181640 97516 182416 97544
rect 181640 97504 181646 97516
rect 182410 97504 182416 97516
rect 182468 97504 182474 97556
rect 23250 97436 23256 97488
rect 23308 97476 23314 97488
rect 24906 97476 24912 97488
rect 23308 97448 24912 97476
rect 23308 97436 23314 97448
rect 24906 97436 24912 97448
rect 24964 97436 24970 97488
rect 27298 97300 27304 97352
rect 27356 97340 27362 97352
rect 29046 97340 29052 97352
rect 27356 97312 29052 97340
rect 27356 97300 27362 97312
rect 29046 97300 29052 97312
rect 29104 97300 29110 97352
rect 105222 97300 105228 97352
rect 105280 97340 105286 97352
rect 107062 97340 107068 97352
rect 105280 97312 107068 97340
rect 105280 97300 105286 97312
rect 107062 97300 107068 97312
rect 107120 97300 107126 97352
rect 163826 97300 163832 97352
rect 163884 97340 163890 97352
rect 167598 97340 167604 97352
rect 163884 97312 167604 97340
rect 163884 97300 163890 97312
rect 167598 97300 167604 97312
rect 167656 97300 167662 97352
rect 169254 97300 169260 97352
rect 169312 97340 169318 97352
rect 170450 97340 170456 97352
rect 169312 97312 170456 97340
rect 169312 97300 169318 97312
rect 170450 97300 170456 97312
rect 170508 97300 170514 97352
rect 23526 97232 23532 97284
rect 23584 97272 23590 97284
rect 23584 97244 25504 97272
rect 23584 97232 23590 97244
rect 24538 97164 24544 97216
rect 24596 97204 24602 97216
rect 24596 97176 25412 97204
rect 24596 97164 24602 97176
rect 25384 97068 25412 97176
rect 25476 97136 25504 97244
rect 28586 97232 28592 97284
rect 28644 97272 28650 97284
rect 30426 97272 30432 97284
rect 28644 97244 30432 97272
rect 28644 97232 28650 97244
rect 30426 97232 30432 97244
rect 30484 97232 30490 97284
rect 30518 97232 30524 97284
rect 30576 97272 30582 97284
rect 31622 97272 31628 97284
rect 30576 97244 31628 97272
rect 30576 97232 30582 97244
rect 31622 97232 31628 97244
rect 31680 97232 31686 97284
rect 37602 97232 37608 97284
rect 37660 97272 37666 97284
rect 39718 97272 39724 97284
rect 37660 97244 39724 97272
rect 37660 97232 37666 97244
rect 39718 97232 39724 97244
rect 39776 97232 39782 97284
rect 40362 97232 40368 97284
rect 40420 97272 40426 97284
rect 42294 97272 42300 97284
rect 40420 97244 42300 97272
rect 40420 97232 40426 97244
rect 42294 97232 42300 97244
rect 42352 97232 42358 97284
rect 103750 97232 103756 97284
rect 103808 97272 103814 97284
rect 105406 97272 105412 97284
rect 103808 97244 105412 97272
rect 103808 97232 103814 97244
rect 105406 97232 105412 97244
rect 105464 97232 105470 97284
rect 106602 97232 106608 97284
rect 106660 97272 106666 97284
rect 108718 97272 108724 97284
rect 106660 97244 108724 97272
rect 106660 97232 106666 97244
rect 108718 97232 108724 97244
rect 108776 97232 108782 97284
rect 163734 97232 163740 97284
rect 163792 97272 163798 97284
rect 165298 97272 165304 97284
rect 163792 97244 165304 97272
rect 163792 97232 163798 97244
rect 165298 97232 165304 97244
rect 165356 97232 165362 97284
rect 169898 97232 169904 97284
rect 169956 97272 169962 97284
rect 170818 97272 170824 97284
rect 169956 97244 170824 97272
rect 169956 97232 169962 97244
rect 170818 97232 170824 97244
rect 170876 97232 170882 97284
rect 184434 97232 184440 97284
rect 184492 97272 184498 97284
rect 186366 97272 186372 97284
rect 184492 97244 186372 97272
rect 184492 97232 184498 97244
rect 186366 97232 186372 97244
rect 186424 97232 186430 97284
rect 26010 97164 26016 97216
rect 26068 97204 26074 97216
rect 26068 97176 27804 97204
rect 26068 97164 26074 97176
rect 27666 97136 27672 97148
rect 25476 97108 27672 97136
rect 27666 97096 27672 97108
rect 27724 97096 27730 97148
rect 27776 97136 27804 97176
rect 29138 97164 29144 97216
rect 29196 97204 29202 97216
rect 29196 97176 30012 97204
rect 29196 97164 29202 97176
rect 28862 97136 28868 97148
rect 27776 97108 28868 97136
rect 28862 97096 28868 97108
rect 28920 97096 28926 97148
rect 29984 97136 30012 97176
rect 30058 97164 30064 97216
rect 30116 97204 30122 97216
rect 31254 97204 31260 97216
rect 30116 97176 31260 97204
rect 30116 97164 30122 97176
rect 31254 97164 31260 97176
rect 31312 97164 31318 97216
rect 31346 97164 31352 97216
rect 31404 97204 31410 97216
rect 37510 97204 37516 97216
rect 31404 97176 32128 97204
rect 31404 97164 31410 97176
rect 30886 97136 30892 97148
rect 29984 97108 30892 97136
rect 30886 97096 30892 97108
rect 30944 97096 30950 97148
rect 32100 97080 32128 97176
rect 36424 97176 37516 97204
rect 36038 97096 36044 97148
rect 36096 97136 36102 97148
rect 36424 97136 36452 97176
rect 37510 97164 37516 97176
rect 37568 97164 37574 97216
rect 38982 97204 38988 97216
rect 38356 97176 38988 97204
rect 36096 97108 36452 97136
rect 36096 97096 36102 97108
rect 36498 97096 36504 97148
rect 36556 97136 36562 97148
rect 38246 97136 38252 97148
rect 36556 97108 38252 97136
rect 36556 97096 36562 97108
rect 38246 97096 38252 97108
rect 38304 97096 38310 97148
rect 28034 97068 28040 97080
rect 25384 97040 28040 97068
rect 28034 97028 28040 97040
rect 28092 97028 28098 97080
rect 32082 97028 32088 97080
rect 32140 97028 32146 97080
rect 35670 97028 35676 97080
rect 35728 97068 35734 97080
rect 36958 97068 36964 97080
rect 35728 97040 36964 97068
rect 35728 97028 35734 97040
rect 36958 97028 36964 97040
rect 37016 97028 37022 97080
rect 37142 97028 37148 97080
rect 37200 97068 37206 97080
rect 38356 97068 38384 97176
rect 38982 97164 38988 97176
rect 39040 97164 39046 97216
rect 41006 97204 41012 97216
rect 39184 97176 41012 97204
rect 38430 97096 38436 97148
rect 38488 97136 38494 97148
rect 39184 97136 39212 97176
rect 41006 97164 41012 97176
rect 41064 97164 41070 97216
rect 92434 97164 92440 97216
rect 92492 97204 92498 97216
rect 93262 97204 93268 97216
rect 92492 97176 93268 97204
rect 92492 97164 92498 97176
rect 93262 97164 93268 97176
rect 93320 97164 93326 97216
rect 105130 97204 105136 97216
rect 103768 97176 105136 97204
rect 38488 97108 39212 97136
rect 38488 97096 38494 97108
rect 40822 97096 40828 97148
rect 40880 97136 40886 97148
rect 45882 97136 45888 97148
rect 40880 97108 45888 97136
rect 40880 97096 40886 97108
rect 45882 97096 45888 97108
rect 45940 97096 45946 97148
rect 85902 97096 85908 97148
rect 85960 97136 85966 97148
rect 87098 97136 87104 97148
rect 85960 97108 87104 97136
rect 85960 97096 85966 97108
rect 87098 97096 87104 97108
rect 87156 97096 87162 97148
rect 103474 97096 103480 97148
rect 103532 97136 103538 97148
rect 103768 97136 103796 97176
rect 105130 97164 105136 97176
rect 105188 97164 105194 97216
rect 106510 97204 106516 97216
rect 105240 97176 106516 97204
rect 103532 97108 103796 97136
rect 103532 97096 103538 97108
rect 104670 97096 104676 97148
rect 104728 97136 104734 97148
rect 105240 97136 105268 97176
rect 106510 97164 106516 97176
rect 106568 97164 106574 97216
rect 108166 97204 108172 97216
rect 106620 97176 108172 97204
rect 104728 97108 105268 97136
rect 104728 97096 104734 97108
rect 105866 97096 105872 97148
rect 105924 97136 105930 97148
rect 106620 97136 106648 97176
rect 108166 97164 108172 97176
rect 108224 97164 108230 97216
rect 109822 97204 109828 97216
rect 108276 97176 109828 97204
rect 105924 97108 106648 97136
rect 105924 97096 105930 97108
rect 107154 97096 107160 97148
rect 107212 97136 107218 97148
rect 108276 97136 108304 97176
rect 109822 97164 109828 97176
rect 109880 97164 109886 97216
rect 111478 97204 111484 97216
rect 110392 97176 111484 97204
rect 107212 97108 108304 97136
rect 107212 97096 107218 97108
rect 108350 97096 108356 97148
rect 108408 97136 108414 97148
rect 110392 97136 110420 97176
rect 111478 97164 111484 97176
rect 111536 97164 111542 97216
rect 165114 97164 165120 97216
rect 165172 97204 165178 97216
rect 165850 97204 165856 97216
rect 165172 97176 165856 97204
rect 165172 97164 165178 97176
rect 165850 97164 165856 97176
rect 165908 97164 165914 97216
rect 168702 97164 168708 97216
rect 168760 97204 168766 97216
rect 170082 97204 170088 97216
rect 168760 97176 170088 97204
rect 168760 97164 168766 97176
rect 170082 97164 170088 97176
rect 170140 97164 170146 97216
rect 176890 97164 176896 97216
rect 176948 97204 176954 97216
rect 178454 97204 178460 97216
rect 176948 97176 178460 97204
rect 176948 97164 176954 97176
rect 178454 97164 178460 97176
rect 178512 97164 178518 97216
rect 180110 97204 180116 97216
rect 178656 97176 180116 97204
rect 108408 97108 110420 97136
rect 108408 97096 108414 97108
rect 123070 97096 123076 97148
rect 123128 97136 123134 97148
rect 124450 97136 124456 97148
rect 123128 97108 124456 97136
rect 123128 97096 123134 97108
rect 124450 97096 124456 97108
rect 124508 97096 124514 97148
rect 127118 97096 127124 97148
rect 127176 97136 127182 97148
rect 127670 97136 127676 97148
rect 127176 97108 127676 97136
rect 127176 97096 127182 97108
rect 127670 97096 127676 97108
rect 127728 97096 127734 97148
rect 154626 97096 154632 97148
rect 154684 97136 154690 97148
rect 160514 97136 160520 97148
rect 154684 97108 160520 97136
rect 154684 97096 154690 97108
rect 160514 97096 160520 97108
rect 160572 97096 160578 97148
rect 176430 97096 176436 97148
rect 176488 97136 176494 97148
rect 177810 97136 177816 97148
rect 176488 97108 177816 97136
rect 176488 97096 176494 97108
rect 177810 97096 177816 97108
rect 177868 97096 177874 97148
rect 178086 97096 178092 97148
rect 178144 97136 178150 97148
rect 178656 97136 178684 97176
rect 180110 97164 180116 97176
rect 180168 97164 180174 97216
rect 182962 97204 182968 97216
rect 182520 97176 182968 97204
rect 178144 97108 178684 97136
rect 178144 97096 178150 97108
rect 179650 97096 179656 97148
rect 179708 97136 179714 97148
rect 181582 97136 181588 97148
rect 179708 97108 181588 97136
rect 179708 97096 179714 97108
rect 181582 97096 181588 97108
rect 181640 97096 181646 97148
rect 182520 97136 182548 97176
rect 182962 97164 182968 97176
rect 183020 97164 183026 97216
rect 184710 97204 184716 97216
rect 183072 97176 184716 97204
rect 181968 97108 182548 97136
rect 37200 97040 38384 97068
rect 37200 97028 37206 97040
rect 38890 97028 38896 97080
rect 38948 97068 38954 97080
rect 40362 97068 40368 97080
rect 38948 97040 40368 97068
rect 38948 97028 38954 97040
rect 40362 97028 40368 97040
rect 40420 97028 40426 97080
rect 40454 97028 40460 97080
rect 40512 97068 40518 97080
rect 45054 97068 45060 97080
rect 40512 97040 45060 97068
rect 40512 97028 40518 97040
rect 45054 97028 45060 97040
rect 45112 97028 45118 97080
rect 50942 97028 50948 97080
rect 51000 97068 51006 97080
rect 57106 97068 57112 97080
rect 51000 97040 57112 97068
rect 51000 97028 51006 97040
rect 57106 97028 57112 97040
rect 57164 97028 57170 97080
rect 105498 97028 105504 97080
rect 105556 97068 105562 97080
rect 107982 97068 107988 97080
rect 105556 97040 107988 97068
rect 105556 97028 105562 97040
rect 107982 97028 107988 97040
rect 108040 97028 108046 97080
rect 126934 97028 126940 97080
rect 126992 97068 126998 97080
rect 129970 97068 129976 97080
rect 126992 97040 129976 97068
rect 126992 97028 126998 97040
rect 129970 97028 129976 97040
rect 130028 97028 130034 97080
rect 176062 97028 176068 97080
rect 176120 97068 176126 97080
rect 177258 97068 177264 97080
rect 176120 97040 177264 97068
rect 176120 97028 176126 97040
rect 177258 97028 177264 97040
rect 177316 97028 177322 97080
rect 177626 97028 177632 97080
rect 177684 97068 177690 97080
rect 179558 97068 179564 97080
rect 177684 97040 179564 97068
rect 177684 97028 177690 97040
rect 179558 97028 179564 97040
rect 179616 97028 179622 97080
rect 180018 97028 180024 97080
rect 180076 97068 180082 97080
rect 181968 97068 181996 97108
rect 180076 97040 181996 97068
rect 180076 97028 180082 97040
rect 20950 96960 20956 97012
rect 21008 97000 21014 97012
rect 26102 97000 26108 97012
rect 21008 96972 26108 97000
rect 21008 96960 21014 96972
rect 26102 96960 26108 96972
rect 26160 96960 26166 97012
rect 26197 97003 26255 97009
rect 26197 96969 26209 97003
rect 26243 97000 26255 97003
rect 26838 97000 26844 97012
rect 26243 96972 26844 97000
rect 26243 96969 26255 96972
rect 26197 96963 26255 96969
rect 26838 96960 26844 96972
rect 26896 96960 26902 97012
rect 37694 96960 37700 97012
rect 37752 97000 37758 97012
rect 40178 97000 40184 97012
rect 37752 96972 40184 97000
rect 37752 96960 37758 96972
rect 40178 96960 40184 96972
rect 40236 96960 40242 97012
rect 107522 96960 107528 97012
rect 107580 97000 107586 97012
rect 110742 97000 110748 97012
rect 107580 96972 110748 97000
rect 107580 96960 107586 96972
rect 110742 96960 110748 96972
rect 110800 96960 110806 97012
rect 178454 96960 178460 97012
rect 178512 97000 178518 97012
rect 180662 97000 180668 97012
rect 178512 96972 180668 97000
rect 178512 96960 178518 96972
rect 180662 96960 180668 96972
rect 180720 96960 180726 97012
rect 181214 96960 181220 97012
rect 181272 97000 181278 97012
rect 183072 97000 183100 97176
rect 184710 97164 184716 97176
rect 184768 97164 184774 97216
rect 184802 97096 184808 97148
rect 184860 97136 184866 97148
rect 189862 97136 189868 97148
rect 184860 97108 189868 97136
rect 184860 97096 184866 97108
rect 189862 97096 189868 97108
rect 189920 97096 189926 97148
rect 185630 97028 185636 97080
rect 185688 97068 185694 97080
rect 190966 97068 190972 97080
rect 185688 97040 190972 97068
rect 185688 97028 185694 97040
rect 190966 97028 190972 97040
rect 191024 97028 191030 97080
rect 181272 96972 183100 97000
rect 181272 96960 181278 96972
rect 184066 96960 184072 97012
rect 184124 97000 184130 97012
rect 188666 97000 188672 97012
rect 184124 96972 188672 97000
rect 184124 96960 184130 96972
rect 188666 96960 188672 96972
rect 188724 96960 188730 97012
rect 41282 96892 41288 96944
rect 41340 96932 41346 96944
rect 46526 96932 46532 96944
rect 41340 96904 46532 96932
rect 41340 96892 41346 96904
rect 46526 96892 46532 96904
rect 46584 96892 46590 96944
rect 107798 96892 107804 96944
rect 107856 96932 107862 96944
rect 110926 96932 110932 96944
rect 107856 96904 110932 96932
rect 107856 96892 107862 96904
rect 110926 96892 110932 96904
rect 110984 96892 110990 96944
rect 165942 96892 165948 96944
rect 166000 96932 166006 96944
rect 166678 96932 166684 96944
rect 166000 96904 166684 96932
rect 166000 96892 166006 96904
rect 166678 96892 166684 96904
rect 166736 96892 166742 96944
rect 177258 96892 177264 96944
rect 177316 96932 177322 96944
rect 179006 96932 179012 96944
rect 177316 96904 179012 96932
rect 177316 96892 177322 96904
rect 179006 96892 179012 96904
rect 179064 96892 179070 96944
rect 182042 96892 182048 96944
rect 182100 96932 182106 96944
rect 185814 96932 185820 96944
rect 182100 96904 185820 96932
rect 182100 96892 182106 96904
rect 185814 96892 185820 96904
rect 185872 96892 185878 96944
rect 24906 96824 24912 96876
rect 24964 96864 24970 96876
rect 27298 96864 27304 96876
rect 24964 96836 27304 96864
rect 24964 96824 24970 96836
rect 27298 96824 27304 96836
rect 27356 96824 27362 96876
rect 27850 96824 27856 96876
rect 27908 96864 27914 96876
rect 30058 96864 30064 96876
rect 27908 96836 30064 96864
rect 27908 96824 27914 96836
rect 30058 96824 30064 96836
rect 30116 96824 30122 96876
rect 41650 96824 41656 96876
rect 41708 96864 41714 96876
rect 47170 96864 47176 96876
rect 41708 96836 47176 96864
rect 41708 96824 41714 96836
rect 47170 96824 47176 96836
rect 47228 96824 47234 96876
rect 51402 96824 51408 96876
rect 51460 96864 51466 96876
rect 53794 96864 53800 96876
rect 51460 96836 53800 96864
rect 51460 96824 51466 96836
rect 53794 96824 53800 96836
rect 53852 96824 53858 96876
rect 84890 96824 84896 96876
rect 84948 96864 84954 96876
rect 88386 96864 88392 96876
rect 84948 96836 88392 96864
rect 84948 96824 84954 96836
rect 88386 96824 88392 96836
rect 88444 96824 88450 96876
rect 127026 96824 127032 96876
rect 127084 96864 127090 96876
rect 128774 96864 128780 96876
rect 127084 96836 128780 96864
rect 127084 96824 127090 96836
rect 128774 96824 128780 96836
rect 128832 96824 128838 96876
rect 185262 96824 185268 96876
rect 185320 96864 185326 96876
rect 190414 96864 190420 96876
rect 185320 96836 190420 96864
rect 185320 96824 185326 96836
rect 190414 96824 190420 96836
rect 190472 96824 190478 96876
rect 22330 96756 22336 96808
rect 22388 96796 22394 96808
rect 26197 96799 26255 96805
rect 26197 96796 26209 96799
rect 22388 96768 26209 96796
rect 22388 96756 22394 96768
rect 26197 96765 26209 96768
rect 26243 96765 26255 96799
rect 26197 96759 26255 96765
rect 38430 96756 38436 96808
rect 38488 96796 38494 96808
rect 41742 96796 41748 96808
rect 38488 96768 41748 96796
rect 38488 96756 38494 96768
rect 41742 96756 41748 96768
rect 41800 96756 41806 96808
rect 108718 96756 108724 96808
rect 108776 96796 108782 96808
rect 112030 96796 112036 96808
rect 108776 96768 112036 96796
rect 108776 96756 108782 96768
rect 112030 96756 112036 96768
rect 112088 96756 112094 96808
rect 175234 96756 175240 96808
rect 175292 96796 175298 96808
rect 176154 96796 176160 96808
rect 175292 96768 176160 96796
rect 175292 96756 175298 96768
rect 176154 96756 176160 96768
rect 176212 96756 176218 96808
rect 180478 96756 180484 96808
rect 180536 96796 180542 96808
rect 182226 96796 182232 96808
rect 180536 96768 182232 96796
rect 180536 96756 180542 96768
rect 182226 96756 182232 96768
rect 182284 96756 182290 96808
rect 182870 96756 182876 96808
rect 182928 96796 182934 96808
rect 187010 96796 187016 96808
rect 182928 96768 187016 96796
rect 182928 96756 182934 96768
rect 187010 96756 187016 96768
rect 187068 96756 187074 96808
rect 84430 96688 84436 96740
rect 84488 96728 84494 96740
rect 88202 96728 88208 96740
rect 84488 96700 88208 96728
rect 84488 96688 84494 96700
rect 88202 96688 88208 96700
rect 88260 96688 88266 96740
rect 108994 96688 109000 96740
rect 109052 96728 109058 96740
rect 112582 96728 112588 96740
rect 109052 96700 112588 96728
rect 109052 96688 109058 96700
rect 112582 96688 112588 96700
rect 112640 96688 112646 96740
rect 181674 96688 181680 96740
rect 181732 96728 181738 96740
rect 185170 96728 185176 96740
rect 181732 96700 185176 96728
rect 181732 96688 181738 96700
rect 185170 96688 185176 96700
rect 185228 96688 185234 96740
rect 175602 96620 175608 96672
rect 175660 96660 175666 96672
rect 176706 96660 176712 96672
rect 175660 96632 176712 96660
rect 175660 96620 175666 96632
rect 176706 96620 176712 96632
rect 176764 96620 176770 96672
rect 83786 96552 83792 96604
rect 83844 96592 83850 96604
rect 88478 96592 88484 96604
rect 83844 96564 88484 96592
rect 83844 96552 83850 96564
rect 88478 96552 88484 96564
rect 88536 96552 88542 96604
rect 180846 96552 180852 96604
rect 180904 96592 180910 96604
rect 184158 96592 184164 96604
rect 180904 96564 184164 96592
rect 180904 96552 180910 96564
rect 184158 96552 184164 96564
rect 184216 96552 184222 96604
rect 50666 96484 50672 96536
rect 50724 96524 50730 96536
rect 58210 96524 58216 96536
rect 50724 96496 58216 96524
rect 50724 96484 50730 96496
rect 58210 96484 58216 96496
rect 58268 96484 58274 96536
rect 82682 96484 82688 96536
rect 82740 96524 82746 96536
rect 89674 96524 89680 96536
rect 82740 96496 89680 96524
rect 82740 96484 82746 96496
rect 89674 96484 89680 96496
rect 89732 96484 89738 96536
rect 109546 96484 109552 96536
rect 109604 96524 109610 96536
rect 113502 96524 113508 96536
rect 109604 96496 113508 96524
rect 109604 96484 109610 96496
rect 113502 96484 113508 96496
rect 113560 96484 113566 96536
rect 182410 96484 182416 96536
rect 182468 96524 182474 96536
rect 184434 96524 184440 96536
rect 182468 96496 184440 96524
rect 182468 96484 182474 96496
rect 184434 96484 184440 96496
rect 184492 96484 184498 96536
rect 39626 96416 39632 96468
rect 39684 96456 39690 96468
rect 43766 96456 43772 96468
rect 39684 96428 43772 96456
rect 39684 96416 39690 96428
rect 43766 96416 43772 96428
rect 43824 96416 43830 96468
rect 53978 96416 53984 96468
rect 54036 96456 54042 96468
rect 77162 96456 77168 96468
rect 54036 96428 77168 96456
rect 54036 96416 54042 96428
rect 77162 96416 77168 96428
rect 77220 96416 77226 96468
rect 79370 96416 79376 96468
rect 79428 96456 79434 96468
rect 88570 96456 88576 96468
rect 79428 96428 88576 96456
rect 79428 96416 79434 96428
rect 88570 96416 88576 96428
rect 88628 96416 88634 96468
rect 109914 96416 109920 96468
rect 109972 96456 109978 96468
rect 113686 96456 113692 96468
rect 109972 96428 113692 96456
rect 109972 96416 109978 96428
rect 113686 96416 113692 96428
rect 113744 96416 113750 96468
rect 113962 96416 113968 96468
rect 114020 96456 114026 96468
rect 119206 96456 119212 96468
rect 114020 96428 119212 96456
rect 114020 96416 114026 96428
rect 119206 96416 119212 96428
rect 119264 96416 119270 96468
rect 125738 96416 125744 96468
rect 125796 96456 125802 96468
rect 148830 96456 148836 96468
rect 125796 96428 148836 96456
rect 125796 96416 125802 96428
rect 148830 96416 148836 96428
rect 148888 96416 148894 96468
rect 151682 96416 151688 96468
rect 151740 96456 151746 96468
rect 160330 96456 160336 96468
rect 151740 96428 160336 96456
rect 151740 96416 151746 96428
rect 160330 96416 160336 96428
rect 160388 96416 160394 96468
rect 23618 96348 23624 96400
rect 23676 96388 23682 96400
rect 26470 96388 26476 96400
rect 23676 96360 26476 96388
rect 23676 96348 23682 96360
rect 26470 96348 26476 96360
rect 26528 96348 26534 96400
rect 110558 96348 110564 96400
rect 110616 96388 110622 96400
rect 114790 96388 114796 96400
rect 110616 96360 114796 96388
rect 110616 96348 110622 96360
rect 114790 96348 114796 96360
rect 114848 96348 114854 96400
rect 25090 96280 25096 96332
rect 25148 96320 25154 96332
rect 28494 96320 28500 96332
rect 25148 96292 28500 96320
rect 25148 96280 25154 96292
rect 28494 96280 28500 96292
rect 28552 96280 28558 96332
rect 40086 96280 40092 96332
rect 40144 96320 40150 96332
rect 44410 96320 44416 96332
rect 40144 96292 44416 96320
rect 40144 96280 40150 96292
rect 44410 96280 44416 96292
rect 44468 96280 44474 96332
rect 110282 96280 110288 96332
rect 110340 96320 110346 96332
rect 114238 96320 114244 96332
rect 110340 96292 114244 96320
rect 110340 96280 110346 96292
rect 114238 96280 114244 96292
rect 114296 96280 114302 96332
rect 156098 96280 156104 96332
rect 156156 96320 156162 96332
rect 160238 96320 160244 96332
rect 156156 96292 160244 96320
rect 156156 96280 156162 96292
rect 160238 96280 160244 96292
rect 160296 96280 160302 96332
rect 39258 96212 39264 96264
rect 39316 96252 39322 96264
rect 43030 96252 43036 96264
rect 39316 96224 43036 96252
rect 39316 96212 39322 96224
rect 43030 96212 43036 96224
rect 43088 96212 43094 96264
rect 111110 96212 111116 96264
rect 111168 96252 111174 96264
rect 115342 96252 115348 96264
rect 111168 96224 115348 96252
rect 111168 96212 111174 96224
rect 115342 96212 115348 96224
rect 115400 96212 115406 96264
rect 157202 96212 157208 96264
rect 157260 96252 157266 96264
rect 160146 96252 160152 96264
rect 157260 96224 160152 96252
rect 157260 96212 157266 96224
rect 160146 96212 160152 96224
rect 160204 96212 160210 96264
rect 35302 96144 35308 96196
rect 35360 96184 35366 96196
rect 36314 96184 36320 96196
rect 35360 96156 36320 96184
rect 35360 96144 35366 96156
rect 36314 96144 36320 96156
rect 36372 96144 36378 96196
rect 111478 96144 111484 96196
rect 111536 96184 111542 96196
rect 116262 96184 116268 96196
rect 111536 96156 116268 96184
rect 111536 96144 111542 96156
rect 116262 96144 116268 96156
rect 116320 96144 116326 96196
rect 111938 96076 111944 96128
rect 111996 96116 112002 96128
rect 116446 96116 116452 96128
rect 111996 96088 116452 96116
rect 111996 96076 112002 96088
rect 116446 96076 116452 96088
rect 116504 96076 116510 96128
rect 184434 96076 184440 96128
rect 184492 96116 184498 96128
rect 189218 96116 189224 96128
rect 184492 96088 189224 96116
rect 184492 96076 184498 96088
rect 189218 96076 189224 96088
rect 189276 96076 189282 96128
rect 102278 96008 102284 96060
rect 102336 96048 102342 96060
rect 103198 96048 103204 96060
rect 102336 96020 103204 96048
rect 102336 96008 102342 96020
rect 103198 96008 103204 96020
rect 103256 96008 103262 96060
rect 112674 96008 112680 96060
rect 112732 96048 112738 96060
rect 117550 96048 117556 96060
rect 112732 96020 117556 96048
rect 112732 96008 112738 96020
rect 117550 96008 117556 96020
rect 117608 96008 117614 96060
rect 100254 95940 100260 95992
rect 100312 95980 100318 95992
rect 100438 95980 100444 95992
rect 100312 95952 100444 95980
rect 100312 95940 100318 95952
rect 100438 95940 100444 95952
rect 100496 95940 100502 95992
rect 101910 95940 101916 95992
rect 101968 95980 101974 95992
rect 102646 95980 102652 95992
rect 101968 95952 102652 95980
rect 101968 95940 101974 95952
rect 102646 95940 102652 95952
rect 102704 95940 102710 95992
rect 103106 95940 103112 95992
rect 103164 95980 103170 95992
rect 104302 95980 104308 95992
rect 103164 95952 104308 95980
rect 103164 95940 103170 95952
rect 104302 95940 104308 95952
rect 104360 95940 104366 95992
rect 113134 95940 113140 95992
rect 113192 95980 113198 95992
rect 118102 95980 118108 95992
rect 113192 95952 118108 95980
rect 113192 95940 113198 95952
rect 118102 95940 118108 95952
rect 118160 95940 118166 95992
rect 159410 95940 159416 95992
rect 159468 95980 159474 95992
rect 161526 95980 161532 95992
rect 159468 95952 161532 95980
rect 159468 95940 159474 95952
rect 161526 95940 161532 95952
rect 161584 95940 161590 95992
rect 183606 95940 183612 95992
rect 183664 95980 183670 95992
rect 188114 95980 188120 95992
rect 183664 95952 188120 95980
rect 183664 95940 183670 95952
rect 188114 95940 188120 95952
rect 188172 95940 188178 95992
rect 101450 95872 101456 95924
rect 101508 95912 101514 95924
rect 102370 95912 102376 95924
rect 101508 95884 102376 95912
rect 101508 95872 101514 95884
rect 102370 95872 102376 95884
rect 102428 95872 102434 95924
rect 102738 95872 102744 95924
rect 102796 95912 102802 95924
rect 103934 95912 103940 95924
rect 102796 95884 103940 95912
rect 102796 95872 102802 95884
rect 103934 95872 103940 95884
rect 103992 95872 103998 95924
rect 112306 95872 112312 95924
rect 112364 95912 112370 95924
rect 116998 95912 117004 95924
rect 112364 95884 117004 95912
rect 112364 95872 112370 95884
rect 116998 95872 117004 95884
rect 117056 95872 117062 95924
rect 178822 95872 178828 95924
rect 178880 95912 178886 95924
rect 180938 95912 180944 95924
rect 178880 95884 180944 95912
rect 178880 95872 178886 95884
rect 180938 95872 180944 95884
rect 180996 95872 181002 95924
rect 183238 95872 183244 95924
rect 183296 95912 183302 95924
rect 187562 95912 187568 95924
rect 183296 95884 187568 95912
rect 183296 95872 183302 95884
rect 187562 95872 187568 95884
rect 187620 95872 187626 95924
rect 26562 95804 26568 95856
rect 26620 95844 26626 95856
rect 29230 95844 29236 95856
rect 26620 95816 29236 95844
rect 26620 95804 26626 95816
rect 29230 95804 29236 95816
rect 29288 95804 29294 95856
rect 101542 95844 101548 95856
rect 100824 95816 101548 95844
rect 100824 95776 100852 95816
rect 101542 95804 101548 95816
rect 101600 95804 101606 95856
rect 104302 95804 104308 95856
rect 104360 95844 104366 95856
rect 105958 95844 105964 95856
rect 104360 95816 105964 95844
rect 104360 95804 104366 95816
rect 105958 95804 105964 95816
rect 106016 95804 106022 95856
rect 106694 95804 106700 95856
rect 106752 95844 106758 95856
rect 109178 95844 109184 95856
rect 106752 95816 109184 95844
rect 106752 95804 106758 95816
rect 109178 95804 109184 95816
rect 109236 95804 109242 95856
rect 113226 95804 113232 95856
rect 113284 95844 113290 95856
rect 118838 95844 118844 95856
rect 113284 95816 118844 95844
rect 113284 95804 113290 95816
rect 118838 95804 118844 95816
rect 118896 95804 118902 95856
rect 179282 95804 179288 95856
rect 179340 95844 179346 95856
rect 179742 95844 179748 95856
rect 179340 95816 179748 95844
rect 179340 95804 179346 95816
rect 179742 95804 179748 95816
rect 179800 95804 179806 95856
rect 100824 95748 101036 95776
rect 101008 95720 101036 95748
rect 100990 95668 100996 95720
rect 101048 95668 101054 95720
rect 164102 94308 164108 94360
rect 164160 94348 164166 94360
rect 168150 94348 168156 94360
rect 164160 94320 168156 94348
rect 164160 94308 164166 94320
rect 168150 94308 168156 94320
rect 168208 94308 168214 94360
rect 91698 94036 91704 94088
rect 91756 94076 91762 94088
rect 95470 94076 95476 94088
rect 91756 94048 95476 94076
rect 91756 94036 91762 94048
rect 95470 94036 95476 94048
rect 95528 94036 95534 94088
rect 91054 92268 91060 92320
rect 91112 92308 91118 92320
rect 118930 92308 118936 92320
rect 91112 92280 118936 92308
rect 91112 92268 91118 92280
rect 118930 92268 118936 92280
rect 118988 92268 118994 92320
rect 91790 91656 91796 91708
rect 91848 91696 91854 91708
rect 95286 91696 95292 91708
rect 91848 91668 95292 91696
rect 91848 91656 91854 91668
rect 95286 91656 95292 91668
rect 95344 91656 95350 91708
rect 188114 91588 188120 91640
rect 188172 91628 188178 91640
rect 198234 91628 198240 91640
rect 188172 91600 198240 91628
rect 188172 91588 188178 91600
rect 198234 91588 198240 91600
rect 198292 91588 198298 91640
rect 91514 91316 91520 91368
rect 91572 91356 91578 91368
rect 93354 91356 93360 91368
rect 91572 91328 93360 91356
rect 91572 91316 91578 91328
rect 93354 91316 93360 91328
rect 93412 91316 93418 91368
rect 163550 91112 163556 91164
rect 163608 91152 163614 91164
rect 165942 91152 165948 91164
rect 163608 91124 165948 91152
rect 163608 91112 163614 91124
rect 165942 91112 165948 91124
rect 166000 91112 166006 91164
rect 188574 90228 188580 90280
rect 188632 90268 188638 90280
rect 197590 90268 197596 90280
rect 188632 90240 197596 90268
rect 188632 90228 188638 90240
rect 197590 90228 197596 90240
rect 197648 90228 197654 90280
rect 18098 90160 18104 90212
rect 18156 90200 18162 90212
rect 22330 90200 22336 90212
rect 18156 90172 22336 90200
rect 18156 90160 18162 90172
rect 22330 90160 22336 90172
rect 22388 90160 22394 90212
rect 163826 90092 163832 90144
rect 163884 90132 163890 90144
rect 166034 90132 166040 90144
rect 163884 90104 166040 90132
rect 163884 90092 163890 90104
rect 166034 90092 166040 90104
rect 166092 90092 166098 90144
rect 92250 88868 92256 88920
rect 92308 88908 92314 88920
rect 95378 88908 95384 88920
rect 92308 88880 95384 88908
rect 92308 88868 92314 88880
rect 95378 88868 95384 88880
rect 95436 88868 95442 88920
rect 163458 88732 163464 88784
rect 163516 88772 163522 88784
rect 165114 88772 165120 88784
rect 163516 88744 165120 88772
rect 163516 88732 163522 88744
rect 165114 88732 165120 88744
rect 165172 88732 165178 88784
rect 92158 87508 92164 87560
rect 92216 87548 92222 87560
rect 95378 87548 95384 87560
rect 92216 87520 95384 87548
rect 92216 87508 92222 87520
rect 95378 87508 95384 87520
rect 95436 87508 95442 87560
rect 188114 84652 188120 84704
rect 188172 84692 188178 84704
rect 196946 84692 196952 84704
rect 188172 84664 196952 84692
rect 188172 84652 188178 84664
rect 196946 84652 196952 84664
rect 197004 84652 197010 84704
rect 163918 84312 163924 84364
rect 163976 84352 163982 84364
rect 167322 84352 167328 84364
rect 163976 84324 167328 84352
rect 163976 84312 163982 84324
rect 167322 84312 167328 84324
rect 167380 84312 167386 84364
rect 116538 83564 116544 83616
rect 116596 83604 116602 83616
rect 119574 83604 119580 83616
rect 116596 83576 119580 83604
rect 116596 83564 116602 83576
rect 119574 83564 119580 83576
rect 119632 83564 119638 83616
rect 163918 82680 163924 82732
rect 163976 82720 163982 82732
rect 167874 82720 167880 82732
rect 163976 82692 167880 82720
rect 163976 82680 163982 82692
rect 167874 82680 167880 82692
rect 167932 82680 167938 82732
rect 13222 82272 13228 82324
rect 13280 82312 13286 82324
rect 15430 82312 15436 82324
rect 13280 82284 15436 82312
rect 13280 82272 13286 82284
rect 15430 82272 15436 82284
rect 15488 82272 15494 82324
rect 13314 81932 13320 81984
rect 13372 81972 13378 81984
rect 22330 81972 22336 81984
rect 13372 81944 22336 81972
rect 13372 81932 13378 81944
rect 22330 81932 22336 81944
rect 22388 81932 22394 81984
rect 163550 81932 163556 81984
rect 163608 81972 163614 81984
rect 167230 81972 167236 81984
rect 163608 81944 167236 81972
rect 163608 81932 163614 81944
rect 167230 81932 167236 81944
rect 167288 81932 167294 81984
rect 91790 80504 91796 80556
rect 91848 80544 91854 80556
rect 94274 80544 94280 80556
rect 91848 80516 94280 80544
rect 91848 80504 91854 80516
rect 94274 80504 94280 80516
rect 94332 80504 94338 80556
rect 164102 80436 164108 80488
rect 164160 80476 164166 80488
rect 167322 80476 167328 80488
rect 164160 80448 167328 80476
rect 164160 80436 164166 80448
rect 167322 80436 167328 80448
rect 167380 80436 167386 80488
rect 164378 78940 164384 78992
rect 164436 78980 164442 78992
rect 167230 78980 167236 78992
rect 164436 78952 167236 78980
rect 164436 78940 164442 78952
rect 167230 78940 167236 78952
rect 167288 78940 167294 78992
rect 91422 78804 91428 78856
rect 91480 78844 91486 78856
rect 95286 78844 95292 78856
rect 91480 78816 95292 78844
rect 91480 78804 91486 78816
rect 95286 78804 95292 78816
rect 95344 78804 95350 78856
rect 167230 77892 167236 77904
rect 164488 77864 167236 77892
rect 164102 77784 164108 77836
rect 164160 77824 164166 77836
rect 164488 77824 164516 77864
rect 167230 77852 167236 77864
rect 167288 77852 167294 77904
rect 164160 77796 164516 77824
rect 164160 77784 164166 77796
rect 91698 77444 91704 77496
rect 91756 77484 91762 77496
rect 95378 77484 95384 77496
rect 91756 77456 95384 77484
rect 91756 77444 91762 77456
rect 95378 77444 95384 77456
rect 95436 77444 95442 77496
rect 167230 76464 167236 76476
rect 164488 76436 167236 76464
rect 163734 76356 163740 76408
rect 163792 76396 163798 76408
rect 164488 76396 164516 76436
rect 167230 76424 167236 76436
rect 167288 76424 167294 76476
rect 163792 76368 164516 76396
rect 163792 76356 163798 76368
rect 91698 76220 91704 76272
rect 91756 76260 91762 76272
rect 94918 76260 94924 76272
rect 91756 76232 94924 76260
rect 91756 76220 91762 76232
rect 94918 76220 94924 76232
rect 94976 76220 94982 76272
rect 15430 74996 15436 75048
rect 15488 75036 15494 75048
rect 22330 75036 22336 75048
rect 15488 75008 22336 75036
rect 15488 74996 15494 75008
rect 22330 74996 22336 75008
rect 22388 74996 22394 75048
rect 45054 74996 45060 75048
rect 45112 75036 45118 75048
rect 47814 75036 47820 75048
rect 45112 75008 47820 75036
rect 45112 74996 45118 75008
rect 47814 74996 47820 75008
rect 47872 74996 47878 75048
rect 164102 74928 164108 74980
rect 164160 74968 164166 74980
rect 167230 74968 167236 74980
rect 164160 74940 167236 74968
rect 164160 74928 164166 74940
rect 167230 74928 167236 74940
rect 167288 74928 167294 74980
rect 164378 73704 164384 73756
rect 164436 73744 164442 73756
rect 167138 73744 167144 73756
rect 164436 73716 167144 73744
rect 164436 73704 164442 73716
rect 167138 73704 167144 73716
rect 167196 73704 167202 73756
rect 91698 72480 91704 72532
rect 91756 72520 91762 72532
rect 95378 72520 95384 72532
rect 91756 72492 95384 72520
rect 91756 72480 91762 72492
rect 95378 72480 95384 72492
rect 95436 72480 95442 72532
rect 164378 72480 164384 72532
rect 164436 72520 164442 72532
rect 167230 72520 167236 72532
rect 164436 72492 167236 72520
rect 164436 72480 164442 72492
rect 167230 72480 167236 72492
rect 167288 72480 167294 72532
rect 91698 71256 91704 71308
rect 91756 71296 91762 71308
rect 95378 71296 95384 71308
rect 91756 71268 95384 71296
rect 91756 71256 91762 71268
rect 95378 71256 95384 71268
rect 95436 71256 95442 71308
rect 164378 71120 164384 71172
rect 164436 71160 164442 71172
rect 167322 71160 167328 71172
rect 164436 71132 167328 71160
rect 164436 71120 164442 71132
rect 167322 71120 167328 71132
rect 167380 71120 167386 71172
rect 163550 69896 163556 69948
rect 163608 69936 163614 69948
rect 167230 69936 167236 69948
rect 163608 69908 167236 69936
rect 163608 69896 163614 69908
rect 167230 69896 167236 69908
rect 167288 69896 167294 69948
rect 91422 69556 91428 69608
rect 91480 69596 91486 69608
rect 93998 69596 94004 69608
rect 91480 69568 94004 69596
rect 91480 69556 91486 69568
rect 93998 69556 94004 69568
rect 94056 69556 94062 69608
rect 91422 68672 91428 68724
rect 91480 68712 91486 68724
rect 93906 68712 93912 68724
rect 91480 68684 93912 68712
rect 91480 68672 91486 68684
rect 93906 68672 93912 68684
rect 93964 68672 93970 68724
rect 163734 68196 163740 68248
rect 163792 68236 163798 68248
rect 167322 68236 167328 68248
rect 163792 68208 167328 68236
rect 163792 68196 163798 68208
rect 167322 68196 167328 68208
rect 167380 68196 167386 68248
rect 189954 67448 189960 67500
rect 190012 67488 190018 67500
rect 190598 67488 190604 67500
rect 190012 67460 190604 67488
rect 190012 67448 190018 67460
rect 190598 67448 190604 67460
rect 190656 67488 190662 67500
rect 197590 67488 197596 67500
rect 190656 67460 197596 67488
rect 190656 67448 190662 67460
rect 197590 67448 197596 67460
rect 197648 67448 197654 67500
rect 91514 66768 91520 66820
rect 91572 66808 91578 66820
rect 93630 66808 93636 66820
rect 91572 66780 93636 66808
rect 91572 66768 91578 66780
rect 93630 66768 93636 66780
rect 93688 66768 93694 66820
rect 164378 66768 164384 66820
rect 164436 66808 164442 66820
rect 167874 66808 167880 66820
rect 164436 66780 167880 66808
rect 164436 66768 164442 66780
rect 167874 66768 167880 66780
rect 167932 66768 167938 66820
rect 44410 65408 44416 65460
rect 44468 65448 44474 65460
rect 47170 65448 47176 65460
rect 44468 65420 47176 65448
rect 44468 65408 44474 65420
rect 47170 65408 47176 65420
rect 47228 65408 47234 65460
rect 164378 65408 164384 65460
rect 164436 65448 164442 65460
rect 167138 65448 167144 65460
rect 164436 65420 167144 65448
rect 164436 65408 164442 65420
rect 167138 65408 167144 65420
rect 167196 65408 167202 65460
rect 164378 64456 164384 64508
rect 164436 64496 164442 64508
rect 167046 64496 167052 64508
rect 164436 64468 167052 64496
rect 164436 64456 164442 64468
rect 167046 64456 167052 64468
rect 167104 64456 167110 64508
rect 92618 64048 92624 64100
rect 92676 64088 92682 64100
rect 93538 64088 93544 64100
rect 92676 64060 93544 64088
rect 92676 64048 92682 64060
rect 93538 64048 93544 64060
rect 93596 64048 93602 64100
rect 164378 64048 164384 64100
rect 164436 64088 164442 64100
rect 166494 64088 166500 64100
rect 164436 64060 166500 64088
rect 164436 64048 164442 64060
rect 166494 64048 166500 64060
rect 166552 64048 166558 64100
rect 117458 62620 117464 62672
rect 117516 62660 117522 62672
rect 119482 62660 119488 62672
rect 117516 62632 119488 62660
rect 117516 62620 117522 62632
rect 119482 62620 119488 62632
rect 119540 62620 119546 62672
rect 13314 62552 13320 62604
rect 13372 62592 13378 62604
rect 22698 62592 22704 62604
rect 13372 62564 22704 62592
rect 13372 62552 13378 62564
rect 22698 62552 22704 62564
rect 22756 62552 22762 62604
rect 91422 61260 91428 61312
rect 91480 61300 91486 61312
rect 93446 61300 93452 61312
rect 91480 61272 93452 61300
rect 91480 61260 91486 61272
rect 93446 61260 93452 61272
rect 93504 61260 93510 61312
rect 92526 59696 92532 59748
rect 92584 59736 92590 59748
rect 94090 59736 94096 59748
rect 92584 59708 94096 59736
rect 92584 59696 92590 59708
rect 94090 59696 94096 59708
rect 94148 59696 94154 59748
rect 91514 58540 91520 58592
rect 91572 58580 91578 58592
rect 93630 58580 93636 58592
rect 91572 58552 93636 58580
rect 91572 58540 91578 58552
rect 93630 58540 93636 58552
rect 93688 58540 93694 58592
rect 164378 58540 164384 58592
rect 164436 58580 164442 58592
rect 166034 58580 166040 58592
rect 164436 58552 166040 58580
rect 164436 58540 164442 58552
rect 166034 58540 166040 58552
rect 166092 58540 166098 58592
rect 92342 58472 92348 58524
rect 92400 58512 92406 58524
rect 95194 58512 95200 58524
rect 92400 58484 95200 58512
rect 92400 58472 92406 58484
rect 95194 58472 95200 58484
rect 95252 58472 95258 58524
rect 187930 57928 187936 57980
rect 187988 57968 187994 57980
rect 189954 57968 189960 57980
rect 187988 57940 189960 57968
rect 187988 57928 187994 57940
rect 189954 57928 189960 57940
rect 190012 57928 190018 57980
rect 164378 57112 164384 57164
rect 164436 57152 164442 57164
rect 165942 57152 165948 57164
rect 164436 57124 165948 57152
rect 164436 57112 164442 57124
rect 165942 57112 165948 57124
rect 166000 57112 166006 57164
rect 74681 51579 74739 51585
rect 74681 51545 74693 51579
rect 74727 51576 74739 51579
rect 82130 51576 82136 51588
rect 74727 51548 82136 51576
rect 74727 51545 74739 51548
rect 74681 51539 74739 51545
rect 82130 51536 82136 51548
rect 82188 51536 82194 51588
rect 84338 51536 84344 51588
rect 84396 51576 84402 51588
rect 145150 51576 145156 51588
rect 84396 51548 145156 51576
rect 84396 51536 84402 51548
rect 145150 51536 145156 51548
rect 145208 51536 145214 51588
rect 173946 51536 173952 51588
rect 174004 51576 174010 51588
rect 174130 51576 174136 51588
rect 174004 51548 174136 51576
rect 174004 51536 174010 51548
rect 174130 51536 174136 51548
rect 174188 51536 174194 51588
rect 175234 51536 175240 51588
rect 175292 51576 175298 51588
rect 176154 51576 176160 51588
rect 175292 51548 176160 51576
rect 175292 51536 175298 51548
rect 176154 51536 176160 51548
rect 176212 51536 176218 51588
rect 98230 51468 98236 51520
rect 98288 51508 98294 51520
rect 98966 51508 98972 51520
rect 98288 51480 98972 51508
rect 98288 51468 98294 51480
rect 98966 51468 98972 51480
rect 99024 51468 99030 51520
rect 103382 51468 103388 51520
rect 103440 51508 103446 51520
rect 103842 51508 103848 51520
rect 103440 51480 103848 51508
rect 103440 51468 103446 51480
rect 103842 51468 103848 51480
rect 103900 51468 103906 51520
rect 105038 51468 105044 51520
rect 105096 51508 105102 51520
rect 106142 51508 106148 51520
rect 105096 51480 106148 51508
rect 105096 51468 105102 51480
rect 106142 51468 106148 51480
rect 106200 51468 106206 51520
rect 106326 51468 106332 51520
rect 106384 51508 106390 51520
rect 107798 51508 107804 51520
rect 106384 51480 107804 51508
rect 106384 51468 106390 51480
rect 107798 51468 107804 51480
rect 107856 51468 107862 51520
rect 111478 51468 111484 51520
rect 111536 51508 111542 51520
rect 112398 51508 112404 51520
rect 111536 51480 112404 51508
rect 111536 51468 111542 51480
rect 112398 51468 112404 51480
rect 112456 51468 112462 51520
rect 113134 51468 113140 51520
rect 113192 51508 113198 51520
rect 114606 51508 114612 51520
rect 113192 51480 114612 51508
rect 113192 51468 113198 51480
rect 114606 51468 114612 51480
rect 114664 51468 114670 51520
rect 174866 51468 174872 51520
rect 174924 51508 174930 51520
rect 175510 51508 175516 51520
rect 174924 51480 175516 51508
rect 174924 51468 174930 51480
rect 175510 51468 175516 51480
rect 175568 51468 175574 51520
rect 72010 51400 72016 51452
rect 72068 51440 72074 51452
rect 73206 51440 73212 51452
rect 72068 51412 73212 51440
rect 72068 51400 72074 51412
rect 73206 51400 73212 51412
rect 73264 51440 73270 51452
rect 83602 51440 83608 51452
rect 73264 51412 83608 51440
rect 73264 51400 73270 51412
rect 83602 51400 83608 51412
rect 83660 51440 83666 51452
rect 84338 51440 84344 51452
rect 83660 51412 84344 51440
rect 83660 51400 83666 51412
rect 84338 51400 84344 51412
rect 84396 51400 84402 51452
rect 96761 51443 96819 51449
rect 96761 51409 96773 51443
rect 96807 51440 96819 51443
rect 96807 51412 99702 51440
rect 96807 51409 96819 51412
rect 96761 51403 96819 51409
rect 66582 51332 66588 51384
rect 66640 51372 66646 51384
rect 74681 51375 74739 51381
rect 74681 51372 74693 51375
rect 66640 51344 74693 51372
rect 66640 51332 66646 51344
rect 74681 51341 74693 51344
rect 74727 51341 74739 51375
rect 74681 51335 74739 51341
rect 82130 51264 82136 51316
rect 82188 51304 82194 51316
rect 87193 51307 87251 51313
rect 87193 51304 87205 51307
rect 82188 51276 87205 51304
rect 82188 51264 82194 51276
rect 87193 51273 87205 51276
rect 87239 51273 87251 51307
rect 87193 51267 87251 51273
rect 87193 51171 87251 51177
rect 87193 51137 87205 51171
rect 87239 51168 87251 51171
rect 96761 51171 96819 51177
rect 96761 51168 96773 51171
rect 87239 51140 96773 51168
rect 87239 51137 87251 51140
rect 87193 51131 87251 51137
rect 96761 51137 96773 51140
rect 96807 51137 96819 51171
rect 99674 51168 99702 51412
rect 105498 51400 105504 51452
rect 105556 51440 105562 51452
rect 106694 51440 106700 51452
rect 105556 51412 106700 51440
rect 105556 51400 105562 51412
rect 106694 51400 106700 51412
rect 106752 51400 106758 51452
rect 107154 51400 107160 51452
rect 107212 51440 107218 51452
rect 108902 51440 108908 51452
rect 107212 51412 108908 51440
rect 107212 51400 107218 51412
rect 108902 51400 108908 51412
rect 108960 51400 108966 51452
rect 110282 51400 110288 51452
rect 110340 51440 110346 51452
rect 111754 51440 111760 51452
rect 110340 51412 111760 51440
rect 110340 51400 110346 51412
rect 111754 51400 111760 51412
rect 111812 51400 111818 51452
rect 112674 51400 112680 51452
rect 112732 51440 112738 51452
rect 114698 51440 114704 51452
rect 112732 51412 114704 51440
rect 112732 51400 112738 51412
rect 114698 51400 114704 51412
rect 114756 51400 114762 51452
rect 116173 51443 116231 51449
rect 116173 51409 116185 51443
rect 116219 51440 116231 51443
rect 125741 51443 125799 51449
rect 125741 51440 125753 51443
rect 116219 51412 125753 51440
rect 116219 51409 116231 51412
rect 116173 51403 116231 51409
rect 125741 51409 125753 51412
rect 125787 51409 125799 51443
rect 125741 51403 125799 51409
rect 105958 51332 105964 51384
rect 106016 51372 106022 51384
rect 107246 51372 107252 51384
rect 106016 51344 107252 51372
rect 106016 51332 106022 51344
rect 107246 51332 107252 51344
rect 107304 51332 107310 51384
rect 128792 51344 138204 51372
rect 106602 51264 106608 51316
rect 106660 51304 106666 51316
rect 108442 51304 108448 51316
rect 106660 51276 108448 51304
rect 106660 51264 106666 51276
rect 108442 51264 108448 51276
rect 108500 51264 108506 51316
rect 125741 51307 125799 51313
rect 125741 51273 125753 51307
rect 125787 51304 125799 51307
rect 128501 51307 128559 51313
rect 128501 51304 128513 51307
rect 125787 51276 128513 51304
rect 125787 51273 125799 51276
rect 125741 51267 125799 51273
rect 128501 51273 128513 51276
rect 128547 51273 128559 51307
rect 128501 51267 128559 51273
rect 128593 51307 128651 51313
rect 128593 51273 128605 51307
rect 128639 51304 128651 51307
rect 128792 51304 128820 51344
rect 128639 51276 128820 51304
rect 138176 51304 138204 51344
rect 138342 51304 138348 51316
rect 138176 51276 138348 51304
rect 128639 51273 128651 51276
rect 128593 51267 128651 51273
rect 138342 51264 138348 51276
rect 138400 51264 138406 51316
rect 116173 51239 116231 51245
rect 106528 51208 116124 51236
rect 106528 51168 106556 51208
rect 99674 51140 106556 51168
rect 116096 51168 116124 51208
rect 116173 51205 116185 51239
rect 116219 51205 116231 51239
rect 116173 51199 116231 51205
rect 116188 51168 116216 51199
rect 116096 51140 116216 51168
rect 96761 51131 96819 51137
rect 40822 50992 40828 51044
rect 40880 51032 40886 51044
rect 42938 51032 42944 51044
rect 40880 51004 42944 51032
rect 40880 50992 40886 51004
rect 42938 50992 42944 51004
rect 42996 50992 43002 51044
rect 109546 50992 109552 51044
rect 109604 51032 109610 51044
rect 111846 51032 111852 51044
rect 109604 51004 111852 51032
rect 109604 50992 109610 51004
rect 111846 50992 111852 51004
rect 111904 50992 111910 51044
rect 112306 50992 112312 51044
rect 112364 51032 112370 51044
rect 114422 51032 114428 51044
rect 112364 51004 114428 51032
rect 112364 50992 112370 51004
rect 114422 50992 114428 51004
rect 114480 50992 114486 51044
rect 64558 50924 64564 50976
rect 64616 50964 64622 50976
rect 86546 50964 86552 50976
rect 64616 50936 86552 50964
rect 64616 50924 64622 50936
rect 86546 50924 86552 50936
rect 86604 50924 86610 50976
rect 13314 50856 13320 50908
rect 13372 50896 13378 50908
rect 72010 50896 72016 50908
rect 13372 50868 72016 50896
rect 13372 50856 13378 50868
rect 72010 50856 72016 50868
rect 72068 50856 72074 50908
rect 138158 50856 138164 50908
rect 138216 50896 138222 50908
rect 151590 50896 151596 50908
rect 138216 50868 151596 50896
rect 138216 50856 138222 50868
rect 151590 50856 151596 50868
rect 151648 50856 151654 50908
rect 36498 50788 36504 50840
rect 36556 50828 36562 50840
rect 38614 50828 38620 50840
rect 36556 50800 38620 50828
rect 36556 50788 36562 50800
rect 38614 50788 38620 50800
rect 38672 50788 38678 50840
rect 104670 50788 104676 50840
rect 104728 50828 104734 50840
rect 105498 50828 105504 50840
rect 104728 50800 105504 50828
rect 104728 50788 104734 50800
rect 105498 50788 105504 50800
rect 105556 50788 105562 50840
rect 36038 50720 36044 50772
rect 36096 50760 36102 50772
rect 37418 50760 37424 50772
rect 36096 50732 37424 50760
rect 36096 50720 36102 50732
rect 37418 50720 37424 50732
rect 37476 50720 37482 50772
rect 175602 50720 175608 50772
rect 175660 50760 175666 50772
rect 176706 50760 176712 50772
rect 175660 50732 176712 50760
rect 175660 50720 175666 50732
rect 176706 50720 176712 50732
rect 176764 50720 176770 50772
rect 182410 50720 182416 50772
rect 182468 50760 182474 50772
rect 184986 50760 184992 50772
rect 182468 50732 184992 50760
rect 182468 50720 182474 50732
rect 184986 50720 184992 50732
rect 185044 50720 185050 50772
rect 35302 50652 35308 50704
rect 35360 50692 35366 50704
rect 36498 50692 36504 50704
rect 35360 50664 36504 50692
rect 35360 50652 35366 50664
rect 36498 50652 36504 50664
rect 36556 50652 36562 50704
rect 180018 50652 180024 50704
rect 180076 50692 180082 50704
rect 182042 50692 182048 50704
rect 180076 50664 182048 50692
rect 180076 50652 180082 50664
rect 182042 50652 182048 50664
rect 182100 50652 182106 50704
rect 39258 50584 39264 50636
rect 39316 50624 39322 50636
rect 41374 50624 41380 50636
rect 39316 50596 41380 50624
rect 39316 50584 39322 50596
rect 41374 50584 41380 50596
rect 41432 50584 41438 50636
rect 178822 50584 178828 50636
rect 178880 50624 178886 50636
rect 180938 50624 180944 50636
rect 178880 50596 180944 50624
rect 178880 50584 178886 50596
rect 180938 50584 180944 50596
rect 180996 50584 181002 50636
rect 184066 50584 184072 50636
rect 184124 50624 184130 50636
rect 186274 50624 186280 50636
rect 184124 50596 186280 50624
rect 184124 50584 184130 50596
rect 186274 50584 186280 50596
rect 186332 50584 186338 50636
rect 38890 50516 38896 50568
rect 38948 50556 38954 50568
rect 40822 50556 40828 50568
rect 38948 50528 40828 50556
rect 38948 50516 38954 50528
rect 40822 50516 40828 50528
rect 40880 50516 40886 50568
rect 179650 50516 179656 50568
rect 179708 50556 179714 50568
rect 182318 50556 182324 50568
rect 179708 50528 182324 50556
rect 179708 50516 179714 50528
rect 182318 50516 182324 50528
rect 182376 50516 182382 50568
rect 183606 50516 183612 50568
rect 183664 50556 183670 50568
rect 188114 50556 188120 50568
rect 183664 50528 188120 50556
rect 183664 50516 183670 50528
rect 188114 50516 188120 50528
rect 188172 50516 188178 50568
rect 38062 50448 38068 50500
rect 38120 50488 38126 50500
rect 39718 50488 39724 50500
rect 38120 50460 39724 50488
rect 38120 50448 38126 50460
rect 39718 50448 39724 50460
rect 39776 50448 39782 50500
rect 111110 50448 111116 50500
rect 111168 50488 111174 50500
rect 112674 50488 112680 50500
rect 111168 50460 112680 50488
rect 111168 50448 111174 50460
rect 112674 50448 112680 50460
rect 112732 50448 112738 50500
rect 177258 50448 177264 50500
rect 177316 50488 177322 50500
rect 179006 50488 179012 50500
rect 177316 50460 179012 50488
rect 177316 50448 177322 50460
rect 179006 50448 179012 50460
rect 179064 50448 179070 50500
rect 181674 50448 181680 50500
rect 181732 50488 181738 50500
rect 183422 50488 183428 50500
rect 181732 50460 183428 50488
rect 181732 50448 181738 50460
rect 183422 50448 183428 50460
rect 183480 50448 183486 50500
rect 184434 50448 184440 50500
rect 184492 50488 184498 50500
rect 186458 50488 186464 50500
rect 184492 50460 186464 50488
rect 184492 50448 184498 50460
rect 186458 50448 186464 50460
rect 186516 50448 186522 50500
rect 37694 50380 37700 50432
rect 37752 50420 37758 50432
rect 40178 50420 40184 50432
rect 37752 50392 40184 50420
rect 37752 50380 37758 50392
rect 40178 50380 40184 50392
rect 40236 50380 40242 50432
rect 41650 50380 41656 50432
rect 41708 50420 41714 50432
rect 44042 50420 44048 50432
rect 41708 50392 44048 50420
rect 41708 50380 41714 50392
rect 44042 50380 44048 50392
rect 44100 50380 44106 50432
rect 109914 50380 109920 50432
rect 109972 50420 109978 50432
rect 109972 50392 111800 50420
rect 109972 50380 109978 50392
rect 27850 50312 27856 50364
rect 27908 50352 27914 50364
rect 30058 50352 30064 50364
rect 27908 50324 30064 50352
rect 27908 50312 27914 50324
rect 30058 50312 30064 50324
rect 30116 50312 30122 50364
rect 36866 50312 36872 50364
rect 36924 50352 36930 50364
rect 36924 50324 38844 50352
rect 36924 50312 36930 50324
rect 26102 50284 26108 50296
rect 23728 50256 26108 50284
rect 20858 50176 20864 50228
rect 20916 50216 20922 50228
rect 23728 50216 23756 50256
rect 26102 50244 26108 50256
rect 26160 50244 26166 50296
rect 26194 50244 26200 50296
rect 26252 50284 26258 50296
rect 26470 50284 26476 50296
rect 26252 50256 26476 50284
rect 26252 50244 26258 50256
rect 26470 50244 26476 50256
rect 26528 50244 26534 50296
rect 28862 50284 28868 50296
rect 27684 50256 28868 50284
rect 20916 50188 23756 50216
rect 20916 50176 20922 50188
rect 25642 50176 25648 50228
rect 25700 50216 25706 50228
rect 27684 50216 27712 50256
rect 28862 50244 28868 50256
rect 28920 50244 28926 50296
rect 30886 50284 30892 50296
rect 29248 50256 30892 50284
rect 25700 50188 27712 50216
rect 25700 50176 25706 50188
rect 29046 50176 29052 50228
rect 29104 50216 29110 50228
rect 29248 50216 29276 50256
rect 30886 50244 30892 50256
rect 30944 50244 30950 50296
rect 36130 50244 36136 50296
rect 36188 50284 36194 50296
rect 37234 50284 37240 50296
rect 36188 50256 37240 50284
rect 36188 50244 36194 50256
rect 37234 50244 37240 50256
rect 37292 50244 37298 50296
rect 37326 50244 37332 50296
rect 37384 50284 37390 50296
rect 37384 50256 38660 50284
rect 37384 50244 37390 50256
rect 29104 50188 29276 50216
rect 29104 50176 29110 50188
rect 22882 50108 22888 50160
rect 22940 50148 22946 50160
rect 27298 50148 27304 50160
rect 22940 50120 27304 50148
rect 22940 50108 22946 50120
rect 27298 50108 27304 50120
rect 27356 50108 27362 50160
rect 38632 50148 38660 50256
rect 38816 50216 38844 50324
rect 40086 50312 40092 50364
rect 40144 50352 40150 50364
rect 44686 50352 44692 50364
rect 40144 50324 44692 50352
rect 40144 50312 40150 50324
rect 44686 50312 44692 50324
rect 44744 50312 44750 50364
rect 108350 50312 108356 50364
rect 108408 50352 108414 50364
rect 110558 50352 110564 50364
rect 108408 50324 110564 50352
rect 108408 50312 108414 50324
rect 110558 50312 110564 50324
rect 110616 50312 110622 50364
rect 39626 50244 39632 50296
rect 39684 50284 39690 50296
rect 39684 50256 40408 50284
rect 39684 50244 39690 50256
rect 39258 50216 39264 50228
rect 38816 50188 39264 50216
rect 39258 50176 39264 50188
rect 39316 50176 39322 50228
rect 39994 50148 40000 50160
rect 38632 50120 40000 50148
rect 39994 50108 40000 50120
rect 40052 50108 40058 50160
rect 27022 50040 27028 50092
rect 27080 50080 27086 50092
rect 29414 50080 29420 50092
rect 27080 50052 29420 50080
rect 27080 50040 27086 50052
rect 29414 50040 29420 50052
rect 29472 50040 29478 50092
rect 30426 50040 30432 50092
rect 30484 50080 30490 50092
rect 31622 50080 31628 50092
rect 30484 50052 31628 50080
rect 30484 50040 30490 50052
rect 31622 50040 31628 50052
rect 31680 50040 31686 50092
rect 40380 50080 40408 50256
rect 40454 50244 40460 50296
rect 40512 50284 40518 50296
rect 40512 50256 41236 50284
rect 40512 50244 40518 50256
rect 41208 50216 41236 50256
rect 41282 50244 41288 50296
rect 41340 50284 41346 50296
rect 41340 50256 42984 50284
rect 41340 50244 41346 50256
rect 42956 50216 42984 50256
rect 107522 50244 107528 50296
rect 107580 50284 107586 50296
rect 107580 50256 108488 50284
rect 107580 50244 107586 50256
rect 46802 50216 46808 50228
rect 41208 50188 42892 50216
rect 42956 50188 46808 50216
rect 42864 50148 42892 50188
rect 46802 50176 46808 50188
rect 46860 50176 46866 50228
rect 93630 50176 93636 50228
rect 93688 50216 93694 50228
rect 94366 50216 94372 50228
rect 93688 50188 94372 50216
rect 93688 50176 93694 50188
rect 94366 50176 94372 50188
rect 94424 50176 94430 50228
rect 97678 50176 97684 50228
rect 97736 50216 97742 50228
rect 98598 50216 98604 50228
rect 97736 50188 98604 50216
rect 97736 50176 97742 50188
rect 98598 50176 98604 50188
rect 98656 50176 98662 50228
rect 108460 50216 108488 50256
rect 108718 50244 108724 50296
rect 108776 50284 108782 50296
rect 111772 50284 111800 50392
rect 176430 50380 176436 50432
rect 176488 50420 176494 50432
rect 177810 50420 177816 50432
rect 176488 50392 177816 50420
rect 176488 50380 176494 50392
rect 177810 50380 177816 50392
rect 177868 50380 177874 50432
rect 178454 50380 178460 50432
rect 178512 50420 178518 50432
rect 180662 50420 180668 50432
rect 178512 50392 180668 50420
rect 178512 50380 178518 50392
rect 180662 50380 180668 50392
rect 180720 50380 180726 50432
rect 182870 50380 182876 50432
rect 182928 50420 182934 50432
rect 184894 50420 184900 50432
rect 182928 50392 184900 50420
rect 182928 50380 182934 50392
rect 184894 50380 184900 50392
rect 184952 50380 184958 50432
rect 185262 50380 185268 50432
rect 185320 50420 185326 50432
rect 187746 50420 187752 50432
rect 185320 50392 187752 50420
rect 185320 50380 185326 50392
rect 187746 50380 187752 50392
rect 187804 50380 187810 50432
rect 176062 50312 176068 50364
rect 176120 50352 176126 50364
rect 177258 50352 177264 50364
rect 176120 50324 177264 50352
rect 176120 50312 176126 50324
rect 177258 50312 177264 50324
rect 177316 50312 177322 50364
rect 177626 50312 177632 50364
rect 177684 50352 177690 50364
rect 179558 50352 179564 50364
rect 177684 50324 179564 50352
rect 177684 50312 177690 50324
rect 179558 50312 179564 50324
rect 179616 50312 179622 50364
rect 180478 50312 180484 50364
rect 180536 50352 180542 50364
rect 180536 50324 182272 50352
rect 180536 50312 180542 50324
rect 108776 50256 110604 50284
rect 111772 50256 111892 50284
rect 108776 50244 108782 50256
rect 109454 50216 109460 50228
rect 108460 50188 109460 50216
rect 109454 50176 109460 50188
rect 109512 50176 109518 50228
rect 110576 50216 110604 50256
rect 111110 50216 111116 50228
rect 110576 50188 111116 50216
rect 111110 50176 111116 50188
rect 111168 50176 111174 50228
rect 111864 50216 111892 50256
rect 111938 50244 111944 50296
rect 111996 50284 112002 50296
rect 111996 50256 112904 50284
rect 111996 50244 112002 50256
rect 112766 50216 112772 50228
rect 111864 50188 112772 50216
rect 112766 50176 112772 50188
rect 112824 50176 112830 50228
rect 112876 50216 112904 50256
rect 113962 50244 113968 50296
rect 114020 50284 114026 50296
rect 114020 50256 116124 50284
rect 114020 50244 114026 50256
rect 115618 50216 115624 50228
rect 112876 50188 115624 50216
rect 115618 50176 115624 50188
rect 115676 50176 115682 50228
rect 116096 50216 116124 50256
rect 176798 50244 176804 50296
rect 176856 50284 176862 50296
rect 176856 50256 178224 50284
rect 176856 50244 176862 50256
rect 118378 50216 118384 50228
rect 116096 50188 118384 50216
rect 118378 50176 118384 50188
rect 118436 50176 118442 50228
rect 165114 50176 165120 50228
rect 165172 50216 165178 50228
rect 167046 50216 167052 50228
rect 165172 50188 167052 50216
rect 165172 50176 165178 50188
rect 167046 50176 167052 50188
rect 167104 50176 167110 50228
rect 169898 50176 169904 50228
rect 169956 50216 169962 50228
rect 170818 50216 170824 50228
rect 169956 50188 170824 50216
rect 169956 50176 169962 50188
rect 170818 50176 170824 50188
rect 170876 50176 170882 50228
rect 171002 50176 171008 50228
rect 171060 50216 171066 50228
rect 171646 50216 171652 50228
rect 171060 50188 171652 50216
rect 171060 50176 171066 50188
rect 171646 50176 171652 50188
rect 171704 50176 171710 50228
rect 178196 50216 178224 50256
rect 179466 50244 179472 50296
rect 179524 50244 179530 50296
rect 181214 50244 181220 50296
rect 181272 50284 181278 50296
rect 181272 50256 182180 50284
rect 181272 50244 181278 50256
rect 178454 50216 178460 50228
rect 178196 50188 178460 50216
rect 178454 50176 178460 50188
rect 178512 50176 178518 50228
rect 179484 50216 179512 50244
rect 181858 50216 181864 50228
rect 179484 50188 181864 50216
rect 181858 50176 181864 50188
rect 181916 50176 181922 50228
rect 45422 50148 45428 50160
rect 42864 50120 45428 50148
rect 45422 50108 45428 50120
rect 45480 50108 45486 50160
rect 93446 50108 93452 50160
rect 93504 50148 93510 50160
rect 95470 50148 95476 50160
rect 93504 50120 95476 50148
rect 93504 50108 93510 50120
rect 95470 50108 95476 50120
rect 95528 50108 95534 50160
rect 97126 50108 97132 50160
rect 97184 50148 97190 50160
rect 98322 50148 98328 50160
rect 97184 50120 98328 50148
rect 97184 50108 97190 50120
rect 98322 50108 98328 50120
rect 98380 50108 98386 50160
rect 98782 50108 98788 50160
rect 98840 50148 98846 50160
rect 99702 50148 99708 50160
rect 98840 50120 99708 50148
rect 98840 50108 98846 50120
rect 99702 50108 99708 50120
rect 99760 50108 99766 50160
rect 107890 50108 107896 50160
rect 107948 50148 107954 50160
rect 110006 50148 110012 50160
rect 107948 50120 110012 50148
rect 107948 50108 107954 50120
rect 110006 50108 110012 50120
rect 110064 50108 110070 50160
rect 110650 50108 110656 50160
rect 110708 50148 110714 50160
rect 113962 50148 113968 50160
rect 110708 50120 113968 50148
rect 110708 50108 110714 50120
rect 113962 50108 113968 50120
rect 114020 50108 114026 50160
rect 163826 50108 163832 50160
rect 163884 50148 163890 50160
rect 167598 50148 167604 50160
rect 163884 50120 167604 50148
rect 163884 50108 163890 50120
rect 167598 50108 167604 50120
rect 167656 50108 167662 50160
rect 168702 50108 168708 50160
rect 168760 50148 168766 50160
rect 170082 50148 170088 50160
rect 168760 50120 170088 50148
rect 168760 50108 168766 50120
rect 170082 50108 170088 50120
rect 170140 50108 170146 50160
rect 178270 50108 178276 50160
rect 178328 50148 178334 50160
rect 180110 50148 180116 50160
rect 178328 50120 180116 50148
rect 178328 50108 178334 50120
rect 180110 50108 180116 50120
rect 180168 50108 180174 50160
rect 182152 50148 182180 50256
rect 182244 50216 182272 50324
rect 184802 50312 184808 50364
rect 184860 50352 184866 50364
rect 189862 50352 189868 50364
rect 184860 50324 189868 50352
rect 184860 50312 184866 50324
rect 189862 50312 189868 50324
rect 189920 50312 189926 50364
rect 183238 50244 183244 50296
rect 183296 50284 183302 50296
rect 183296 50256 185124 50284
rect 183296 50244 183302 50256
rect 183514 50216 183520 50228
rect 182244 50188 183520 50216
rect 183514 50176 183520 50188
rect 183572 50176 183578 50228
rect 185096 50216 185124 50256
rect 185630 50244 185636 50296
rect 185688 50284 185694 50296
rect 185688 50256 187884 50284
rect 185688 50244 185694 50256
rect 187562 50216 187568 50228
rect 185096 50188 187568 50216
rect 187562 50176 187568 50188
rect 187620 50176 187626 50228
rect 184710 50148 184716 50160
rect 182152 50120 184716 50148
rect 184710 50108 184716 50120
rect 184768 50108 184774 50160
rect 184986 50108 184992 50160
rect 185044 50148 185050 50160
rect 186366 50148 186372 50160
rect 185044 50120 186372 50148
rect 185044 50108 185050 50120
rect 186366 50108 186372 50120
rect 186424 50108 186430 50160
rect 43766 50080 43772 50092
rect 40380 50052 43772 50080
rect 43766 50040 43772 50052
rect 43824 50040 43830 50092
rect 93354 50040 93360 50092
rect 93412 50080 93418 50092
rect 96022 50080 96028 50092
rect 93412 50052 96028 50080
rect 93412 50040 93418 50052
rect 96022 50040 96028 50052
rect 96080 50040 96086 50092
rect 109270 50040 109276 50092
rect 109328 50080 109334 50092
rect 111662 50080 111668 50092
rect 109328 50052 111668 50080
rect 109328 50040 109334 50052
rect 111662 50040 111668 50052
rect 111720 50040 111726 50092
rect 169254 50040 169260 50092
rect 169312 50080 169318 50092
rect 170450 50080 170456 50092
rect 169312 50052 170456 50080
rect 169312 50040 169318 50052
rect 170450 50040 170456 50052
rect 170508 50040 170514 50092
rect 184894 50040 184900 50092
rect 184952 50080 184958 50092
rect 187010 50080 187016 50092
rect 184952 50052 187016 50080
rect 184952 50040 184958 50052
rect 187010 50040 187016 50052
rect 187068 50040 187074 50092
rect 24262 49972 24268 50024
rect 24320 50012 24326 50024
rect 28034 50012 28040 50024
rect 24320 49984 28040 50012
rect 24320 49972 24326 49984
rect 28034 49972 28040 49984
rect 28092 49972 28098 50024
rect 28310 49972 28316 50024
rect 28368 50012 28374 50024
rect 30150 50012 30156 50024
rect 28368 49984 30156 50012
rect 28368 49972 28374 49984
rect 30150 49972 30156 49984
rect 30208 49972 30214 50024
rect 31070 49972 31076 50024
rect 31128 50012 31134 50024
rect 32082 50012 32088 50024
rect 31128 49984 32088 50012
rect 31128 49972 31134 49984
rect 32082 49972 32088 49984
rect 32140 49972 32146 50024
rect 40822 49972 40828 50024
rect 40880 50012 40886 50024
rect 42662 50012 42668 50024
rect 40880 49984 42668 50012
rect 40880 49972 40886 49984
rect 42662 49972 42668 49984
rect 42720 49972 42726 50024
rect 42938 49972 42944 50024
rect 42996 50012 43002 50024
rect 46066 50012 46072 50024
rect 42996 49984 46072 50012
rect 42996 49972 43002 49984
rect 46066 49972 46072 49984
rect 46124 49972 46130 50024
rect 112674 49972 112680 50024
rect 112732 50012 112738 50024
rect 114514 50012 114520 50024
rect 112732 49984 114520 50012
rect 112732 49972 112738 49984
rect 114514 49972 114520 49984
rect 114572 49972 114578 50024
rect 181122 49972 181128 50024
rect 181180 50012 181186 50024
rect 184158 50012 184164 50024
rect 181180 49984 184164 50012
rect 181180 49972 181186 49984
rect 184158 49972 184164 49984
rect 184216 49972 184222 50024
rect 187856 50012 187884 50256
rect 190966 50012 190972 50024
rect 187856 49984 190972 50012
rect 190966 49972 190972 49984
rect 191024 49972 191030 50024
rect 23618 49904 23624 49956
rect 23676 49944 23682 49956
rect 27666 49944 27672 49956
rect 23676 49916 27672 49944
rect 23676 49904 23682 49916
rect 27666 49904 27672 49916
rect 27724 49904 27730 49956
rect 29690 49904 29696 49956
rect 29748 49944 29754 49956
rect 31254 49944 31260 49956
rect 29748 49916 31260 49944
rect 29748 49904 29754 49916
rect 31254 49904 31260 49916
rect 31312 49904 31318 49956
rect 41374 49904 41380 49956
rect 41432 49944 41438 49956
rect 43398 49944 43404 49956
rect 41432 49916 43404 49944
rect 41432 49904 41438 49916
rect 43398 49904 43404 49916
rect 43456 49904 43462 49956
rect 183422 49904 183428 49956
rect 183480 49944 183486 49956
rect 185262 49944 185268 49956
rect 183480 49916 185268 49944
rect 183480 49904 183486 49916
rect 185262 49904 185268 49916
rect 185320 49904 185326 49956
rect 187746 49904 187752 49956
rect 187804 49944 187810 49956
rect 190414 49944 190420 49956
rect 187804 49916 190420 49944
rect 187804 49904 187810 49916
rect 190414 49904 190420 49916
rect 190472 49904 190478 49956
rect 38890 49836 38896 49888
rect 38948 49876 38954 49888
rect 42018 49876 42024 49888
rect 38948 49848 42024 49876
rect 38948 49836 38954 49848
rect 42018 49836 42024 49848
rect 42076 49836 42082 49888
rect 182502 49836 182508 49888
rect 182560 49876 182566 49888
rect 185814 49876 185820 49888
rect 182560 49848 185820 49876
rect 182560 49836 182566 49848
rect 185814 49836 185820 49848
rect 185872 49836 185878 49888
rect 44042 49768 44048 49820
rect 44100 49808 44106 49820
rect 47446 49808 47452 49820
rect 44100 49780 47452 49808
rect 44100 49768 44106 49780
rect 47446 49768 47452 49780
rect 47504 49768 47510 49820
rect 112398 49768 112404 49820
rect 112456 49808 112462 49820
rect 115066 49808 115072 49820
rect 112456 49780 115072 49808
rect 112456 49768 112462 49780
rect 115066 49768 115072 49780
rect 115124 49768 115130 49820
rect 186458 49768 186464 49820
rect 186516 49808 186522 49820
rect 189218 49808 189224 49820
rect 186516 49780 189224 49808
rect 186516 49768 186522 49780
rect 189218 49768 189224 49780
rect 189276 49768 189282 49820
rect 26286 49700 26292 49752
rect 26344 49740 26350 49752
rect 29230 49740 29236 49752
rect 26344 49712 29236 49740
rect 26344 49700 26350 49712
rect 29230 49700 29236 49712
rect 29288 49700 29294 49752
rect 163734 49700 163740 49752
rect 163792 49740 163798 49752
rect 168150 49740 168156 49752
rect 163792 49712 168156 49740
rect 163792 49700 163798 49712
rect 168150 49700 168156 49712
rect 168208 49700 168214 49752
rect 24906 49632 24912 49684
rect 24964 49672 24970 49684
rect 28494 49672 28500 49684
rect 24964 49644 28500 49672
rect 24964 49632 24970 49644
rect 28494 49632 28500 49644
rect 28552 49632 28558 49684
rect 39718 49632 39724 49684
rect 39776 49672 39782 49684
rect 41282 49672 41288 49684
rect 39776 49644 41288 49672
rect 39776 49632 39782 49644
rect 41282 49632 41288 49644
rect 41340 49632 41346 49684
rect 186274 49632 186280 49684
rect 186332 49672 186338 49684
rect 188666 49672 188672 49684
rect 186332 49644 188672 49672
rect 186332 49632 186338 49644
rect 188666 49632 188672 49644
rect 188724 49632 188730 49684
rect 113502 49564 113508 49616
rect 113560 49604 113566 49616
rect 117826 49604 117832 49616
rect 113560 49576 117832 49604
rect 113560 49564 113566 49576
rect 117826 49564 117832 49576
rect 117884 49564 117890 49616
rect 20214 49496 20220 49548
rect 20272 49536 20278 49548
rect 44410 49536 44416 49548
rect 20272 49508 44416 49536
rect 20272 49496 20278 49508
rect 44410 49496 44416 49508
rect 44468 49496 44474 49548
rect 114698 49496 114704 49548
rect 114756 49536 114762 49548
rect 116722 49536 116728 49548
rect 114756 49508 116728 49536
rect 114756 49496 114762 49508
rect 116722 49496 116728 49508
rect 116780 49496 116786 49548
rect 168518 49496 168524 49548
rect 168576 49536 168582 49548
rect 191518 49536 191524 49548
rect 168576 49508 191524 49536
rect 168576 49496 168582 49508
rect 191518 49496 191524 49508
rect 191576 49496 191582 49548
rect 111754 49360 111760 49412
rect 111812 49400 111818 49412
rect 113410 49400 113416 49412
rect 111812 49372 113416 49400
rect 111812 49360 111818 49372
rect 113410 49360 113416 49372
rect 113468 49360 113474 49412
rect 91422 49224 91428 49276
rect 91480 49264 91486 49276
rect 92894 49264 92900 49276
rect 91480 49236 92900 49264
rect 91480 49224 91486 49236
rect 92894 49224 92900 49236
rect 92952 49224 92958 49276
rect 96574 49088 96580 49140
rect 96632 49128 96638 49140
rect 97770 49128 97776 49140
rect 96632 49100 97776 49128
rect 96632 49088 96638 49100
rect 97770 49088 97776 49100
rect 97828 49088 97834 49140
rect 114606 49088 114612 49140
rect 114664 49128 114670 49140
rect 117274 49128 117280 49140
rect 114664 49100 117280 49128
rect 114664 49088 114670 49100
rect 117274 49088 117280 49100
rect 117332 49088 117338 49140
rect 21502 48952 21508 49004
rect 21560 48992 21566 49004
rect 26194 48992 26200 49004
rect 21560 48964 26200 48992
rect 21560 48952 21566 48964
rect 26194 48952 26200 48964
rect 26252 48952 26258 49004
rect 114422 48952 114428 49004
rect 114480 48992 114486 49004
rect 116170 48992 116176 49004
rect 114480 48964 116176 48992
rect 114480 48952 114486 48964
rect 116170 48952 116176 48964
rect 116228 48952 116234 49004
rect 182042 48952 182048 49004
rect 182100 48992 182106 49004
rect 182962 48992 182968 49004
rect 182100 48964 182968 48992
rect 182100 48952 182106 48964
rect 182962 48952 182968 48964
rect 183020 48952 183026 49004
rect 22238 48884 22244 48936
rect 22296 48924 22302 48936
rect 26378 48924 26384 48936
rect 22296 48896 26384 48924
rect 22296 48884 22302 48896
rect 26378 48884 26384 48896
rect 26436 48884 26442 48936
rect 103934 47728 103940 47780
rect 103992 47768 103998 47780
rect 104394 47768 104400 47780
rect 103992 47740 104400 47768
rect 103992 47728 103998 47740
rect 104394 47728 104400 47740
rect 104452 47728 104458 47780
rect 50758 46504 50764 46556
rect 50816 46544 50822 46556
rect 61614 46544 61620 46556
rect 50816 46516 61620 46544
rect 50816 46504 50822 46516
rect 61614 46504 61620 46516
rect 61672 46504 61678 46556
rect 122794 46504 122800 46556
rect 122852 46544 122858 46556
rect 129142 46544 129148 46556
rect 122852 46516 129148 46544
rect 122852 46504 122858 46516
rect 129142 46504 129148 46516
rect 129200 46504 129206 46556
rect 51034 46436 51040 46488
rect 51092 46476 51098 46488
rect 63086 46476 63092 46488
rect 51092 46448 63092 46476
rect 51092 46436 51098 46448
rect 63086 46436 63092 46448
rect 63144 46436 63150 46488
rect 122334 46436 122340 46488
rect 122392 46476 122398 46488
rect 127670 46476 127676 46488
rect 122392 46448 127676 46476
rect 122392 46436 122398 46448
rect 127670 46436 127676 46448
rect 127728 46436 127734 46488
rect 51126 46368 51132 46420
rect 51184 46408 51190 46420
rect 60050 46408 60056 46420
rect 51184 46380 60056 46408
rect 51184 46368 51190 46380
rect 60050 46368 60056 46380
rect 60108 46368 60114 46420
rect 122426 46368 122432 46420
rect 122484 46408 122490 46420
rect 130614 46408 130620 46420
rect 122484 46380 130620 46408
rect 122484 46368 122490 46380
rect 130614 46368 130620 46380
rect 130672 46368 130678 46420
rect 148646 46368 148652 46420
rect 148704 46408 148710 46420
rect 158214 46408 158220 46420
rect 148704 46380 158220 46408
rect 148704 46368 148710 46380
rect 158214 46368 158220 46380
rect 158272 46368 158278 46420
rect 50942 46300 50948 46352
rect 51000 46340 51006 46352
rect 58578 46340 58584 46352
rect 51000 46312 58584 46340
rect 51000 46300 51006 46312
rect 58578 46300 58584 46312
rect 58636 46300 58642 46352
rect 76610 46300 76616 46352
rect 76668 46340 76674 46352
rect 87834 46340 87840 46352
rect 76668 46312 87840 46340
rect 76668 46300 76674 46312
rect 87834 46300 87840 46312
rect 87892 46300 87898 46352
rect 122518 46300 122524 46352
rect 122576 46340 122582 46352
rect 132086 46340 132092 46352
rect 122576 46312 132092 46340
rect 122576 46300 122582 46312
rect 132086 46300 132092 46312
rect 132144 46300 132150 46352
rect 150118 46300 150124 46352
rect 150176 46340 150182 46352
rect 159594 46340 159600 46352
rect 150176 46312 159600 46340
rect 150176 46300 150182 46312
rect 159594 46300 159600 46312
rect 159652 46300 159658 46352
rect 50666 46232 50672 46284
rect 50724 46272 50730 46284
rect 55634 46272 55640 46284
rect 50724 46244 55640 46272
rect 50724 46232 50730 46244
rect 55634 46232 55640 46244
rect 55692 46232 55698 46284
rect 81118 46232 81124 46284
rect 81176 46272 81182 46284
rect 87926 46272 87932 46284
rect 81176 46244 87932 46272
rect 81176 46232 81182 46244
rect 87926 46232 87932 46244
rect 87984 46232 87990 46284
rect 126474 46232 126480 46284
rect 126532 46272 126538 46284
rect 136594 46272 136600 46284
rect 126532 46244 136600 46272
rect 126532 46232 126538 46244
rect 136594 46232 136600 46244
rect 136652 46232 136658 46284
rect 151590 46232 151596 46284
rect 151648 46272 151654 46284
rect 159686 46272 159692 46284
rect 151648 46244 159692 46272
rect 151648 46232 151654 46244
rect 159686 46232 159692 46244
rect 159744 46232 159750 46284
rect 50850 46164 50856 46216
rect 50908 46204 50914 46216
rect 57106 46204 57112 46216
rect 50908 46176 57112 46204
rect 50908 46164 50914 46176
rect 57106 46164 57112 46176
rect 57164 46164 57170 46216
rect 78082 46164 78088 46216
rect 78140 46204 78146 46216
rect 86454 46204 86460 46216
rect 78140 46176 86460 46204
rect 78140 46164 78146 46176
rect 86454 46164 86460 46176
rect 86512 46164 86518 46216
rect 122702 46164 122708 46216
rect 122760 46204 122766 46216
rect 133650 46204 133656 46216
rect 122760 46176 133656 46204
rect 122760 46164 122766 46176
rect 133650 46164 133656 46176
rect 133708 46164 133714 46216
rect 54070 46096 54076 46148
rect 54128 46136 54134 46148
rect 67594 46136 67600 46148
rect 54128 46108 67600 46136
rect 54128 46096 54134 46108
rect 67594 46096 67600 46108
rect 67652 46096 67658 46148
rect 79554 46096 79560 46148
rect 79612 46136 79618 46148
rect 85074 46136 85080 46148
rect 79612 46108 85080 46136
rect 79612 46096 79618 46108
rect 85074 46096 85080 46108
rect 85132 46096 85138 46148
rect 122886 46096 122892 46148
rect 122944 46136 122950 46148
rect 135122 46136 135128 46148
rect 122944 46108 135128 46136
rect 122944 46096 122950 46108
rect 135122 46096 135128 46108
rect 135180 46096 135186 46148
rect 153154 46096 153160 46148
rect 153212 46136 153218 46148
rect 158306 46136 158312 46148
rect 153212 46108 158312 46136
rect 153212 46096 153218 46108
rect 158306 46096 158312 46108
rect 158364 46096 158370 46148
rect 121690 44872 121696 44924
rect 121748 44912 121754 44924
rect 123530 44912 123536 44924
rect 121748 44884 123536 44912
rect 121748 44872 121754 44884
rect 123530 44872 123536 44884
rect 123588 44872 123594 44924
rect 121690 44736 121696 44788
rect 121748 44776 121754 44788
rect 123346 44776 123352 44788
rect 121748 44748 123352 44776
rect 121748 44736 121754 44748
rect 123346 44736 123352 44748
rect 123404 44736 123410 44788
rect 154718 44736 154724 44788
rect 154776 44776 154782 44788
rect 156834 44776 156840 44788
rect 154776 44748 156840 44776
rect 154776 44736 154782 44748
rect 156834 44736 156840 44748
rect 156892 44736 156898 44788
rect 84338 44396 84344 44448
rect 84396 44436 84402 44448
rect 85166 44436 85172 44448
rect 84396 44408 85172 44436
rect 84396 44396 84402 44408
rect 85166 44396 85172 44408
rect 85224 44396 85230 44448
rect 159778 43648 159784 43700
rect 159836 43688 159842 43700
rect 160054 43688 160060 43700
rect 159836 43660 160060 43688
rect 159836 43648 159842 43660
rect 160054 43648 160060 43660
rect 160112 43648 160118 43700
rect 121690 43376 121696 43428
rect 121748 43416 121754 43428
rect 124358 43416 124364 43428
rect 121748 43388 124364 43416
rect 121748 43376 121754 43388
rect 124358 43376 124364 43388
rect 124416 43376 124422 43428
rect 121690 42016 121696 42068
rect 121748 42056 121754 42068
rect 124266 42056 124272 42068
rect 121748 42028 124272 42056
rect 121748 42016 121754 42028
rect 124266 42016 124272 42028
rect 124324 42016 124330 42068
rect 121690 40656 121696 40708
rect 121748 40696 121754 40708
rect 124358 40696 124364 40708
rect 121748 40668 124364 40696
rect 121748 40656 121754 40668
rect 124358 40656 124364 40668
rect 124416 40656 124422 40708
rect 14694 40520 14700 40572
rect 14752 40560 14758 40572
rect 18006 40560 18012 40572
rect 14752 40532 18012 40560
rect 14752 40520 14758 40532
rect 18006 40520 18012 40532
rect 18064 40520 18070 40572
rect 156466 39704 156472 39756
rect 156524 39744 156530 39756
rect 156926 39744 156932 39756
rect 156524 39716 156932 39744
rect 156524 39704 156530 39716
rect 156926 39704 156932 39716
rect 156984 39704 156990 39756
rect 122518 39160 122524 39212
rect 122576 39200 122582 39212
rect 122794 39200 122800 39212
rect 122576 39172 122800 39200
rect 122576 39160 122582 39172
rect 122794 39160 122800 39172
rect 122852 39160 122858 39212
rect 159042 38548 159048 38600
rect 159100 38588 159106 38600
rect 160514 38588 160520 38600
rect 159100 38560 160520 38588
rect 159100 38548 159106 38560
rect 160514 38548 160520 38560
rect 160572 38548 160578 38600
rect 121782 38412 121788 38464
rect 121840 38452 121846 38464
rect 123898 38452 123904 38464
rect 121840 38424 123904 38452
rect 121840 38412 121846 38424
rect 123898 38412 123904 38424
rect 123956 38412 123962 38464
rect 121690 38208 121696 38260
rect 121748 38248 121754 38260
rect 123438 38248 123444 38260
rect 121748 38220 123444 38248
rect 121748 38208 121754 38220
rect 123438 38208 123444 38220
rect 123496 38208 123502 38260
rect 121690 37800 121696 37852
rect 121748 37840 121754 37852
rect 124358 37840 124364 37852
rect 121748 37812 124364 37840
rect 121748 37800 121754 37812
rect 124358 37800 124364 37812
rect 124416 37800 124422 37852
rect 88202 37324 88208 37376
rect 88260 37364 88266 37376
rect 88754 37364 88760 37376
rect 88260 37336 88760 37364
rect 88260 37324 88266 37336
rect 88754 37324 88760 37336
rect 88812 37324 88818 37376
rect 121690 35080 121696 35132
rect 121748 35120 121754 35132
rect 123622 35120 123628 35132
rect 121748 35092 123628 35120
rect 121748 35080 121754 35092
rect 123622 35080 123628 35092
rect 123680 35080 123686 35132
rect 121690 33992 121696 34044
rect 121748 34032 121754 34044
rect 124358 34032 124364 34044
rect 121748 34004 124364 34032
rect 121748 33992 121754 34004
rect 124358 33992 124364 34004
rect 124416 33992 124422 34044
rect 121690 33720 121696 33772
rect 121748 33760 121754 33772
rect 124266 33760 124272 33772
rect 121748 33732 124272 33760
rect 121748 33720 121754 33732
rect 124266 33720 124272 33732
rect 124324 33720 124330 33772
rect 121690 32360 121696 32412
rect 121748 32400 121754 32412
rect 123990 32400 123996 32412
rect 121748 32372 123996 32400
rect 121748 32360 121754 32372
rect 123990 32360 123996 32372
rect 124048 32360 124054 32412
rect 121690 31000 121696 31052
rect 121748 31040 121754 31052
rect 124358 31040 124364 31052
rect 121748 31012 124364 31040
rect 121748 31000 121754 31012
rect 124358 31000 124364 31012
rect 124416 31000 124422 31052
rect 121690 28824 121696 28876
rect 121748 28864 121754 28876
rect 123530 28864 123536 28876
rect 121748 28836 123536 28864
rect 121748 28824 121754 28836
rect 123530 28824 123536 28836
rect 123588 28824 123594 28876
rect 121690 28484 121696 28536
rect 121748 28524 121754 28536
rect 124358 28524 124364 28536
rect 121748 28496 124364 28524
rect 121748 28484 121754 28496
rect 124358 28484 124364 28496
rect 124416 28484 124422 28536
rect 121690 28144 121696 28196
rect 121748 28184 121754 28196
rect 124082 28184 124088 28196
rect 121748 28156 124088 28184
rect 121748 28144 121754 28156
rect 124082 28144 124088 28156
rect 124140 28144 124146 28196
rect 159042 28144 159048 28196
rect 159100 28184 159106 28196
rect 160698 28184 160704 28196
rect 159100 28156 160704 28184
rect 159100 28144 159106 28156
rect 160698 28144 160704 28156
rect 160756 28144 160762 28196
rect 88294 27668 88300 27720
rect 88352 27708 88358 27720
rect 88754 27708 88760 27720
rect 88352 27680 88760 27708
rect 88352 27668 88358 27680
rect 88754 27668 88760 27680
rect 88812 27668 88818 27720
rect 158950 25152 158956 25204
rect 159008 25192 159014 25204
rect 160330 25192 160336 25204
rect 159008 25164 160336 25192
rect 159008 25152 159014 25164
rect 160330 25152 160336 25164
rect 160388 25152 160394 25204
rect 50574 24472 50580 24524
rect 50632 24512 50638 24524
rect 50850 24512 50856 24524
rect 50632 24484 50856 24512
rect 50632 24472 50638 24484
rect 50850 24472 50856 24484
rect 50908 24472 50914 24524
rect 121690 24200 121696 24252
rect 121748 24240 121754 24252
rect 123438 24240 123444 24252
rect 121748 24212 123444 24240
rect 121748 24200 121754 24212
rect 123438 24200 123444 24212
rect 123496 24200 123502 24252
rect 51034 24064 51040 24116
rect 51092 24104 51098 24116
rect 51310 24104 51316 24116
rect 51092 24076 51316 24104
rect 51092 24064 51098 24076
rect 51310 24064 51316 24076
rect 51368 24064 51374 24116
rect 159042 22636 159048 22688
rect 159100 22676 159106 22688
rect 160698 22676 160704 22688
rect 159100 22648 160704 22676
rect 159100 22636 159106 22648
rect 160698 22636 160704 22648
rect 160756 22636 160762 22688
rect 85166 22568 85172 22620
rect 85224 22608 85230 22620
rect 88754 22608 88760 22620
rect 85224 22580 88760 22608
rect 85224 22568 85230 22580
rect 88754 22568 88760 22580
rect 88812 22568 88818 22620
rect 156926 22568 156932 22620
rect 156984 22608 156990 22620
rect 160422 22608 160428 22620
rect 156984 22580 160428 22608
rect 156984 22568 156990 22580
rect 160422 22568 160428 22580
rect 160480 22568 160486 22620
rect 156834 22500 156840 22552
rect 156892 22540 156898 22552
rect 160514 22540 160520 22552
rect 156892 22512 160520 22540
rect 156892 22500 156898 22512
rect 160514 22500 160520 22512
rect 160572 22500 160578 22552
rect 85074 21208 85080 21260
rect 85132 21248 85138 21260
rect 88570 21248 88576 21260
rect 85132 21220 88576 21248
rect 85132 21208 85138 21220
rect 88570 21208 88576 21220
rect 88628 21208 88634 21260
rect 158306 21208 158312 21260
rect 158364 21248 158370 21260
rect 160330 21248 160336 21260
rect 158364 21220 160336 21248
rect 158364 21208 158370 21220
rect 160330 21208 160336 21220
rect 160388 21208 160394 21260
rect 86454 19780 86460 19832
rect 86512 19820 86518 19832
rect 88570 19820 88576 19832
rect 86512 19792 88576 19820
rect 86512 19780 86518 19792
rect 88570 19780 88576 19792
rect 88628 19780 88634 19832
rect 158214 19780 158220 19832
rect 158272 19820 158278 19832
rect 160330 19820 160336 19832
rect 158272 19792 160336 19820
rect 158272 19780 158278 19792
rect 160330 19780 160336 19792
rect 160388 19780 160394 19832
rect 13130 19100 13136 19152
rect 13188 19140 13194 19152
rect 66490 19140 66496 19152
rect 13188 19112 66496 19140
rect 13188 19100 13194 19112
rect 66490 19100 66496 19112
rect 66548 19100 66554 19152
rect 18098 18420 18104 18472
rect 18156 18460 18162 18472
rect 62534 18460 62540 18472
rect 18156 18432 62540 18460
rect 18156 18420 18162 18432
rect 62534 18420 62540 18432
rect 62592 18420 62598 18472
rect 69986 18420 69992 18472
rect 70044 18460 70050 18472
rect 73942 18460 73948 18472
rect 70044 18432 73948 18460
rect 70044 18420 70050 18432
rect 73942 18420 73948 18432
rect 74000 18420 74006 18472
rect 74037 18463 74095 18469
rect 74037 18429 74049 18463
rect 74083 18460 74095 18463
rect 119666 18460 119672 18472
rect 74083 18432 119672 18460
rect 74083 18429 74095 18432
rect 74037 18423 74095 18429
rect 119666 18420 119672 18432
rect 119724 18420 119730 18472
rect 50390 18352 50396 18404
rect 50448 18392 50454 18404
rect 63546 18392 63552 18404
rect 50448 18364 63552 18392
rect 50448 18352 50454 18364
rect 63546 18352 63552 18364
rect 63604 18392 63610 18404
rect 94642 18392 94648 18404
rect 63604 18364 94648 18392
rect 63604 18352 63610 18364
rect 94642 18352 94648 18364
rect 94700 18392 94706 18404
rect 95378 18392 95384 18404
rect 94700 18364 95384 18392
rect 94700 18352 94706 18364
rect 95378 18352 95384 18364
rect 95436 18352 95442 18404
rect 100162 18352 100168 18404
rect 100220 18392 100226 18404
rect 134570 18392 134576 18404
rect 100220 18364 134576 18392
rect 100220 18352 100226 18364
rect 134570 18352 134576 18364
rect 134628 18352 134634 18404
rect 55082 18284 55088 18336
rect 55140 18324 55146 18336
rect 75966 18324 75972 18336
rect 55140 18296 75972 18324
rect 55140 18284 55146 18296
rect 75966 18284 75972 18296
rect 76024 18284 76030 18336
rect 81762 18284 81768 18336
rect 81820 18324 81826 18336
rect 83234 18324 83240 18336
rect 81820 18296 83240 18324
rect 81820 18284 81826 18296
rect 83234 18284 83240 18296
rect 83292 18284 83298 18336
rect 143770 18284 143776 18336
rect 143828 18324 143834 18336
rect 144966 18324 144972 18336
rect 143828 18296 144972 18324
rect 143828 18284 143834 18296
rect 144966 18284 144972 18296
rect 145024 18284 145030 18336
rect 145150 18284 145156 18336
rect 145208 18324 145214 18336
rect 145978 18324 145984 18336
rect 145208 18296 145984 18324
rect 145208 18284 145214 18296
rect 145978 18284 145984 18296
rect 146036 18284 146042 18336
rect 39074 18216 39080 18268
rect 39132 18256 39138 18268
rect 66674 18256 66680 18268
rect 39132 18228 66680 18256
rect 39132 18216 39138 18228
rect 66674 18216 66680 18228
rect 66732 18216 66738 18268
rect 71090 18216 71096 18268
rect 71148 18256 71154 18268
rect 72930 18256 72936 18268
rect 71148 18228 72936 18256
rect 71148 18216 71154 18228
rect 72930 18216 72936 18228
rect 72988 18216 72994 18268
rect 82222 18216 82228 18268
rect 82280 18256 82286 18268
rect 84338 18256 84344 18268
rect 82280 18228 84344 18256
rect 82280 18216 82286 18228
rect 84338 18216 84344 18228
rect 84396 18216 84402 18268
rect 49746 18148 49752 18200
rect 49804 18188 49810 18200
rect 77070 18188 77076 18200
rect 49804 18160 77076 18188
rect 49804 18148 49810 18160
rect 77070 18148 77076 18160
rect 77128 18148 77134 18200
rect 80290 18148 80296 18200
rect 80348 18188 80354 18200
rect 84246 18188 84252 18200
rect 80348 18160 84252 18188
rect 80348 18148 80354 18160
rect 84246 18148 84252 18160
rect 84304 18148 84310 18200
rect 44410 18080 44416 18132
rect 44468 18120 44474 18132
rect 78082 18120 78088 18132
rect 44468 18092 78088 18120
rect 44468 18080 44474 18092
rect 78082 18080 78088 18092
rect 78140 18080 78146 18132
rect 33738 18012 33744 18064
rect 33796 18052 33802 18064
rect 33796 18024 65616 18052
rect 33796 18012 33802 18024
rect 28402 17944 28408 17996
rect 28460 17984 28466 17996
rect 65588 17984 65616 18024
rect 65662 18012 65668 18064
rect 65720 18052 65726 18064
rect 74037 18055 74095 18061
rect 74037 18052 74049 18055
rect 65720 18024 74049 18052
rect 65720 18012 65726 18024
rect 74037 18021 74049 18024
rect 74083 18021 74095 18055
rect 74037 18015 74095 18021
rect 145794 18012 145800 18064
rect 145852 18052 145858 18064
rect 149106 18052 149112 18064
rect 145852 18024 149112 18052
rect 145852 18012 145858 18024
rect 149106 18012 149112 18024
rect 149164 18012 149170 18064
rect 67686 17984 67692 17996
rect 28460 17956 65524 17984
rect 65588 17956 67692 17984
rect 28460 17944 28466 17956
rect 17730 17876 17736 17928
rect 17788 17916 17794 17928
rect 65496 17916 65524 17956
rect 67686 17944 67692 17956
rect 67744 17944 67750 17996
rect 124450 17944 124456 17996
rect 124508 17984 124514 17996
rect 140826 17984 140832 17996
rect 124508 17956 140832 17984
rect 124508 17944 124514 17956
rect 140826 17944 140832 17956
rect 140884 17944 140890 17996
rect 68790 17916 68796 17928
rect 17788 17888 65432 17916
rect 65496 17888 68796 17916
rect 17788 17876 17794 17888
rect 23066 17808 23072 17860
rect 23124 17848 23130 17860
rect 65404 17848 65432 17888
rect 68790 17876 68796 17888
rect 68848 17876 68854 17928
rect 119114 17876 119120 17928
rect 119172 17916 119178 17928
rect 141838 17916 141844 17928
rect 119172 17888 141844 17916
rect 119172 17876 119178 17888
rect 141838 17876 141844 17888
rect 141896 17876 141902 17928
rect 70814 17848 70820 17860
rect 23124 17820 65340 17848
rect 65404 17820 70820 17848
rect 23124 17808 23130 17820
rect 12486 17740 12492 17792
rect 12544 17780 12550 17792
rect 65205 17783 65263 17789
rect 65205 17780 65217 17783
rect 12544 17752 65217 17780
rect 12544 17740 12550 17752
rect 65205 17749 65217 17752
rect 65251 17749 65263 17783
rect 65312 17780 65340 17820
rect 70814 17808 70820 17820
rect 70872 17808 70878 17860
rect 113778 17808 113784 17860
rect 113836 17848 113842 17860
rect 142850 17848 142856 17860
rect 113836 17820 142856 17848
rect 113836 17808 113842 17820
rect 142850 17808 142856 17820
rect 142908 17808 142914 17860
rect 69802 17780 69808 17792
rect 65312 17752 69808 17780
rect 65205 17743 65263 17749
rect 69802 17740 69808 17752
rect 69860 17740 69866 17792
rect 81210 17740 81216 17792
rect 81268 17780 81274 17792
rect 92434 17780 92440 17792
rect 81268 17752 92440 17780
rect 81268 17740 81274 17752
rect 92434 17740 92440 17752
rect 92492 17740 92498 17792
rect 108442 17740 108448 17792
rect 108500 17780 108506 17792
rect 143862 17780 143868 17792
rect 108500 17752 143868 17780
rect 108500 17740 108506 17752
rect 143862 17740 143868 17752
rect 143920 17740 143926 17792
rect 146990 17740 146996 17792
rect 147048 17780 147054 17792
rect 154810 17780 154816 17792
rect 147048 17752 154816 17780
rect 147048 17740 147054 17752
rect 154810 17740 154816 17752
rect 154868 17740 154874 17792
rect 60418 17672 60424 17724
rect 60476 17712 60482 17724
rect 74954 17712 74960 17724
rect 60476 17684 74960 17712
rect 60476 17672 60482 17684
rect 74954 17672 74960 17684
rect 75012 17672 75018 17724
rect 65205 17647 65263 17653
rect 65205 17613 65217 17647
rect 65251 17644 65263 17647
rect 71826 17644 71832 17656
rect 65251 17616 71832 17644
rect 65251 17613 65263 17616
rect 65205 17607 65263 17613
rect 71826 17604 71832 17616
rect 71884 17604 71890 17656
rect 79186 17468 79192 17520
rect 79244 17508 79250 17520
rect 80106 17508 80112 17520
rect 79244 17480 80112 17508
rect 79244 17468 79250 17480
rect 80106 17468 80112 17480
rect 80164 17468 80170 17520
rect 148002 17128 148008 17180
rect 148060 17168 148066 17180
rect 150578 17168 150584 17180
rect 148060 17140 150584 17168
rect 148060 17128 148066 17140
rect 150578 17128 150584 17140
rect 150636 17128 150642 17180
rect 61522 17060 61528 17112
rect 61580 17100 61586 17112
rect 105774 17100 105780 17112
rect 61580 17072 105780 17100
rect 61580 17060 61586 17072
rect 105774 17060 105780 17072
rect 105832 17060 105838 17112
rect 116998 17060 117004 17112
rect 117056 17100 117062 17112
rect 126474 17100 126480 17112
rect 117056 17072 126480 17100
rect 117056 17060 117062 17072
rect 126474 17060 126480 17072
rect 126532 17060 126538 17112
rect 133558 17060 133564 17112
rect 133616 17100 133622 17112
rect 187102 17100 187108 17112
rect 133616 17072 187108 17100
rect 133616 17060 133622 17072
rect 187102 17060 187108 17072
rect 187160 17060 187166 17112
rect 95378 16992 95384 17044
rect 95436 17032 95442 17044
rect 135582 17032 135588 17044
rect 95436 17004 135588 17032
rect 95436 16992 95442 17004
rect 135582 16992 135588 17004
rect 135640 17032 135646 17044
rect 168518 17032 168524 17044
rect 135640 17004 168524 17032
rect 135640 16992 135646 17004
rect 168518 16992 168524 17004
rect 168576 16992 168582 17044
rect 154810 12912 154816 12964
rect 154868 12952 154874 12964
rect 156466 12952 156472 12964
rect 154868 12924 156472 12952
rect 154868 12912 154874 12924
rect 156466 12912 156472 12924
rect 156524 12912 156530 12964
rect 84338 12844 84344 12896
rect 84396 12884 84402 12896
rect 87098 12884 87104 12896
rect 84396 12856 87104 12884
rect 84396 12844 84402 12856
rect 87098 12844 87104 12856
rect 87156 12844 87162 12896
rect 156282 12708 156288 12760
rect 156340 12748 156346 12760
rect 172474 12748 172480 12760
rect 156340 12720 172480 12748
rect 156340 12708 156346 12720
rect 172474 12708 172480 12720
rect 172532 12708 172538 12760
rect 145150 12640 145156 12692
rect 145208 12680 145214 12692
rect 161802 12680 161808 12692
rect 145208 12652 161808 12680
rect 145208 12640 145214 12652
rect 161802 12640 161808 12652
rect 161860 12640 161866 12692
rect 155270 12572 155276 12624
rect 155328 12612 155334 12624
rect 177810 12612 177816 12624
rect 155328 12584 177816 12612
rect 155328 12572 155334 12584
rect 177810 12572 177816 12584
rect 177868 12572 177874 12624
rect 143770 12504 143776 12556
rect 143828 12544 143834 12556
rect 167138 12544 167144 12556
rect 143828 12516 167144 12544
rect 143828 12504 143834 12516
rect 167138 12504 167144 12516
rect 167196 12504 167202 12556
rect 154258 12436 154264 12488
rect 154316 12476 154322 12488
rect 183146 12476 183152 12488
rect 154316 12448 183152 12476
rect 154316 12436 154322 12448
rect 183146 12436 183152 12448
rect 183204 12436 183210 12488
rect 153246 12368 153252 12420
rect 153304 12408 153310 12420
rect 188482 12408 188488 12420
rect 153304 12380 188488 12408
rect 153304 12368 153310 12380
rect 188482 12368 188488 12380
rect 188540 12368 188546 12420
rect 79186 12300 79192 12352
rect 79244 12340 79250 12352
rect 97770 12340 97776 12352
rect 79244 12312 97776 12340
rect 79244 12300 79250 12312
rect 97770 12300 97776 12312
rect 97828 12300 97834 12352
rect 135122 12300 135128 12352
rect 135180 12340 135186 12352
rect 138250 12340 138256 12352
rect 135180 12312 138256 12340
rect 135180 12300 135186 12312
rect 138250 12300 138256 12312
rect 138308 12300 138314 12352
rect 140458 12300 140464 12352
rect 140516 12340 140522 12352
rect 150118 12340 150124 12352
rect 140516 12312 150124 12340
rect 140516 12300 140522 12312
rect 150118 12300 150124 12312
rect 150176 12300 150182 12352
rect 152142 12300 152148 12352
rect 152200 12340 152206 12352
rect 193818 12340 193824 12352
rect 152200 12312 193824 12340
rect 152200 12300 152206 12312
rect 193818 12300 193824 12312
rect 193876 12300 193882 12352
rect 78910 12232 78916 12284
rect 78968 12272 78974 12284
rect 103106 12272 103112 12284
rect 78968 12244 103112 12272
rect 78968 12232 78974 12244
rect 103106 12232 103112 12244
rect 103164 12232 103170 12284
rect 129786 12232 129792 12284
rect 129844 12272 129850 12284
rect 139814 12272 139820 12284
rect 129844 12244 139820 12272
rect 129844 12232 129850 12244
rect 139814 12232 139820 12244
rect 139872 12232 139878 12284
rect 151130 12232 151136 12284
rect 151188 12272 151194 12284
rect 199154 12272 199160 12284
rect 151188 12244 199160 12272
rect 151188 12232 151194 12244
rect 199154 12232 199160 12244
rect 199212 12232 199218 12284
rect 76426 12096 76432 12148
rect 76484 12136 76490 12148
rect 80290 12136 80296 12148
rect 76484 12108 80296 12136
rect 76484 12096 76490 12108
rect 80290 12096 80296 12108
rect 80348 12096 80354 12148
rect 150578 12096 150584 12148
rect 150636 12136 150642 12148
rect 151130 12136 151136 12148
rect 150636 12108 151136 12136
rect 150636 12096 150642 12108
rect 151130 12096 151136 12108
rect 151188 12096 151194 12148
rect 65754 11688 65760 11740
rect 65812 11728 65818 11740
rect 69986 11728 69992 11740
rect 65812 11700 69992 11728
rect 65812 11688 65818 11700
rect 69986 11688 69992 11700
rect 70044 11688 70050 11740
<< via1 >>
rect 80204 216504 80256 216556
rect 89772 216504 89824 216556
rect 83148 216436 83200 216488
rect 153804 216436 153856 216488
rect 155552 216436 155604 216488
rect 185820 216436 185872 216488
rect 22704 213104 22756 213156
rect 56744 213104 56796 213156
rect 66496 213104 66548 213156
rect 115072 213104 115124 213156
rect 56192 211676 56244 211728
rect 56744 211676 56796 211728
rect 96488 211676 96540 211728
rect 128872 211676 128924 211728
rect 25832 210996 25884 211048
rect 76524 210996 76576 211048
rect 121788 210996 121840 211048
rect 151596 210996 151648 211048
rect 57664 210928 57716 210980
rect 148284 210928 148336 210980
rect 28132 210588 28184 210640
rect 105964 210588 106016 210640
rect 47268 210384 47320 210436
rect 59872 210384 59924 210436
rect 69808 210316 69860 210368
rect 128872 210384 128924 210436
rect 192076 210384 192128 210436
rect 141476 210316 141528 210368
rect 156840 210316 156892 210368
rect 160336 210316 160388 210368
rect 13320 209568 13372 209620
rect 191708 209568 191760 209620
rect 88576 208956 88628 209008
rect 159048 207188 159100 207240
rect 160520 207188 160572 207240
rect 159048 206780 159100 206832
rect 160612 206780 160664 206832
rect 122156 205352 122208 205404
rect 124364 205352 124416 205404
rect 49292 204672 49344 204724
rect 50488 204672 50540 204724
rect 159048 203380 159100 203432
rect 160520 203380 160572 203432
rect 84988 202199 85040 202208
rect 84988 202165 84997 202199
rect 84997 202165 85031 202199
rect 85031 202165 85040 202199
rect 84988 202156 85040 202165
rect 120868 202020 120920 202072
rect 122432 202020 122484 202072
rect 84988 201952 85040 202004
rect 158956 201884 159008 201936
rect 160612 201884 160664 201936
rect 87196 201272 87248 201324
rect 88944 201272 88996 201324
rect 87196 199300 87248 199352
rect 88944 199300 88996 199352
rect 158956 198688 159008 198740
rect 160520 198688 160572 198740
rect 87196 197532 87248 197584
rect 88944 197532 88996 197584
rect 121788 196512 121840 196564
rect 124180 196512 124232 196564
rect 158956 195356 159008 195408
rect 160520 195356 160572 195408
rect 122248 194132 122300 194184
rect 123352 194132 123404 194184
rect 50304 192364 50356 192416
rect 50488 192364 50540 192416
rect 84528 192407 84580 192416
rect 84528 192373 84537 192407
rect 84537 192373 84571 192407
rect 84571 192373 84580 192407
rect 84528 192364 84580 192373
rect 122524 192339 122576 192348
rect 122524 192305 122533 192339
rect 122533 192305 122567 192339
rect 122567 192305 122576 192339
rect 122524 192296 122576 192305
rect 87196 192092 87248 192144
rect 88852 192092 88904 192144
rect 122156 191480 122208 191532
rect 123352 191480 123404 191532
rect 194744 191004 194796 191056
rect 196860 191004 196912 191056
rect 158956 190868 159008 190920
rect 160612 190868 160664 190920
rect 121972 188760 122024 188812
rect 123352 188760 123404 188812
rect 87196 188216 87248 188268
rect 88668 188216 88720 188268
rect 87104 186856 87156 186908
rect 88576 186856 88628 186908
rect 122892 185972 122944 186024
rect 126480 185972 126532 186024
rect 87012 185904 87064 185956
rect 88576 185904 88628 185956
rect 122984 185700 123036 185752
rect 126572 185700 126624 185752
rect 85724 185632 85776 185684
rect 88576 185632 88628 185684
rect 157484 185564 157536 185616
rect 160612 185564 160664 185616
rect 49936 185496 49988 185548
rect 52052 185496 52104 185548
rect 158864 185496 158916 185548
rect 160520 185496 160572 185548
rect 84528 185292 84580 185344
rect 84252 185224 84304 185276
rect 122892 184204 122944 184256
rect 124456 184204 124508 184256
rect 86460 184136 86512 184188
rect 88668 184136 88720 184188
rect 122340 184136 122392 184188
rect 125468 184136 125520 184188
rect 85172 184068 85224 184120
rect 88576 184068 88628 184120
rect 122984 184068 123036 184120
rect 124548 184068 124600 184120
rect 158220 184068 158272 184120
rect 160336 184068 160388 184120
rect 122616 182776 122668 182828
rect 50396 182572 50448 182624
rect 86552 182708 86604 182760
rect 88576 182708 88628 182760
rect 158312 182708 158364 182760
rect 160336 182708 160388 182760
rect 55456 182640 55508 182692
rect 122616 182640 122668 182692
rect 127584 182640 127636 182692
rect 67140 182436 67192 182488
rect 69808 182436 69860 182488
rect 70452 182436 70504 182488
rect 74040 182436 74092 182488
rect 143684 182436 143736 182488
rect 147548 182436 147600 182488
rect 66036 182368 66088 182420
rect 68336 182368 68388 182420
rect 69348 182368 69400 182420
rect 72660 182368 72712 182420
rect 137244 182368 137296 182420
rect 138992 182368 139044 182420
rect 139452 182368 139504 182420
rect 141844 182368 141896 182420
rect 142764 182368 142816 182420
rect 146076 182368 146128 182420
rect 68244 182300 68296 182352
rect 71188 182300 71240 182352
rect 144880 182300 144932 182352
rect 148928 182300 148980 182352
rect 146076 182232 146128 182284
rect 150400 182232 150452 182284
rect 134944 182164 134996 182216
rect 136140 182164 136192 182216
rect 73764 182028 73816 182080
rect 78364 182028 78416 182080
rect 136140 182028 136192 182080
rect 137520 182028 137572 182080
rect 138164 181960 138216 182012
rect 140372 181960 140424 182012
rect 61528 181892 61580 181944
rect 62632 181892 62684 181944
rect 147180 181824 147232 181876
rect 151780 181824 151832 181876
rect 62632 181756 62684 181808
rect 64104 181756 64156 181808
rect 74868 181756 74920 181808
rect 79744 181756 79796 181808
rect 64932 181416 64984 181468
rect 66956 181416 67008 181468
rect 72660 181416 72712 181468
rect 76892 181416 76944 181468
rect 140556 181416 140608 181468
rect 143224 181416 143276 181468
rect 148284 181416 148336 181468
rect 153252 181416 153304 181468
rect 63828 181348 63880 181400
rect 65484 181348 65536 181400
rect 71556 181348 71608 181400
rect 75512 181348 75564 181400
rect 141660 181348 141712 181400
rect 144696 181348 144748 181400
rect 175700 181348 175752 181400
rect 176436 181348 176488 181400
rect 20864 181280 20916 181332
rect 26108 181280 26160 181332
rect 29972 181280 30024 181332
rect 31352 181280 31404 181332
rect 31904 181280 31956 181332
rect 32824 181280 32876 181332
rect 33192 181280 33244 181332
rect 33652 181280 33704 181332
rect 36872 181280 36924 181332
rect 37700 181280 37752 181332
rect 38896 181280 38948 181332
rect 41012 181280 41064 181332
rect 106700 181280 106752 181332
rect 107988 181280 108040 181332
rect 108356 181280 108408 181332
rect 109828 181280 109880 181332
rect 130436 181280 130488 181332
rect 190972 181280 191024 181332
rect 27764 181212 27816 181264
rect 30432 181212 30484 181264
rect 37424 181212 37476 181264
rect 38436 181212 38488 181264
rect 107160 181212 107212 181264
rect 108172 181212 108224 181264
rect 168984 181212 169036 181264
rect 170456 181212 170508 181264
rect 176436 181212 176488 181264
rect 177264 181212 177316 181264
rect 177540 181212 177592 181264
rect 178276 181212 178328 181264
rect 179104 181212 179156 181264
rect 180484 181212 180536 181264
rect 182876 181212 182928 181264
rect 186004 181212 186056 181264
rect 37700 181144 37752 181196
rect 39080 181144 39132 181196
rect 40460 181144 40512 181196
rect 43588 181144 43640 181196
rect 106240 181144 106292 181196
rect 107068 181144 107120 181196
rect 107528 181144 107580 181196
rect 108724 181144 108776 181196
rect 109092 181144 109144 181196
rect 110932 181144 110984 181196
rect 168432 181144 168484 181196
rect 170088 181144 170140 181196
rect 176804 181144 176856 181196
rect 177816 181144 177868 181196
rect 178092 181144 178144 181196
rect 179380 181144 179432 181196
rect 182416 181144 182468 181196
rect 185452 181144 185504 181196
rect 38436 181076 38488 181128
rect 40368 181076 40420 181128
rect 177632 181076 177684 181128
rect 178828 181076 178880 181128
rect 181220 181076 181272 181128
rect 183796 181076 183848 181128
rect 28592 181008 28644 181060
rect 30892 181008 30944 181060
rect 40092 181008 40144 181060
rect 43036 181008 43088 181060
rect 108724 181008 108776 181060
rect 110748 181008 110800 181060
rect 183612 181008 183664 181060
rect 187108 181008 187160 181060
rect 163188 180940 163240 180992
rect 167880 180940 167932 180992
rect 180852 180940 180904 180992
rect 183244 180940 183296 180992
rect 27304 180872 27356 180924
rect 30064 180872 30116 180924
rect 39632 180872 39684 180924
rect 42300 180872 42352 180924
rect 99340 180872 99392 180924
rect 99800 180872 99852 180924
rect 181680 180872 181732 180924
rect 184348 180872 184400 180924
rect 183244 180804 183296 180856
rect 186556 180804 186608 180856
rect 105964 180736 106016 180788
rect 106516 180736 106568 180788
rect 182048 180736 182100 180788
rect 184900 180736 184952 180788
rect 39264 180600 39316 180652
rect 41748 180600 41800 180652
rect 168524 180600 168576 180652
rect 190420 180600 190472 180652
rect 26384 180532 26436 180584
rect 27856 180532 27908 180584
rect 178460 180532 178512 180584
rect 179932 180532 179984 180584
rect 30524 180464 30576 180516
rect 32088 180464 32140 180516
rect 24728 180396 24780 180448
rect 26568 180396 26620 180448
rect 25372 180328 25424 180380
rect 28868 180328 28920 180380
rect 31260 180328 31312 180380
rect 32456 180328 32508 180380
rect 22796 180260 22848 180312
rect 26384 180260 26436 180312
rect 92164 180260 92216 180312
rect 94372 180260 94424 180312
rect 110564 180260 110616 180312
rect 113508 180260 113560 180312
rect 23440 180192 23492 180244
rect 25372 180192 25424 180244
rect 26016 180192 26068 180244
rect 27948 180192 28000 180244
rect 29144 180192 29196 180244
rect 31260 180192 31312 180244
rect 92440 180192 92492 180244
rect 93268 180192 93320 180244
rect 98880 180192 98932 180244
rect 99616 180192 99668 180244
rect 107804 180192 107856 180244
rect 109368 180192 109420 180244
rect 111116 180192 111168 180244
rect 113692 180192 113744 180244
rect 24084 180124 24136 180176
rect 27764 180124 27816 180176
rect 21508 180056 21560 180108
rect 26476 180056 26528 180108
rect 38068 180056 38120 180108
rect 39724 180056 39776 180108
rect 92716 180124 92768 180176
rect 111576 180124 111628 180176
rect 114244 180124 114296 180176
rect 169536 180124 169588 180176
rect 170824 180124 170876 180176
rect 179288 180124 179340 180176
rect 181036 180124 181088 180176
rect 92348 180056 92400 180108
rect 94924 180056 94976 180108
rect 97776 180056 97828 180108
rect 98696 180056 98748 180108
rect 110288 180056 110340 180108
rect 112588 180056 112640 180108
rect 180760 180056 180812 180108
rect 182692 180056 182744 180108
rect 184072 180056 184124 180108
rect 187660 180056 187712 180108
rect 22152 179988 22204 180040
rect 26844 179988 26896 180040
rect 91980 179988 92032 180040
rect 92072 179988 92124 180040
rect 92440 179988 92492 180040
rect 92624 179988 92676 180040
rect 95476 179988 95528 180040
rect 97224 179988 97276 180040
rect 98236 179988 98288 180040
rect 109920 179988 109972 180040
rect 112036 179988 112088 180040
rect 112220 179988 112272 180040
rect 115348 179988 115400 180040
rect 170640 179988 170692 180040
rect 171652 179988 171704 180040
rect 179656 179988 179708 180040
rect 181588 179988 181640 180040
rect 36228 179920 36280 179972
rect 92256 179920 92308 179972
rect 94096 179920 94148 179972
rect 96672 179920 96724 179972
rect 97776 179920 97828 179972
rect 98144 179920 98196 179972
rect 98972 179920 99024 179972
rect 100720 179920 100772 179972
rect 100996 179920 101048 179972
rect 105044 179920 105096 179972
rect 105504 179920 105556 179972
rect 109552 179920 109604 179972
rect 111484 179920 111536 179972
rect 111944 179920 111996 179972
rect 114796 179920 114848 179972
rect 171192 179920 171244 179972
rect 172020 179920 172072 179972
rect 180024 179920 180076 179972
rect 182140 179920 182192 179972
rect 36044 179852 36096 179904
rect 163096 179852 163148 179904
rect 163280 179852 163332 179904
rect 113048 178492 113100 178544
rect 116452 178492 116504 178544
rect 126572 178492 126624 178544
rect 127676 178492 127728 178544
rect 25372 178424 25424 178476
rect 27672 178424 27724 178476
rect 81584 178424 81636 178476
rect 85172 178424 85224 178476
rect 113508 178424 113560 178476
rect 117004 178424 117056 178476
rect 112680 178356 112732 178408
rect 116268 178356 116320 178408
rect 124456 178356 124508 178408
rect 126664 178356 126716 178408
rect 52052 178288 52104 178340
rect 56008 178288 56060 178340
rect 26384 178152 26436 178204
rect 27304 178152 27356 178204
rect 83792 178152 83844 178204
rect 86460 178152 86512 178204
rect 80480 178016 80532 178068
rect 87840 178016 87892 178068
rect 113968 178016 114020 178068
rect 117556 178016 117608 178068
rect 153896 178016 153948 178068
rect 161072 178016 161124 178068
rect 82688 177948 82740 178000
rect 89220 177948 89272 178000
rect 151688 177948 151740 178000
rect 158312 177948 158364 178000
rect 122432 177880 122484 177932
rect 129976 177880 130028 177932
rect 50672 177812 50724 177864
rect 58216 177812 58268 177864
rect 58308 177812 58360 177864
rect 88208 177812 88260 177864
rect 128596 177812 128648 177864
rect 161072 177812 161124 177864
rect 41656 177744 41708 177796
rect 45796 177744 45848 177796
rect 154632 177744 154684 177796
rect 161256 177744 161308 177796
rect 27856 177676 27908 177728
rect 29696 177676 29748 177728
rect 50120 177676 50172 177728
rect 53800 177676 53852 177728
rect 126480 177676 126532 177728
rect 128780 177676 128832 177728
rect 159416 177676 159468 177728
rect 160980 177676 161032 177728
rect 185268 177676 185320 177728
rect 189316 177676 189368 177728
rect 27948 177608 28000 177660
rect 29236 177608 29288 177660
rect 33376 177608 33428 177660
rect 34112 177608 34164 177660
rect 41288 177608 41340 177660
rect 44876 177608 44928 177660
rect 50028 177608 50080 177660
rect 52696 177608 52748 177660
rect 75972 177608 76024 177660
rect 80296 177608 80348 177660
rect 84896 177608 84948 177660
rect 85724 177608 85776 177660
rect 99708 177608 99760 177660
rect 100168 177608 100220 177660
rect 100260 177608 100312 177660
rect 100720 177608 100772 177660
rect 104216 177608 104268 177660
rect 104676 177608 104728 177660
rect 156104 177608 156156 177660
rect 158220 177608 158272 177660
rect 158312 177608 158364 177660
rect 158864 177608 158916 177660
rect 169996 177608 170048 177660
rect 171284 177608 171336 177660
rect 172848 177608 172900 177660
rect 173216 177608 173268 177660
rect 175608 177608 175660 177660
rect 176160 177608 176212 177660
rect 184440 177608 184492 177660
rect 188212 177608 188264 177660
rect 152792 177540 152844 177592
rect 159600 177540 159652 177592
rect 185636 177540 185688 177592
rect 189868 177540 189920 177592
rect 50212 177472 50264 177524
rect 54904 177472 54956 177524
rect 86000 177472 86052 177524
rect 87012 177472 87064 177524
rect 105504 177472 105556 177524
rect 106148 177472 106200 177524
rect 26568 177404 26620 177456
rect 28500 177404 28552 177456
rect 79376 177404 79428 177456
rect 86552 177404 86604 177456
rect 184808 177404 184860 177456
rect 188764 177404 188816 177456
rect 40828 177336 40880 177388
rect 44416 177336 44468 177388
rect 51960 177336 52012 177388
rect 57112 177336 57164 177388
rect 31996 177268 32048 177320
rect 33284 177268 33336 177320
rect 171744 177200 171796 177252
rect 172480 177200 172532 177252
rect 164384 174004 164436 174056
rect 167144 174004 167196 174056
rect 188028 172984 188080 173036
rect 196952 172984 197004 173036
rect 164292 172780 164344 172832
rect 166776 172780 166828 172832
rect 92624 171692 92676 171744
rect 95016 171692 95068 171744
rect 164016 171556 164068 171608
rect 166224 171556 166276 171608
rect 163372 170332 163424 170384
rect 165672 170332 165724 170384
rect 163188 169108 163240 169160
rect 165120 169108 165172 169160
rect 91704 168904 91756 168956
rect 94832 168904 94884 168956
rect 114060 168904 114112 168956
rect 118936 168904 118988 168956
rect 13320 167544 13372 167596
rect 22244 167544 22296 167596
rect 163188 165912 163240 165964
rect 167512 165912 167564 165964
rect 91980 165844 92032 165896
rect 94556 165844 94608 165896
rect 116544 164756 116596 164808
rect 119580 164756 119632 164808
rect 188028 164756 188080 164808
rect 197596 164756 197648 164808
rect 164292 164348 164344 164400
rect 167328 164348 167380 164400
rect 164292 163124 164344 163176
rect 167236 163124 167288 163176
rect 164476 162104 164528 162156
rect 168432 162104 168484 162156
rect 92624 161900 92676 161952
rect 95384 161900 95436 161952
rect 164292 161900 164344 161952
rect 167972 161900 168024 161952
rect 91980 161152 92032 161204
rect 94188 161152 94240 161204
rect 91980 160540 92032 160592
rect 94096 160540 94148 160592
rect 164292 160540 164344 160592
rect 168524 160608 168576 160660
rect 91980 159180 92032 159232
rect 94004 159180 94056 159232
rect 164292 158228 164344 158280
rect 168524 158228 168576 158280
rect 91796 157208 91848 157260
rect 94004 157208 94056 157260
rect 164292 156936 164344 156988
rect 168524 156936 168576 156988
rect 45060 156392 45112 156444
rect 47820 156392 47872 156444
rect 164384 155304 164436 155356
rect 167144 155304 167196 155356
rect 13412 155100 13464 155152
rect 22336 155100 22388 155152
rect 163372 154488 163424 154540
rect 167144 154488 167196 154540
rect 91428 154080 91480 154132
rect 94740 154080 94792 154132
rect 91796 152516 91848 152568
rect 95384 152516 95436 152568
rect 164384 152380 164436 152432
rect 167236 152380 167288 152432
rect 91704 151564 91756 151616
rect 94188 151564 94240 151616
rect 164384 151496 164436 151548
rect 167328 151496 167380 151548
rect 164384 149728 164436 149780
rect 167144 149728 167196 149780
rect 91428 149592 91480 149644
rect 94004 149592 94056 149644
rect 163924 149592 163976 149644
rect 167236 149592 167288 149644
rect 164384 148504 164436 148556
rect 167052 148504 167104 148556
rect 13320 146804 13372 146856
rect 22336 146804 22388 146856
rect 91428 146804 91480 146856
rect 93544 146804 93596 146856
rect 164384 146804 164436 146856
rect 167880 146804 167932 146856
rect 164384 145444 164436 145496
rect 167972 145444 168024 145496
rect 91336 143540 91388 143592
rect 94372 143540 94424 143592
rect 91796 142724 91848 142776
rect 95660 142724 95712 142776
rect 91704 142656 91756 142708
rect 95384 142656 95436 142708
rect 116820 142588 116872 142640
rect 118936 142588 118988 142640
rect 164384 141568 164436 141620
rect 167052 141568 167104 141620
rect 91704 141475 91756 141484
rect 91704 141441 91713 141475
rect 91713 141441 91747 141475
rect 91747 141441 91756 141475
rect 91704 141432 91756 141441
rect 91796 141296 91848 141348
rect 95016 141296 95068 141348
rect 92532 140004 92584 140056
rect 93452 140004 93504 140056
rect 164292 140004 164344 140056
rect 166408 140004 166460 140056
rect 92624 139936 92676 139988
rect 93912 139936 93964 139988
rect 164384 139936 164436 139988
rect 165856 139936 165908 139988
rect 188028 139188 188080 139240
rect 192076 139188 192128 139240
rect 193456 139188 193508 139240
rect 48464 134700 48516 134752
rect 82136 134360 82188 134412
rect 84344 134360 84396 134412
rect 145156 134360 145208 134412
rect 23624 134224 23676 134276
rect 27672 134224 27724 134276
rect 73212 134224 73264 134276
rect 83608 134224 83660 134276
rect 84344 134224 84396 134276
rect 66588 134156 66640 134208
rect 82136 134088 82188 134140
rect 138256 134156 138308 134208
rect 182416 134020 182468 134072
rect 186372 134020 186424 134072
rect 27028 133952 27080 134004
rect 29696 133952 29748 134004
rect 38436 133952 38488 134004
rect 41564 133952 41616 134004
rect 26292 133884 26344 133936
rect 29236 133884 29288 133936
rect 37700 133884 37752 133936
rect 40644 133884 40696 133936
rect 28316 133816 28368 133868
rect 30432 133816 30484 133868
rect 31076 133816 31128 133868
rect 32088 133816 32140 133868
rect 37240 133816 37292 133868
rect 40000 133816 40052 133868
rect 40828 133816 40880 133868
rect 43588 133816 43640 133868
rect 29696 133748 29748 133800
rect 31260 133748 31312 133800
rect 34848 133748 34900 133800
rect 35860 133748 35912 133800
rect 36504 133748 36556 133800
rect 38620 133748 38672 133800
rect 41288 133748 41340 133800
rect 44324 133748 44376 133800
rect 27672 133680 27724 133732
rect 30064 133680 30116 133732
rect 40460 133680 40512 133732
rect 43036 133680 43088 133732
rect 62356 133680 62408 133732
rect 86552 133680 86604 133732
rect 38068 133612 38120 133664
rect 41012 133612 41064 133664
rect 114060 133952 114112 134004
rect 182876 133952 182928 134004
rect 186464 133952 186516 134004
rect 107528 133884 107580 133936
rect 110196 133884 110248 133936
rect 169260 133884 169312 133936
rect 170456 133884 170508 133936
rect 178460 133884 178512 133936
rect 180668 133884 180720 133936
rect 181220 133884 181272 133936
rect 184716 133884 184768 133936
rect 169904 133816 169956 133868
rect 170824 133816 170876 133868
rect 175608 133816 175660 133868
rect 176712 133816 176764 133868
rect 177264 133816 177316 133868
rect 179012 133816 179064 133868
rect 184440 133816 184492 133868
rect 186832 133816 186884 133868
rect 109000 133748 109052 133800
rect 110840 133748 110892 133800
rect 113968 133748 114020 133800
rect 119488 133748 119540 133800
rect 168708 133748 168760 133800
rect 170088 133748 170140 133800
rect 170456 133748 170508 133800
rect 171284 133748 171336 133800
rect 175240 133748 175292 133800
rect 176160 133748 176212 133800
rect 176436 133748 176488 133800
rect 177816 133748 177868 133800
rect 183612 133748 183664 133800
rect 185544 133748 185596 133800
rect 110288 133680 110340 133732
rect 113232 133680 113284 133732
rect 113324 133680 113376 133732
rect 118936 133680 118988 133732
rect 174872 133680 174924 133732
rect 175608 133680 175660 133732
rect 176804 133680 176856 133732
rect 178460 133680 178512 133732
rect 184072 133680 184124 133732
rect 186648 133680 186700 133732
rect 108356 133612 108408 133664
rect 111392 133612 111444 133664
rect 181680 133612 181732 133664
rect 185084 133612 185136 133664
rect 39264 133544 39316 133596
rect 42944 133544 42996 133596
rect 109920 133544 109972 133596
rect 113324 133544 113376 133596
rect 149664 133544 149716 133596
rect 151596 133544 151648 133596
rect 184808 133544 184860 133596
rect 187292 133544 187344 133596
rect 39632 133476 39684 133528
rect 41840 133476 41892 133528
rect 108724 133476 108776 133528
rect 111944 133476 111996 133528
rect 177632 133476 177684 133528
rect 179564 133476 179616 133528
rect 180852 133476 180904 133528
rect 182508 133476 182560 133528
rect 29052 133408 29104 133460
rect 30892 133408 30944 133460
rect 34480 133408 34532 133460
rect 35216 133408 35268 133460
rect 36872 133408 36924 133460
rect 39264 133408 39316 133460
rect 40092 133408 40144 133460
rect 42300 133408 42352 133460
rect 107160 133408 107212 133460
rect 109644 133408 109696 133460
rect 183244 133408 183296 133460
rect 185728 133408 185780 133460
rect 25004 133340 25056 133392
rect 26108 133340 26160 133392
rect 38896 133340 38948 133392
rect 42668 133340 42720 133392
rect 107804 133340 107856 133392
rect 110564 133340 110616 133392
rect 111484 133340 111536 133392
rect 114428 133340 114480 133392
rect 180024 133340 180076 133392
rect 182968 133340 183020 133392
rect 30432 133272 30484 133324
rect 31628 133272 31680 133324
rect 106700 133272 106752 133324
rect 109000 133272 109052 133324
rect 111116 133272 111168 133324
rect 113416 133272 113468 133324
rect 176068 133272 176120 133324
rect 177264 133272 177316 133324
rect 178092 133272 178144 133324
rect 180116 133272 180168 133324
rect 182048 133272 182100 133324
rect 184808 133272 184860 133324
rect 24912 133204 24964 133256
rect 28500 133204 28552 133256
rect 105504 133204 105556 133256
rect 107252 133204 107304 133256
rect 111852 133204 111904 133256
rect 114704 133204 114756 133256
rect 179288 133204 179340 133256
rect 181864 133204 181916 133256
rect 185268 133204 185320 133256
rect 190420 133204 190472 133256
rect 24268 133136 24320 133188
rect 28040 133136 28092 133188
rect 35676 133136 35728 133188
rect 37240 133136 37292 133188
rect 103572 133136 103624 133188
rect 104952 133136 105004 133188
rect 105044 133136 105096 133188
rect 106700 133136 106752 133188
rect 110472 133136 110524 133188
rect 112588 133136 112640 133188
rect 112680 133136 112732 133188
rect 116084 133136 116136 133188
rect 178828 133136 178880 133188
rect 181312 133136 181364 133188
rect 25648 133068 25700 133120
rect 28868 133068 28920 133120
rect 35308 133068 35360 133120
rect 36504 133068 36556 133120
rect 41656 133068 41708 133120
rect 47452 133068 47504 133120
rect 96764 133068 96816 133120
rect 97776 133068 97828 133120
rect 97960 133068 98012 133120
rect 98604 133068 98656 133120
rect 103480 133068 103532 133120
rect 104400 133068 104452 133120
rect 104676 133068 104728 133120
rect 106148 133068 106200 133120
rect 106332 133068 106384 133120
rect 108448 133068 108500 133120
rect 112312 133068 112364 133120
rect 114796 133068 114848 133120
rect 180484 133068 180536 133120
rect 183520 133068 183572 133120
rect 22888 133000 22940 133052
rect 27304 133000 27356 133052
rect 36044 133000 36096 133052
rect 37884 133000 37936 133052
rect 97408 133000 97460 133052
rect 98236 133000 98288 133052
rect 103112 133000 103164 133052
rect 103756 133000 103808 133052
rect 104308 133000 104360 133052
rect 105504 133000 105556 133052
rect 105964 133000 106016 133052
rect 107896 133000 107948 133052
rect 109552 133000 109604 133052
rect 112772 133000 112824 133052
rect 113140 133000 113192 133052
rect 115716 133000 115768 133052
rect 179656 133000 179708 133052
rect 182416 133000 182468 133052
rect 185636 133000 185688 133052
rect 190972 133000 191024 133052
rect 92072 131572 92124 131624
rect 92716 131572 92768 131624
rect 93452 131572 93504 131624
rect 94464 131572 94516 131624
rect 110840 131572 110892 131624
rect 112496 131572 112548 131624
rect 116084 131572 116136 131624
rect 117740 131572 117792 131624
rect 114428 131504 114480 131556
rect 115992 131504 116044 131556
rect 21508 131368 21560 131420
rect 26476 131368 26528 131420
rect 43588 131368 43640 131420
rect 46072 131368 46124 131420
rect 114704 131368 114756 131420
rect 116636 131368 116688 131420
rect 22244 131232 22296 131284
rect 26844 131232 26896 131284
rect 113232 131232 113284 131284
rect 114244 131232 114296 131284
rect 114796 131232 114848 131284
rect 117188 131232 117240 131284
rect 44324 131096 44376 131148
rect 46808 131096 46860 131148
rect 91980 131096 92032 131148
rect 96212 131096 96264 131148
rect 113416 131096 113468 131148
rect 115440 131096 115492 131148
rect 115716 130960 115768 131012
rect 118384 130960 118436 131012
rect 20220 130892 20272 130944
rect 44416 130892 44468 130944
rect 168524 130892 168576 130944
rect 191524 130892 191576 130944
rect 112588 130688 112640 130740
rect 114888 130688 114940 130740
rect 185636 130552 185688 130604
rect 188120 130552 188172 130604
rect 185728 130484 185780 130536
rect 187568 130484 187620 130536
rect 43036 130416 43088 130468
rect 45428 130416 45480 130468
rect 163740 130416 163792 130468
rect 168156 130416 168208 130468
rect 186832 130416 186884 130468
rect 189224 130416 189276 130468
rect 42300 130348 42352 130400
rect 44692 130348 44744 130400
rect 163832 130348 163884 130400
rect 167604 130348 167656 130400
rect 186648 130348 186700 130400
rect 188672 130348 188724 130400
rect 20864 130280 20916 130332
rect 25004 130280 25056 130332
rect 41840 130280 41892 130332
rect 44048 130280 44100 130332
rect 163924 130280 163976 130332
rect 165304 130280 165356 130332
rect 182508 130280 182560 130332
rect 184164 130280 184216 130332
rect 184808 130280 184860 130332
rect 185820 130280 185872 130332
rect 187292 130280 187344 130332
rect 189868 130280 189920 130332
rect 121696 126880 121748 126932
rect 123996 126880 124048 126932
rect 121788 126200 121840 126252
rect 124364 126200 124416 126252
rect 121696 126132 121748 126184
rect 123904 126132 123956 126184
rect 121696 125112 121748 125164
rect 123720 125112 123772 125164
rect 87748 124568 87800 124620
rect 88760 124568 88812 124620
rect 121696 123480 121748 123532
rect 123536 123480 123588 123532
rect 121696 122120 121748 122172
rect 123444 122120 123496 122172
rect 121696 121984 121748 122036
rect 123352 121984 123404 122036
rect 121696 120896 121748 120948
rect 124364 120896 124416 120948
rect 121696 119332 121748 119384
rect 124272 119332 124324 119384
rect 51132 119264 51184 119316
rect 51592 119264 51644 119316
rect 121696 118176 121748 118228
rect 124364 118176 124416 118228
rect 123076 116544 123128 116596
rect 124272 116544 124324 116596
rect 50580 116476 50632 116528
rect 51592 116476 51644 116528
rect 121696 115660 121748 115712
rect 124364 115660 124416 115712
rect 121696 115388 121748 115440
rect 123996 115388 124048 115440
rect 121696 115116 121748 115168
rect 124272 115116 124324 115168
rect 159048 115116 159100 115168
rect 160612 115116 160664 115168
rect 121696 113960 121748 114012
rect 123444 113960 123496 114012
rect 121696 112328 121748 112380
rect 123352 112328 123404 112380
rect 51224 111240 51276 111292
rect 51592 111240 51644 111292
rect 51224 111104 51276 111156
rect 51684 111104 51736 111156
rect 121696 110968 121748 111020
rect 124272 110968 124324 111020
rect 121696 109744 121748 109796
rect 124364 109744 124416 109796
rect 121696 108724 121748 108776
rect 123444 108724 123496 108776
rect 51224 108520 51276 108572
rect 51592 108520 51644 108572
rect 85172 106863 85224 106872
rect 85172 106829 85181 106863
rect 85181 106829 85215 106863
rect 85215 106829 85224 106863
rect 85172 106820 85224 106829
rect 121696 106820 121748 106872
rect 124272 106820 124324 106872
rect 121696 105868 121748 105920
rect 124364 105868 124416 105920
rect 121696 105596 121748 105648
rect 124180 105596 124232 105648
rect 91060 104687 91112 104696
rect 91060 104653 91069 104687
rect 91069 104653 91103 104687
rect 91103 104653 91112 104687
rect 91060 104644 91112 104653
rect 85908 104100 85960 104152
rect 88668 104100 88720 104152
rect 121788 104100 121840 104152
rect 126940 104100 126992 104152
rect 85816 104032 85868 104084
rect 88576 104032 88628 104084
rect 121696 104032 121748 104084
rect 127032 104032 127084 104084
rect 157576 104032 157628 104084
rect 160336 104032 160388 104084
rect 50764 103012 50816 103064
rect 54076 103012 54128 103064
rect 121696 102808 121748 102860
rect 124548 102808 124600 102860
rect 51224 102740 51276 102792
rect 55364 102740 55416 102792
rect 121788 102740 121840 102792
rect 125928 102740 125980 102792
rect 127124 102740 127176 102792
rect 121880 102672 121932 102724
rect 81584 101380 81636 101432
rect 88668 101380 88720 101432
rect 152792 101380 152844 101432
rect 160428 101380 160480 101432
rect 51224 101312 51276 101364
rect 52604 101312 52656 101364
rect 80480 101312 80532 101364
rect 88576 101312 88628 101364
rect 153896 101312 153948 101364
rect 160336 101312 160388 101364
rect 18012 101244 18064 101296
rect 58400 101244 58452 101296
rect 128964 101244 129016 101296
rect 193548 101244 193600 101296
rect 116360 101040 116412 101092
rect 127584 101040 127636 101092
rect 73764 100768 73816 100820
rect 78364 100768 78416 100820
rect 127584 100564 127636 100616
rect 190604 100564 190656 100616
rect 193456 100564 193508 100616
rect 71556 100360 71608 100412
rect 69348 100156 69400 100208
rect 72660 100156 72712 100208
rect 75512 100156 75564 100208
rect 64932 100088 64984 100140
rect 66956 100088 67008 100140
rect 68244 100088 68296 100140
rect 71188 100088 71240 100140
rect 145984 100156 146036 100208
rect 150400 100156 150452 100208
rect 75972 100088 76024 100140
rect 81216 100088 81268 100140
rect 95936 100088 95988 100140
rect 116360 100088 116412 100140
rect 144972 100088 145024 100140
rect 148928 100088 148980 100140
rect 56744 100020 56796 100072
rect 67140 100020 67192 100072
rect 69808 100020 69860 100072
rect 70452 100020 70504 100072
rect 74040 100020 74092 100072
rect 74868 100020 74920 100072
rect 79744 100020 79796 100072
rect 141660 100020 141712 100072
rect 144696 100020 144748 100072
rect 148284 100020 148336 100072
rect 153252 100020 153304 100072
rect 63828 99952 63880 100004
rect 65484 99952 65536 100004
rect 66036 99952 66088 100004
rect 68336 99952 68388 100004
rect 72660 99952 72712 100004
rect 76892 99952 76944 100004
rect 136048 99952 136100 100004
rect 137520 99952 137572 100004
rect 138164 99952 138216 100004
rect 140372 99952 140424 100004
rect 140556 99952 140608 100004
rect 143224 99952 143276 100004
rect 143684 99952 143736 100004
rect 147548 99952 147600 100004
rect 59320 99884 59372 99936
rect 59780 99884 59832 99936
rect 60424 99884 60476 99936
rect 61252 99884 61304 99936
rect 61528 99884 61580 99936
rect 62632 99884 62684 99936
rect 63000 99884 63052 99936
rect 64104 99884 64156 99936
rect 95936 99884 95988 99936
rect 97040 99884 97092 99936
rect 130436 99884 130488 99936
rect 131264 99884 131316 99936
rect 131816 99884 131868 99936
rect 132552 99884 132604 99936
rect 133288 99884 133340 99936
rect 133840 99884 133892 99936
rect 134668 99884 134720 99936
rect 134944 99884 134996 99936
rect 136140 99884 136192 99936
rect 137244 99884 137296 99936
rect 138992 99884 139044 99936
rect 139452 99884 139504 99936
rect 141844 99884 141896 99936
rect 142764 99884 142816 99936
rect 146076 99884 146128 99936
rect 147180 99884 147232 99936
rect 151780 99884 151832 99936
rect 154632 99884 154684 99936
rect 160980 99884 161032 99936
rect 56928 98456 56980 98508
rect 97132 98456 97184 98508
rect 93360 98252 93412 98304
rect 94372 98252 94424 98304
rect 92164 98116 92216 98168
rect 94096 98116 94148 98168
rect 171008 98116 171060 98168
rect 171652 98116 171704 98168
rect 182232 98116 182284 98168
rect 183520 98116 183572 98168
rect 92348 98048 92400 98100
rect 94924 98048 94976 98100
rect 21784 97776 21836 97828
rect 23624 97776 23676 97828
rect 168524 97776 168576 97828
rect 191524 97776 191576 97828
rect 179748 97640 179800 97692
rect 181864 97640 181916 97692
rect 181588 97504 181640 97556
rect 182416 97504 182468 97556
rect 23256 97436 23308 97488
rect 24912 97436 24964 97488
rect 27304 97300 27356 97352
rect 29052 97300 29104 97352
rect 105228 97300 105280 97352
rect 107068 97300 107120 97352
rect 163832 97300 163884 97352
rect 167604 97300 167656 97352
rect 169260 97300 169312 97352
rect 170456 97300 170508 97352
rect 23532 97232 23584 97284
rect 24544 97164 24596 97216
rect 28592 97232 28644 97284
rect 30432 97232 30484 97284
rect 30524 97232 30576 97284
rect 31628 97232 31680 97284
rect 37608 97232 37660 97284
rect 39724 97232 39776 97284
rect 40368 97232 40420 97284
rect 42300 97232 42352 97284
rect 103756 97232 103808 97284
rect 105412 97232 105464 97284
rect 106608 97232 106660 97284
rect 108724 97232 108776 97284
rect 163740 97232 163792 97284
rect 165304 97232 165356 97284
rect 169904 97232 169956 97284
rect 170824 97232 170876 97284
rect 184440 97232 184492 97284
rect 186372 97232 186424 97284
rect 26016 97164 26068 97216
rect 27672 97096 27724 97148
rect 29144 97164 29196 97216
rect 28868 97096 28920 97148
rect 30064 97164 30116 97216
rect 31260 97164 31312 97216
rect 31352 97164 31404 97216
rect 30892 97096 30944 97148
rect 36044 97096 36096 97148
rect 37516 97164 37568 97216
rect 36504 97096 36556 97148
rect 38252 97096 38304 97148
rect 28040 97028 28092 97080
rect 32088 97028 32140 97080
rect 35676 97028 35728 97080
rect 36964 97028 37016 97080
rect 37148 97028 37200 97080
rect 38988 97164 39040 97216
rect 38436 97096 38488 97148
rect 41012 97164 41064 97216
rect 92440 97164 92492 97216
rect 93268 97164 93320 97216
rect 40828 97096 40880 97148
rect 45888 97096 45940 97148
rect 85908 97096 85960 97148
rect 87104 97096 87156 97148
rect 103480 97096 103532 97148
rect 105136 97164 105188 97216
rect 104676 97096 104728 97148
rect 106516 97164 106568 97216
rect 105872 97096 105924 97148
rect 108172 97164 108224 97216
rect 107160 97096 107212 97148
rect 109828 97164 109880 97216
rect 108356 97096 108408 97148
rect 111484 97164 111536 97216
rect 165120 97164 165172 97216
rect 165856 97164 165908 97216
rect 168708 97164 168760 97216
rect 170088 97164 170140 97216
rect 176896 97164 176948 97216
rect 178460 97164 178512 97216
rect 123076 97096 123128 97148
rect 124456 97096 124508 97148
rect 127124 97096 127176 97148
rect 127676 97096 127728 97148
rect 154632 97096 154684 97148
rect 160520 97096 160572 97148
rect 176436 97096 176488 97148
rect 177816 97096 177868 97148
rect 178092 97096 178144 97148
rect 180116 97164 180168 97216
rect 179656 97096 179708 97148
rect 181588 97096 181640 97148
rect 182968 97164 183020 97216
rect 38896 97028 38948 97080
rect 40368 97028 40420 97080
rect 40460 97028 40512 97080
rect 45060 97028 45112 97080
rect 50948 97028 51000 97080
rect 57112 97028 57164 97080
rect 105504 97028 105556 97080
rect 107988 97028 108040 97080
rect 126940 97028 126992 97080
rect 129976 97028 130028 97080
rect 176068 97028 176120 97080
rect 177264 97028 177316 97080
rect 177632 97028 177684 97080
rect 179564 97028 179616 97080
rect 180024 97028 180076 97080
rect 20956 96960 21008 97012
rect 26108 96960 26160 97012
rect 26844 96960 26896 97012
rect 37700 96960 37752 97012
rect 40184 96960 40236 97012
rect 107528 96960 107580 97012
rect 110748 96960 110800 97012
rect 178460 96960 178512 97012
rect 180668 96960 180720 97012
rect 181220 96960 181272 97012
rect 184716 97164 184768 97216
rect 184808 97096 184860 97148
rect 189868 97096 189920 97148
rect 185636 97028 185688 97080
rect 190972 97028 191024 97080
rect 184072 96960 184124 97012
rect 188672 96960 188724 97012
rect 41288 96892 41340 96944
rect 46532 96892 46584 96944
rect 107804 96892 107856 96944
rect 110932 96892 110984 96944
rect 165948 96892 166000 96944
rect 166684 96892 166736 96944
rect 177264 96892 177316 96944
rect 179012 96892 179064 96944
rect 182048 96892 182100 96944
rect 185820 96892 185872 96944
rect 24912 96824 24964 96876
rect 27304 96824 27356 96876
rect 27856 96824 27908 96876
rect 30064 96824 30116 96876
rect 41656 96824 41708 96876
rect 47176 96824 47228 96876
rect 51408 96824 51460 96876
rect 53800 96824 53852 96876
rect 84896 96824 84948 96876
rect 88392 96824 88444 96876
rect 127032 96824 127084 96876
rect 128780 96824 128832 96876
rect 185268 96824 185320 96876
rect 190420 96824 190472 96876
rect 22336 96756 22388 96808
rect 38436 96756 38488 96808
rect 41748 96756 41800 96808
rect 108724 96756 108776 96808
rect 112036 96756 112088 96808
rect 175240 96756 175292 96808
rect 176160 96756 176212 96808
rect 180484 96756 180536 96808
rect 182232 96756 182284 96808
rect 182876 96756 182928 96808
rect 187016 96756 187068 96808
rect 84436 96688 84488 96740
rect 88208 96688 88260 96740
rect 109000 96688 109052 96740
rect 112588 96688 112640 96740
rect 181680 96688 181732 96740
rect 185176 96688 185228 96740
rect 175608 96620 175660 96672
rect 176712 96620 176764 96672
rect 83792 96552 83844 96604
rect 88484 96552 88536 96604
rect 180852 96552 180904 96604
rect 184164 96552 184216 96604
rect 50672 96484 50724 96536
rect 58216 96484 58268 96536
rect 82688 96484 82740 96536
rect 89680 96484 89732 96536
rect 109552 96484 109604 96536
rect 113508 96484 113560 96536
rect 182416 96484 182468 96536
rect 184440 96484 184492 96536
rect 39632 96416 39684 96468
rect 43772 96416 43824 96468
rect 53984 96416 54036 96468
rect 77168 96416 77220 96468
rect 79376 96416 79428 96468
rect 88576 96416 88628 96468
rect 109920 96416 109972 96468
rect 113692 96416 113744 96468
rect 113968 96416 114020 96468
rect 119212 96416 119264 96468
rect 125744 96416 125796 96468
rect 148836 96416 148888 96468
rect 151688 96416 151740 96468
rect 160336 96416 160388 96468
rect 23624 96348 23676 96400
rect 26476 96348 26528 96400
rect 110564 96348 110616 96400
rect 114796 96348 114848 96400
rect 25096 96280 25148 96332
rect 28500 96280 28552 96332
rect 40092 96280 40144 96332
rect 44416 96280 44468 96332
rect 110288 96280 110340 96332
rect 114244 96280 114296 96332
rect 156104 96280 156156 96332
rect 160244 96280 160296 96332
rect 39264 96212 39316 96264
rect 43036 96212 43088 96264
rect 111116 96212 111168 96264
rect 115348 96212 115400 96264
rect 157208 96212 157260 96264
rect 160152 96212 160204 96264
rect 35308 96144 35360 96196
rect 36320 96144 36372 96196
rect 111484 96144 111536 96196
rect 116268 96144 116320 96196
rect 111944 96076 111996 96128
rect 116452 96076 116504 96128
rect 184440 96076 184492 96128
rect 189224 96076 189276 96128
rect 102284 96008 102336 96060
rect 103204 96008 103256 96060
rect 112680 96008 112732 96060
rect 117556 96008 117608 96060
rect 100260 95940 100312 95992
rect 100444 95940 100496 95992
rect 101916 95940 101968 95992
rect 102652 95940 102704 95992
rect 103112 95940 103164 95992
rect 104308 95940 104360 95992
rect 113140 95940 113192 95992
rect 118108 95940 118160 95992
rect 159416 95940 159468 95992
rect 161532 95940 161584 95992
rect 183612 95940 183664 95992
rect 188120 95940 188172 95992
rect 101456 95872 101508 95924
rect 102376 95872 102428 95924
rect 102744 95872 102796 95924
rect 103940 95872 103992 95924
rect 112312 95872 112364 95924
rect 117004 95872 117056 95924
rect 178828 95872 178880 95924
rect 180944 95872 180996 95924
rect 183244 95872 183296 95924
rect 187568 95872 187620 95924
rect 26568 95804 26620 95856
rect 29236 95804 29288 95856
rect 101548 95804 101600 95856
rect 104308 95804 104360 95856
rect 105964 95804 106016 95856
rect 106700 95804 106752 95856
rect 109184 95804 109236 95856
rect 113232 95804 113284 95856
rect 118844 95804 118896 95856
rect 179288 95804 179340 95856
rect 179748 95804 179800 95856
rect 100996 95668 101048 95720
rect 164108 94308 164160 94360
rect 168156 94308 168208 94360
rect 91704 94036 91756 94088
rect 95476 94036 95528 94088
rect 91060 92268 91112 92320
rect 118936 92268 118988 92320
rect 91796 91656 91848 91708
rect 95292 91656 95344 91708
rect 188120 91588 188172 91640
rect 198240 91588 198292 91640
rect 91520 91316 91572 91368
rect 93360 91316 93412 91368
rect 163556 91112 163608 91164
rect 165948 91112 166000 91164
rect 188580 90228 188632 90280
rect 197596 90228 197648 90280
rect 18104 90160 18156 90212
rect 22336 90160 22388 90212
rect 163832 90092 163884 90144
rect 166040 90092 166092 90144
rect 92256 88868 92308 88920
rect 95384 88868 95436 88920
rect 163464 88732 163516 88784
rect 165120 88732 165172 88784
rect 92164 87508 92216 87560
rect 95384 87508 95436 87560
rect 188120 84652 188172 84704
rect 196952 84652 197004 84704
rect 163924 84312 163976 84364
rect 167328 84312 167380 84364
rect 116544 83564 116596 83616
rect 119580 83564 119632 83616
rect 163924 82680 163976 82732
rect 167880 82680 167932 82732
rect 13228 82272 13280 82324
rect 15436 82272 15488 82324
rect 13320 81932 13372 81984
rect 22336 81932 22388 81984
rect 163556 81932 163608 81984
rect 167236 81932 167288 81984
rect 91796 80504 91848 80556
rect 94280 80504 94332 80556
rect 164108 80436 164160 80488
rect 167328 80436 167380 80488
rect 164384 78940 164436 78992
rect 167236 78940 167288 78992
rect 91428 78804 91480 78856
rect 95292 78804 95344 78856
rect 164108 77784 164160 77836
rect 167236 77852 167288 77904
rect 91704 77444 91756 77496
rect 95384 77444 95436 77496
rect 163740 76356 163792 76408
rect 167236 76424 167288 76476
rect 91704 76220 91756 76272
rect 94924 76220 94976 76272
rect 15436 74996 15488 75048
rect 22336 74996 22388 75048
rect 45060 74996 45112 75048
rect 47820 74996 47872 75048
rect 164108 74928 164160 74980
rect 167236 74928 167288 74980
rect 164384 73704 164436 73756
rect 167144 73704 167196 73756
rect 91704 72480 91756 72532
rect 95384 72480 95436 72532
rect 164384 72480 164436 72532
rect 167236 72480 167288 72532
rect 91704 71256 91756 71308
rect 95384 71256 95436 71308
rect 164384 71120 164436 71172
rect 167328 71120 167380 71172
rect 163556 69896 163608 69948
rect 167236 69896 167288 69948
rect 91428 69556 91480 69608
rect 94004 69556 94056 69608
rect 91428 68672 91480 68724
rect 93912 68672 93964 68724
rect 163740 68196 163792 68248
rect 167328 68196 167380 68248
rect 189960 67448 190012 67500
rect 190604 67448 190656 67500
rect 197596 67448 197648 67500
rect 91520 66768 91572 66820
rect 93636 66768 93688 66820
rect 164384 66768 164436 66820
rect 167880 66768 167932 66820
rect 44416 65408 44468 65460
rect 47176 65408 47228 65460
rect 164384 65408 164436 65460
rect 167144 65408 167196 65460
rect 164384 64456 164436 64508
rect 167052 64456 167104 64508
rect 92624 64048 92676 64100
rect 93544 64048 93596 64100
rect 164384 64048 164436 64100
rect 166500 64048 166552 64100
rect 117464 62620 117516 62672
rect 119488 62620 119540 62672
rect 13320 62552 13372 62604
rect 22704 62552 22756 62604
rect 91428 61260 91480 61312
rect 93452 61260 93504 61312
rect 92532 59696 92584 59748
rect 94096 59696 94148 59748
rect 91520 58540 91572 58592
rect 93636 58540 93688 58592
rect 164384 58540 164436 58592
rect 166040 58540 166092 58592
rect 92348 58472 92400 58524
rect 95200 58472 95252 58524
rect 187936 57928 187988 57980
rect 189960 57928 190012 57980
rect 164384 57112 164436 57164
rect 165948 57112 166000 57164
rect 82136 51536 82188 51588
rect 84344 51536 84396 51588
rect 145156 51536 145208 51588
rect 173952 51536 174004 51588
rect 174136 51536 174188 51588
rect 175240 51536 175292 51588
rect 176160 51536 176212 51588
rect 98236 51468 98288 51520
rect 98972 51468 99024 51520
rect 103388 51468 103440 51520
rect 103848 51468 103900 51520
rect 105044 51468 105096 51520
rect 106148 51468 106200 51520
rect 106332 51468 106384 51520
rect 107804 51468 107856 51520
rect 111484 51468 111536 51520
rect 112404 51468 112456 51520
rect 113140 51468 113192 51520
rect 114612 51468 114664 51520
rect 174872 51468 174924 51520
rect 175516 51468 175568 51520
rect 72016 51400 72068 51452
rect 73212 51400 73264 51452
rect 83608 51400 83660 51452
rect 84344 51400 84396 51452
rect 66588 51332 66640 51384
rect 82136 51264 82188 51316
rect 105504 51400 105556 51452
rect 106700 51400 106752 51452
rect 107160 51400 107212 51452
rect 108908 51400 108960 51452
rect 110288 51400 110340 51452
rect 111760 51400 111812 51452
rect 112680 51400 112732 51452
rect 114704 51400 114756 51452
rect 105964 51332 106016 51384
rect 107252 51332 107304 51384
rect 106608 51264 106660 51316
rect 108448 51264 108500 51316
rect 138348 51264 138400 51316
rect 40828 50992 40880 51044
rect 42944 50992 42996 51044
rect 109552 50992 109604 51044
rect 111852 50992 111904 51044
rect 112312 50992 112364 51044
rect 114428 50992 114480 51044
rect 64564 50924 64616 50976
rect 86552 50924 86604 50976
rect 13320 50856 13372 50908
rect 72016 50856 72068 50908
rect 138164 50856 138216 50908
rect 151596 50856 151648 50908
rect 36504 50788 36556 50840
rect 38620 50788 38672 50840
rect 104676 50788 104728 50840
rect 105504 50788 105556 50840
rect 36044 50720 36096 50772
rect 37424 50720 37476 50772
rect 175608 50720 175660 50772
rect 176712 50720 176764 50772
rect 182416 50720 182468 50772
rect 184992 50720 185044 50772
rect 35308 50652 35360 50704
rect 36504 50652 36556 50704
rect 180024 50652 180076 50704
rect 182048 50652 182100 50704
rect 39264 50584 39316 50636
rect 41380 50584 41432 50636
rect 178828 50584 178880 50636
rect 180944 50584 180996 50636
rect 184072 50584 184124 50636
rect 186280 50584 186332 50636
rect 38896 50516 38948 50568
rect 40828 50516 40880 50568
rect 179656 50516 179708 50568
rect 182324 50516 182376 50568
rect 183612 50516 183664 50568
rect 188120 50516 188172 50568
rect 38068 50448 38120 50500
rect 39724 50448 39776 50500
rect 111116 50448 111168 50500
rect 112680 50448 112732 50500
rect 177264 50448 177316 50500
rect 179012 50448 179064 50500
rect 181680 50448 181732 50500
rect 183428 50448 183480 50500
rect 184440 50448 184492 50500
rect 186464 50448 186516 50500
rect 37700 50380 37752 50432
rect 40184 50380 40236 50432
rect 41656 50380 41708 50432
rect 44048 50380 44100 50432
rect 109920 50380 109972 50432
rect 27856 50312 27908 50364
rect 30064 50312 30116 50364
rect 36872 50312 36924 50364
rect 20864 50176 20916 50228
rect 26108 50244 26160 50296
rect 26200 50244 26252 50296
rect 26476 50244 26528 50296
rect 25648 50176 25700 50228
rect 28868 50244 28920 50296
rect 29052 50176 29104 50228
rect 30892 50244 30944 50296
rect 36136 50244 36188 50296
rect 37240 50244 37292 50296
rect 37332 50244 37384 50296
rect 22888 50108 22940 50160
rect 27304 50108 27356 50160
rect 40092 50312 40144 50364
rect 44692 50312 44744 50364
rect 108356 50312 108408 50364
rect 110564 50312 110616 50364
rect 39632 50244 39684 50296
rect 39264 50176 39316 50228
rect 40000 50108 40052 50160
rect 27028 50040 27080 50092
rect 29420 50040 29472 50092
rect 30432 50040 30484 50092
rect 31628 50040 31680 50092
rect 40460 50244 40512 50296
rect 41288 50244 41340 50296
rect 107528 50244 107580 50296
rect 46808 50176 46860 50228
rect 93636 50176 93688 50228
rect 94372 50176 94424 50228
rect 97684 50176 97736 50228
rect 98604 50176 98656 50228
rect 108724 50244 108776 50296
rect 176436 50380 176488 50432
rect 177816 50380 177868 50432
rect 178460 50380 178512 50432
rect 180668 50380 180720 50432
rect 182876 50380 182928 50432
rect 184900 50380 184952 50432
rect 185268 50380 185320 50432
rect 187752 50380 187804 50432
rect 176068 50312 176120 50364
rect 177264 50312 177316 50364
rect 177632 50312 177684 50364
rect 179564 50312 179616 50364
rect 180484 50312 180536 50364
rect 109460 50176 109512 50228
rect 111116 50176 111168 50228
rect 111944 50244 111996 50296
rect 112772 50176 112824 50228
rect 113968 50244 114020 50296
rect 115624 50176 115676 50228
rect 176804 50244 176856 50296
rect 118384 50176 118436 50228
rect 165120 50176 165172 50228
rect 167052 50176 167104 50228
rect 169904 50176 169956 50228
rect 170824 50176 170876 50228
rect 171008 50176 171060 50228
rect 171652 50176 171704 50228
rect 179472 50244 179524 50296
rect 181220 50244 181272 50296
rect 178460 50176 178512 50228
rect 181864 50176 181916 50228
rect 45428 50108 45480 50160
rect 93452 50108 93504 50160
rect 95476 50108 95528 50160
rect 97132 50108 97184 50160
rect 98328 50108 98380 50160
rect 98788 50108 98840 50160
rect 99708 50108 99760 50160
rect 107896 50108 107948 50160
rect 110012 50108 110064 50160
rect 110656 50108 110708 50160
rect 113968 50108 114020 50160
rect 163832 50108 163884 50160
rect 167604 50108 167656 50160
rect 168708 50108 168760 50160
rect 170088 50108 170140 50160
rect 178276 50108 178328 50160
rect 180116 50108 180168 50160
rect 184808 50312 184860 50364
rect 189868 50312 189920 50364
rect 183244 50244 183296 50296
rect 183520 50176 183572 50228
rect 185636 50244 185688 50296
rect 187568 50176 187620 50228
rect 184716 50108 184768 50160
rect 184992 50108 185044 50160
rect 186372 50108 186424 50160
rect 43772 50040 43824 50092
rect 93360 50040 93412 50092
rect 96028 50040 96080 50092
rect 109276 50040 109328 50092
rect 111668 50040 111720 50092
rect 169260 50040 169312 50092
rect 170456 50040 170508 50092
rect 184900 50040 184952 50092
rect 187016 50040 187068 50092
rect 24268 49972 24320 50024
rect 28040 49972 28092 50024
rect 28316 49972 28368 50024
rect 30156 49972 30208 50024
rect 31076 49972 31128 50024
rect 32088 49972 32140 50024
rect 40828 49972 40880 50024
rect 42668 49972 42720 50024
rect 42944 49972 42996 50024
rect 46072 49972 46124 50024
rect 112680 49972 112732 50024
rect 114520 49972 114572 50024
rect 181128 49972 181180 50024
rect 184164 49972 184216 50024
rect 190972 49972 191024 50024
rect 23624 49904 23676 49956
rect 27672 49904 27724 49956
rect 29696 49904 29748 49956
rect 31260 49904 31312 49956
rect 41380 49904 41432 49956
rect 43404 49904 43456 49956
rect 183428 49904 183480 49956
rect 185268 49904 185320 49956
rect 187752 49904 187804 49956
rect 190420 49904 190472 49956
rect 38896 49836 38948 49888
rect 42024 49836 42076 49888
rect 182508 49836 182560 49888
rect 185820 49836 185872 49888
rect 44048 49768 44100 49820
rect 47452 49768 47504 49820
rect 112404 49768 112456 49820
rect 115072 49768 115124 49820
rect 186464 49768 186516 49820
rect 189224 49768 189276 49820
rect 26292 49700 26344 49752
rect 29236 49700 29288 49752
rect 163740 49700 163792 49752
rect 168156 49700 168208 49752
rect 24912 49632 24964 49684
rect 28500 49632 28552 49684
rect 39724 49632 39776 49684
rect 41288 49632 41340 49684
rect 186280 49632 186332 49684
rect 188672 49632 188724 49684
rect 113508 49564 113560 49616
rect 117832 49564 117884 49616
rect 20220 49496 20272 49548
rect 44416 49496 44468 49548
rect 114704 49496 114756 49548
rect 116728 49496 116780 49548
rect 168524 49496 168576 49548
rect 191524 49496 191576 49548
rect 111760 49360 111812 49412
rect 113416 49360 113468 49412
rect 91428 49224 91480 49276
rect 92900 49224 92952 49276
rect 96580 49088 96632 49140
rect 97776 49088 97828 49140
rect 114612 49088 114664 49140
rect 117280 49088 117332 49140
rect 21508 48952 21560 49004
rect 26200 48952 26252 49004
rect 114428 48952 114480 49004
rect 116176 48952 116228 49004
rect 182048 48952 182100 49004
rect 182968 48952 183020 49004
rect 22244 48884 22296 48936
rect 26384 48884 26436 48936
rect 103940 47728 103992 47780
rect 104400 47728 104452 47780
rect 50764 46504 50816 46556
rect 61620 46504 61672 46556
rect 122800 46504 122852 46556
rect 129148 46504 129200 46556
rect 51040 46436 51092 46488
rect 63092 46436 63144 46488
rect 122340 46436 122392 46488
rect 127676 46436 127728 46488
rect 51132 46368 51184 46420
rect 60056 46368 60108 46420
rect 122432 46368 122484 46420
rect 130620 46368 130672 46420
rect 148652 46368 148704 46420
rect 158220 46368 158272 46420
rect 50948 46300 51000 46352
rect 58584 46300 58636 46352
rect 76616 46300 76668 46352
rect 87840 46300 87892 46352
rect 122524 46300 122576 46352
rect 132092 46300 132144 46352
rect 150124 46300 150176 46352
rect 159600 46300 159652 46352
rect 50672 46232 50724 46284
rect 55640 46232 55692 46284
rect 81124 46232 81176 46284
rect 87932 46232 87984 46284
rect 126480 46232 126532 46284
rect 136600 46232 136652 46284
rect 151596 46232 151648 46284
rect 159692 46232 159744 46284
rect 50856 46164 50908 46216
rect 57112 46164 57164 46216
rect 78088 46164 78140 46216
rect 86460 46164 86512 46216
rect 122708 46164 122760 46216
rect 133656 46164 133708 46216
rect 54076 46096 54128 46148
rect 67600 46096 67652 46148
rect 79560 46096 79612 46148
rect 85080 46096 85132 46148
rect 122892 46096 122944 46148
rect 135128 46096 135180 46148
rect 153160 46096 153212 46148
rect 158312 46096 158364 46148
rect 121696 44872 121748 44924
rect 123536 44872 123588 44924
rect 121696 44736 121748 44788
rect 123352 44736 123404 44788
rect 154724 44736 154776 44788
rect 156840 44736 156892 44788
rect 84344 44396 84396 44448
rect 85172 44396 85224 44448
rect 159784 43648 159836 43700
rect 160060 43648 160112 43700
rect 121696 43376 121748 43428
rect 124364 43376 124416 43428
rect 121696 42016 121748 42068
rect 124272 42016 124324 42068
rect 121696 40656 121748 40708
rect 124364 40656 124416 40708
rect 14700 40520 14752 40572
rect 18012 40520 18064 40572
rect 156472 39704 156524 39756
rect 156932 39704 156984 39756
rect 122524 39160 122576 39212
rect 122800 39160 122852 39212
rect 159048 38548 159100 38600
rect 160520 38548 160572 38600
rect 121788 38412 121840 38464
rect 123904 38412 123956 38464
rect 121696 38208 121748 38260
rect 123444 38208 123496 38260
rect 121696 37800 121748 37852
rect 124364 37800 124416 37852
rect 88208 37324 88260 37376
rect 88760 37324 88812 37376
rect 121696 35080 121748 35132
rect 123628 35080 123680 35132
rect 121696 33992 121748 34044
rect 124364 33992 124416 34044
rect 121696 33720 121748 33772
rect 124272 33720 124324 33772
rect 121696 32360 121748 32412
rect 123996 32360 124048 32412
rect 121696 31000 121748 31052
rect 124364 31000 124416 31052
rect 121696 28824 121748 28876
rect 123536 28824 123588 28876
rect 121696 28484 121748 28536
rect 124364 28484 124416 28536
rect 121696 28144 121748 28196
rect 124088 28144 124140 28196
rect 159048 28144 159100 28196
rect 160704 28144 160756 28196
rect 88300 27668 88352 27720
rect 88760 27668 88812 27720
rect 158956 25152 159008 25204
rect 160336 25152 160388 25204
rect 50580 24472 50632 24524
rect 50856 24472 50908 24524
rect 121696 24200 121748 24252
rect 123444 24200 123496 24252
rect 51040 24064 51092 24116
rect 51316 24064 51368 24116
rect 159048 22636 159100 22688
rect 160704 22636 160756 22688
rect 85172 22568 85224 22620
rect 88760 22568 88812 22620
rect 156932 22568 156984 22620
rect 160428 22568 160480 22620
rect 156840 22500 156892 22552
rect 160520 22500 160572 22552
rect 85080 21208 85132 21260
rect 88576 21208 88628 21260
rect 158312 21208 158364 21260
rect 160336 21208 160388 21260
rect 86460 19780 86512 19832
rect 88576 19780 88628 19832
rect 158220 19780 158272 19832
rect 160336 19780 160388 19832
rect 13136 19100 13188 19152
rect 66496 19100 66548 19152
rect 18104 18420 18156 18472
rect 62540 18420 62592 18472
rect 69992 18420 70044 18472
rect 73948 18420 74000 18472
rect 119672 18420 119724 18472
rect 50396 18352 50448 18404
rect 63552 18352 63604 18404
rect 94648 18352 94700 18404
rect 95384 18352 95436 18404
rect 100168 18352 100220 18404
rect 134576 18352 134628 18404
rect 55088 18284 55140 18336
rect 75972 18284 76024 18336
rect 81768 18284 81820 18336
rect 83240 18284 83292 18336
rect 143776 18284 143828 18336
rect 144972 18284 145024 18336
rect 145156 18284 145208 18336
rect 145984 18284 146036 18336
rect 39080 18216 39132 18268
rect 66680 18216 66732 18268
rect 71096 18216 71148 18268
rect 72936 18216 72988 18268
rect 82228 18216 82280 18268
rect 84344 18216 84396 18268
rect 49752 18148 49804 18200
rect 77076 18148 77128 18200
rect 80296 18148 80348 18200
rect 84252 18148 84304 18200
rect 44416 18080 44468 18132
rect 78088 18080 78140 18132
rect 33744 18012 33796 18064
rect 28408 17944 28460 17996
rect 65668 18012 65720 18064
rect 145800 18012 145852 18064
rect 149112 18012 149164 18064
rect 17736 17876 17788 17928
rect 67692 17944 67744 17996
rect 124456 17944 124508 17996
rect 140832 17944 140884 17996
rect 23072 17808 23124 17860
rect 68796 17876 68848 17928
rect 119120 17876 119172 17928
rect 141844 17876 141896 17928
rect 12492 17740 12544 17792
rect 70820 17808 70872 17860
rect 113784 17808 113836 17860
rect 142856 17808 142908 17860
rect 69808 17740 69860 17792
rect 81216 17740 81268 17792
rect 92440 17740 92492 17792
rect 108448 17740 108500 17792
rect 143868 17740 143920 17792
rect 146996 17740 147048 17792
rect 154816 17740 154868 17792
rect 60424 17672 60476 17724
rect 74960 17672 75012 17724
rect 71832 17604 71884 17656
rect 79192 17468 79244 17520
rect 80112 17468 80164 17520
rect 148008 17128 148060 17180
rect 150584 17128 150636 17180
rect 61528 17060 61580 17112
rect 105780 17060 105832 17112
rect 117004 17060 117056 17112
rect 126480 17060 126532 17112
rect 133564 17060 133616 17112
rect 187108 17060 187160 17112
rect 95384 16992 95436 17044
rect 135588 16992 135640 17044
rect 168524 16992 168576 17044
rect 154816 12912 154868 12964
rect 156472 12912 156524 12964
rect 84344 12844 84396 12896
rect 87104 12844 87156 12896
rect 156288 12708 156340 12760
rect 172480 12708 172532 12760
rect 145156 12640 145208 12692
rect 161808 12640 161860 12692
rect 155276 12572 155328 12624
rect 177816 12572 177868 12624
rect 143776 12504 143828 12556
rect 167144 12504 167196 12556
rect 154264 12436 154316 12488
rect 183152 12436 183204 12488
rect 153252 12368 153304 12420
rect 188488 12368 188540 12420
rect 79192 12300 79244 12352
rect 97776 12300 97828 12352
rect 135128 12300 135180 12352
rect 138256 12300 138308 12352
rect 140464 12300 140516 12352
rect 150124 12300 150176 12352
rect 152148 12300 152200 12352
rect 193824 12300 193876 12352
rect 78916 12232 78968 12284
rect 103112 12232 103164 12284
rect 129792 12232 129844 12284
rect 139820 12232 139872 12284
rect 151136 12232 151188 12284
rect 199160 12232 199212 12284
rect 76432 12096 76484 12148
rect 80296 12096 80348 12148
rect 150584 12096 150636 12148
rect 151136 12096 151188 12148
rect 65760 11688 65812 11740
rect 69992 11688 70044 11740
<< metal2 >>
rect 25830 220344 25886 220824
rect 57754 220344 57810 220824
rect 89770 220344 89826 220824
rect 121786 220344 121842 220824
rect 153802 220344 153858 220824
rect 185818 220344 185874 220824
rect 22704 213156 22756 213162
rect 22704 213098 22756 213104
rect 22716 210730 22744 213098
rect 25844 211054 25872 220344
rect 57768 220250 57796 220344
rect 57676 220222 57796 220250
rect 33374 213192 33430 213201
rect 33374 213127 33430 213136
rect 39446 213192 39502 213201
rect 39446 213127 39502 213136
rect 56744 213156 56796 213162
rect 25832 211048 25884 211054
rect 25832 210990 25884 210996
rect 22408 210702 22744 210730
rect 33388 210730 33416 213127
rect 39460 210730 39488 213127
rect 56744 213098 56796 213104
rect 56756 211734 56784 213098
rect 56192 211728 56244 211734
rect 56192 211670 56244 211676
rect 56744 211728 56796 211734
rect 56744 211670 56796 211676
rect 33388 210702 33540 210730
rect 39152 210702 39488 210730
rect 28132 210640 28184 210646
rect 27928 210588 28132 210594
rect 27928 210582 28184 210588
rect 27928 210566 28172 210582
rect 49290 210472 49346 210481
rect 47268 210436 47320 210442
rect 49290 210407 49346 210416
rect 47268 210378 47320 210384
rect 13318 210200 13374 210209
rect 13318 210135 13374 210144
rect 13332 209626 13360 210135
rect 13320 209620 13372 209626
rect 13320 209562 13372 209568
rect 14698 188984 14754 188993
rect 14698 188919 14754 188928
rect 13318 167768 13374 167777
rect 13318 167703 13374 167712
rect 13332 167602 13360 167703
rect 13320 167596 13372 167602
rect 13320 167538 13372 167544
rect 13412 155152 13464 155158
rect 13412 155094 13464 155100
rect 13320 146856 13372 146862
rect 13320 146798 13372 146804
rect 13332 125345 13360 146798
rect 13424 146561 13452 155094
rect 13410 146552 13466 146561
rect 13410 146487 13466 146496
rect 13318 125336 13374 125345
rect 13318 125271 13374 125280
rect 13318 104120 13374 104129
rect 13318 104055 13374 104064
rect 13226 82904 13282 82913
rect 13226 82839 13282 82848
rect 13240 82330 13268 82839
rect 13228 82324 13280 82330
rect 13228 82266 13280 82272
rect 13332 81990 13360 104055
rect 13320 81984 13372 81990
rect 13320 81926 13372 81932
rect 13320 62604 13372 62610
rect 13320 62546 13372 62552
rect 13332 61697 13360 62546
rect 13318 61688 13374 61697
rect 13318 61623 13374 61632
rect 13320 50908 13372 50914
rect 13320 50850 13372 50856
rect 13332 40481 13360 50850
rect 14712 40578 14740 188919
rect 47280 183258 47308 210378
rect 49304 204730 49332 210407
rect 49934 209928 49990 209937
rect 49934 209863 49990 209872
rect 49948 208985 49976 209863
rect 51314 209384 51370 209393
rect 51314 209319 51370 209328
rect 49934 208976 49990 208985
rect 49934 208911 49990 208920
rect 51328 208305 51356 209319
rect 56204 208826 56232 211670
rect 57676 210986 57704 220222
rect 89784 216562 89812 220344
rect 80204 216556 80256 216562
rect 80204 216498 80256 216504
rect 89772 216556 89824 216562
rect 89772 216498 89824 216504
rect 66496 213156 66548 213162
rect 66496 213098 66548 213104
rect 57664 210980 57716 210986
rect 57664 210922 57716 210928
rect 59872 210436 59924 210442
rect 59872 210378 59924 210384
rect 56204 208798 56586 208826
rect 59884 208812 59912 210378
rect 66508 208812 66536 213098
rect 76524 211048 76576 211054
rect 76524 210990 76576 210996
rect 69808 210368 69860 210374
rect 69808 210310 69860 210316
rect 73210 210336 73266 210345
rect 69820 208812 69848 210310
rect 73210 210271 73266 210280
rect 73224 208812 73252 210271
rect 76536 208812 76564 210990
rect 80216 208826 80244 216498
rect 83148 216488 83200 216494
rect 83148 216430 83200 216436
rect 79862 208798 80244 208826
rect 83160 208812 83188 216430
rect 115072 213156 115124 213162
rect 115072 213098 115124 213104
rect 96488 211728 96540 211734
rect 96488 211670 96540 211676
rect 96500 210716 96528 211670
rect 115084 210716 115112 213098
rect 121800 211054 121828 220344
rect 153816 216494 153844 220344
rect 185832 216494 185860 220344
rect 153804 216488 153856 216494
rect 153804 216430 153856 216436
rect 155552 216488 155604 216494
rect 155552 216430 155604 216436
rect 185820 216488 185872 216494
rect 185820 216430 185872 216436
rect 128872 211728 128924 211734
rect 128872 211670 128924 211676
rect 121788 211048 121840 211054
rect 121788 210990 121840 210996
rect 105964 210640 106016 210646
rect 105806 210588 105964 210594
rect 105806 210582 106016 210588
rect 105806 210566 106004 210582
rect 120866 210472 120922 210481
rect 128884 210442 128912 211670
rect 151596 211048 151648 211054
rect 151596 210990 151648 210996
rect 148284 210980 148336 210986
rect 148284 210922 148336 210928
rect 138806 210744 138862 210753
rect 138806 210679 138862 210688
rect 120866 210407 120922 210416
rect 128872 210436 128924 210442
rect 88574 209928 88630 209937
rect 88574 209863 88630 209872
rect 88588 209014 88616 209863
rect 88576 209008 88628 209014
rect 88576 208950 88628 208956
rect 88666 208840 88722 208849
rect 88666 208775 88722 208784
rect 51498 208432 51554 208441
rect 51498 208367 51554 208376
rect 51314 208296 51370 208305
rect 51314 208231 51370 208240
rect 51314 208160 51370 208169
rect 51314 208095 51370 208104
rect 51328 207081 51356 208095
rect 51406 207616 51462 207625
rect 51406 207551 51462 207560
rect 51314 207072 51370 207081
rect 51314 207007 51370 207016
rect 51314 206800 51370 206809
rect 51314 206735 51370 206744
rect 51328 205993 51356 206735
rect 51420 206129 51448 207551
rect 51512 207489 51540 208367
rect 88574 208296 88630 208305
rect 88574 208231 88630 208240
rect 51498 207480 51554 207489
rect 51498 207415 51554 207424
rect 88482 207208 88538 207217
rect 88588 207194 88616 208231
rect 88680 207897 88708 208775
rect 88666 207888 88722 207897
rect 88666 207823 88722 207832
rect 88666 207752 88722 207761
rect 88666 207687 88722 207696
rect 88538 207166 88616 207194
rect 88482 207143 88538 207152
rect 88482 206664 88538 206673
rect 88680 206650 88708 207687
rect 88758 207208 88814 207217
rect 88758 207143 88814 207152
rect 88538 206622 88708 206650
rect 88482 206599 88538 206608
rect 51498 206528 51554 206537
rect 51498 206463 51554 206472
rect 51406 206120 51462 206129
rect 51406 206055 51462 206064
rect 51314 205984 51370 205993
rect 51314 205919 51370 205928
rect 51512 205313 51540 206463
rect 88772 206265 88800 207143
rect 88850 206664 88906 206673
rect 88850 206599 88906 206608
rect 88758 206256 88814 206265
rect 88758 206191 88814 206200
rect 87194 205984 87250 205993
rect 87194 205919 87250 205928
rect 51590 205576 51646 205585
rect 51590 205511 51646 205520
rect 51314 205304 51370 205313
rect 51314 205239 51370 205248
rect 51498 205304 51554 205313
rect 51498 205239 51554 205248
rect 49292 204724 49344 204730
rect 49292 204666 49344 204672
rect 50488 204724 50540 204730
rect 50488 204666 50540 204672
rect 50500 202049 50528 204666
rect 51328 204089 51356 205239
rect 51604 204769 51632 205511
rect 87208 204905 87236 205919
rect 88482 205848 88538 205857
rect 88864 205834 88892 206599
rect 88538 205806 88892 205834
rect 88482 205783 88538 205792
rect 87194 204896 87250 204905
rect 88666 204896 88722 204905
rect 87194 204831 87250 204840
rect 88588 204854 88666 204882
rect 51406 204760 51462 204769
rect 51406 204695 51462 204704
rect 51590 204760 51646 204769
rect 51590 204695 51646 204704
rect 51314 204080 51370 204089
rect 51314 204015 51370 204024
rect 51314 203944 51370 203953
rect 51314 203879 51370 203888
rect 51328 203001 51356 203879
rect 51420 203409 51448 204695
rect 51498 203672 51554 203681
rect 51498 203607 51554 203616
rect 88482 203672 88538 203681
rect 88588 203658 88616 204854
rect 88666 204831 88722 204840
rect 88666 204352 88722 204361
rect 88666 204287 88722 204296
rect 88538 203630 88616 203658
rect 88482 203607 88538 203616
rect 51406 203400 51462 203409
rect 51406 203335 51462 203344
rect 51406 203128 51462 203137
rect 51406 203063 51462 203072
rect 51314 202992 51370 203001
rect 51314 202927 51370 202936
rect 51314 202448 51370 202457
rect 51314 202383 51370 202392
rect 50302 202040 50358 202049
rect 50302 201975 50358 201984
rect 50486 202040 50542 202049
rect 50486 201975 50542 201984
rect 50316 192422 50344 201975
rect 51222 201904 51278 201913
rect 51222 201839 51278 201848
rect 51236 200666 51264 201839
rect 51328 201097 51356 202383
rect 51420 201777 51448 203063
rect 51512 201913 51540 203607
rect 88680 203545 88708 204287
rect 88758 203808 88814 203817
rect 88758 203743 88814 203752
rect 88666 203536 88722 203545
rect 88666 203471 88722 203480
rect 88482 202448 88538 202457
rect 88772 202434 88800 203743
rect 88850 203264 88906 203273
rect 88850 203199 88906 203208
rect 88538 202406 88800 202434
rect 88482 202383 88538 202392
rect 88574 202312 88630 202321
rect 88574 202247 88630 202256
rect 84988 202208 85040 202214
rect 84988 202150 85040 202156
rect 85000 202010 85028 202150
rect 84988 202004 85040 202010
rect 84988 201946 85040 201952
rect 51498 201904 51554 201913
rect 51498 201839 51554 201848
rect 51406 201768 51462 201777
rect 51406 201703 51462 201712
rect 88588 201618 88616 202247
rect 88864 202185 88892 203199
rect 88942 202720 88998 202729
rect 88942 202655 88998 202664
rect 88850 202176 88906 202185
rect 88850 202111 88906 202120
rect 88496 201590 88616 201618
rect 51498 201360 51554 201369
rect 51498 201295 51554 201304
rect 87196 201324 87248 201330
rect 51314 201088 51370 201097
rect 51314 201023 51370 201032
rect 51406 200816 51462 200825
rect 51406 200751 51462 200760
rect 51236 200638 51356 200666
rect 51328 200553 51356 200638
rect 51314 200544 51370 200553
rect 51314 200479 51370 200488
rect 51314 200272 51370 200281
rect 51314 200207 51370 200216
rect 51328 198785 51356 200207
rect 51420 199057 51448 200751
rect 51512 200009 51540 201295
rect 87196 201266 87248 201272
rect 87208 201233 87236 201266
rect 87194 201224 87250 201233
rect 87194 201159 87250 201168
rect 88496 200689 88524 201590
rect 88574 201496 88630 201505
rect 88574 201431 88630 201440
rect 88482 200680 88538 200689
rect 88482 200615 88538 200624
rect 88482 200136 88538 200145
rect 88588 200122 88616 201431
rect 88956 201330 88984 202655
rect 120880 202078 120908 210407
rect 128872 210378 128924 210384
rect 122982 209928 123038 209937
rect 123038 209886 123116 209914
rect 122982 209863 123038 209872
rect 122982 209384 123038 209393
rect 122982 209319 123038 209328
rect 122996 208690 123024 209319
rect 123088 208849 123116 209886
rect 123074 208840 123130 208849
rect 123074 208775 123130 208784
rect 128884 208690 128912 210378
rect 138820 208690 138848 210679
rect 141476 210368 141528 210374
rect 141476 210310 141528 210316
rect 145614 210336 145670 210345
rect 141488 208826 141516 210310
rect 145614 210271 145670 210280
rect 141488 208798 141870 208826
rect 145628 208690 145656 210271
rect 148296 208826 148324 210922
rect 151608 208826 151636 210990
rect 148296 208798 148586 208826
rect 151608 208798 151898 208826
rect 155564 208690 155592 216430
rect 160334 210472 160390 210481
rect 160334 210407 160390 210416
rect 192076 210436 192128 210442
rect 160348 210374 160376 210407
rect 192076 210378 192128 210384
rect 156840 210368 156892 210374
rect 156840 210310 156892 210316
rect 160336 210368 160388 210374
rect 160336 210310 160388 210316
rect 122996 208662 123116 208690
rect 128622 208662 128912 208690
rect 138558 208662 138848 208690
rect 145274 208662 145656 208690
rect 155210 208662 155592 208690
rect 123088 208305 123116 208662
rect 123258 208432 123314 208441
rect 123258 208367 123314 208376
rect 123074 208296 123130 208305
rect 123074 208231 123130 208240
rect 122982 208160 123038 208169
rect 123038 208118 123116 208146
rect 122982 208095 123038 208104
rect 123088 207081 123116 208118
rect 123166 207616 123222 207625
rect 123166 207551 123222 207560
rect 123074 207072 123130 207081
rect 123074 207007 123130 207016
rect 122982 206800 123038 206809
rect 123038 206758 123116 206786
rect 122982 206735 123038 206744
rect 122982 206528 123038 206537
rect 122982 206463 123038 206472
rect 122154 205984 122210 205993
rect 122154 205919 122210 205928
rect 122168 205410 122196 205919
rect 122996 205834 123024 206463
rect 123088 205993 123116 206758
rect 123180 206129 123208 207551
rect 123272 207489 123300 208367
rect 123258 207480 123314 207489
rect 123258 207415 123314 207424
rect 123166 206120 123222 206129
rect 123166 206055 123222 206064
rect 123074 205984 123130 205993
rect 123074 205919 123130 205928
rect 122996 205806 123116 205834
rect 122156 205404 122208 205410
rect 122156 205346 122208 205352
rect 123088 205177 123116 205806
rect 124364 205404 124416 205410
rect 124364 205346 124416 205352
rect 123258 205304 123314 205313
rect 123258 205239 123314 205248
rect 123074 205168 123130 205177
rect 123074 205103 123130 205112
rect 122982 204760 123038 204769
rect 123038 204718 123116 204746
rect 122982 204695 123038 204704
rect 122982 204216 123038 204225
rect 122982 204151 123038 204160
rect 122996 203250 123024 204151
rect 123088 203409 123116 204718
rect 123272 204089 123300 205239
rect 124376 204497 124404 205346
rect 124362 204488 124418 204497
rect 124362 204423 124418 204432
rect 123258 204080 123314 204089
rect 123258 204015 123314 204024
rect 123166 203672 123222 203681
rect 123166 203607 123222 203616
rect 123074 203400 123130 203409
rect 123074 203335 123130 203344
rect 122996 203222 123116 203250
rect 123088 203001 123116 203222
rect 123074 202992 123130 203001
rect 123074 202927 123130 202936
rect 122982 202448 123038 202457
rect 123038 202406 123116 202434
rect 122982 202383 123038 202392
rect 120868 202072 120920 202078
rect 120868 202014 120920 202020
rect 122432 202072 122484 202078
rect 122432 202014 122484 202020
rect 88944 201324 88996 201330
rect 88944 201266 88996 201272
rect 88666 200952 88722 200961
rect 88666 200887 88722 200896
rect 88538 200094 88616 200122
rect 88482 200071 88538 200080
rect 51498 200000 51554 200009
rect 51498 199935 51554 199944
rect 51498 199592 51554 199601
rect 51498 199527 51554 199536
rect 51406 199048 51462 199057
rect 51406 198983 51462 198992
rect 51406 198912 51462 198921
rect 51406 198847 51462 198856
rect 51314 198776 51370 198785
rect 51314 198711 51370 198720
rect 51314 198504 51370 198513
rect 51314 198439 51370 198448
rect 51328 196473 51356 198439
rect 51420 197561 51448 198847
rect 51512 197697 51540 199527
rect 88482 199456 88538 199465
rect 88680 199442 88708 200887
rect 88758 200408 88814 200417
rect 88758 200343 88814 200352
rect 88538 199414 88708 199442
rect 88482 199391 88538 199400
rect 87196 199352 87248 199358
rect 88772 199329 88800 200343
rect 88850 199864 88906 199873
rect 88850 199799 88906 199808
rect 87196 199294 87248 199300
rect 88758 199320 88814 199329
rect 51590 197960 51646 197969
rect 51590 197895 51646 197904
rect 51498 197688 51554 197697
rect 51498 197623 51554 197632
rect 51406 197552 51462 197561
rect 51406 197487 51462 197496
rect 51498 197416 51554 197425
rect 51498 197351 51554 197360
rect 51406 196736 51462 196745
rect 51406 196671 51462 196680
rect 51314 196464 51370 196473
rect 51314 196399 51370 196408
rect 51314 196192 51370 196201
rect 51314 196127 51370 196136
rect 51328 194569 51356 196127
rect 51420 195113 51448 196671
rect 51512 195793 51540 197351
rect 51604 196337 51632 197895
rect 87208 197697 87236 199294
rect 88758 199255 88814 199264
rect 88864 198354 88892 199799
rect 88944 199352 88996 199358
rect 88942 199320 88944 199329
rect 88996 199320 88998 199329
rect 88942 199255 88998 199264
rect 88942 198776 88998 198785
rect 88942 198711 88998 198720
rect 88496 198326 88892 198354
rect 88496 198241 88524 198326
rect 88482 198232 88538 198241
rect 88666 198232 88722 198241
rect 88482 198167 88538 198176
rect 88588 198190 88666 198218
rect 88588 197946 88616 198190
rect 88666 198167 88722 198176
rect 88496 197918 88616 197946
rect 87194 197688 87250 197697
rect 87194 197623 87250 197632
rect 87196 197584 87248 197590
rect 87196 197526 87248 197532
rect 87208 197153 87236 197526
rect 87194 197144 87250 197153
rect 87194 197079 87250 197088
rect 88496 196473 88524 197918
rect 88574 197688 88630 197697
rect 88574 197623 88630 197632
rect 88482 196464 88538 196473
rect 88482 196399 88538 196408
rect 51590 196328 51646 196337
rect 51590 196263 51646 196272
rect 88482 196328 88538 196337
rect 88588 196314 88616 197623
rect 88956 197590 88984 198711
rect 88944 197584 88996 197590
rect 88944 197526 88996 197532
rect 88666 197144 88722 197153
rect 88666 197079 88722 197088
rect 88538 196286 88616 196314
rect 88482 196263 88538 196272
rect 88680 196042 88708 197079
rect 121786 196736 121842 196745
rect 121786 196671 121842 196680
rect 121800 196570 121828 196671
rect 121788 196564 121840 196570
rect 121788 196506 121840 196512
rect 89218 196464 89274 196473
rect 89218 196399 89274 196408
rect 88496 196014 88708 196042
rect 88496 195793 88524 196014
rect 88574 195920 88630 195929
rect 88574 195855 88630 195864
rect 51498 195784 51554 195793
rect 51498 195719 51554 195728
rect 88482 195784 88538 195793
rect 88482 195719 88538 195728
rect 51498 195648 51554 195657
rect 51498 195583 51554 195592
rect 51406 195104 51462 195113
rect 51406 195039 51462 195048
rect 51406 194832 51462 194841
rect 51406 194767 51462 194776
rect 51314 194560 51370 194569
rect 51314 194495 51370 194504
rect 51314 193880 51370 193889
rect 51314 193815 51370 193824
rect 51328 193186 51356 193815
rect 51420 193345 51448 194767
rect 51512 193753 51540 195583
rect 88390 195376 88446 195385
rect 88390 195311 88446 195320
rect 88298 194288 88354 194297
rect 88298 194223 88354 194232
rect 51590 194152 51646 194161
rect 51590 194087 51646 194096
rect 51498 193744 51554 193753
rect 51498 193679 51554 193688
rect 51406 193336 51462 193345
rect 51406 193271 51462 193280
rect 51328 193158 51448 193186
rect 51314 193064 51370 193073
rect 51314 192999 51370 193008
rect 50500 192422 50528 192453
rect 50304 192416 50356 192422
rect 50488 192416 50540 192422
rect 50304 192358 50356 192364
rect 50408 192364 50488 192370
rect 50408 192358 50540 192364
rect 50408 192342 50528 192358
rect 49934 185992 49990 186001
rect 49934 185927 49990 185936
rect 49948 185554 49976 185927
rect 49936 185548 49988 185554
rect 49936 185490 49988 185496
rect 50210 185312 50266 185321
rect 50210 185247 50266 185256
rect 50118 184768 50174 184777
rect 50118 184703 50174 184712
rect 50026 184224 50082 184233
rect 50026 184159 50082 184168
rect 47156 183230 47308 183258
rect 49934 183136 49990 183145
rect 49934 183071 49990 183080
rect 19924 182822 20260 182850
rect 20568 182822 20904 182850
rect 21212 182822 21548 182850
rect 21856 182822 22192 182850
rect 22500 182822 22836 182850
rect 23144 182822 23480 182850
rect 23788 182822 24124 182850
rect 24432 182822 24768 182850
rect 25076 182822 25412 182850
rect 25720 182822 26056 182850
rect 26364 182822 26424 182850
rect 27008 182822 27344 182850
rect 27652 182822 27804 182850
rect 28296 182822 28632 182850
rect 28940 182822 29184 182850
rect 29676 182822 30012 182850
rect 30320 182822 30564 182850
rect 30964 182822 31300 182850
rect 31608 182822 31944 182850
rect 20232 180561 20260 182822
rect 20876 181338 20904 182822
rect 20864 181332 20916 181338
rect 20864 181274 20916 181280
rect 20218 180552 20274 180561
rect 20218 180487 20274 180496
rect 21520 180114 21548 182822
rect 21508 180108 21560 180114
rect 21508 180050 21560 180056
rect 22164 180046 22192 182822
rect 22808 180318 22836 182822
rect 22796 180312 22848 180318
rect 22796 180254 22848 180260
rect 23452 180250 23480 182822
rect 23440 180244 23492 180250
rect 23440 180186 23492 180192
rect 24096 180182 24124 182822
rect 24740 180454 24768 182822
rect 24728 180448 24780 180454
rect 24728 180390 24780 180396
rect 25384 180386 25412 182822
rect 25372 180380 25424 180386
rect 25372 180322 25424 180328
rect 26028 180250 26056 182822
rect 26108 181332 26160 181338
rect 26108 181274 26160 181280
rect 25372 180244 25424 180250
rect 25372 180186 25424 180192
rect 26016 180244 26068 180250
rect 26016 180186 26068 180192
rect 24084 180176 24136 180182
rect 24084 180118 24136 180124
rect 22152 180040 22204 180046
rect 22152 179982 22204 179988
rect 25384 178482 25412 180186
rect 25372 178476 25424 178482
rect 25372 178418 25424 178424
rect 26120 175764 26148 181274
rect 26396 180590 26424 182822
rect 27316 180930 27344 182822
rect 27776 181270 27804 182822
rect 27764 181264 27816 181270
rect 27764 181206 27816 181212
rect 28604 181066 28632 182822
rect 28592 181060 28644 181066
rect 28592 181002 28644 181008
rect 27304 180924 27356 180930
rect 27304 180866 27356 180872
rect 26384 180584 26436 180590
rect 26384 180526 26436 180532
rect 27856 180584 27908 180590
rect 27856 180526 27908 180532
rect 26568 180448 26620 180454
rect 26568 180390 26620 180396
rect 26384 180312 26436 180318
rect 26384 180254 26436 180260
rect 26396 178210 26424 180254
rect 26476 180108 26528 180114
rect 26476 180050 26528 180056
rect 26384 178204 26436 178210
rect 26384 178146 26436 178152
rect 26488 175764 26516 180050
rect 26580 177462 26608 180390
rect 27764 180176 27816 180182
rect 27764 180118 27816 180124
rect 26844 180040 26896 180046
rect 26844 179982 26896 179988
rect 26568 177456 26620 177462
rect 26568 177398 26620 177404
rect 26856 175764 26884 179982
rect 27672 178476 27724 178482
rect 27672 178418 27724 178424
rect 27304 178204 27356 178210
rect 27304 178146 27356 178152
rect 27316 175764 27344 178146
rect 27684 175764 27712 178418
rect 27776 177274 27804 180118
rect 27868 177734 27896 180526
rect 28868 180380 28920 180386
rect 28868 180322 28920 180328
rect 27948 180244 28000 180250
rect 27948 180186 28000 180192
rect 27856 177728 27908 177734
rect 27856 177670 27908 177676
rect 27960 177666 27988 180186
rect 27948 177660 28000 177666
rect 27948 177602 28000 177608
rect 28500 177456 28552 177462
rect 28500 177398 28552 177404
rect 27776 177246 27896 177274
rect 27868 175778 27896 177246
rect 27868 175750 28066 175778
rect 28512 175764 28540 177398
rect 28880 175764 28908 180322
rect 29156 180250 29184 182822
rect 29984 181338 30012 182822
rect 29972 181332 30024 181338
rect 29972 181274 30024 181280
rect 30432 181264 30484 181270
rect 30432 181206 30484 181212
rect 30064 180924 30116 180930
rect 30064 180866 30116 180872
rect 29144 180244 29196 180250
rect 29144 180186 29196 180192
rect 29696 177728 29748 177734
rect 29696 177670 29748 177676
rect 29236 177660 29288 177666
rect 29236 177602 29288 177608
rect 29248 175764 29276 177602
rect 29708 175764 29736 177670
rect 30076 175764 30104 180866
rect 30444 175764 30472 181206
rect 30536 180522 30564 182822
rect 30892 181060 30944 181066
rect 30892 181002 30944 181008
rect 30524 180516 30576 180522
rect 30524 180458 30576 180464
rect 30904 175764 30932 181002
rect 31272 180386 31300 182822
rect 31916 181338 31944 182822
rect 32008 182822 32252 182850
rect 32896 182822 33232 182850
rect 31352 181332 31404 181338
rect 31352 181274 31404 181280
rect 31904 181332 31956 181338
rect 31904 181274 31956 181280
rect 31260 180380 31312 180386
rect 31260 180322 31312 180328
rect 31260 180244 31312 180250
rect 31260 180186 31312 180192
rect 31272 175764 31300 180186
rect 31364 175778 31392 181274
rect 32008 177326 32036 182822
rect 33204 181338 33232 182822
rect 33388 182822 33540 182850
rect 34184 182822 34244 182850
rect 34828 182822 34888 182850
rect 35472 182822 35532 182850
rect 36116 182822 36176 182850
rect 32824 181332 32876 181338
rect 32824 181274 32876 181280
rect 33192 181332 33244 181338
rect 33192 181274 33244 181280
rect 32088 180516 32140 180522
rect 32088 180458 32140 180464
rect 31996 177320 32048 177326
rect 31996 177262 32048 177268
rect 31364 175750 31654 175778
rect 32100 175764 32128 180458
rect 32456 180380 32508 180386
rect 32456 180322 32508 180328
rect 32468 175764 32496 180322
rect 32836 175764 32864 181274
rect 33388 177666 33416 182822
rect 33652 181332 33704 181338
rect 33652 181274 33704 181280
rect 33376 177660 33428 177666
rect 33376 177602 33428 177608
rect 33284 177320 33336 177326
rect 33284 177262 33336 177268
rect 33296 175764 33324 177262
rect 33664 175764 33692 181274
rect 34112 177660 34164 177666
rect 34112 177602 34164 177608
rect 34124 175764 34152 177602
rect 34216 175778 34244 182822
rect 34216 175750 34506 175778
rect 34860 175764 34888 182822
rect 35504 175778 35532 182822
rect 36148 179994 36176 182822
rect 35964 179966 36176 179994
rect 36240 182822 36760 182850
rect 36884 182822 37404 182850
rect 37712 182822 38048 182850
rect 38448 182822 38784 182850
rect 39092 182822 39428 182850
rect 39736 182822 40072 182850
rect 40380 182822 40716 182850
rect 41024 182822 41360 182850
rect 41760 182822 42004 182850
rect 42312 182822 42648 182850
rect 43048 182822 43292 182850
rect 43600 182822 43936 182850
rect 44428 182822 44580 182850
rect 44888 182822 45224 182850
rect 45808 182822 45868 182850
rect 36240 179978 36268 182822
rect 36884 181490 36912 182822
rect 36332 181462 36912 181490
rect 36228 179972 36280 179978
rect 35964 175778 35992 179966
rect 36228 179914 36280 179920
rect 36044 179904 36096 179910
rect 36044 179846 36096 179852
rect 35334 175750 35532 175778
rect 35702 175750 35992 175778
rect 36056 175764 36084 179846
rect 36332 175778 36360 181462
rect 37712 181338 37740 182822
rect 36872 181332 36924 181338
rect 36872 181274 36924 181280
rect 37700 181332 37752 181338
rect 37700 181274 37752 181280
rect 36332 175750 36530 175778
rect 36884 175764 36912 181274
rect 38448 181270 38476 182822
rect 38896 181332 38948 181338
rect 38896 181274 38948 181280
rect 37424 181264 37476 181270
rect 37424 181206 37476 181212
rect 38436 181264 38488 181270
rect 38436 181206 38488 181212
rect 37436 175778 37464 181206
rect 37700 181196 37752 181202
rect 37700 181138 37752 181144
rect 37266 175750 37464 175778
rect 37712 175764 37740 181138
rect 38436 181128 38488 181134
rect 38436 181070 38488 181076
rect 38068 180108 38120 180114
rect 38068 180050 38120 180056
rect 38080 175764 38108 180050
rect 38448 175764 38476 181070
rect 38908 175764 38936 181274
rect 39092 181202 39120 182822
rect 39080 181196 39132 181202
rect 39080 181138 39132 181144
rect 39632 180924 39684 180930
rect 39632 180866 39684 180872
rect 39264 180652 39316 180658
rect 39264 180594 39316 180600
rect 39276 175764 39304 180594
rect 39644 175764 39672 180866
rect 39736 180114 39764 182822
rect 40380 181134 40408 182822
rect 41024 181338 41052 182822
rect 41012 181332 41064 181338
rect 41012 181274 41064 181280
rect 40460 181196 40512 181202
rect 40460 181138 40512 181144
rect 40368 181128 40420 181134
rect 40368 181070 40420 181076
rect 40092 181060 40144 181066
rect 40092 181002 40144 181008
rect 39724 180108 39776 180114
rect 39724 180050 39776 180056
rect 40104 175764 40132 181002
rect 40472 175764 40500 181138
rect 41760 180658 41788 182822
rect 42312 180930 42340 182822
rect 43048 181066 43076 182822
rect 43600 181202 43628 182822
rect 43588 181196 43640 181202
rect 43588 181138 43640 181144
rect 43036 181060 43088 181066
rect 43036 181002 43088 181008
rect 42300 180924 42352 180930
rect 42300 180866 42352 180872
rect 41748 180652 41800 180658
rect 41748 180594 41800 180600
rect 41656 177796 41708 177802
rect 41656 177738 41708 177744
rect 41288 177660 41340 177666
rect 41288 177602 41340 177608
rect 40828 177388 40880 177394
rect 40828 177330 40880 177336
rect 40840 175764 40868 177330
rect 41300 175764 41328 177602
rect 41668 175764 41696 177738
rect 44428 177394 44456 182822
rect 44888 177666 44916 182822
rect 45808 177802 45836 182822
rect 45796 177796 45848 177802
rect 45796 177738 45848 177744
rect 44876 177660 44928 177666
rect 44876 177602 44928 177608
rect 44416 177388 44468 177394
rect 44416 177330 44468 177336
rect 49948 175642 49976 183071
rect 50040 177666 50068 184159
rect 50132 177734 50160 184703
rect 50120 177728 50172 177734
rect 50120 177670 50172 177676
rect 50028 177660 50080 177666
rect 50028 177602 50080 177608
rect 50224 177530 50252 185247
rect 50408 182630 50436 192342
rect 51328 191577 51356 192999
rect 51420 192121 51448 193158
rect 51498 192792 51554 192801
rect 51498 192727 51554 192736
rect 51406 192112 51462 192121
rect 51406 192047 51462 192056
rect 51406 191704 51462 191713
rect 51406 191639 51462 191648
rect 51314 191568 51370 191577
rect 51314 191503 51370 191512
rect 51314 190480 51370 190489
rect 51314 190415 51370 190424
rect 51328 188177 51356 190415
rect 51420 189265 51448 191639
rect 51512 190897 51540 192727
rect 51604 192393 51632 194087
rect 84528 192416 84580 192422
rect 51590 192384 51646 192393
rect 84528 192358 84580 192364
rect 51590 192319 51646 192328
rect 51682 192248 51738 192257
rect 51682 192183 51738 192192
rect 51590 191024 51646 191033
rect 51590 190959 51646 190968
rect 51498 190888 51554 190897
rect 51498 190823 51554 190832
rect 51498 189936 51554 189945
rect 51498 189871 51554 189880
rect 51406 189256 51462 189265
rect 51406 189191 51462 189200
rect 51406 189120 51462 189129
rect 51406 189055 51462 189064
rect 51314 188168 51370 188177
rect 51314 188103 51370 188112
rect 51314 187896 51370 187905
rect 51314 187831 51370 187840
rect 50670 187080 50726 187089
rect 50670 187015 50726 187024
rect 50396 182624 50448 182630
rect 50396 182566 50448 182572
rect 50684 177870 50712 187015
rect 51328 186137 51356 187831
rect 51420 187361 51448 189055
rect 51512 188041 51540 189871
rect 51604 189129 51632 190959
rect 51696 190353 51724 192183
rect 51682 190344 51738 190353
rect 51682 190279 51738 190288
rect 51590 189120 51646 189129
rect 51590 189055 51646 189064
rect 51590 188848 51646 188857
rect 51590 188783 51646 188792
rect 51498 188032 51554 188041
rect 51498 187967 51554 187976
rect 51498 187624 51554 187633
rect 51498 187559 51554 187568
rect 51406 187352 51462 187361
rect 51406 187287 51462 187296
rect 51314 186128 51370 186137
rect 51314 186063 51370 186072
rect 51512 185457 51540 187559
rect 51604 186817 51632 188783
rect 51590 186808 51646 186817
rect 51590 186743 51646 186752
rect 51958 186536 52014 186545
rect 51958 186471 52014 186480
rect 51498 185448 51554 185457
rect 51498 185383 51554 185392
rect 51314 183680 51370 183689
rect 51314 183615 51370 183624
rect 50672 177864 50724 177870
rect 50672 177806 50724 177812
rect 50212 177524 50264 177530
rect 50212 177466 50264 177472
rect 51328 175778 51356 183615
rect 51972 177394 52000 186471
rect 52052 185548 52104 185554
rect 52052 185490 52104 185496
rect 52064 178346 52092 185490
rect 84540 185350 84568 192358
rect 88312 192257 88340 194223
rect 88404 193481 88432 195311
rect 88482 194152 88538 194161
rect 88588 194138 88616 195855
rect 89232 195249 89260 196399
rect 89218 195240 89274 195249
rect 89218 195175 89274 195184
rect 88666 194832 88722 194841
rect 88666 194767 88722 194776
rect 88538 194110 88616 194138
rect 88482 194087 88538 194096
rect 88390 193472 88446 193481
rect 88390 193407 88446 193416
rect 88680 193050 88708 194767
rect 122246 194560 122302 194569
rect 122246 194495 122302 194504
rect 122260 194190 122288 194495
rect 122248 194184 122300 194190
rect 122248 194126 122300 194132
rect 88758 193744 88814 193753
rect 88758 193679 88814 193688
rect 88496 193022 88708 193050
rect 88496 192937 88524 193022
rect 88482 192928 88538 192937
rect 88482 192863 88538 192872
rect 88390 192656 88446 192665
rect 88390 192591 88446 192600
rect 88298 192248 88354 192257
rect 88298 192183 88354 192192
rect 87196 192144 87248 192150
rect 87196 192086 87248 192092
rect 87208 191169 87236 192086
rect 88298 191432 88354 191441
rect 88298 191367 88354 191376
rect 87194 191160 87250 191169
rect 87194 191095 87250 191104
rect 88206 189800 88262 189809
rect 88206 189735 88262 189744
rect 87196 188268 87248 188274
rect 87196 188210 87248 188216
rect 87104 186908 87156 186914
rect 87104 186850 87156 186856
rect 87012 185956 87064 185962
rect 87012 185898 87064 185904
rect 85724 185684 85776 185690
rect 85724 185626 85776 185632
rect 84528 185344 84580 185350
rect 84528 185286 84580 185292
rect 84252 185276 84304 185282
rect 84252 185218 84304 185224
rect 84264 185162 84292 185218
rect 84094 185134 84292 185162
rect 82226 185040 82282 185049
rect 82282 184998 82622 185026
rect 82226 184975 82282 184984
rect 55468 184862 55574 184890
rect 58320 184862 58426 184890
rect 59608 184862 59806 184890
rect 60988 184862 61278 184890
rect 55468 182698 55496 184862
rect 55456 182692 55508 182698
rect 55456 182634 55508 182640
rect 52052 178340 52104 178346
rect 52052 178282 52104 178288
rect 56008 178340 56060 178346
rect 56008 178282 56060 178288
rect 53800 177728 53852 177734
rect 53800 177670 53852 177676
rect 52696 177660 52748 177666
rect 52696 177602 52748 177608
rect 51960 177388 52012 177394
rect 51960 177330 52012 177336
rect 51328 175750 51618 175778
rect 52708 175764 52736 177602
rect 53812 175764 53840 177670
rect 54904 177524 54956 177530
rect 54904 177466 54956 177472
rect 54916 175764 54944 177466
rect 56020 175764 56048 178282
rect 58320 177870 58348 184862
rect 59608 182442 59636 184862
rect 60988 182442 61016 184862
rect 59516 182414 59636 182442
rect 60896 182414 61016 182442
rect 58216 177864 58268 177870
rect 58216 177806 58268 177812
rect 58308 177864 58360 177870
rect 58308 177806 58360 177812
rect 57112 177388 57164 177394
rect 57112 177330 57164 177336
rect 57124 175764 57152 177330
rect 58228 175764 58256 177806
rect 59516 175778 59544 182414
rect 60896 175778 60924 182414
rect 62644 181950 62672 184876
rect 61528 181944 61580 181950
rect 61528 181886 61580 181892
rect 62632 181944 62684 181950
rect 62632 181886 62684 181892
rect 59346 175750 59544 175778
rect 60450 175750 60924 175778
rect 61540 175764 61568 181886
rect 64116 181814 64144 184876
rect 62632 181808 62684 181814
rect 62632 181750 62684 181756
rect 64104 181808 64156 181814
rect 64104 181750 64156 181756
rect 62644 175764 62672 181750
rect 64932 181468 64984 181474
rect 64932 181410 64984 181416
rect 63828 181400 63880 181406
rect 63828 181342 63880 181348
rect 63840 175764 63868 181342
rect 64944 175764 64972 181410
rect 65496 181406 65524 184876
rect 66036 182420 66088 182426
rect 66036 182362 66088 182368
rect 65484 181400 65536 181406
rect 65484 181342 65536 181348
rect 66048 175764 66076 182362
rect 66968 181474 66996 184876
rect 67140 182488 67192 182494
rect 67140 182430 67192 182436
rect 66956 181468 67008 181474
rect 66956 181410 67008 181416
rect 67152 175764 67180 182430
rect 68348 182426 68376 184876
rect 69820 182494 69848 184876
rect 69808 182488 69860 182494
rect 69808 182430 69860 182436
rect 70452 182488 70504 182494
rect 70452 182430 70504 182436
rect 68336 182420 68388 182426
rect 68336 182362 68388 182368
rect 69348 182420 69400 182426
rect 69348 182362 69400 182368
rect 68244 182352 68296 182358
rect 68244 182294 68296 182300
rect 68256 175764 68284 182294
rect 69360 175764 69388 182362
rect 70464 175764 70492 182430
rect 71200 182358 71228 184876
rect 72672 182426 72700 184876
rect 74052 182494 74080 184876
rect 74040 182488 74092 182494
rect 74040 182430 74092 182436
rect 72660 182420 72712 182426
rect 72660 182362 72712 182368
rect 71188 182352 71240 182358
rect 71188 182294 71240 182300
rect 73764 182080 73816 182086
rect 73764 182022 73816 182028
rect 72660 181468 72712 181474
rect 72660 181410 72712 181416
rect 71556 181400 71608 181406
rect 71556 181342 71608 181348
rect 71568 175764 71596 181342
rect 72672 175764 72700 181410
rect 73776 175764 73804 182022
rect 74868 181808 74920 181814
rect 74868 181750 74920 181756
rect 74880 175764 74908 181750
rect 75524 181406 75552 184876
rect 76904 181474 76932 184876
rect 78376 182086 78404 184876
rect 78364 182080 78416 182086
rect 78364 182022 78416 182028
rect 79756 181814 79784 184876
rect 80308 184862 81242 184890
rect 79744 181808 79796 181814
rect 79744 181750 79796 181756
rect 76892 181468 76944 181474
rect 76892 181410 76944 181416
rect 75512 181400 75564 181406
rect 75512 181342 75564 181348
rect 80308 177666 80336 184862
rect 85172 184120 85224 184126
rect 85172 184062 85224 184068
rect 85184 178482 85212 184062
rect 81584 178476 81636 178482
rect 81584 178418 81636 178424
rect 85172 178476 85224 178482
rect 85172 178418 85224 178424
rect 80480 178068 80532 178074
rect 80480 178010 80532 178016
rect 75972 177660 76024 177666
rect 75972 177602 76024 177608
rect 80296 177660 80348 177666
rect 80296 177602 80348 177608
rect 75984 175764 76012 177602
rect 79376 177456 79428 177462
rect 79376 177398 79428 177404
rect 77166 177288 77222 177297
rect 77166 177223 77222 177232
rect 77180 175764 77208 177223
rect 79388 175764 79416 177398
rect 80492 175764 80520 178010
rect 81596 175764 81624 178418
rect 83792 178204 83844 178210
rect 83792 178146 83844 178152
rect 82688 178000 82740 178006
rect 82688 177942 82740 177948
rect 82700 175764 82728 177942
rect 83804 175764 83832 178146
rect 85736 177666 85764 185626
rect 86460 184188 86512 184194
rect 86460 184130 86512 184136
rect 86472 178210 86500 184130
rect 86552 182760 86604 182766
rect 86552 182702 86604 182708
rect 86460 178204 86512 178210
rect 86460 178146 86512 178152
rect 84896 177660 84948 177666
rect 84896 177602 84948 177608
rect 85724 177660 85776 177666
rect 85724 177602 85776 177608
rect 84908 175764 84936 177602
rect 86000 177524 86052 177530
rect 86000 177466 86052 177472
rect 86012 175764 86040 177466
rect 86564 177462 86592 182702
rect 87024 177530 87052 185898
rect 87012 177524 87064 177530
rect 87012 177466 87064 177472
rect 86552 177456 86604 177462
rect 86552 177398 86604 177404
rect 87116 175764 87144 186850
rect 87208 186273 87236 188210
rect 88220 187497 88248 189735
rect 88312 189265 88340 191367
rect 88404 190489 88432 192591
rect 88772 192098 88800 193679
rect 88850 193200 88906 193209
rect 88850 193135 88906 193144
rect 88864 192150 88892 193135
rect 122444 193050 122472 202014
rect 122982 201904 123038 201913
rect 122982 201839 123038 201848
rect 122996 200938 123024 201839
rect 123088 201097 123116 202406
rect 123180 201913 123208 203607
rect 123258 203128 123314 203137
rect 123258 203063 123314 203072
rect 123166 201904 123222 201913
rect 123166 201839 123222 201848
rect 123272 201777 123300 203063
rect 123258 201768 123314 201777
rect 123258 201703 123314 201712
rect 123166 201360 123222 201369
rect 123166 201295 123222 201304
rect 123074 201088 123130 201097
rect 123074 201023 123130 201032
rect 122996 200910 123116 200938
rect 122982 200816 123038 200825
rect 122982 200751 123038 200760
rect 122996 200394 123024 200751
rect 123088 200553 123116 200910
rect 123074 200544 123130 200553
rect 123074 200479 123130 200488
rect 122996 200366 123116 200394
rect 122982 199592 123038 199601
rect 122982 199527 123038 199536
rect 122996 199034 123024 199527
rect 123088 199193 123116 200366
rect 123180 200009 123208 201295
rect 123166 200000 123222 200009
rect 123166 199935 123222 199944
rect 123166 199864 123222 199873
rect 123166 199799 123222 199808
rect 123074 199184 123130 199193
rect 123074 199119 123130 199128
rect 122996 199006 123116 199034
rect 122982 198776 123038 198785
rect 122982 198711 123038 198720
rect 122996 197674 123024 198711
rect 123088 197833 123116 199006
rect 123180 198785 123208 199799
rect 123166 198776 123222 198785
rect 123166 198711 123222 198720
rect 123166 198504 123222 198513
rect 123166 198439 123222 198448
rect 123074 197824 123130 197833
rect 123074 197759 123130 197768
rect 122996 197646 123116 197674
rect 123088 197561 123116 197646
rect 123074 197552 123130 197561
rect 123074 197487 123130 197496
rect 122982 197416 123038 197425
rect 123038 197374 123116 197402
rect 122982 197351 123038 197360
rect 123088 196314 123116 197374
rect 123180 196473 123208 198439
rect 123258 197960 123314 197969
rect 123258 197895 123314 197904
rect 123166 196464 123222 196473
rect 123166 196399 123222 196408
rect 123272 196337 123300 197895
rect 124180 196564 124232 196570
rect 124180 196506 124232 196512
rect 123258 196328 123314 196337
rect 123088 196286 123208 196314
rect 123074 196192 123130 196201
rect 123074 196127 123130 196136
rect 122982 195104 123038 195113
rect 122982 195039 123038 195048
rect 122996 194410 123024 195039
rect 123088 194569 123116 196127
rect 123180 195793 123208 196286
rect 123258 196263 123314 196272
rect 123166 195784 123222 195793
rect 123166 195719 123222 195728
rect 123166 195648 123222 195657
rect 123166 195583 123222 195592
rect 123074 194560 123130 194569
rect 123074 194495 123130 194504
rect 122996 194382 123116 194410
rect 123088 193345 123116 194382
rect 123180 193753 123208 195583
rect 124192 194977 124220 196506
rect 124178 194968 124234 194977
rect 124178 194903 124234 194912
rect 123352 194184 123404 194190
rect 123352 194126 123404 194132
rect 123258 193880 123314 193889
rect 123258 193815 123314 193824
rect 123166 193744 123222 193753
rect 123166 193679 123222 193688
rect 123074 193336 123130 193345
rect 123074 193271 123130 193280
rect 122982 193064 123038 193073
rect 122444 193022 122564 193050
rect 122536 192354 122564 193022
rect 123038 193022 123116 193050
rect 122982 192999 123038 193008
rect 122524 192348 122576 192354
rect 122524 192290 122576 192296
rect 88496 192070 88800 192098
rect 88852 192144 88904 192150
rect 88852 192086 88904 192092
rect 88496 191713 88524 192070
rect 88574 191976 88630 191985
rect 88574 191911 88630 191920
rect 88482 191704 88538 191713
rect 88482 191639 88538 191648
rect 88390 190480 88446 190489
rect 88390 190415 88446 190424
rect 88390 190344 88446 190353
rect 88390 190279 88446 190288
rect 88298 189256 88354 189265
rect 88298 189191 88354 189200
rect 88404 188177 88432 190279
rect 88482 189936 88538 189945
rect 88588 189922 88616 191911
rect 122154 191704 122210 191713
rect 122154 191639 122210 191648
rect 122168 191538 122196 191639
rect 123088 191577 123116 193022
rect 123166 192792 123222 192801
rect 123166 192727 123222 192736
rect 123074 191568 123130 191577
rect 122156 191532 122208 191538
rect 123074 191503 123130 191512
rect 122156 191474 122208 191480
rect 122982 191024 123038 191033
rect 123038 190982 123116 191010
rect 122982 190959 123038 190968
rect 88666 190888 88722 190897
rect 88666 190823 88722 190832
rect 88538 189894 88616 189922
rect 88482 189871 88538 189880
rect 88680 188834 88708 190823
rect 122982 189392 123038 189401
rect 122982 189327 123038 189336
rect 88758 189256 88814 189265
rect 88758 189191 88814 189200
rect 88496 188806 88708 188834
rect 88496 188721 88524 188806
rect 88482 188712 88538 188721
rect 88482 188647 88538 188656
rect 88666 188712 88722 188721
rect 88666 188647 88722 188656
rect 88680 188274 88708 188647
rect 88668 188268 88720 188274
rect 88668 188210 88720 188216
rect 88390 188168 88446 188177
rect 88390 188103 88446 188112
rect 88206 187488 88262 187497
rect 88206 187423 88262 187432
rect 88390 187488 88446 187497
rect 88390 187423 88446 187432
rect 87194 186264 87250 186273
rect 87194 186199 87250 186208
rect 88404 185185 88432 187423
rect 88482 187352 88538 187361
rect 88772 187338 88800 189191
rect 122996 188970 123024 189327
rect 123088 189129 123116 190982
rect 123180 190897 123208 192727
rect 123272 192121 123300 193815
rect 123364 192257 123392 194126
rect 123350 192248 123406 192257
rect 123350 192183 123406 192192
rect 123258 192112 123314 192121
rect 123258 192047 123314 192056
rect 123258 191976 123314 191985
rect 123258 191911 123314 191920
rect 123166 190888 123222 190897
rect 123166 190823 123222 190832
rect 123166 190480 123222 190489
rect 123166 190415 123222 190424
rect 123074 189120 123130 189129
rect 123074 189055 123130 189064
rect 122996 188942 123116 188970
rect 121970 188848 122026 188857
rect 121970 188783 121972 188792
rect 122024 188783 122026 188792
rect 121972 188754 122024 188760
rect 88850 188168 88906 188177
rect 88850 188103 88906 188112
rect 122982 188168 123038 188177
rect 122982 188103 123038 188112
rect 88538 187310 88800 187338
rect 88482 187287 88538 187296
rect 88574 186944 88630 186953
rect 88574 186879 88576 186888
rect 88628 186879 88630 186888
rect 88576 186850 88628 186856
rect 88864 186522 88892 188103
rect 122996 187202 123024 188103
rect 123088 187361 123116 188942
rect 123180 188177 123208 190415
rect 123272 190353 123300 191911
rect 123352 191532 123404 191538
rect 123352 191474 123404 191480
rect 123258 190344 123314 190353
rect 123258 190279 123314 190288
rect 123258 189936 123314 189945
rect 123258 189871 123314 189880
rect 123166 188168 123222 188177
rect 123166 188103 123222 188112
rect 123272 188041 123300 189871
rect 123364 189537 123392 191474
rect 123350 189528 123406 189537
rect 123350 189463 123406 189472
rect 123352 188812 123404 188818
rect 123352 188754 123404 188760
rect 123258 188032 123314 188041
rect 123258 187967 123314 187976
rect 123074 187352 123130 187361
rect 123074 187287 123130 187296
rect 122996 187174 123116 187202
rect 122430 187080 122486 187089
rect 122430 187015 122486 187024
rect 88496 186494 88892 186522
rect 88496 185729 88524 186494
rect 88574 186400 88630 186409
rect 88574 186335 88630 186344
rect 88588 185962 88616 186335
rect 88576 185956 88628 185962
rect 88576 185898 88628 185904
rect 88574 185856 88630 185865
rect 88574 185791 88630 185800
rect 88482 185720 88538 185729
rect 88588 185690 88616 185791
rect 88482 185655 88538 185664
rect 88576 185684 88628 185690
rect 88576 185626 88628 185632
rect 88666 185312 88722 185321
rect 88666 185247 88722 185256
rect 88390 185176 88446 185185
rect 88390 185111 88446 185120
rect 88574 184224 88630 184233
rect 88680 184194 88708 185247
rect 89218 184768 89274 184777
rect 89218 184703 89274 184712
rect 122338 184768 122394 184777
rect 122338 184703 122394 184712
rect 88574 184159 88630 184168
rect 88668 184188 88720 184194
rect 88588 184126 88616 184159
rect 88668 184130 88720 184136
rect 88576 184120 88628 184126
rect 88576 184062 88628 184068
rect 87838 183680 87894 183689
rect 87838 183615 87894 183624
rect 87852 178074 87880 183615
rect 88574 183136 88630 183145
rect 88574 183071 88630 183080
rect 88588 182766 88616 183071
rect 88576 182760 88628 182766
rect 88576 182702 88628 182708
rect 87840 178068 87892 178074
rect 87840 178010 87892 178016
rect 89232 178006 89260 184703
rect 122352 184194 122380 184703
rect 122340 184188 122392 184194
rect 122340 184130 122392 184136
rect 122154 183136 122210 183145
rect 122154 183071 122210 183080
rect 91348 182958 92098 182986
rect 92268 182958 92558 182986
rect 92728 182958 93110 182986
rect 93280 182958 93662 182986
rect 94108 182958 94214 182986
rect 94384 182958 94766 182986
rect 94936 182958 95318 182986
rect 95488 182958 95870 182986
rect 100180 182958 100286 182986
rect 100732 182958 100838 182986
rect 101284 182958 101390 182986
rect 101836 182958 101942 182986
rect 102388 182958 102494 182986
rect 102940 182958 103046 182986
rect 103952 182958 104150 182986
rect 105148 182958 105254 182986
rect 105516 182958 105806 182986
rect 106160 182958 106266 182986
rect 106528 182958 106818 182986
rect 107080 182958 107370 182986
rect 108184 182958 108474 182986
rect 108736 182958 109026 182986
rect 109380 182958 109578 182986
rect 109840 182958 110130 182986
rect 110944 182958 111234 182986
rect 111496 182958 111786 182986
rect 112048 182958 112338 182986
rect 112600 182958 112890 182986
rect 113704 182958 113994 182986
rect 114256 182958 114546 182986
rect 114808 182958 115098 182986
rect 115360 182958 115650 182986
rect 116464 182958 116754 182986
rect 117016 182958 117306 182986
rect 117568 182958 117858 182986
rect 89220 178000 89272 178006
rect 89220 177942 89272 177948
rect 88208 177864 88260 177870
rect 88208 177806 88260 177812
rect 88220 175764 88248 177806
rect 49948 175614 50514 175642
rect 45058 171848 45114 171857
rect 45058 171783 45114 171792
rect 22244 167596 22296 167602
rect 22244 167538 22296 167544
rect 22256 163833 22284 167538
rect 22242 163824 22298 163833
rect 22242 163759 22298 163768
rect 45072 156450 45100 171783
rect 48462 169264 48518 169273
rect 48462 169199 48518 169208
rect 45060 156444 45112 156450
rect 45060 156386 45112 156392
rect 47820 156444 47872 156450
rect 47820 156386 47872 156392
rect 47832 155945 47860 156386
rect 47818 155936 47874 155945
rect 47818 155871 47874 155880
rect 22334 155800 22390 155809
rect 22334 155735 22390 155744
rect 22348 155158 22376 155735
rect 22336 155152 22388 155158
rect 22336 155094 22388 155100
rect 22334 147776 22390 147785
rect 22334 147711 22390 147720
rect 45794 147776 45850 147785
rect 45794 147711 45850 147720
rect 22348 146862 22376 147711
rect 22336 146856 22388 146862
rect 22336 146798 22388 146804
rect 45808 142617 45836 147711
rect 45794 142608 45850 142617
rect 45794 142543 45850 142552
rect 44414 139888 44470 139897
rect 44414 139823 44470 139832
rect 23624 134276 23676 134282
rect 23624 134218 23676 134224
rect 22888 133052 22940 133058
rect 22888 132994 22940 133000
rect 21508 131420 21560 131426
rect 21508 131362 21560 131368
rect 20220 130944 20272 130950
rect 20220 130886 20272 130892
rect 20232 128708 20260 130886
rect 20864 130332 20916 130338
rect 20864 130274 20916 130280
rect 20876 128708 20904 130274
rect 21520 128708 21548 131362
rect 22244 131284 22296 131290
rect 22244 131226 22296 131232
rect 22256 128708 22284 131226
rect 22900 128708 22928 132994
rect 23636 128708 23664 134218
rect 26120 133398 26148 135916
rect 26292 133936 26344 133942
rect 26292 133878 26344 133884
rect 25004 133392 25056 133398
rect 25004 133334 25056 133340
rect 26108 133392 26160 133398
rect 26108 133334 26160 133340
rect 24912 133256 24964 133262
rect 24912 133198 24964 133204
rect 24268 133188 24320 133194
rect 24268 133130 24320 133136
rect 24280 128708 24308 133130
rect 24924 128708 24952 133198
rect 25016 130338 25044 133334
rect 25648 133120 25700 133126
rect 25648 133062 25700 133068
rect 25004 130332 25056 130338
rect 25004 130274 25056 130280
rect 25660 128708 25688 133062
rect 26304 128708 26332 133878
rect 26488 131426 26516 135916
rect 26476 131420 26528 131426
rect 26476 131362 26528 131368
rect 26856 131290 26884 135916
rect 27028 134004 27080 134010
rect 27028 133946 27080 133952
rect 26844 131284 26896 131290
rect 26844 131226 26896 131232
rect 27040 128708 27068 133946
rect 27316 133058 27344 135916
rect 27684 134282 27712 135916
rect 27672 134276 27724 134282
rect 27672 134218 27724 134224
rect 27672 133732 27724 133738
rect 27672 133674 27724 133680
rect 27304 133052 27356 133058
rect 27304 132994 27356 133000
rect 27684 128708 27712 133674
rect 28052 133194 28080 135916
rect 28316 133868 28368 133874
rect 28316 133810 28368 133816
rect 28040 133188 28092 133194
rect 28040 133130 28092 133136
rect 28328 128708 28356 133810
rect 28512 133262 28540 135916
rect 28500 133256 28552 133262
rect 28500 133198 28552 133204
rect 28880 133126 28908 135916
rect 29248 133942 29276 135916
rect 29708 134010 29736 135916
rect 29696 134004 29748 134010
rect 29696 133946 29748 133952
rect 29236 133936 29288 133942
rect 29236 133878 29288 133884
rect 29696 133800 29748 133806
rect 29696 133742 29748 133748
rect 29052 133460 29104 133466
rect 29052 133402 29104 133408
rect 28868 133120 28920 133126
rect 28868 133062 28920 133068
rect 29064 128708 29092 133402
rect 29708 128708 29736 133742
rect 30076 133738 30104 135916
rect 30444 133874 30472 135916
rect 30432 133868 30484 133874
rect 30432 133810 30484 133816
rect 30064 133732 30116 133738
rect 30064 133674 30116 133680
rect 30904 133466 30932 135916
rect 31076 133868 31128 133874
rect 31076 133810 31128 133816
rect 30892 133460 30944 133466
rect 30892 133402 30944 133408
rect 30432 133324 30484 133330
rect 30432 133266 30484 133272
rect 30444 128708 30472 133266
rect 31088 128708 31116 133810
rect 31272 133806 31300 135916
rect 31260 133800 31312 133806
rect 31260 133742 31312 133748
rect 31640 133330 31668 135916
rect 32100 133874 32128 135916
rect 32192 135902 32482 135930
rect 32088 133868 32140 133874
rect 32088 133810 32140 133816
rect 32192 133754 32220 135902
rect 31824 133726 32220 133754
rect 31628 133324 31680 133330
rect 31628 133266 31680 133272
rect 31824 128708 31852 133726
rect 32836 128722 32864 135916
rect 33296 128722 33324 135916
rect 32482 128694 32864 128722
rect 33126 128694 33324 128722
rect 33664 128722 33692 135916
rect 34124 128722 34152 135916
rect 34492 133466 34520 135916
rect 34860 133806 34888 135916
rect 34848 133800 34900 133806
rect 34848 133742 34900 133748
rect 34480 133460 34532 133466
rect 34480 133402 34532 133408
rect 35216 133460 35268 133466
rect 35216 133402 35268 133408
rect 33664 128694 33862 128722
rect 34124 128694 34506 128722
rect 35228 128708 35256 133402
rect 35320 133126 35348 135916
rect 35688 133194 35716 135916
rect 35860 133800 35912 133806
rect 35860 133742 35912 133748
rect 35676 133188 35728 133194
rect 35676 133130 35728 133136
rect 35308 133120 35360 133126
rect 35308 133062 35360 133068
rect 35872 128708 35900 133742
rect 36056 133058 36084 135916
rect 36516 133806 36544 135916
rect 36504 133800 36556 133806
rect 36504 133742 36556 133748
rect 36884 133466 36912 135916
rect 37252 133874 37280 135916
rect 37712 133942 37740 135916
rect 37700 133936 37752 133942
rect 37700 133878 37752 133884
rect 37240 133868 37292 133874
rect 37240 133810 37292 133816
rect 38080 133670 38108 135916
rect 38448 134010 38476 135916
rect 38436 134004 38488 134010
rect 38436 133946 38488 133952
rect 38620 133800 38672 133806
rect 38620 133742 38672 133748
rect 38068 133664 38120 133670
rect 38068 133606 38120 133612
rect 36872 133460 36924 133466
rect 36872 133402 36924 133408
rect 37240 133188 37292 133194
rect 37240 133130 37292 133136
rect 36504 133120 36556 133126
rect 36504 133062 36556 133068
rect 36044 133052 36096 133058
rect 36044 132994 36096 133000
rect 36516 128708 36544 133062
rect 37252 128708 37280 133130
rect 37884 133052 37936 133058
rect 37884 132994 37936 133000
rect 37896 128708 37924 132994
rect 38632 128708 38660 133742
rect 38908 133398 38936 135916
rect 39276 133602 39304 135916
rect 39264 133596 39316 133602
rect 39264 133538 39316 133544
rect 39644 133534 39672 135916
rect 40000 133868 40052 133874
rect 40000 133810 40052 133816
rect 39632 133528 39684 133534
rect 39632 133470 39684 133476
rect 39264 133460 39316 133466
rect 39264 133402 39316 133408
rect 38896 133392 38948 133398
rect 38896 133334 38948 133340
rect 39276 128708 39304 133402
rect 40012 128708 40040 133810
rect 40104 133466 40132 135916
rect 40472 133738 40500 135916
rect 40644 133936 40696 133942
rect 40644 133878 40696 133884
rect 40460 133732 40512 133738
rect 40460 133674 40512 133680
rect 40092 133460 40144 133466
rect 40092 133402 40144 133408
rect 40656 128708 40684 133878
rect 40840 133874 40868 135916
rect 40828 133868 40880 133874
rect 40828 133810 40880 133816
rect 41300 133806 41328 135916
rect 41564 134004 41616 134010
rect 41564 133946 41616 133952
rect 41288 133800 41340 133806
rect 41288 133742 41340 133748
rect 41012 133664 41064 133670
rect 41012 133606 41064 133612
rect 41024 128722 41052 133606
rect 41576 130354 41604 133946
rect 41668 133126 41696 135916
rect 43588 133868 43640 133874
rect 43588 133810 43640 133816
rect 43036 133732 43088 133738
rect 43036 133674 43088 133680
rect 42944 133596 42996 133602
rect 42944 133538 42996 133544
rect 41840 133528 41892 133534
rect 41840 133470 41892 133476
rect 41656 133120 41708 133126
rect 41656 133062 41708 133068
rect 41576 130326 41788 130354
rect 41852 130338 41880 133470
rect 42300 133460 42352 133466
rect 42300 133402 42352 133408
rect 42312 130406 42340 133402
rect 42668 133392 42720 133398
rect 42668 133334 42720 133340
rect 42300 130400 42352 130406
rect 42300 130342 42352 130348
rect 41760 128722 41788 130326
rect 41840 130332 41892 130338
rect 41840 130274 41892 130280
rect 41024 128694 41314 128722
rect 41760 128694 42050 128722
rect 42680 128708 42708 133334
rect 42956 130354 42984 133538
rect 43048 130474 43076 133674
rect 43600 131426 43628 133810
rect 44324 133800 44376 133806
rect 44324 133742 44376 133748
rect 43588 131420 43640 131426
rect 43588 131362 43640 131368
rect 44336 131154 44364 133742
rect 44324 131148 44376 131154
rect 44324 131090 44376 131096
rect 44428 130950 44456 139823
rect 48476 134758 48504 169199
rect 91348 166689 91376 182958
rect 92268 180538 92296 182958
rect 91532 180510 92296 180538
rect 91532 179314 91560 180510
rect 92164 180312 92216 180318
rect 92164 180254 92216 180260
rect 91980 180040 92032 180046
rect 91980 179982 92032 179988
rect 92072 180040 92124 180046
rect 92072 179982 92124 179988
rect 91440 179286 91560 179314
rect 91440 167913 91468 179286
rect 91992 169137 92020 179982
rect 92084 170361 92112 179982
rect 92176 172809 92204 180254
rect 92440 180244 92492 180250
rect 92440 180186 92492 180192
rect 92348 180108 92400 180114
rect 92348 180050 92400 180056
rect 92256 179972 92308 179978
rect 92256 179914 92308 179920
rect 92162 172800 92218 172809
rect 92162 172735 92218 172744
rect 92268 171585 92296 179914
rect 92360 174033 92388 180050
rect 92452 180046 92480 180186
rect 92728 180182 92756 182958
rect 93280 180250 93308 182958
rect 93268 180244 93320 180250
rect 93268 180186 93320 180192
rect 92716 180176 92768 180182
rect 92716 180118 92768 180124
rect 92440 180040 92492 180046
rect 92440 179982 92492 179988
rect 92624 180040 92676 180046
rect 92624 179982 92676 179988
rect 92636 175257 92664 179982
rect 94108 179978 94136 182958
rect 94384 180318 94412 182958
rect 94372 180312 94424 180318
rect 94372 180254 94424 180260
rect 94936 180114 94964 182958
rect 94924 180108 94976 180114
rect 94924 180050 94976 180056
rect 95488 180046 95516 182958
rect 96422 182822 96712 182850
rect 96974 182822 97264 182850
rect 97526 182822 97816 182850
rect 98078 182822 98184 182850
rect 98630 182822 98920 182850
rect 99182 182822 99380 182850
rect 99734 182822 99840 182850
rect 95476 180040 95528 180046
rect 95476 179982 95528 179988
rect 96684 179978 96712 182822
rect 97236 180046 97264 182822
rect 97788 180114 97816 182822
rect 97776 180108 97828 180114
rect 97776 180050 97828 180056
rect 97224 180040 97276 180046
rect 97224 179982 97276 179988
rect 98156 179978 98184 182822
rect 98892 180250 98920 182822
rect 99352 180930 99380 182822
rect 99812 181354 99840 182822
rect 99720 181326 99840 181354
rect 100180 181354 100208 182958
rect 100180 181326 100300 181354
rect 99340 180924 99392 180930
rect 99340 180866 99392 180872
rect 98880 180244 98932 180250
rect 98880 180186 98932 180192
rect 99616 180244 99668 180250
rect 99616 180186 99668 180192
rect 98696 180108 98748 180114
rect 98696 180050 98748 180056
rect 98236 180040 98288 180046
rect 98236 179982 98288 179988
rect 94096 179972 94148 179978
rect 94096 179914 94148 179920
rect 96672 179972 96724 179978
rect 96672 179914 96724 179920
rect 97776 179972 97828 179978
rect 97776 179914 97828 179920
rect 98144 179972 98196 179978
rect 98144 179914 98196 179920
rect 97788 175778 97816 179914
rect 98248 175778 98276 179982
rect 98708 175778 98736 180050
rect 98972 179972 99024 179978
rect 98972 179914 99024 179920
rect 98984 175778 99012 179914
rect 99628 176050 99656 180186
rect 99720 177666 99748 181326
rect 99800 180924 99852 180930
rect 99800 180866 99852 180872
rect 99708 177660 99760 177666
rect 99708 177602 99760 177608
rect 99628 176022 99702 176050
rect 97788 175750 98124 175778
rect 98248 175750 98492 175778
rect 98708 175750 98860 175778
rect 98984 175750 99320 175778
rect 99674 175764 99702 176022
rect 99812 175778 99840 180866
rect 100272 177666 100300 181326
rect 100732 179978 100760 182958
rect 101284 181354 101312 182958
rect 101836 181354 101864 182958
rect 102388 181354 102416 182958
rect 102940 181354 102968 182958
rect 103598 182822 103704 182850
rect 103676 181354 103704 182822
rect 101284 181326 101404 181354
rect 101836 181326 101956 181354
rect 102388 181326 102508 181354
rect 102940 181326 103060 181354
rect 100720 179972 100772 179978
rect 100720 179914 100772 179920
rect 100996 179972 101048 179978
rect 100996 179914 101048 179920
rect 100168 177660 100220 177666
rect 100168 177602 100220 177608
rect 100260 177660 100312 177666
rect 100260 177602 100312 177608
rect 100720 177660 100772 177666
rect 100720 177602 100772 177608
rect 100180 175778 100208 177602
rect 100732 175778 100760 177602
rect 101008 175778 101036 179914
rect 101376 175778 101404 181326
rect 101928 175778 101956 181326
rect 102480 176050 102508 181326
rect 102434 176022 102508 176050
rect 99812 175750 100056 175778
rect 100180 175750 100516 175778
rect 100732 175750 100884 175778
rect 101008 175750 101252 175778
rect 101376 175750 101712 175778
rect 101928 175750 102080 175778
rect 102434 175764 102462 176022
rect 103032 175778 103060 181326
rect 103584 181326 103704 181354
rect 103584 175914 103612 181326
rect 103492 175886 103612 175914
rect 103492 175778 103520 175886
rect 102908 175750 103060 175778
rect 103276 175750 103520 175778
rect 103952 175642 103980 182958
rect 104702 182822 104808 182850
rect 104780 181354 104808 182822
rect 104688 181326 104808 181354
rect 104688 177666 104716 181326
rect 105148 181218 105176 182958
rect 104780 181190 105176 181218
rect 104216 177660 104268 177666
rect 104216 177602 104268 177608
rect 104676 177660 104728 177666
rect 104676 177602 104728 177608
rect 104228 175778 104256 177602
rect 104780 176050 104808 181190
rect 105516 179978 105544 182958
rect 105964 180788 106016 180794
rect 105964 180730 106016 180736
rect 105044 179972 105096 179978
rect 105044 179914 105096 179920
rect 105504 179972 105556 179978
rect 105504 179914 105556 179920
rect 104688 176022 104808 176050
rect 104688 175778 104716 176022
rect 105056 175778 105084 179914
rect 105504 177524 105556 177530
rect 105504 177466 105556 177472
rect 105516 175778 105544 177466
rect 105976 175778 106004 180730
rect 106160 177530 106188 182958
rect 106240 181196 106292 181202
rect 106240 181138 106292 181144
rect 106148 177524 106200 177530
rect 106148 177466 106200 177472
rect 106252 175778 106280 181138
rect 106528 180794 106556 182958
rect 106700 181332 106752 181338
rect 106700 181274 106752 181280
rect 106516 180788 106568 180794
rect 106516 180730 106568 180736
rect 106712 175778 106740 181274
rect 107080 181202 107108 182958
rect 107922 182822 108028 182850
rect 108000 181338 108028 182822
rect 107988 181332 108040 181338
rect 107988 181274 108040 181280
rect 108184 181270 108212 182958
rect 108356 181332 108408 181338
rect 108356 181274 108408 181280
rect 107160 181264 107212 181270
rect 107160 181206 107212 181212
rect 108172 181264 108224 181270
rect 108172 181206 108224 181212
rect 107068 181196 107120 181202
rect 107068 181138 107120 181144
rect 107172 175778 107200 181206
rect 107528 181196 107580 181202
rect 107528 181138 107580 181144
rect 107540 175778 107568 181138
rect 107804 180244 107856 180250
rect 107804 180186 107856 180192
rect 107816 175778 107844 180186
rect 108368 175778 108396 181274
rect 108736 181202 108764 182958
rect 108724 181196 108776 181202
rect 108724 181138 108776 181144
rect 109092 181196 109144 181202
rect 109092 181138 109144 181144
rect 108724 181060 108776 181066
rect 108724 181002 108776 181008
rect 108736 175778 108764 181002
rect 109104 175778 109132 181138
rect 109380 180250 109408 182958
rect 109840 181338 109868 182958
rect 110682 182822 110788 182850
rect 109828 181332 109880 181338
rect 109828 181274 109880 181280
rect 110760 181066 110788 182822
rect 110944 181202 110972 182958
rect 110932 181196 110984 181202
rect 110932 181138 110984 181144
rect 110748 181060 110800 181066
rect 110748 181002 110800 181008
rect 110564 180312 110616 180318
rect 110564 180254 110616 180260
rect 109368 180244 109420 180250
rect 109368 180186 109420 180192
rect 110288 180108 110340 180114
rect 110288 180050 110340 180056
rect 109920 180040 109972 180046
rect 109920 179982 109972 179988
rect 109552 179972 109604 179978
rect 109552 179914 109604 179920
rect 109564 175778 109592 179914
rect 109932 175778 109960 179982
rect 110300 175778 110328 180050
rect 110576 175778 110604 180254
rect 111116 180244 111168 180250
rect 111116 180186 111168 180192
rect 111128 175778 111156 180186
rect 111496 179978 111524 182958
rect 111576 180176 111628 180182
rect 111576 180118 111628 180124
rect 111484 179972 111536 179978
rect 111484 179914 111536 179920
rect 111588 179314 111616 180118
rect 112048 180046 112076 182958
rect 112600 180114 112628 182958
rect 113442 182822 113548 182850
rect 113520 180318 113548 182822
rect 113508 180312 113560 180318
rect 113508 180254 113560 180260
rect 113704 180250 113732 182958
rect 113692 180244 113744 180250
rect 113692 180186 113744 180192
rect 114256 180182 114284 182958
rect 114244 180176 114296 180182
rect 114244 180118 114296 180124
rect 112588 180108 112640 180114
rect 112588 180050 112640 180056
rect 112036 180040 112088 180046
rect 112036 179982 112088 179988
rect 112220 180040 112272 180046
rect 112220 179982 112272 179988
rect 111944 179972 111996 179978
rect 111944 179914 111996 179920
rect 111496 179286 111616 179314
rect 111496 175778 111524 179286
rect 111956 175778 111984 179914
rect 112232 175778 112260 179982
rect 114808 179978 114836 182958
rect 115360 180046 115388 182958
rect 116202 182822 116308 182850
rect 115348 180040 115400 180046
rect 115348 179982 115400 179988
rect 114796 179972 114848 179978
rect 114796 179914 114848 179920
rect 113048 178544 113100 178550
rect 113048 178486 113100 178492
rect 112680 178408 112732 178414
rect 112680 178350 112732 178356
rect 112692 175778 112720 178350
rect 113060 175778 113088 178486
rect 113508 178476 113560 178482
rect 113508 178418 113560 178424
rect 104104 175750 104256 175778
rect 104472 175750 104716 175778
rect 104840 175750 105084 175778
rect 105300 175750 105544 175778
rect 105668 175750 106004 175778
rect 106128 175750 106280 175778
rect 106496 175750 106740 175778
rect 106864 175750 107200 175778
rect 107324 175750 107568 175778
rect 107692 175750 107844 175778
rect 108060 175750 108396 175778
rect 108520 175750 108764 175778
rect 108888 175750 109132 175778
rect 109256 175750 109592 175778
rect 109716 175750 109960 175778
rect 110084 175750 110328 175778
rect 110452 175750 110604 175778
rect 110912 175750 111156 175778
rect 111280 175750 111524 175778
rect 111648 175750 111984 175778
rect 112108 175750 112260 175778
rect 112476 175750 112720 175778
rect 112844 175750 113088 175778
rect 113520 175642 113548 178418
rect 116280 178414 116308 182822
rect 116464 178550 116492 182958
rect 116452 178544 116504 178550
rect 116452 178486 116504 178492
rect 117016 178482 117044 182958
rect 117004 178476 117056 178482
rect 117004 178418 117056 178424
rect 116268 178408 116320 178414
rect 116268 178350 116320 178356
rect 117568 178074 117596 182958
rect 113968 178068 114020 178074
rect 113968 178010 114020 178016
rect 117556 178068 117608 178074
rect 117556 178010 117608 178016
rect 113980 175778 114008 178010
rect 113672 175750 114008 175778
rect 122168 175778 122196 183071
rect 122444 177938 122472 187015
rect 122890 186536 122946 186545
rect 122890 186471 122946 186480
rect 122904 186030 122932 186471
rect 123088 186137 123116 187174
rect 123364 186817 123392 188754
rect 123534 187624 123590 187633
rect 123534 187559 123590 187568
rect 123350 186808 123406 186817
rect 123350 186743 123406 186752
rect 123074 186128 123130 186137
rect 123074 186063 123130 186072
rect 122892 186024 122944 186030
rect 122892 185966 122944 185972
rect 122982 185992 123038 186001
rect 122982 185927 123038 185936
rect 122996 185758 123024 185927
rect 122984 185752 123036 185758
rect 122984 185694 123036 185700
rect 122890 185312 122946 185321
rect 122890 185247 122946 185256
rect 122904 184262 122932 185247
rect 123548 185185 123576 187559
rect 126480 186024 126532 186030
rect 126480 185966 126532 185972
rect 123534 185176 123590 185185
rect 123534 185111 123590 185120
rect 122892 184256 122944 184262
rect 124456 184256 124508 184262
rect 122892 184198 122944 184204
rect 122982 184224 123038 184233
rect 124456 184198 124508 184204
rect 122982 184159 123038 184168
rect 122996 184126 123024 184159
rect 122984 184120 123036 184126
rect 122984 184062 123036 184068
rect 123074 183680 123130 183689
rect 123074 183615 123130 183624
rect 122616 182828 122668 182834
rect 122616 182770 122668 182776
rect 122628 182698 122656 182770
rect 122616 182692 122668 182698
rect 122616 182634 122668 182640
rect 122432 177932 122484 177938
rect 122432 177874 122484 177880
rect 122168 175750 122504 175778
rect 103644 175614 103980 175642
rect 113304 175614 113548 175642
rect 123088 175642 123116 183615
rect 124468 178414 124496 184198
rect 125468 184188 125520 184194
rect 125468 184130 125520 184136
rect 124548 184120 124600 184126
rect 124548 184062 124600 184068
rect 124456 178408 124508 178414
rect 124456 178350 124508 178356
rect 124560 175778 124588 184062
rect 125480 175778 125508 184130
rect 126492 177734 126520 185966
rect 126572 185752 126624 185758
rect 126572 185694 126624 185700
rect 126584 178550 126612 185694
rect 156852 185298 156880 210310
rect 160334 209928 160390 209937
rect 160334 209863 160390 209872
rect 160242 208432 160298 208441
rect 160348 208418 160376 209863
rect 191708 209620 191760 209626
rect 191708 209562 191760 209568
rect 160426 209384 160482 209393
rect 160426 209319 160482 209328
rect 160298 208390 160376 208418
rect 160242 208367 160298 208376
rect 160242 207888 160298 207897
rect 160440 207874 160468 209319
rect 191720 208985 191748 209562
rect 191706 208976 191762 208985
rect 191706 208911 191762 208920
rect 160518 208840 160574 208849
rect 160518 208775 160574 208784
rect 160298 207846 160468 207874
rect 160242 207823 160298 207832
rect 160150 207616 160206 207625
rect 160150 207551 160206 207560
rect 159048 207240 159100 207246
rect 159046 207208 159048 207217
rect 159100 207208 159102 207217
rect 159046 207143 159102 207152
rect 159048 206832 159100 206838
rect 159048 206774 159100 206780
rect 159060 206673 159088 206774
rect 159046 206664 159102 206673
rect 159046 206599 159102 206608
rect 160164 206129 160192 207551
rect 160532 207246 160560 208775
rect 160610 207888 160666 207897
rect 160610 207823 160666 207832
rect 160520 207240 160572 207246
rect 160520 207182 160572 207188
rect 160426 207072 160482 207081
rect 160426 207007 160482 207016
rect 160334 206528 160390 206537
rect 160334 206463 160390 206472
rect 160150 206120 160206 206129
rect 160150 206055 160206 206064
rect 160348 205698 160376 206463
rect 160164 205670 160376 205698
rect 160164 204905 160192 205670
rect 160440 205562 160468 207007
rect 160624 206838 160652 207823
rect 160612 206832 160664 206838
rect 160612 206774 160664 206780
rect 160518 205984 160574 205993
rect 160518 205919 160574 205928
rect 160256 205534 160468 205562
rect 160256 205449 160284 205534
rect 160242 205440 160298 205449
rect 160242 205375 160298 205384
rect 160334 205304 160390 205313
rect 160334 205239 160390 205248
rect 160150 204896 160206 204905
rect 160150 204831 160206 204840
rect 160348 204066 160376 205239
rect 160532 204905 160560 205919
rect 160518 204896 160574 204905
rect 160518 204831 160574 204840
rect 160426 204760 160482 204769
rect 160426 204695 160482 204704
rect 160256 204038 160376 204066
rect 160256 203681 160284 204038
rect 160334 203944 160390 203953
rect 160334 203879 160390 203888
rect 160242 203672 160298 203681
rect 160242 203607 160298 203616
rect 159048 203432 159100 203438
rect 159048 203374 159100 203380
rect 158956 201936 159008 201942
rect 159060 201913 159088 203374
rect 160242 202448 160298 202457
rect 160348 202434 160376 203879
rect 160440 203545 160468 204695
rect 160518 203672 160574 203681
rect 160518 203607 160574 203616
rect 160426 203536 160482 203545
rect 160426 203471 160482 203480
rect 160532 203438 160560 203607
rect 160520 203432 160572 203438
rect 160520 203374 160572 203380
rect 160610 203128 160666 203137
rect 160610 203063 160666 203072
rect 160298 202406 160376 202434
rect 160426 202448 160482 202457
rect 160242 202383 160298 202392
rect 160426 202383 160482 202392
rect 158956 201878 159008 201884
rect 159046 201904 159102 201913
rect 158968 201233 158996 201878
rect 159046 201839 159102 201848
rect 160440 201482 160468 202383
rect 160624 201942 160652 203063
rect 160612 201936 160664 201942
rect 160518 201904 160574 201913
rect 160612 201878 160664 201884
rect 160518 201839 160574 201848
rect 160256 201454 160468 201482
rect 158954 201224 159010 201233
rect 158954 201159 159010 201168
rect 160150 200816 160206 200825
rect 160150 200751 160206 200760
rect 160164 198921 160192 200751
rect 160256 200689 160284 201454
rect 160334 201360 160390 201369
rect 160334 201295 160390 201304
rect 160242 200680 160298 200689
rect 160242 200615 160298 200624
rect 160242 199456 160298 199465
rect 160348 199442 160376 201295
rect 160532 200689 160560 201839
rect 160518 200680 160574 200689
rect 160518 200615 160574 200624
rect 160518 200272 160574 200281
rect 160518 200207 160574 200216
rect 160298 199414 160376 199442
rect 160242 199391 160298 199400
rect 160242 199320 160298 199329
rect 160242 199255 160298 199264
rect 160150 198912 160206 198921
rect 160150 198847 160206 198856
rect 158956 198740 159008 198746
rect 158956 198682 159008 198688
rect 158968 198241 158996 198682
rect 160058 198504 160114 198513
rect 160058 198439 160114 198448
rect 158954 198232 159010 198241
rect 158954 198167 159010 198176
rect 160072 196473 160100 198439
rect 160256 198354 160284 199255
rect 160426 199048 160482 199057
rect 160426 198983 160482 198992
rect 160164 198326 160284 198354
rect 160164 197697 160192 198326
rect 160242 197960 160298 197969
rect 160242 197895 160298 197904
rect 160150 197688 160206 197697
rect 160150 197623 160206 197632
rect 160256 197266 160284 197895
rect 160164 197238 160284 197266
rect 160058 196464 160114 196473
rect 160058 196399 160114 196408
rect 160164 195929 160192 197238
rect 160242 197144 160298 197153
rect 160440 197130 160468 198983
rect 160532 198746 160560 200207
rect 160520 198740 160572 198746
rect 160520 198682 160572 198688
rect 160518 197416 160574 197425
rect 160518 197351 160574 197360
rect 160298 197102 160468 197130
rect 160242 197079 160298 197088
rect 160242 196736 160298 196745
rect 160242 196671 160298 196680
rect 160150 195920 160206 195929
rect 160150 195855 160206 195864
rect 160150 195648 160206 195657
rect 160150 195583 160206 195592
rect 158956 195408 159008 195414
rect 158956 195350 159008 195356
rect 158968 195249 158996 195350
rect 158954 195240 159010 195249
rect 158954 195175 159010 195184
rect 159966 194560 160022 194569
rect 159966 194495 160022 194504
rect 159980 192257 160008 194495
rect 160058 193880 160114 193889
rect 160058 193815 160114 193824
rect 159966 192248 160022 192257
rect 159966 192183 160022 192192
rect 160072 192121 160100 193815
rect 160164 193481 160192 195583
rect 160256 194705 160284 196671
rect 160334 196192 160390 196201
rect 160334 196127 160390 196136
rect 160242 194696 160298 194705
rect 160242 194631 160298 194640
rect 160242 194152 160298 194161
rect 160348 194138 160376 196127
rect 160532 195414 160560 197351
rect 160520 195408 160572 195414
rect 160520 195350 160572 195356
rect 160426 195104 160482 195113
rect 160426 195039 160482 195048
rect 160298 194110 160376 194138
rect 160242 194087 160298 194096
rect 160150 193472 160206 193481
rect 160150 193407 160206 193416
rect 160440 193050 160468 195039
rect 160518 193336 160574 193345
rect 160518 193271 160574 193280
rect 160256 193022 160468 193050
rect 160256 192937 160284 193022
rect 160242 192928 160298 192937
rect 160242 192863 160298 192872
rect 160150 192792 160206 192801
rect 160150 192727 160206 192736
rect 160058 192112 160114 192121
rect 160058 192047 160114 192056
rect 160058 191704 160114 191713
rect 160058 191639 160114 191648
rect 158956 190920 159008 190926
rect 158956 190862 159008 190868
rect 158968 189945 158996 190862
rect 158954 189936 159010 189945
rect 158954 189871 159010 189880
rect 159966 189664 160022 189673
rect 159966 189599 160022 189608
rect 159980 187497 160008 189599
rect 160072 189265 160100 191639
rect 160164 190897 160192 192727
rect 160242 191160 160298 191169
rect 160532 191146 160560 193271
rect 160610 192248 160666 192257
rect 160610 192183 160666 192192
rect 160298 191118 160560 191146
rect 160242 191095 160298 191104
rect 160242 191024 160298 191033
rect 160242 190959 160298 190968
rect 160150 190888 160206 190897
rect 160150 190823 160206 190832
rect 160150 190480 160206 190489
rect 160150 190415 160206 190424
rect 160058 189256 160114 189265
rect 160058 189191 160114 189200
rect 160058 188848 160114 188857
rect 160058 188783 160114 188792
rect 159966 187488 160022 187497
rect 159966 187423 160022 187432
rect 160072 186273 160100 188783
rect 160164 188177 160192 190415
rect 160256 188721 160284 190959
rect 160624 190926 160652 192183
rect 160612 190920 160664 190926
rect 160612 190862 160664 190868
rect 160334 189392 160390 189401
rect 160334 189327 160390 189336
rect 160242 188712 160298 188721
rect 160242 188647 160298 188656
rect 160150 188168 160206 188177
rect 160150 188103 160206 188112
rect 160150 187624 160206 187633
rect 160150 187559 160206 187568
rect 160058 186264 160114 186273
rect 160058 186199 160114 186208
rect 157484 185616 157536 185622
rect 157484 185558 157536 185564
rect 156130 185270 156880 185298
rect 154354 185040 154410 185049
rect 154410 184998 154658 185026
rect 154354 184975 154410 184984
rect 127596 182698 127624 184876
rect 128608 184862 128990 184890
rect 127584 182692 127636 182698
rect 127584 182634 127636 182640
rect 126572 178544 126624 178550
rect 126572 178486 126624 178492
rect 127676 178544 127728 178550
rect 127676 178486 127728 178492
rect 126664 178408 126716 178414
rect 126664 178350 126716 178356
rect 126480 177728 126532 177734
rect 126480 177670 126532 177676
rect 126676 175778 126704 178350
rect 127688 175778 127716 178486
rect 128608 177870 128636 184862
rect 130448 181338 130476 184876
rect 131368 184862 131842 184890
rect 132840 184862 133314 184890
rect 134128 184862 134694 184890
rect 131368 182442 131396 184862
rect 131276 182414 131396 182442
rect 130436 181332 130488 181338
rect 130436 181274 130488 181280
rect 129976 177932 130028 177938
rect 129976 177874 130028 177880
rect 128596 177864 128648 177870
rect 128596 177806 128648 177812
rect 128780 177728 128832 177734
rect 128780 177670 128832 177676
rect 128792 175778 128820 177670
rect 129988 175778 130016 177874
rect 131276 175778 131304 182414
rect 132840 181354 132868 184862
rect 134128 182442 134156 184862
rect 132656 181326 132868 181354
rect 133944 182414 134156 182442
rect 132656 175778 132684 181326
rect 133944 175778 133972 182414
rect 136152 182222 136180 184876
rect 137244 182420 137296 182426
rect 137244 182362 137296 182368
rect 134944 182216 134996 182222
rect 134944 182158 134996 182164
rect 136140 182216 136192 182222
rect 136140 182158 136192 182164
rect 134956 175778 134984 182158
rect 136140 182080 136192 182086
rect 136140 182022 136192 182028
rect 136152 175778 136180 182022
rect 137256 175778 137284 182362
rect 137532 182086 137560 184876
rect 139004 182426 139032 184876
rect 138992 182420 139044 182426
rect 138992 182362 139044 182368
rect 139452 182420 139504 182426
rect 139452 182362 139504 182368
rect 137520 182080 137572 182086
rect 137520 182022 137572 182028
rect 138164 182012 138216 182018
rect 138164 181954 138216 181960
rect 138176 175778 138204 181954
rect 139464 175778 139492 182362
rect 140384 182018 140412 184876
rect 141856 182426 141884 184876
rect 141844 182420 141896 182426
rect 141844 182362 141896 182368
rect 142764 182420 142816 182426
rect 142764 182362 142816 182368
rect 140372 182012 140424 182018
rect 140372 181954 140424 181960
rect 140556 181468 140608 181474
rect 140556 181410 140608 181416
rect 140568 175778 140596 181410
rect 141660 181400 141712 181406
rect 141660 181342 141712 181348
rect 141672 175778 141700 181342
rect 142776 175778 142804 182362
rect 143236 181474 143264 184876
rect 143684 182488 143736 182494
rect 143684 182430 143736 182436
rect 143224 181468 143276 181474
rect 143224 181410 143276 181416
rect 143696 175778 143724 182430
rect 144708 181406 144736 184876
rect 146088 182426 146116 184876
rect 147560 182494 147588 184876
rect 147548 182488 147600 182494
rect 147548 182430 147600 182436
rect 146076 182420 146128 182426
rect 146076 182362 146128 182368
rect 148940 182358 148968 184876
rect 144880 182352 144932 182358
rect 144880 182294 144932 182300
rect 148928 182352 148980 182358
rect 148928 182294 148980 182300
rect 144696 181400 144748 181406
rect 144696 181342 144748 181348
rect 144892 175778 144920 182294
rect 150412 182290 150440 184876
rect 146076 182284 146128 182290
rect 146076 182226 146128 182232
rect 150400 182284 150452 182290
rect 150400 182226 150452 182232
rect 146088 175778 146116 182226
rect 151792 181882 151820 184876
rect 147180 181876 147232 181882
rect 147180 181818 147232 181824
rect 151780 181876 151832 181882
rect 151780 181818 151832 181824
rect 147192 175778 147220 181818
rect 153264 181474 153292 184876
rect 148284 181468 148336 181474
rect 148284 181410 148336 181416
rect 153252 181468 153304 181474
rect 153252 181410 153304 181416
rect 148296 175778 148324 181410
rect 153896 178068 153948 178074
rect 153896 178010 153948 178016
rect 151688 178000 151740 178006
rect 151688 177942 151740 177948
rect 148834 177288 148890 177297
rect 148834 177223 148890 177232
rect 124560 175750 124712 175778
rect 125480 175750 125816 175778
rect 126676 175750 126920 175778
rect 127688 175750 128024 175778
rect 128792 175750 129128 175778
rect 129988 175750 130232 175778
rect 131276 175750 131336 175778
rect 132440 175750 132684 175778
rect 133544 175750 133972 175778
rect 134648 175750 134984 175778
rect 135844 175750 136180 175778
rect 136948 175750 137284 175778
rect 138052 175750 138204 175778
rect 139156 175750 139492 175778
rect 140260 175750 140596 175778
rect 141364 175750 141700 175778
rect 142468 175750 142804 175778
rect 143572 175750 143724 175778
rect 144676 175750 144920 175778
rect 145780 175750 146116 175778
rect 146884 175750 147220 175778
rect 147988 175750 148324 175778
rect 148848 175778 148876 177223
rect 151700 175778 151728 177942
rect 152792 177592 152844 177598
rect 152792 177534 152844 177540
rect 152804 175778 152832 177534
rect 153908 175778 153936 178010
rect 154632 177796 154684 177802
rect 154632 177738 154684 177744
rect 148848 175750 149184 175778
rect 151392 175750 151728 175778
rect 152496 175750 152832 175778
rect 153600 175750 153936 175778
rect 154644 175778 154672 177738
rect 156104 177660 156156 177666
rect 156104 177602 156156 177608
rect 156116 175778 156144 177602
rect 154644 175750 154704 175778
rect 155808 175750 156144 175778
rect 157496 175642 157524 185558
rect 158864 185548 158916 185554
rect 158864 185490 158916 185496
rect 158220 184120 158272 184126
rect 158220 184062 158272 184068
rect 158232 177666 158260 184062
rect 158312 182760 158364 182766
rect 158312 182702 158364 182708
rect 158324 178006 158352 182702
rect 158312 178000 158364 178006
rect 158312 177942 158364 177948
rect 158876 177666 158904 185490
rect 160164 185185 160192 187559
rect 160242 186944 160298 186953
rect 160348 186930 160376 189327
rect 160426 188168 160482 188177
rect 160426 188103 160482 188112
rect 160298 186902 160376 186930
rect 160242 186879 160298 186888
rect 160440 185842 160468 188103
rect 160978 187080 161034 187089
rect 160978 187015 161034 187024
rect 160518 186536 160574 186545
rect 160518 186471 160574 186480
rect 160256 185814 160468 185842
rect 160256 185729 160284 185814
rect 160242 185720 160298 185729
rect 160242 185655 160298 185664
rect 160532 185554 160560 186471
rect 160610 185992 160666 186001
rect 160610 185927 160666 185936
rect 160624 185622 160652 185927
rect 160612 185616 160664 185622
rect 160612 185558 160664 185564
rect 160520 185548 160572 185554
rect 160520 185490 160572 185496
rect 160334 185312 160390 185321
rect 160334 185247 160390 185256
rect 160150 185176 160206 185185
rect 160150 185111 160206 185120
rect 160348 184126 160376 185247
rect 160336 184120 160388 184126
rect 160336 184062 160388 184068
rect 159598 183680 159654 183689
rect 159598 183615 159654 183624
rect 159416 177728 159468 177734
rect 159416 177670 159468 177676
rect 158220 177660 158272 177666
rect 158220 177602 158272 177608
rect 158312 177660 158364 177666
rect 158312 177602 158364 177608
rect 158864 177660 158916 177666
rect 158864 177602 158916 177608
rect 158324 175778 158352 177602
rect 159428 175778 159456 177670
rect 159612 177598 159640 183615
rect 160334 183136 160390 183145
rect 160334 183071 160390 183080
rect 160348 182766 160376 183071
rect 160336 182760 160388 182766
rect 160336 182702 160388 182708
rect 160992 177734 161020 187015
rect 192088 185593 192116 210378
rect 196950 208976 197006 208985
rect 196950 208911 197006 208920
rect 194742 191160 194798 191169
rect 194742 191095 194798 191104
rect 194756 191062 194784 191095
rect 194744 191056 194796 191062
rect 194744 190998 194796 191004
rect 196860 191056 196912 191062
rect 196860 190998 196912 191004
rect 192074 185584 192130 185593
rect 192074 185519 192130 185528
rect 161254 184768 161310 184777
rect 161254 184703 161310 184712
rect 161070 184224 161126 184233
rect 161070 184159 161126 184168
rect 161084 178074 161112 184159
rect 161072 178068 161124 178074
rect 161072 178010 161124 178016
rect 161072 177864 161124 177870
rect 161072 177806 161124 177812
rect 160980 177728 161032 177734
rect 160980 177670 161032 177676
rect 159600 177592 159652 177598
rect 159600 177534 159652 177540
rect 158016 175750 158352 175778
rect 159120 175750 159456 175778
rect 161084 175778 161112 177806
rect 161268 177802 161296 184703
rect 163108 182822 164134 182850
rect 163108 179910 163136 182822
rect 163188 180992 163240 180998
rect 163188 180934 163240 180940
rect 163096 179904 163148 179910
rect 163096 179846 163148 179852
rect 161256 177796 161308 177802
rect 161256 177738 161308 177744
rect 161084 175750 161328 175778
rect 123088 175614 123608 175642
rect 156912 175614 157524 175642
rect 163200 175257 163228 180934
rect 163280 179904 163332 179910
rect 163280 179846 163332 179852
rect 92622 175248 92678 175257
rect 92622 175183 92678 175192
rect 163186 175248 163242 175257
rect 163186 175183 163242 175192
rect 94554 174568 94610 174577
rect 94554 174503 94610 174512
rect 92346 174024 92402 174033
rect 92346 173959 92402 173968
rect 92624 171744 92676 171750
rect 92624 171686 92676 171692
rect 92254 171576 92310 171585
rect 92254 171511 92310 171520
rect 92070 170352 92126 170361
rect 92070 170287 92126 170296
rect 91978 169128 92034 169137
rect 91978 169063 92034 169072
rect 91704 168956 91756 168962
rect 91704 168898 91756 168904
rect 91426 167904 91482 167913
rect 91426 167839 91482 167848
rect 91334 166680 91390 166689
rect 91334 166615 91390 166624
rect 91716 163153 91744 168898
rect 91980 165896 92032 165902
rect 91980 165838 92032 165844
rect 91992 165465 92020 165838
rect 91978 165456 92034 165465
rect 91978 165391 92034 165400
rect 92636 164241 92664 171686
rect 94568 165902 94596 174503
rect 95014 172256 95070 172265
rect 95014 172191 95070 172200
rect 95028 171750 95056 172191
rect 95016 171744 95068 171750
rect 95016 171686 95068 171692
rect 94830 169944 94886 169953
rect 94830 169879 94886 169888
rect 94844 168962 94872 169879
rect 163188 169160 163240 169166
rect 163186 169128 163188 169137
rect 163240 169128 163242 169137
rect 163186 169063 163242 169072
rect 118934 168992 118990 169001
rect 94832 168956 94884 168962
rect 94832 168898 94884 168904
rect 114060 168956 114112 168962
rect 118934 168927 118936 168936
rect 114060 168898 114112 168904
rect 118988 168927 118990 168936
rect 118936 168898 118988 168904
rect 95382 167496 95438 167505
rect 95382 167431 95438 167440
rect 94556 165896 94608 165902
rect 94556 165838 94608 165844
rect 94186 165184 94242 165193
rect 94186 165119 94242 165128
rect 92622 164232 92678 164241
rect 92622 164167 92678 164176
rect 91702 163144 91758 163153
rect 91702 163079 91758 163088
rect 94094 162872 94150 162881
rect 94094 162807 94150 162816
rect 92624 161952 92676 161958
rect 92622 161920 92624 161929
rect 92676 161920 92678 161929
rect 92622 161855 92678 161864
rect 91980 161204 92032 161210
rect 91980 161146 92032 161152
rect 91992 160705 92020 161146
rect 91978 160696 92034 160705
rect 91978 160631 92034 160640
rect 94108 160598 94136 162807
rect 94200 161210 94228 165119
rect 95396 161958 95424 167431
rect 95384 161952 95436 161958
rect 95384 161894 95436 161900
rect 94188 161204 94240 161210
rect 94188 161146 94240 161152
rect 91980 160592 92032 160598
rect 91980 160534 92032 160540
rect 94096 160592 94148 160598
rect 94096 160534 94148 160540
rect 91992 159481 92020 160534
rect 94002 160424 94058 160433
rect 94002 160359 94058 160368
rect 91978 159472 92034 159481
rect 91978 159407 92034 159416
rect 94016 159238 94044 160359
rect 91980 159232 92032 159238
rect 91980 159174 92032 159180
rect 94004 159232 94056 159238
rect 94004 159174 94056 159180
rect 91992 158257 92020 159174
rect 91978 158248 92034 158257
rect 91978 158183 92034 158192
rect 94002 158112 94058 158121
rect 94002 158047 94058 158056
rect 94016 157266 94044 158047
rect 91796 157260 91848 157266
rect 91796 157202 91848 157208
rect 94004 157260 94056 157266
rect 94004 157202 94056 157208
rect 91808 157033 91836 157202
rect 91794 157024 91850 157033
rect 91794 156959 91850 156968
rect 91426 154576 91482 154585
rect 91426 154511 91482 154520
rect 91440 154138 91468 154511
rect 91428 154132 91480 154138
rect 91428 154074 91480 154080
rect 94740 154132 94792 154138
rect 94740 154074 94792 154080
rect 94752 153497 94780 154074
rect 94738 153488 94794 153497
rect 94738 153423 94794 153432
rect 91794 153352 91850 153361
rect 91794 153287 91850 153296
rect 91808 152574 91836 153287
rect 91796 152568 91848 152574
rect 91796 152510 91848 152516
rect 95384 152568 95436 152574
rect 95384 152510 95436 152516
rect 91702 152128 91758 152137
rect 91702 152063 91758 152072
rect 91716 151622 91744 152063
rect 91704 151616 91756 151622
rect 91704 151558 91756 151564
rect 94188 151616 94240 151622
rect 94188 151558 94240 151564
rect 91426 150904 91482 150913
rect 91426 150839 91482 150848
rect 91334 149816 91390 149825
rect 91334 149751 91390 149760
rect 91348 143598 91376 149751
rect 91440 149650 91468 150839
rect 91428 149644 91480 149650
rect 91428 149586 91480 149592
rect 94004 149644 94056 149650
rect 94004 149586 94056 149592
rect 91702 148592 91758 148601
rect 91702 148527 91758 148536
rect 91426 147368 91482 147377
rect 91426 147303 91482 147312
rect 91440 146862 91468 147303
rect 91428 146856 91480 146862
rect 91428 146798 91480 146804
rect 91336 143592 91388 143598
rect 91336 143534 91388 143540
rect 91716 142714 91744 148527
rect 93544 146856 93596 146862
rect 93544 146798 93596 146804
rect 93358 146144 93414 146153
rect 93358 146079 93414 146088
rect 91978 144920 92034 144929
rect 91978 144855 92034 144864
rect 91794 143696 91850 143705
rect 91794 143631 91850 143640
rect 91808 142782 91836 143631
rect 91796 142776 91848 142782
rect 91796 142718 91848 142724
rect 91704 142708 91756 142714
rect 91704 142650 91756 142656
rect 91794 142472 91850 142481
rect 91794 142407 91850 142416
rect 91702 141792 91758 141801
rect 91702 141727 91758 141736
rect 91716 141490 91744 141727
rect 91704 141484 91756 141490
rect 91704 141426 91756 141432
rect 91808 141354 91836 142407
rect 91796 141348 91848 141354
rect 91796 141290 91848 141296
rect 53274 135902 54024 135930
rect 48464 134752 48516 134758
rect 48464 134694 48516 134700
rect 47452 133120 47504 133126
rect 47452 133062 47504 133068
rect 46072 131420 46124 131426
rect 46072 131362 46124 131368
rect 44416 130944 44468 130950
rect 44416 130886 44468 130892
rect 43036 130468 43088 130474
rect 43036 130410 43088 130416
rect 45428 130468 45480 130474
rect 45428 130410 45480 130416
rect 44692 130400 44744 130406
rect 42956 130326 43076 130354
rect 44692 130342 44744 130348
rect 43048 128722 43076 130326
rect 44048 130332 44100 130338
rect 44048 130274 44100 130280
rect 43048 128694 43430 128722
rect 44060 128708 44088 130274
rect 44704 128708 44732 130342
rect 45440 128708 45468 130410
rect 46084 128708 46112 131362
rect 46808 131148 46860 131154
rect 46808 131090 46860 131096
rect 46820 128708 46848 131090
rect 47464 128708 47492 133062
rect 51222 128192 51278 128201
rect 51278 128150 51356 128178
rect 51222 128127 51278 128136
rect 51328 127113 51356 128150
rect 51406 127648 51462 127657
rect 51406 127583 51462 127592
rect 51314 127104 51370 127113
rect 51314 127039 51370 127048
rect 51222 126968 51278 126977
rect 51278 126926 51356 126954
rect 51222 126903 51278 126912
rect 51222 126152 51278 126161
rect 51222 126087 51278 126096
rect 51236 125594 51264 126087
rect 51328 125753 51356 126926
rect 51420 125889 51448 127583
rect 51498 126424 51554 126433
rect 51498 126359 51554 126368
rect 51406 125880 51462 125889
rect 51406 125815 51462 125824
rect 51314 125744 51370 125753
rect 51314 125679 51370 125688
rect 51236 125566 51356 125594
rect 51222 125200 51278 125209
rect 51222 125135 51278 125144
rect 51236 124370 51264 125135
rect 51328 124529 51356 125566
rect 51406 124792 51462 124801
rect 51406 124727 51462 124736
rect 51314 124520 51370 124529
rect 51314 124455 51370 124464
rect 51236 124342 51356 124370
rect 51222 124112 51278 124121
rect 51222 124047 51278 124056
rect 51236 123826 51264 124047
rect 51328 123985 51356 124342
rect 51314 123976 51370 123985
rect 51314 123911 51370 123920
rect 51236 123798 51356 123826
rect 18102 123568 18158 123577
rect 18102 123503 18158 123512
rect 18010 114184 18066 114193
rect 18010 114119 18066 114128
rect 18024 101302 18052 114119
rect 18012 101296 18064 101302
rect 18012 101238 18064 101244
rect 18116 90218 18144 123503
rect 51328 123146 51356 123798
rect 51420 123305 51448 124727
rect 51512 124665 51540 126359
rect 51498 124656 51554 124665
rect 51498 124591 51554 124600
rect 51498 123568 51554 123577
rect 51498 123503 51554 123512
rect 51406 123296 51462 123305
rect 51406 123231 51462 123240
rect 51328 123118 51448 123146
rect 51314 122888 51370 122897
rect 51314 122823 51370 122832
rect 51328 121537 51356 122823
rect 51420 122761 51448 123118
rect 51406 122752 51462 122761
rect 51406 122687 51462 122696
rect 51406 122072 51462 122081
rect 51406 122007 51462 122016
rect 51314 121528 51370 121537
rect 51314 121463 51370 121472
rect 51222 120712 51278 120721
rect 51278 120670 51356 120698
rect 51222 120647 51278 120656
rect 51222 120032 51278 120041
rect 51222 119967 51278 119976
rect 51130 119352 51186 119361
rect 51130 119287 51132 119296
rect 51184 119287 51186 119296
rect 51132 119258 51184 119264
rect 51236 118930 51264 119967
rect 51328 119089 51356 120670
rect 51420 120313 51448 122007
rect 51512 121673 51540 123503
rect 51774 122344 51830 122353
rect 51774 122279 51830 122288
rect 51498 121664 51554 121673
rect 51498 121599 51554 121608
rect 51498 121120 51554 121129
rect 51498 121055 51554 121064
rect 51406 120304 51462 120313
rect 51406 120239 51462 120248
rect 51406 119488 51462 119497
rect 51406 119423 51462 119432
rect 51314 119080 51370 119089
rect 51314 119015 51370 119024
rect 51236 118902 51356 118930
rect 51328 118545 51356 118902
rect 51314 118536 51370 118545
rect 51314 118471 51370 118480
rect 51222 118264 51278 118273
rect 51278 118222 51356 118250
rect 51222 118199 51278 118208
rect 51328 117706 51356 118222
rect 51420 117865 51448 119423
rect 51512 119225 51540 121055
rect 51788 120449 51816 122279
rect 51774 120440 51830 120449
rect 51774 120375 51830 120384
rect 51592 119316 51644 119322
rect 51592 119258 51644 119264
rect 51498 119216 51554 119225
rect 51498 119151 51554 119160
rect 51498 117992 51554 118001
rect 51498 117927 51554 117936
rect 51406 117856 51462 117865
rect 51406 117791 51462 117800
rect 51328 117678 51448 117706
rect 50578 117040 50634 117049
rect 50578 116975 50634 116984
rect 50592 116534 50620 116975
rect 50580 116528 50632 116534
rect 50580 116470 50632 116476
rect 51222 116496 51278 116505
rect 51278 116454 51356 116482
rect 51222 116431 51278 116440
rect 51222 115952 51278 115961
rect 51222 115887 51278 115896
rect 51236 114850 51264 115887
rect 51328 115009 51356 116454
rect 51420 116233 51448 117678
rect 51406 116224 51462 116233
rect 51406 116159 51462 116168
rect 51512 116097 51540 117927
rect 51604 117321 51632 119258
rect 51590 117312 51646 117321
rect 51590 117247 51646 117256
rect 51592 116528 51644 116534
rect 51592 116470 51644 116476
rect 51498 116088 51554 116097
rect 51498 116023 51554 116032
rect 51604 115553 51632 116470
rect 51590 115544 51646 115553
rect 51590 115479 51646 115488
rect 51406 115408 51462 115417
rect 51406 115343 51462 115352
rect 51314 115000 51370 115009
rect 51314 114935 51370 114944
rect 51236 114822 51356 114850
rect 51328 114329 51356 114822
rect 51314 114320 51370 114329
rect 51314 114255 51370 114264
rect 51314 114184 51370 114193
rect 51314 114119 51370 114128
rect 51222 112960 51278 112969
rect 51222 112895 51278 112904
rect 51236 112130 51264 112895
rect 51328 112289 51356 114119
rect 51420 113649 51448 115343
rect 51498 115136 51554 115145
rect 51498 115071 51554 115080
rect 51406 113640 51462 113649
rect 51406 113575 51462 113584
rect 51512 113105 51540 115071
rect 51590 113776 51646 113785
rect 51590 113711 51646 113720
rect 51498 113096 51554 113105
rect 51498 113031 51554 113040
rect 51498 112552 51554 112561
rect 51498 112487 51554 112496
rect 51314 112280 51370 112289
rect 51314 112215 51370 112224
rect 51236 112102 51356 112130
rect 51222 111872 51278 111881
rect 51222 111807 51278 111816
rect 51236 111298 51264 111807
rect 51224 111292 51276 111298
rect 51224 111234 51276 111240
rect 51222 111192 51278 111201
rect 51222 111127 51224 111136
rect 51276 111127 51278 111136
rect 51224 111098 51276 111104
rect 51222 111056 51278 111065
rect 51222 110991 51278 111000
rect 51236 110770 51264 110991
rect 51328 110929 51356 112102
rect 51314 110920 51370 110929
rect 51314 110855 51370 110864
rect 51512 110793 51540 112487
rect 51604 112017 51632 113711
rect 51590 112008 51646 112017
rect 51590 111943 51646 111952
rect 51592 111292 51644 111298
rect 51592 111234 51644 111240
rect 51498 110784 51554 110793
rect 51236 110742 51356 110770
rect 51328 109025 51356 110742
rect 51498 110719 51554 110728
rect 51604 110113 51632 111234
rect 51684 111156 51736 111162
rect 51684 111098 51736 111104
rect 51406 110104 51462 110113
rect 51406 110039 51462 110048
rect 51590 110104 51646 110113
rect 51590 110039 51646 110048
rect 51314 109016 51370 109025
rect 51314 108951 51370 108960
rect 51222 108880 51278 108889
rect 51222 108815 51278 108824
rect 51236 108578 51264 108815
rect 51224 108572 51276 108578
rect 51224 108514 51276 108520
rect 51222 108336 51278 108345
rect 51278 108294 51356 108322
rect 51222 108271 51278 108280
rect 51222 107112 51278 107121
rect 51222 107047 51278 107056
rect 51236 106418 51264 107047
rect 51328 106577 51356 108294
rect 51420 108209 51448 110039
rect 51498 109696 51554 109705
rect 51498 109631 51554 109640
rect 51406 108200 51462 108209
rect 51406 108135 51462 108144
rect 51406 107928 51462 107937
rect 51406 107863 51462 107872
rect 51314 106568 51370 106577
rect 51314 106503 51370 106512
rect 51236 106390 51356 106418
rect 51222 106024 51278 106033
rect 51222 105959 51278 105968
rect 51236 105194 51264 105959
rect 51328 105353 51356 106390
rect 51420 106033 51448 107863
rect 51512 107801 51540 109631
rect 51696 109569 51724 111098
rect 51682 109560 51738 109569
rect 51682 109495 51738 109504
rect 51592 108572 51644 108578
rect 51592 108514 51644 108520
rect 51498 107792 51554 107801
rect 51498 107727 51554 107736
rect 51498 106840 51554 106849
rect 51498 106775 51554 106784
rect 51406 106024 51462 106033
rect 51406 105959 51462 105968
rect 51406 105480 51462 105489
rect 51406 105415 51462 105424
rect 51314 105344 51370 105353
rect 51314 105279 51370 105288
rect 51236 105166 51356 105194
rect 50670 104800 50726 104809
rect 50670 104735 50726 104744
rect 50486 101128 50542 101137
rect 50486 101063 50542 101072
rect 20246 100950 20536 100978
rect 21534 100950 21824 100978
rect 22914 100950 23296 100978
rect 24294 100950 24584 100978
rect 24938 100950 25044 100978
rect 25674 100950 26056 100978
rect 26318 100950 26424 100978
rect 27054 100950 27344 100978
rect 27698 100950 27804 100978
rect 28342 100950 28632 100978
rect 29078 100950 29184 100978
rect 29722 100950 30104 100978
rect 30458 100950 30564 100978
rect 31102 100950 31392 100978
rect 31838 100950 31944 100978
rect 32482 100950 32864 100978
rect 33126 100950 33324 100978
rect 20508 97873 20536 100950
rect 20784 100814 20890 100842
rect 20494 97864 20550 97873
rect 20494 97799 20550 97808
rect 20784 97306 20812 100814
rect 21796 97834 21824 100950
rect 22164 100814 22270 100842
rect 21784 97828 21836 97834
rect 21784 97770 21836 97776
rect 20784 97278 20996 97306
rect 20968 97018 20996 97278
rect 22164 97170 22192 100814
rect 23268 97494 23296 100950
rect 23544 100814 23650 100842
rect 23256 97488 23308 97494
rect 23256 97430 23308 97436
rect 23544 97290 23572 100814
rect 23624 97828 23676 97834
rect 23624 97770 23676 97776
rect 23532 97284 23584 97290
rect 23532 97226 23584 97232
rect 22164 97142 22376 97170
rect 20956 97012 21008 97018
rect 20956 96954 21008 96960
rect 22348 96814 22376 97142
rect 22336 96808 22388 96814
rect 22336 96750 22388 96756
rect 23636 96406 23664 97770
rect 24556 97222 24584 100950
rect 24912 97488 24964 97494
rect 24912 97430 24964 97436
rect 24544 97216 24596 97222
rect 24544 97158 24596 97164
rect 24924 96882 24952 97430
rect 25016 97170 25044 100950
rect 26028 97222 26056 100950
rect 26016 97216 26068 97222
rect 25016 97142 25136 97170
rect 26016 97158 26068 97164
rect 26396 97170 26424 100950
rect 27316 97358 27344 100950
rect 27304 97352 27356 97358
rect 27304 97294 27356 97300
rect 27776 97170 27804 100950
rect 28604 97290 28632 100950
rect 29052 97352 29104 97358
rect 29052 97294 29104 97300
rect 28592 97284 28644 97290
rect 28592 97226 28644 97232
rect 26396 97142 26608 97170
rect 24912 96876 24964 96882
rect 24912 96818 24964 96824
rect 23624 96400 23676 96406
rect 23624 96342 23676 96348
rect 25108 96338 25136 97142
rect 26108 97012 26160 97018
rect 26108 96954 26160 96960
rect 25096 96332 25148 96338
rect 25096 96274 25148 96280
rect 26120 93756 26148 96954
rect 26476 96400 26528 96406
rect 26476 96342 26528 96348
rect 26488 93756 26516 96342
rect 26580 95862 26608 97142
rect 27672 97148 27724 97154
rect 27776 97142 27896 97170
rect 27672 97090 27724 97096
rect 26844 97012 26896 97018
rect 26844 96954 26896 96960
rect 26568 95856 26620 95862
rect 26568 95798 26620 95804
rect 26856 93756 26884 96954
rect 27304 96876 27356 96882
rect 27304 96818 27356 96824
rect 27316 93756 27344 96818
rect 27684 93756 27712 97090
rect 27868 96882 27896 97142
rect 28868 97148 28920 97154
rect 28868 97090 28920 97096
rect 28040 97080 28092 97086
rect 28040 97022 28092 97028
rect 27856 96876 27908 96882
rect 27856 96818 27908 96824
rect 28052 93756 28080 97022
rect 28500 96332 28552 96338
rect 28500 96274 28552 96280
rect 28512 93756 28540 96274
rect 28880 93756 28908 97090
rect 29064 95946 29092 97294
rect 29156 97222 29184 100950
rect 30076 97222 30104 100950
rect 30536 97290 30564 100950
rect 30432 97284 30484 97290
rect 30432 97226 30484 97232
rect 30524 97284 30576 97290
rect 30524 97226 30576 97232
rect 29144 97216 29196 97222
rect 29144 97158 29196 97164
rect 30064 97216 30116 97222
rect 30064 97158 30116 97164
rect 30064 96876 30116 96882
rect 30064 96818 30116 96824
rect 29064 95918 29368 95946
rect 29236 95856 29288 95862
rect 29236 95798 29288 95804
rect 29248 93756 29276 95798
rect 29340 93770 29368 95918
rect 29340 93742 29722 93770
rect 30076 93756 30104 96818
rect 30444 93756 30472 97226
rect 31364 97222 31392 100950
rect 31628 97284 31680 97290
rect 31628 97226 31680 97232
rect 31260 97216 31312 97222
rect 31260 97158 31312 97164
rect 31352 97216 31404 97222
rect 31352 97158 31404 97164
rect 30892 97148 30944 97154
rect 30892 97090 30944 97096
rect 30904 93756 30932 97090
rect 31272 93756 31300 97158
rect 31640 93756 31668 97226
rect 31916 97170 31944 100950
rect 31916 97142 32220 97170
rect 32088 97080 32140 97086
rect 32088 97022 32140 97028
rect 32100 93756 32128 97022
rect 32192 93770 32220 97142
rect 32192 93742 32482 93770
rect 32836 93756 32864 100950
rect 33296 93756 33324 100950
rect 33664 100814 33862 100842
rect 34308 100814 34506 100842
rect 34768 100814 35242 100842
rect 35320 100814 35886 100842
rect 36332 100814 36530 100842
rect 36976 100814 37266 100842
rect 37528 100814 37910 100842
rect 38264 100814 38646 100842
rect 39000 100814 39290 100842
rect 39736 100814 40026 100842
rect 40288 100814 40670 100842
rect 41024 100814 41314 100842
rect 41760 100814 42050 100842
rect 42312 100814 42694 100842
rect 43048 100814 43430 100842
rect 43784 100814 44074 100842
rect 44428 100814 44718 100842
rect 45072 100814 45454 100842
rect 45900 100814 46098 100842
rect 46544 100814 46834 100842
rect 47188 100814 47478 100842
rect 33664 93756 33692 100814
rect 34308 93770 34336 100814
rect 34768 95810 34796 100814
rect 35320 96354 35348 100814
rect 36044 97148 36096 97154
rect 36044 97090 36096 97096
rect 35676 97080 35728 97086
rect 35676 97022 35728 97028
rect 34676 95782 34796 95810
rect 35228 96326 35348 96354
rect 34676 93770 34704 95782
rect 35228 93770 35256 96326
rect 35308 96196 35360 96202
rect 35308 96138 35360 96144
rect 34138 93742 34336 93770
rect 34506 93742 34704 93770
rect 34874 93742 35256 93770
rect 35320 93756 35348 96138
rect 35688 93756 35716 97022
rect 36056 93756 36084 97090
rect 36332 96202 36360 100814
rect 36504 97148 36556 97154
rect 36504 97090 36556 97096
rect 36320 96196 36372 96202
rect 36320 96138 36372 96144
rect 36516 93756 36544 97090
rect 36976 97086 37004 100814
rect 37528 97222 37556 100814
rect 37608 97284 37660 97290
rect 37608 97226 37660 97232
rect 37516 97216 37568 97222
rect 37516 97158 37568 97164
rect 36964 97080 37016 97086
rect 36964 97022 37016 97028
rect 37148 97080 37200 97086
rect 37148 97022 37200 97028
rect 37160 93770 37188 97022
rect 37620 95946 37648 97226
rect 38264 97154 38292 100814
rect 39000 97222 39028 100814
rect 39736 97290 39764 100814
rect 39724 97284 39776 97290
rect 39724 97226 39776 97232
rect 38988 97216 39040 97222
rect 40288 97170 40316 100814
rect 40368 97284 40420 97290
rect 40368 97226 40420 97232
rect 38988 97158 39040 97164
rect 38252 97148 38304 97154
rect 38436 97148 38488 97154
rect 38252 97090 38304 97096
rect 38356 97108 38436 97136
rect 37700 97012 37752 97018
rect 37700 96954 37752 96960
rect 37436 95918 37648 95946
rect 37436 93770 37464 95918
rect 36898 93742 37188 93770
rect 37266 93742 37464 93770
rect 37712 93756 37740 96954
rect 38356 93770 38384 97108
rect 38436 97090 38488 97096
rect 40196 97142 40316 97170
rect 38896 97080 38948 97086
rect 38896 97022 38948 97028
rect 38436 96808 38488 96814
rect 38436 96750 38488 96756
rect 38094 93742 38384 93770
rect 38448 93756 38476 96750
rect 38908 93756 38936 97022
rect 40196 97018 40224 97142
rect 40380 97086 40408 97226
rect 41024 97222 41052 100814
rect 41012 97216 41064 97222
rect 41012 97158 41064 97164
rect 40828 97148 40880 97154
rect 40828 97090 40880 97096
rect 40368 97080 40420 97086
rect 40368 97022 40420 97028
rect 40460 97080 40512 97086
rect 40460 97022 40512 97028
rect 40184 97012 40236 97018
rect 40184 96954 40236 96960
rect 39632 96468 39684 96474
rect 39632 96410 39684 96416
rect 39264 96264 39316 96270
rect 39264 96206 39316 96212
rect 39276 93756 39304 96206
rect 39644 93756 39672 96410
rect 40092 96332 40144 96338
rect 40092 96274 40144 96280
rect 40104 93756 40132 96274
rect 40472 93756 40500 97022
rect 40840 93756 40868 97090
rect 41288 96944 41340 96950
rect 41288 96886 41340 96892
rect 41300 93756 41328 96886
rect 41656 96876 41708 96882
rect 41656 96818 41708 96824
rect 41668 93756 41696 96818
rect 41760 96814 41788 100814
rect 42312 97290 42340 100814
rect 42300 97284 42352 97290
rect 42300 97226 42352 97232
rect 41748 96808 41800 96814
rect 41748 96750 41800 96756
rect 43048 96270 43076 100814
rect 43784 96474 43812 100814
rect 43772 96468 43824 96474
rect 43772 96410 43824 96416
rect 44428 96338 44456 100814
rect 45072 97086 45100 100814
rect 45900 97154 45928 100814
rect 45888 97148 45940 97154
rect 45888 97090 45940 97096
rect 45060 97080 45112 97086
rect 45060 97022 45112 97028
rect 46544 96950 46572 100814
rect 46532 96944 46584 96950
rect 46532 96886 46584 96892
rect 47188 96882 47216 100814
rect 47176 96876 47228 96882
rect 47176 96818 47228 96824
rect 44416 96332 44468 96338
rect 44416 96274 44468 96280
rect 43036 96264 43088 96270
rect 43036 96206 43088 96212
rect 50500 93756 50528 101063
rect 50684 96542 50712 104735
rect 50946 104256 51002 104265
rect 50946 104191 51002 104200
rect 50762 103168 50818 103177
rect 50762 103103 50818 103112
rect 50776 103070 50804 103103
rect 50764 103064 50816 103070
rect 50764 103006 50816 103012
rect 50960 97086 50988 104191
rect 51328 103993 51356 105166
rect 51314 103984 51370 103993
rect 51314 103919 51370 103928
rect 51222 103712 51278 103721
rect 51222 103647 51278 103656
rect 51236 102798 51264 103647
rect 51420 103585 51448 105415
rect 51512 104809 51540 106775
rect 51604 106713 51632 108514
rect 51590 106704 51646 106713
rect 51590 106639 51646 106648
rect 51498 104800 51554 104809
rect 51498 104735 51554 104744
rect 51406 103576 51462 103585
rect 51406 103511 51462 103520
rect 51224 102792 51276 102798
rect 51224 102734 51276 102740
rect 51406 102760 51462 102769
rect 51406 102695 51462 102704
rect 51222 101944 51278 101953
rect 51222 101879 51278 101888
rect 51236 101370 51264 101879
rect 51314 101400 51370 101409
rect 51224 101364 51276 101370
rect 51314 101335 51370 101344
rect 51224 101306 51276 101312
rect 50948 97080 51000 97086
rect 50948 97022 51000 97028
rect 50672 96536 50724 96542
rect 50672 96478 50724 96484
rect 51328 93770 51356 101335
rect 51420 96882 51448 102695
rect 52604 101364 52656 101370
rect 52604 101306 52656 101312
rect 52616 97034 52644 101306
rect 52616 97006 52736 97034
rect 51408 96876 51460 96882
rect 51408 96818 51460 96824
rect 51328 93742 51618 93770
rect 52708 93756 52736 97006
rect 53800 96876 53852 96882
rect 53800 96818 53852 96824
rect 53812 93756 53840 96818
rect 53996 96474 54024 135902
rect 66600 134214 66628 135916
rect 73224 134282 73252 135916
rect 82136 134412 82188 134418
rect 82136 134354 82188 134360
rect 84344 134412 84396 134418
rect 84344 134354 84396 134360
rect 73212 134276 73264 134282
rect 73212 134218 73264 134224
rect 66588 134208 66640 134214
rect 66588 134150 66640 134156
rect 82148 134146 82176 134354
rect 84356 134282 84384 134354
rect 83608 134276 83660 134282
rect 83608 134218 83660 134224
rect 84344 134276 84396 134282
rect 84344 134218 84396 134224
rect 82136 134140 82188 134146
rect 82136 134082 82188 134088
rect 62356 133732 62408 133738
rect 62356 133674 62408 133680
rect 62368 126804 62396 133674
rect 82148 133097 82176 134082
rect 83620 133097 83648 134218
rect 86564 133738 86592 135916
rect 86552 133732 86604 133738
rect 86552 133674 86604 133680
rect 82134 133088 82190 133097
rect 82134 133023 82190 133032
rect 83606 133088 83662 133097
rect 83606 133023 83662 133032
rect 91992 131154 92020 144855
rect 92530 141248 92586 141257
rect 92530 141183 92586 141192
rect 92544 140062 92572 141183
rect 92532 140056 92584 140062
rect 92532 139998 92584 140004
rect 92622 140024 92678 140033
rect 92622 139959 92624 139968
rect 92676 139959 92678 139968
rect 92624 139930 92676 139936
rect 93266 138800 93322 138809
rect 93266 138735 93322 138744
rect 92070 137576 92126 137585
rect 92070 137511 92126 137520
rect 92084 131630 92112 137511
rect 92162 136488 92218 136497
rect 92162 136423 92218 136432
rect 92072 131624 92124 131630
rect 92072 131566 92124 131572
rect 91980 131148 92032 131154
rect 91980 131090 92032 131096
rect 92176 128708 92204 136423
rect 92716 131624 92768 131630
rect 92716 131566 92768 131572
rect 92728 128708 92756 131566
rect 93280 128708 93308 138735
rect 93372 137041 93400 146079
rect 93452 140056 93504 140062
rect 93452 139998 93504 140004
rect 93358 137032 93414 137041
rect 93358 136967 93414 136976
rect 93464 131630 93492 139998
rect 93556 138673 93584 146798
rect 94016 145609 94044 149586
rect 94200 148737 94228 151558
rect 95396 151049 95424 152510
rect 95382 151040 95438 151049
rect 95382 150975 95438 150984
rect 94186 148728 94242 148737
rect 94186 148663 94242 148672
rect 94002 145600 94058 145609
rect 94002 145535 94058 145544
rect 94370 143968 94426 143977
rect 94370 143903 94426 143912
rect 94384 143598 94412 143903
rect 94372 143592 94424 143598
rect 94372 143534 94424 143540
rect 95660 142776 95712 142782
rect 95660 142718 95712 142724
rect 95384 142708 95436 142714
rect 95384 142650 95436 142656
rect 95396 141665 95424 142650
rect 95382 141656 95438 141665
rect 95382 141591 95438 141600
rect 95016 141348 95068 141354
rect 95016 141290 95068 141296
rect 93912 139988 93964 139994
rect 93912 139930 93964 139936
rect 93542 138664 93598 138673
rect 93542 138599 93598 138608
rect 93452 131624 93504 131630
rect 93452 131566 93504 131572
rect 93924 128708 93952 139930
rect 94464 131624 94516 131630
rect 94464 131566 94516 131572
rect 94476 128708 94504 131566
rect 95028 128708 95056 141290
rect 95672 128708 95700 142718
rect 97788 135902 98124 135930
rect 98248 135902 98492 135930
rect 98616 135902 98860 135930
rect 98984 135902 99320 135930
rect 97788 133126 97816 135902
rect 96764 133120 96816 133126
rect 96764 133062 96816 133068
rect 97776 133120 97828 133126
rect 97776 133062 97828 133068
rect 97960 133120 98012 133126
rect 97960 133062 98012 133068
rect 96212 131148 96264 131154
rect 96212 131090 96264 131096
rect 96224 128708 96252 131090
rect 96776 128708 96804 133062
rect 97408 133052 97460 133058
rect 97408 132994 97460 133000
rect 97420 128708 97448 132994
rect 97972 128708 98000 133062
rect 98248 133058 98276 135902
rect 98616 133126 98644 135902
rect 98604 133120 98656 133126
rect 98604 133062 98656 133068
rect 98236 133052 98288 133058
rect 98236 132994 98288 133000
rect 98984 128722 99012 135902
rect 99674 135658 99702 135916
rect 99628 135630 99702 135658
rect 99904 135902 100056 135930
rect 100272 135902 100516 135930
rect 99628 133754 99656 135630
rect 99536 133726 99656 133754
rect 99536 128722 99564 133726
rect 99904 128722 99932 135902
rect 98538 128694 99012 128722
rect 99182 128694 99564 128722
rect 99734 128694 99932 128722
rect 100272 128708 100300 135902
rect 100870 135658 100898 135916
rect 101252 135902 101496 135930
rect 101712 135902 101864 135930
rect 102080 135902 102324 135930
rect 102448 135902 102784 135930
rect 102908 135902 103152 135930
rect 103276 135902 103520 135930
rect 100870 135630 100944 135658
rect 100916 128708 100944 135630
rect 101468 128708 101496 135902
rect 101836 128722 101864 135902
rect 102296 133074 102324 135902
rect 102296 133046 102416 133074
rect 102388 128722 102416 133046
rect 102756 128994 102784 135902
rect 103124 133058 103152 135902
rect 103492 133126 103520 135902
rect 103630 135658 103658 135916
rect 104104 135902 104348 135930
rect 104472 135902 104716 135930
rect 104840 135902 105084 135930
rect 105300 135902 105544 135930
rect 105668 135902 106004 135930
rect 106128 135902 106372 135930
rect 106496 135902 106740 135930
rect 106864 135902 107200 135930
rect 107324 135902 107568 135930
rect 107692 135902 107844 135930
rect 108060 135902 108396 135930
rect 108520 135902 108764 135930
rect 108888 135902 109040 135930
rect 109256 135902 109592 135930
rect 109716 135902 109960 135930
rect 110084 135902 110328 135930
rect 103584 135630 103658 135658
rect 103584 133194 103612 135630
rect 103572 133188 103624 133194
rect 103572 133130 103624 133136
rect 103480 133120 103532 133126
rect 103480 133062 103532 133068
rect 104320 133058 104348 135902
rect 104688 133126 104716 135902
rect 105056 133194 105084 135902
rect 105516 133262 105544 135902
rect 105504 133256 105556 133262
rect 105504 133198 105556 133204
rect 104952 133188 105004 133194
rect 104952 133130 105004 133136
rect 105044 133188 105096 133194
rect 105044 133130 105096 133136
rect 104400 133120 104452 133126
rect 104400 133062 104452 133068
rect 104676 133120 104728 133126
rect 104676 133062 104728 133068
rect 103112 133052 103164 133058
rect 103112 132994 103164 133000
rect 103756 133052 103808 133058
rect 103756 132994 103808 133000
rect 104308 133052 104360 133058
rect 104308 132994 104360 133000
rect 102756 128966 102876 128994
rect 102848 128722 102876 128966
rect 101836 128694 102034 128722
rect 102388 128694 102678 128722
rect 102848 128694 103230 128722
rect 103768 128708 103796 132994
rect 104412 128708 104440 133062
rect 104964 128708 104992 133130
rect 105976 133058 106004 135902
rect 106344 133126 106372 135902
rect 106712 133330 106740 135902
rect 107172 133466 107200 135902
rect 107540 133942 107568 135902
rect 107528 133936 107580 133942
rect 107528 133878 107580 133884
rect 107160 133460 107212 133466
rect 107160 133402 107212 133408
rect 107816 133398 107844 135902
rect 108368 133670 108396 135902
rect 108356 133664 108408 133670
rect 108356 133606 108408 133612
rect 108736 133534 108764 135902
rect 109012 133806 109040 135902
rect 109000 133800 109052 133806
rect 109000 133742 109052 133748
rect 108724 133528 108776 133534
rect 108724 133470 108776 133476
rect 107804 133392 107856 133398
rect 107804 133334 107856 133340
rect 106700 133324 106752 133330
rect 106700 133266 106752 133272
rect 109000 133324 109052 133330
rect 109000 133266 109052 133272
rect 107252 133256 107304 133262
rect 107252 133198 107304 133204
rect 106700 133188 106752 133194
rect 106700 133130 106752 133136
rect 106148 133120 106200 133126
rect 106148 133062 106200 133068
rect 106332 133120 106384 133126
rect 106332 133062 106384 133068
rect 105504 133052 105556 133058
rect 105504 132994 105556 133000
rect 105964 133052 106016 133058
rect 105964 132994 106016 133000
rect 105516 128708 105544 132994
rect 106160 128708 106188 133062
rect 106712 128708 106740 133130
rect 107264 128708 107292 133198
rect 108448 133120 108500 133126
rect 108448 133062 108500 133068
rect 107896 133052 107948 133058
rect 107896 132994 107948 133000
rect 107908 128708 107936 132994
rect 108460 128708 108488 133062
rect 109012 128708 109040 133266
rect 109564 133058 109592 135902
rect 109932 133602 109960 135902
rect 110196 133936 110248 133942
rect 110196 133878 110248 133884
rect 109920 133596 109972 133602
rect 109920 133538 109972 133544
rect 109644 133460 109696 133466
rect 109644 133402 109696 133408
rect 109552 133052 109604 133058
rect 109552 132994 109604 133000
rect 109656 128708 109684 133402
rect 110208 128708 110236 133878
rect 110300 133738 110328 135902
rect 110438 135658 110466 135916
rect 110912 135902 111156 135930
rect 111280 135902 111524 135930
rect 111648 135902 111892 135930
rect 112108 135902 112352 135930
rect 112476 135902 112720 135930
rect 112844 135902 113180 135930
rect 110438 135630 110512 135658
rect 110288 133732 110340 133738
rect 110288 133674 110340 133680
rect 110484 133194 110512 135630
rect 110840 133800 110892 133806
rect 110840 133742 110892 133748
rect 110564 133392 110616 133398
rect 110564 133334 110616 133340
rect 110472 133188 110524 133194
rect 110472 133130 110524 133136
rect 110576 131578 110604 133334
rect 110852 131630 110880 133742
rect 111128 133330 111156 135902
rect 111392 133664 111444 133670
rect 111392 133606 111444 133612
rect 111116 133324 111168 133330
rect 111116 133266 111168 133272
rect 110840 131624 110892 131630
rect 110576 131550 110696 131578
rect 110840 131566 110892 131572
rect 110668 128722 110696 131550
rect 110668 128694 110774 128722
rect 111404 128708 111432 133606
rect 111496 133398 111524 135902
rect 111484 133392 111536 133398
rect 111484 133334 111536 133340
rect 111864 133262 111892 135902
rect 111944 133528 111996 133534
rect 111944 133470 111996 133476
rect 111852 133256 111904 133262
rect 111852 133198 111904 133204
rect 111956 128708 111984 133470
rect 112324 133126 112352 135902
rect 112692 133194 112720 135902
rect 112588 133188 112640 133194
rect 112588 133130 112640 133136
rect 112680 133188 112732 133194
rect 112680 133130 112732 133136
rect 112312 133120 112364 133126
rect 112312 133062 112364 133068
rect 112496 131624 112548 131630
rect 112496 131566 112548 131572
rect 112508 128708 112536 131566
rect 112600 130746 112628 133130
rect 113152 133058 113180 135902
rect 113290 135658 113318 135916
rect 113672 135902 114008 135930
rect 113290 135630 113364 135658
rect 113336 133738 113364 135630
rect 113980 133806 114008 135902
rect 114072 134010 114100 168898
rect 163292 166689 163320 179846
rect 164384 174056 164436 174062
rect 164382 174024 164384 174033
rect 164436 174024 164438 174033
rect 164382 173959 164438 173968
rect 164292 172832 164344 172838
rect 164290 172800 164292 172809
rect 164344 172800 164346 172809
rect 164290 172735 164346 172744
rect 164016 171608 164068 171614
rect 164014 171576 164016 171585
rect 164068 171576 164070 171585
rect 164014 171511 164070 171520
rect 163372 170384 163424 170390
rect 163370 170352 163372 170361
rect 163424 170352 163426 170361
rect 163370 170287 163426 170296
rect 164580 168026 164608 182836
rect 165132 169166 165160 182836
rect 165684 170390 165712 182836
rect 166236 171614 166264 182836
rect 166788 172838 166816 182836
rect 167248 182822 167354 182850
rect 167248 181218 167276 182822
rect 167156 181190 167276 181218
rect 167156 174062 167184 181190
rect 167892 180998 167920 182836
rect 168444 181202 168472 182836
rect 168996 181270 169024 182836
rect 168984 181264 169036 181270
rect 168984 181206 169036 181212
rect 168432 181196 168484 181202
rect 168432 181138 168484 181144
rect 167880 180992 167932 180998
rect 167880 180934 167932 180940
rect 168524 180652 168576 180658
rect 168524 180594 168576 180600
rect 168536 174849 168564 180594
rect 169548 180182 169576 182836
rect 170008 182822 170114 182850
rect 169536 180176 169588 180182
rect 169536 180118 169588 180124
rect 170008 177666 170036 182822
rect 170456 181264 170508 181270
rect 170456 181206 170508 181212
rect 170088 181196 170140 181202
rect 170088 181138 170140 181144
rect 169996 177660 170048 177666
rect 169996 177602 170048 177608
rect 170100 175764 170128 181138
rect 170468 175764 170496 181206
rect 170652 180046 170680 182836
rect 170824 180176 170876 180182
rect 170824 180118 170876 180124
rect 170640 180040 170692 180046
rect 170640 179982 170692 179988
rect 170836 175764 170864 180118
rect 171204 179978 171232 182836
rect 171652 180040 171704 180046
rect 171652 179982 171704 179988
rect 171192 179972 171244 179978
rect 171192 179914 171244 179920
rect 171284 177660 171336 177666
rect 171284 177602 171336 177608
rect 171296 175764 171324 177602
rect 171664 175764 171692 179982
rect 171756 177258 171784 182836
rect 172322 182822 172612 182850
rect 172584 181218 172612 182822
rect 172584 181190 172796 181218
rect 172020 179972 172072 179978
rect 172020 179914 172072 179920
rect 171744 177252 171796 177258
rect 171744 177194 171796 177200
rect 172032 175764 172060 179914
rect 172480 177252 172532 177258
rect 172480 177194 172532 177200
rect 172492 175764 172520 177194
rect 172768 175778 172796 181190
rect 172860 177666 172888 182836
rect 172848 177660 172900 177666
rect 172848 177602 172900 177608
rect 173216 177660 173268 177666
rect 173216 177602 173268 177608
rect 172768 175750 172874 175778
rect 173228 175764 173256 177602
rect 173412 175778 173440 182836
rect 173964 175778 173992 182836
rect 174516 175778 174544 182836
rect 175068 175778 175096 182836
rect 175620 181218 175648 182836
rect 175700 181400 175752 181406
rect 175700 181342 175752 181348
rect 175436 181190 175648 181218
rect 175436 175778 175464 181190
rect 175608 177660 175660 177666
rect 175608 177602 175660 177608
rect 173412 175750 173702 175778
rect 173964 175750 174070 175778
rect 174438 175750 174544 175778
rect 174898 175750 175096 175778
rect 175266 175750 175464 175778
rect 175620 175764 175648 177602
rect 175712 175778 175740 181342
rect 176172 177666 176200 182836
rect 176448 182822 176738 182850
rect 176448 181406 176476 182822
rect 176436 181400 176488 181406
rect 176436 181342 176488 181348
rect 177276 181270 177304 182836
rect 176436 181264 176488 181270
rect 176436 181206 176488 181212
rect 177264 181264 177316 181270
rect 177264 181206 177316 181212
rect 177540 181264 177592 181270
rect 177540 181206 177592 181212
rect 176160 177660 176212 177666
rect 176160 177602 176212 177608
rect 175712 175750 176094 175778
rect 176448 175764 176476 181206
rect 176804 181196 176856 181202
rect 176804 181138 176856 181144
rect 176816 175764 176844 181138
rect 177552 175778 177580 181206
rect 177828 181202 177856 182836
rect 178288 181270 178316 182836
rect 178276 181264 178328 181270
rect 178276 181206 178328 181212
rect 177816 181196 177868 181202
rect 177816 181138 177868 181144
rect 178092 181196 178144 181202
rect 178092 181138 178144 181144
rect 177632 181128 177684 181134
rect 177632 181070 177684 181076
rect 177290 175750 177580 175778
rect 177644 175764 177672 181070
rect 178104 175764 178132 181138
rect 178840 181134 178868 182836
rect 179104 181264 179156 181270
rect 179104 181206 179156 181212
rect 178828 181128 178880 181134
rect 178828 181070 178880 181076
rect 178460 180584 178512 180590
rect 178460 180526 178512 180532
rect 178472 175764 178500 180526
rect 179116 175778 179144 181206
rect 179392 181202 179420 182836
rect 179380 181196 179432 181202
rect 179380 181138 179432 181144
rect 179944 180590 179972 182836
rect 180496 181270 180524 182836
rect 180484 181264 180536 181270
rect 180484 181206 180536 181212
rect 180852 180992 180904 180998
rect 180852 180934 180904 180940
rect 179932 180584 179984 180590
rect 179932 180526 179984 180532
rect 179288 180176 179340 180182
rect 179288 180118 179340 180124
rect 178854 175750 179144 175778
rect 179300 175764 179328 180118
rect 180760 180108 180812 180114
rect 180760 180050 180812 180056
rect 179656 180040 179708 180046
rect 179656 179982 179708 179988
rect 179668 175764 179696 179982
rect 180024 179972 180076 179978
rect 180024 179914 180076 179920
rect 180036 175764 180064 179914
rect 180772 175778 180800 180050
rect 180510 175750 180800 175778
rect 180864 175764 180892 180934
rect 181048 180182 181076 182836
rect 181220 181128 181272 181134
rect 181220 181070 181272 181076
rect 181036 180176 181088 180182
rect 181036 180118 181088 180124
rect 181232 175764 181260 181070
rect 181600 180046 181628 182836
rect 181680 180924 181732 180930
rect 181680 180866 181732 180872
rect 181588 180040 181640 180046
rect 181588 179982 181640 179988
rect 181692 175764 181720 180866
rect 182048 180788 182100 180794
rect 182048 180730 182100 180736
rect 182060 175764 182088 180730
rect 182152 179978 182180 182836
rect 182416 181196 182468 181202
rect 182416 181138 182468 181144
rect 182140 179972 182192 179978
rect 182140 179914 182192 179920
rect 182428 175764 182456 181138
rect 182704 180114 182732 182836
rect 182876 181264 182928 181270
rect 182876 181206 182928 181212
rect 182692 180108 182744 180114
rect 182692 180050 182744 180056
rect 182888 175764 182916 181206
rect 183256 180998 183284 182836
rect 183808 181134 183836 182836
rect 183796 181128 183848 181134
rect 183796 181070 183848 181076
rect 183612 181060 183664 181066
rect 183612 181002 183664 181008
rect 183244 180992 183296 180998
rect 183244 180934 183296 180940
rect 183244 180856 183296 180862
rect 183244 180798 183296 180804
rect 183256 175764 183284 180798
rect 183624 175764 183652 181002
rect 184360 180930 184388 182836
rect 184348 180924 184400 180930
rect 184348 180866 184400 180872
rect 184912 180794 184940 182836
rect 185464 181202 185492 182836
rect 186016 181270 186044 182836
rect 186004 181264 186056 181270
rect 186004 181206 186056 181212
rect 185452 181196 185504 181202
rect 185452 181138 185504 181144
rect 186568 180862 186596 182836
rect 187120 181066 187148 182836
rect 187108 181060 187160 181066
rect 187108 181002 187160 181008
rect 186556 180856 186608 180862
rect 186556 180798 186608 180804
rect 184900 180788 184952 180794
rect 184900 180730 184952 180736
rect 187672 180114 187700 182836
rect 184072 180108 184124 180114
rect 184072 180050 184124 180056
rect 187660 180108 187712 180114
rect 187660 180050 187712 180056
rect 184084 175764 184112 180050
rect 185268 177728 185320 177734
rect 185268 177670 185320 177676
rect 184440 177660 184492 177666
rect 184440 177602 184492 177608
rect 184452 175764 184480 177602
rect 184808 177456 184860 177462
rect 184808 177398 184860 177404
rect 184820 175764 184848 177398
rect 185280 175764 185308 177670
rect 188224 177666 188252 182836
rect 188212 177660 188264 177666
rect 188212 177602 188264 177608
rect 185636 177592 185688 177598
rect 185636 177534 185688 177540
rect 185648 175764 185676 177534
rect 188776 177462 188804 182836
rect 189328 177734 189356 182836
rect 189316 177728 189368 177734
rect 189316 177670 189368 177676
rect 189880 177598 189908 182836
rect 190432 180658 190460 182836
rect 190984 181338 191012 182836
rect 190972 181332 191024 181338
rect 190972 181274 191024 181280
rect 190420 180652 190472 180658
rect 190420 180594 190472 180600
rect 189868 177592 189920 177598
rect 189868 177534 189920 177540
rect 188764 177456 188816 177462
rect 188764 177398 188816 177404
rect 168522 174840 168578 174849
rect 168522 174775 168578 174784
rect 167144 174056 167196 174062
rect 167144 173998 167196 174004
rect 188028 173036 188080 173042
rect 188028 172978 188080 172984
rect 166776 172832 166828 172838
rect 166776 172774 166828 172780
rect 188040 172537 188068 172978
rect 188026 172528 188082 172537
rect 188026 172463 188082 172472
rect 166224 171608 166276 171614
rect 166224 171550 166276 171556
rect 167510 170488 167566 170497
rect 167510 170423 167566 170432
rect 165672 170384 165724 170390
rect 165672 170326 165724 170332
rect 165120 169160 165172 169166
rect 165120 169102 165172 169108
rect 167326 168176 167382 168185
rect 167326 168111 167382 168120
rect 164396 167998 164608 168026
rect 164396 167913 164424 167998
rect 164382 167904 164438 167913
rect 164382 167839 164438 167848
rect 163278 166680 163334 166689
rect 163278 166615 163334 166624
rect 167234 166272 167290 166281
rect 167234 166207 167290 166216
rect 163188 165964 163240 165970
rect 163188 165906 163240 165912
rect 163200 165465 163228 165906
rect 163186 165456 163242 165465
rect 163186 165391 163242 165400
rect 116542 165184 116598 165193
rect 116542 165119 116598 165128
rect 116556 164814 116584 165119
rect 116544 164808 116596 164814
rect 116544 164750 116596 164756
rect 119580 164808 119632 164814
rect 119580 164750 119632 164756
rect 119592 155945 119620 164750
rect 164292 164400 164344 164406
rect 164292 164342 164344 164348
rect 164304 164241 164332 164342
rect 164290 164232 164346 164241
rect 164290 164167 164346 164176
rect 167248 163182 167276 166207
rect 167340 164406 167368 168111
rect 167524 165970 167552 170423
rect 167512 165964 167564 165970
rect 167512 165906 167564 165912
rect 188026 165864 188082 165873
rect 188026 165799 188082 165808
rect 188040 164814 188068 165799
rect 188028 164808 188080 164814
rect 188028 164750 188080 164756
rect 167328 164400 167380 164406
rect 167328 164342 167380 164348
rect 167970 164096 168026 164105
rect 167970 164031 168026 164040
rect 164292 163176 164344 163182
rect 164290 163144 164292 163153
rect 167236 163176 167288 163182
rect 164344 163144 164346 163153
rect 167236 163118 167288 163124
rect 164290 163079 164346 163088
rect 164476 162156 164528 162162
rect 164476 162098 164528 162104
rect 164292 161952 164344 161958
rect 164290 161920 164292 161929
rect 164344 161920 164346 161929
rect 164290 161855 164346 161864
rect 164382 160696 164438 160705
rect 164488 160682 164516 162098
rect 167984 161958 168012 164031
rect 168430 162192 168486 162201
rect 168430 162127 168432 162136
rect 168484 162127 168486 162136
rect 168432 162098 168484 162104
rect 167972 161952 168024 161958
rect 167972 161894 168024 161900
rect 168522 160832 168578 160841
rect 168522 160767 168578 160776
rect 164438 160654 164516 160682
rect 168536 160666 168564 160767
rect 168524 160660 168576 160666
rect 164382 160631 164438 160640
rect 168524 160602 168576 160608
rect 164292 160592 164344 160598
rect 164292 160534 164344 160540
rect 164304 159481 164332 160534
rect 164290 159472 164346 159481
rect 164290 159407 164346 159416
rect 168522 158520 168578 158529
rect 168522 158455 168578 158464
rect 168536 158286 168564 158455
rect 164292 158280 164344 158286
rect 164290 158248 164292 158257
rect 168524 158280 168576 158286
rect 164344 158248 164346 158257
rect 168524 158222 168576 158228
rect 164290 158183 164346 158192
rect 164290 157024 164346 157033
rect 164290 156959 164292 156968
rect 164344 156959 164346 156968
rect 168524 156988 168576 156994
rect 164292 156930 164344 156936
rect 168524 156930 168576 156936
rect 168536 156897 168564 156930
rect 168522 156888 168578 156897
rect 168522 156823 168578 156832
rect 119578 155936 119634 155945
rect 119578 155871 119634 155880
rect 164382 155800 164438 155809
rect 164382 155735 164438 155744
rect 164396 155362 164424 155735
rect 164384 155356 164436 155362
rect 164384 155298 164436 155304
rect 167144 155356 167196 155362
rect 167144 155298 167196 155304
rect 167156 154857 167184 155298
rect 167142 154848 167198 154857
rect 167142 154783 167198 154792
rect 163370 154576 163426 154585
rect 163370 154511 163372 154520
rect 163424 154511 163426 154520
rect 167144 154540 167196 154546
rect 163372 154482 163424 154488
rect 167144 154482 167196 154488
rect 164382 153352 164438 153361
rect 164382 153287 164438 153296
rect 164396 152438 164424 153287
rect 167156 152817 167184 154482
rect 167142 152808 167198 152817
rect 167142 152743 167198 152752
rect 164384 152432 164436 152438
rect 164384 152374 164436 152380
rect 167236 152432 167288 152438
rect 167236 152374 167288 152380
rect 164382 152128 164438 152137
rect 164382 152063 164438 152072
rect 164396 151554 164424 152063
rect 164384 151548 164436 151554
rect 164384 151490 164436 151496
rect 163922 150904 163978 150913
rect 163922 150839 163978 150848
rect 163936 149650 163964 150839
rect 167248 150777 167276 152374
rect 167328 151548 167380 151554
rect 167328 151490 167380 151496
rect 167234 150768 167290 150777
rect 167234 150703 167290 150712
rect 164382 149816 164438 149825
rect 164382 149751 164384 149760
rect 164436 149751 164438 149760
rect 167144 149780 167196 149786
rect 164384 149722 164436 149728
rect 167144 149722 167196 149728
rect 163924 149644 163976 149650
rect 163924 149586 163976 149592
rect 164382 148592 164438 148601
rect 164382 148527 164384 148536
rect 164436 148527 164438 148536
rect 167052 148556 167104 148562
rect 164384 148498 164436 148504
rect 167052 148498 167104 148504
rect 164382 147368 164438 147377
rect 164382 147303 164438 147312
rect 164396 146862 164424 147303
rect 164384 146856 164436 146862
rect 164384 146798 164436 146804
rect 164382 146144 164438 146153
rect 164382 146079 164438 146088
rect 116818 145600 116874 145609
rect 116818 145535 116874 145544
rect 116832 142646 116860 145535
rect 164396 145502 164424 146079
rect 164384 145496 164436 145502
rect 164384 145438 164436 145444
rect 163738 144920 163794 144929
rect 163738 144855 163794 144864
rect 116820 142640 116872 142646
rect 116818 142608 116820 142617
rect 118936 142640 118988 142646
rect 116872 142608 116874 142617
rect 116818 142543 116874 142552
rect 118934 142608 118936 142617
rect 118988 142608 118990 142617
rect 118934 142543 118990 142552
rect 116832 142517 116860 142543
rect 163094 136488 163150 136497
rect 163094 136423 163150 136432
rect 125264 135902 125784 135930
rect 114060 134004 114112 134010
rect 114060 133946 114112 133952
rect 113968 133800 114020 133806
rect 113968 133742 114020 133748
rect 119488 133800 119540 133806
rect 119488 133742 119540 133748
rect 113232 133732 113284 133738
rect 113232 133674 113284 133680
rect 113324 133732 113376 133738
rect 113324 133674 113376 133680
rect 118936 133732 118988 133738
rect 118936 133674 118988 133680
rect 112772 133052 112824 133058
rect 112772 132994 112824 133000
rect 113140 133052 113192 133058
rect 113140 132994 113192 133000
rect 112588 130740 112640 130746
rect 112588 130682 112640 130688
rect 112784 128722 112812 132994
rect 113244 131290 113272 133674
rect 113324 133596 113376 133602
rect 113324 133538 113376 133544
rect 113232 131284 113284 131290
rect 113232 131226 113284 131232
rect 113336 130354 113364 133538
rect 114428 133392 114480 133398
rect 114428 133334 114480 133340
rect 113416 133324 113468 133330
rect 113416 133266 113468 133272
rect 113428 131154 113456 133266
rect 114440 131562 114468 133334
rect 114704 133256 114756 133262
rect 114704 133198 114756 133204
rect 114428 131556 114480 131562
rect 114428 131498 114480 131504
rect 114716 131426 114744 133198
rect 116084 133188 116136 133194
rect 116084 133130 116136 133136
rect 114796 133120 114848 133126
rect 114796 133062 114848 133068
rect 114704 131420 114756 131426
rect 114704 131362 114756 131368
rect 114808 131290 114836 133062
rect 115716 133052 115768 133058
rect 115716 132994 115768 133000
rect 114244 131284 114296 131290
rect 114244 131226 114296 131232
rect 114796 131284 114848 131290
rect 114796 131226 114848 131232
rect 113416 131148 113468 131154
rect 113416 131090 113468 131096
rect 113336 130326 113456 130354
rect 113428 128722 113456 130326
rect 112784 128694 113166 128722
rect 113428 128694 113718 128722
rect 114256 128708 114284 131226
rect 115440 131148 115492 131154
rect 115440 131090 115492 131096
rect 114888 130740 114940 130746
rect 114888 130682 114940 130688
rect 114900 128708 114928 130682
rect 115452 128708 115480 131090
rect 115728 131018 115756 132994
rect 116096 131630 116124 133130
rect 116084 131624 116136 131630
rect 116084 131566 116136 131572
rect 117740 131624 117792 131630
rect 117740 131566 117792 131572
rect 115992 131556 116044 131562
rect 115992 131498 116044 131504
rect 115716 131012 115768 131018
rect 115716 130954 115768 130960
rect 116004 128708 116032 131498
rect 116636 131420 116688 131426
rect 116636 131362 116688 131368
rect 116648 128708 116676 131362
rect 117188 131284 117240 131290
rect 117188 131226 117240 131232
rect 117200 128708 117228 131226
rect 117752 128708 117780 131566
rect 118384 131012 118436 131018
rect 118384 130954 118436 130960
rect 118396 128708 118424 130954
rect 118948 128708 118976 133674
rect 119500 128708 119528 133742
rect 88574 128464 88630 128473
rect 88574 128399 88630 128408
rect 88390 127920 88446 127929
rect 88390 127855 88446 127864
rect 88298 126696 88354 126705
rect 88298 126631 88354 126640
rect 88312 124665 88340 126631
rect 88404 125889 88432 127855
rect 88482 126424 88538 126433
rect 88588 126410 88616 128399
rect 123074 128192 123130 128201
rect 123074 128127 123130 128136
rect 88666 127376 88722 127385
rect 88666 127311 88722 127320
rect 88538 126382 88616 126410
rect 88482 126359 88538 126368
rect 88482 126152 88538 126161
rect 88482 126087 88538 126096
rect 88390 125880 88446 125889
rect 88390 125815 88446 125824
rect 88496 125458 88524 126087
rect 88404 125430 88524 125458
rect 88298 124656 88354 124665
rect 87748 124620 87800 124626
rect 88298 124591 88354 124600
rect 87748 124562 87800 124568
rect 87760 123441 87788 124562
rect 88404 124121 88432 125430
rect 88680 125322 88708 127311
rect 121694 127240 121750 127249
rect 121694 127175 121750 127184
rect 121708 126938 121736 127175
rect 123088 127113 123116 128127
rect 123166 127784 123222 127793
rect 123166 127719 123222 127728
rect 123074 127104 123130 127113
rect 123074 127039 123130 127048
rect 121696 126932 121748 126938
rect 121696 126874 121748 126880
rect 121786 126560 121842 126569
rect 121786 126495 121842 126504
rect 121800 126258 121828 126495
rect 121788 126252 121840 126258
rect 121788 126194 121840 126200
rect 121696 126184 121748 126190
rect 121694 126152 121696 126161
rect 121748 126152 121750 126161
rect 121694 126087 121750 126096
rect 123180 125889 123208 127719
rect 123996 126932 124048 126938
rect 123996 126874 124048 126880
rect 123904 126184 123956 126190
rect 123904 126126 123956 126132
rect 123166 125880 123222 125889
rect 123166 125815 123222 125824
rect 88758 125608 88814 125617
rect 88758 125543 88814 125552
rect 88496 125294 88708 125322
rect 88496 125209 88524 125294
rect 88482 125200 88538 125209
rect 88482 125135 88538 125144
rect 88482 124928 88538 124937
rect 88482 124863 88538 124872
rect 88390 124112 88446 124121
rect 88390 124047 88446 124056
rect 88390 123840 88446 123849
rect 88390 123775 88446 123784
rect 87746 123432 87802 123441
rect 87746 123367 87802 123376
rect 88206 122616 88262 122625
rect 88206 122551 88262 122560
rect 88220 120449 88248 122551
rect 88298 122072 88354 122081
rect 88298 122007 88354 122016
rect 88206 120440 88262 120449
rect 88206 120375 88262 120384
rect 88312 119905 88340 122007
rect 88404 121673 88432 123775
rect 88496 122897 88524 124863
rect 88772 124626 88800 125543
rect 121694 125472 121750 125481
rect 121694 125407 121750 125416
rect 121708 125170 121736 125407
rect 121696 125164 121748 125170
rect 121696 125106 121748 125112
rect 123720 125164 123772 125170
rect 123720 125106 123772 125112
rect 123166 124928 123222 124937
rect 123166 124863 123222 124872
rect 88760 124620 88812 124626
rect 88760 124562 88812 124568
rect 88666 124384 88722 124393
rect 88666 124319 88722 124328
rect 88574 123296 88630 123305
rect 88574 123231 88630 123240
rect 88482 122888 88538 122897
rect 88482 122823 88538 122832
rect 88390 121664 88446 121673
rect 88390 121599 88446 121608
rect 88390 121528 88446 121537
rect 88390 121463 88446 121472
rect 88298 119896 88354 119905
rect 88298 119831 88354 119840
rect 88298 119760 88354 119769
rect 88298 119695 88354 119704
rect 88206 119352 88262 119361
rect 88206 119287 88262 119296
rect 88114 117992 88170 118001
rect 88114 117927 88170 117936
rect 88128 115689 88156 117927
rect 88220 116913 88248 119287
rect 88312 117457 88340 119695
rect 88404 119225 88432 121463
rect 88482 121120 88538 121129
rect 88588 121106 88616 123231
rect 88680 122217 88708 124319
rect 122982 124112 123038 124121
rect 123038 124070 123116 124098
rect 122982 124047 123038 124056
rect 121694 123704 121750 123713
rect 121694 123639 121750 123648
rect 121708 123538 121736 123639
rect 121696 123532 121748 123538
rect 121696 123474 121748 123480
rect 122982 122888 123038 122897
rect 122982 122823 123038 122832
rect 121694 122480 121750 122489
rect 121694 122415 121750 122424
rect 88666 122208 88722 122217
rect 121708 122178 121736 122415
rect 88666 122143 88722 122152
rect 121696 122172 121748 122178
rect 121696 122114 121748 122120
rect 121694 122072 121750 122081
rect 122996 122058 123024 122823
rect 123088 122761 123116 124070
rect 123180 123305 123208 124863
rect 123732 123985 123760 125106
rect 123916 124529 123944 126126
rect 124008 125753 124036 126874
rect 124364 126252 124416 126258
rect 124364 126194 124416 126200
rect 123994 125744 124050 125753
rect 123994 125679 124050 125688
rect 124376 124665 124404 126194
rect 124362 124656 124418 124665
rect 124362 124591 124418 124600
rect 123902 124520 123958 124529
rect 123902 124455 123958 124464
rect 123718 123976 123774 123985
rect 123718 123911 123774 123920
rect 123536 123532 123588 123538
rect 123536 123474 123588 123480
rect 123166 123296 123222 123305
rect 123166 123231 123222 123240
rect 123074 122752 123130 122761
rect 123074 122687 123130 122696
rect 123444 122172 123496 122178
rect 123444 122114 123496 122120
rect 122996 122030 123116 122058
rect 121694 122007 121696 122016
rect 121748 122007 121750 122016
rect 121696 121978 121748 121984
rect 123088 121537 123116 122030
rect 123352 122036 123404 122042
rect 123352 121978 123404 121984
rect 123074 121528 123130 121537
rect 123074 121463 123130 121472
rect 121694 121256 121750 121265
rect 121694 121191 121750 121200
rect 88538 121078 88616 121106
rect 88482 121055 88538 121064
rect 121708 120954 121736 121191
rect 121696 120948 121748 120954
rect 121696 120890 121748 120896
rect 88482 120848 88538 120857
rect 88482 120783 88538 120792
rect 88390 119216 88446 119225
rect 88390 119151 88446 119160
rect 88496 118681 88524 120783
rect 122982 120712 123038 120721
rect 123038 120670 123208 120698
rect 122982 120647 123038 120656
rect 88574 120304 88630 120313
rect 88574 120239 88630 120248
rect 88482 118672 88538 118681
rect 88482 118607 88538 118616
rect 88390 118536 88446 118545
rect 88390 118471 88446 118480
rect 88298 117448 88354 117457
rect 88298 117383 88354 117392
rect 88206 116904 88262 116913
rect 88206 116839 88262 116848
rect 88404 116233 88432 118471
rect 88482 118128 88538 118137
rect 88588 118114 88616 120239
rect 122982 120032 123038 120041
rect 123038 119990 123116 120018
rect 122982 119967 123038 119976
rect 121694 119624 121750 119633
rect 121694 119559 121750 119568
rect 121708 119390 121736 119559
rect 121696 119384 121748 119390
rect 121696 119326 121748 119332
rect 123088 118545 123116 119990
rect 123180 119089 123208 120670
rect 123364 120313 123392 121978
rect 123456 120449 123484 122114
rect 123548 121673 123576 123474
rect 123534 121664 123590 121673
rect 123534 121599 123590 121608
rect 124364 120948 124416 120954
rect 124364 120890 124416 120896
rect 123442 120440 123498 120449
rect 123442 120375 123498 120384
rect 123350 120304 123406 120313
rect 123350 120239 123406 120248
rect 124272 119384 124324 119390
rect 123258 119352 123314 119361
rect 124272 119326 124324 119332
rect 123258 119287 123314 119296
rect 123166 119080 123222 119089
rect 123166 119015 123222 119024
rect 123074 118536 123130 118545
rect 123074 118471 123130 118480
rect 121694 118400 121750 118409
rect 121694 118335 121750 118344
rect 121708 118234 121736 118335
rect 121696 118228 121748 118234
rect 121696 118170 121748 118176
rect 88538 118086 88616 118114
rect 88482 118063 88538 118072
rect 123166 117992 123222 118001
rect 123166 117927 123222 117936
rect 88666 117448 88722 117457
rect 88666 117383 88722 117392
rect 88482 116768 88538 116777
rect 88482 116703 88538 116712
rect 88390 116224 88446 116233
rect 88390 116159 88446 116168
rect 88114 115680 88170 115689
rect 88114 115615 88170 115624
rect 88390 115680 88446 115689
rect 88390 115615 88446 115624
rect 88206 115272 88262 115281
rect 88206 115207 88262 115216
rect 88114 113912 88170 113921
rect 88114 113847 88170 113856
rect 88022 113368 88078 113377
rect 88022 113303 88078 113312
rect 88036 110929 88064 113303
rect 88128 111473 88156 113847
rect 88220 112697 88248 115207
rect 88298 114456 88354 114465
rect 88298 114391 88354 114400
rect 88206 112688 88262 112697
rect 88206 112623 88262 112632
rect 88312 112153 88340 114391
rect 88404 113241 88432 115615
rect 88496 115009 88524 116703
rect 88574 116224 88630 116233
rect 88574 116159 88630 116168
rect 88482 115000 88538 115009
rect 88482 114935 88538 114944
rect 88482 114320 88538 114329
rect 88588 114306 88616 116159
rect 88680 115145 88708 117383
rect 122982 117040 123038 117049
rect 123038 116998 123116 117026
rect 122982 116975 123038 116984
rect 123088 116602 123116 116998
rect 123076 116596 123128 116602
rect 123076 116538 123128 116544
rect 123074 116496 123130 116505
rect 123074 116431 123130 116440
rect 121694 115952 121750 115961
rect 121694 115887 121750 115896
rect 121708 115718 121736 115887
rect 121696 115712 121748 115718
rect 121696 115654 121748 115660
rect 121694 115544 121750 115553
rect 121694 115479 121750 115488
rect 121708 115446 121736 115479
rect 121696 115440 121748 115446
rect 121696 115382 121748 115388
rect 121696 115168 121748 115174
rect 88666 115136 88722 115145
rect 88666 115071 88722 115080
rect 121694 115136 121696 115145
rect 121748 115136 121750 115145
rect 121694 115071 121750 115080
rect 123088 115009 123116 116431
rect 123180 116097 123208 117927
rect 123272 117321 123300 119287
rect 124284 117865 124312 119326
rect 124376 119225 124404 120890
rect 124362 119216 124418 119225
rect 124362 119151 124418 119160
rect 124364 118228 124416 118234
rect 124364 118170 124416 118176
rect 124270 117856 124326 117865
rect 124270 117791 124326 117800
rect 123258 117312 123314 117321
rect 123258 117247 123314 117256
rect 124272 116596 124324 116602
rect 124272 116538 124324 116544
rect 123166 116088 123222 116097
rect 123166 116023 123222 116032
rect 124284 115553 124312 116538
rect 124376 116233 124404 118170
rect 124362 116224 124418 116233
rect 124362 116159 124418 116168
rect 124364 115712 124416 115718
rect 124364 115654 124416 115660
rect 124270 115544 124326 115553
rect 124270 115479 124326 115488
rect 123996 115440 124048 115446
rect 123996 115382 124048 115388
rect 123074 115000 123130 115009
rect 123074 114935 123130 114944
rect 88538 114278 88616 114306
rect 121694 114320 121750 114329
rect 88482 114255 88538 114264
rect 121694 114255 121750 114264
rect 121708 114018 121736 114255
rect 121696 114012 121748 114018
rect 121696 113954 121748 113960
rect 123444 114012 123496 114018
rect 123444 113954 123496 113960
rect 122982 113776 123038 113785
rect 123038 113734 123208 113762
rect 122982 113711 123038 113720
rect 88390 113232 88446 113241
rect 88390 113167 88446 113176
rect 88482 112688 88538 112697
rect 88482 112623 88538 112632
rect 88298 112144 88354 112153
rect 88298 112079 88354 112088
rect 88298 111600 88354 111609
rect 88298 111535 88354 111544
rect 88114 111464 88170 111473
rect 88114 111399 88170 111408
rect 88022 110920 88078 110929
rect 88022 110855 88078 110864
rect 88206 109832 88262 109841
rect 88206 109767 88262 109776
rect 88114 109288 88170 109297
rect 88114 109223 88170 109232
rect 88022 107520 88078 107529
rect 88022 107455 88078 107464
rect 85172 106872 85224 106878
rect 85170 106840 85172 106849
rect 85224 106840 85226 106849
rect 85170 106775 85226 106784
rect 88036 104945 88064 107455
rect 88128 106713 88156 109223
rect 88220 107257 88248 109767
rect 88312 109161 88340 111535
rect 88390 111056 88446 111065
rect 88390 110991 88446 111000
rect 88298 109152 88354 109161
rect 88298 109087 88354 109096
rect 88298 108608 88354 108617
rect 88298 108543 88354 108552
rect 88206 107248 88262 107257
rect 88206 107183 88262 107192
rect 88114 106704 88170 106713
rect 88114 106639 88170 106648
rect 88312 106169 88340 108543
rect 88404 108481 88432 110991
rect 88496 110249 88524 112623
rect 121694 112552 121750 112561
rect 121694 112487 121750 112496
rect 121708 112386 121736 112487
rect 121696 112380 121748 112386
rect 121696 112322 121748 112328
rect 88666 112144 88722 112153
rect 88666 112079 88722 112088
rect 88574 110376 88630 110385
rect 88574 110311 88630 110320
rect 88482 110240 88538 110249
rect 88482 110175 88538 110184
rect 88588 109682 88616 110311
rect 88680 109705 88708 112079
rect 123180 111881 123208 113734
rect 123258 112960 123314 112969
rect 123258 112895 123314 112904
rect 122982 111872 123038 111881
rect 123166 111872 123222 111881
rect 123038 111830 123116 111858
rect 122982 111807 123038 111816
rect 121694 111328 121750 111337
rect 121694 111263 121750 111272
rect 121708 111026 121736 111263
rect 121696 111020 121748 111026
rect 121696 110962 121748 110968
rect 123088 110113 123116 111830
rect 123166 111807 123222 111816
rect 123166 111056 123222 111065
rect 123166 110991 123222 111000
rect 123180 110770 123208 110991
rect 123272 110929 123300 112895
rect 123352 112380 123404 112386
rect 123352 112322 123404 112328
rect 123258 110920 123314 110929
rect 123258 110855 123314 110864
rect 123364 110793 123392 112322
rect 123456 112153 123484 113954
rect 124008 113649 124036 115382
rect 124272 115168 124324 115174
rect 124272 115110 124324 115116
rect 123994 113640 124050 113649
rect 123994 113575 124050 113584
rect 124284 113105 124312 115110
rect 124376 114329 124404 115654
rect 124362 114320 124418 114329
rect 124362 114255 124418 114264
rect 124270 113096 124326 113105
rect 124270 113031 124326 113040
rect 123442 112144 123498 112153
rect 123442 112079 123498 112088
rect 124272 111020 124324 111026
rect 124272 110962 124324 110968
rect 123350 110784 123406 110793
rect 123180 110742 123300 110770
rect 121694 110104 121750 110113
rect 121694 110039 121750 110048
rect 123074 110104 123130 110113
rect 123074 110039 123130 110048
rect 121708 109802 121736 110039
rect 121696 109796 121748 109802
rect 121696 109738 121748 109744
rect 88496 109654 88616 109682
rect 88666 109696 88722 109705
rect 88390 108472 88446 108481
rect 88390 108407 88446 108416
rect 88496 107937 88524 109654
rect 88666 109631 88722 109640
rect 122982 109696 123038 109705
rect 122982 109631 123038 109640
rect 122996 109546 123024 109631
rect 122996 109518 123208 109546
rect 121694 109016 121750 109025
rect 121694 108951 121750 108960
rect 121708 108782 121736 108951
rect 121696 108776 121748 108782
rect 121696 108718 121748 108724
rect 88574 108064 88630 108073
rect 88574 107999 88630 108008
rect 88482 107928 88538 107937
rect 88482 107863 88538 107872
rect 88482 106840 88538 106849
rect 88482 106775 88538 106784
rect 88390 106296 88446 106305
rect 88390 106231 88446 106240
rect 88298 106160 88354 106169
rect 88298 106095 88354 106104
rect 88298 105752 88354 105761
rect 88298 105687 88354 105696
rect 88022 104936 88078 104945
rect 88022 104871 88078 104880
rect 85908 104152 85960 104158
rect 85908 104094 85960 104100
rect 85816 104084 85868 104090
rect 85816 104026 85868 104032
rect 54076 103064 54128 103070
rect 54076 103006 54128 103012
rect 53984 96468 54036 96474
rect 53984 96410 54036 96416
rect 54088 93906 54116 103006
rect 55364 102792 55416 102798
rect 55364 102734 55416 102740
rect 55376 95810 55404 102734
rect 55560 101001 55588 102868
rect 55546 100992 55602 101001
rect 55546 100927 55602 100936
rect 56742 100992 56798 101001
rect 56742 100927 56798 100936
rect 56756 100078 56784 100927
rect 56744 100072 56796 100078
rect 56744 100014 56796 100020
rect 56940 98514 56968 102868
rect 58412 101302 58440 102868
rect 58400 101296 58452 101302
rect 58400 101238 58452 101244
rect 59792 99942 59820 102868
rect 61264 99942 61292 102868
rect 62644 99942 62672 102868
rect 63828 100004 63880 100010
rect 63828 99946 63880 99952
rect 59320 99936 59372 99942
rect 59320 99878 59372 99884
rect 59780 99936 59832 99942
rect 59780 99878 59832 99884
rect 60424 99936 60476 99942
rect 60424 99878 60476 99884
rect 61252 99936 61304 99942
rect 61252 99878 61304 99884
rect 61528 99936 61580 99942
rect 61528 99878 61580 99884
rect 62632 99936 62684 99942
rect 62632 99878 62684 99884
rect 63000 99936 63052 99942
rect 63000 99878 63052 99884
rect 56928 98508 56980 98514
rect 56928 98450 56980 98456
rect 57112 97080 57164 97086
rect 57112 97022 57164 97028
rect 55376 95782 55496 95810
rect 54088 93878 54392 93906
rect 54364 93770 54392 93878
rect 55468 93770 55496 95782
rect 54364 93742 54930 93770
rect 55468 93742 56034 93770
rect 57124 93756 57152 97022
rect 58216 96536 58268 96542
rect 58216 96478 58268 96484
rect 58228 93756 58256 96478
rect 59332 93756 59360 99878
rect 60436 93756 60464 99878
rect 61540 93756 61568 99878
rect 63012 93770 63040 99878
rect 62658 93742 63040 93770
rect 63840 93756 63868 99946
rect 64116 99942 64144 102868
rect 64932 100140 64984 100146
rect 64932 100082 64984 100088
rect 64104 99936 64156 99942
rect 64104 99878 64156 99884
rect 64944 93756 64972 100082
rect 65496 100010 65524 102868
rect 66968 100146 66996 102868
rect 66956 100140 67008 100146
rect 66956 100082 67008 100088
rect 68244 100140 68296 100146
rect 68244 100082 68296 100088
rect 67140 100072 67192 100078
rect 67140 100014 67192 100020
rect 65484 100004 65536 100010
rect 65484 99946 65536 99952
rect 66036 100004 66088 100010
rect 66036 99946 66088 99952
rect 66048 93756 66076 99946
rect 67152 93756 67180 100014
rect 68256 93756 68284 100082
rect 68348 100010 68376 102868
rect 69348 100208 69400 100214
rect 69348 100150 69400 100156
rect 68336 100004 68388 100010
rect 68336 99946 68388 99952
rect 69360 93756 69388 100150
rect 69820 100078 69848 102868
rect 71200 100146 71228 102868
rect 71556 100412 71608 100418
rect 71556 100354 71608 100360
rect 71188 100140 71240 100146
rect 71188 100082 71240 100088
rect 69808 100072 69860 100078
rect 69808 100014 69860 100020
rect 70452 100072 70504 100078
rect 70452 100014 70504 100020
rect 70464 93756 70492 100014
rect 71568 93756 71596 100354
rect 72672 100214 72700 102868
rect 73764 100820 73816 100826
rect 73764 100762 73816 100768
rect 72660 100208 72712 100214
rect 72660 100150 72712 100156
rect 72660 100004 72712 100010
rect 72660 99946 72712 99952
rect 72672 93756 72700 99946
rect 73776 93756 73804 100762
rect 74052 100078 74080 102868
rect 75524 100214 75552 102868
rect 75512 100208 75564 100214
rect 75512 100150 75564 100156
rect 75972 100140 76024 100146
rect 75972 100082 76024 100088
rect 74040 100072 74092 100078
rect 74040 100014 74092 100020
rect 74868 100072 74920 100078
rect 74868 100014 74920 100020
rect 74880 93756 74908 100014
rect 75984 93756 76012 100082
rect 76904 100010 76932 102868
rect 78376 100826 78404 102868
rect 78364 100820 78416 100826
rect 78364 100762 78416 100768
rect 79756 100078 79784 102868
rect 80480 101364 80532 101370
rect 80480 101306 80532 101312
rect 79744 100072 79796 100078
rect 79744 100014 79796 100020
rect 76892 100004 76944 100010
rect 76892 99946 76944 99952
rect 77168 96468 77220 96474
rect 77168 96410 77220 96416
rect 79376 96468 79428 96474
rect 79376 96410 79428 96416
rect 77180 93756 77208 96410
rect 79388 93756 79416 96410
rect 80492 93756 80520 101306
rect 81228 100146 81256 102868
rect 84094 102854 84384 102882
rect 81584 101432 81636 101438
rect 81584 101374 81636 101380
rect 81216 100140 81268 100146
rect 81216 100082 81268 100088
rect 81596 93756 81624 101374
rect 84356 100706 84384 102854
rect 84356 100678 84476 100706
rect 84448 96746 84476 100678
rect 84896 96876 84948 96882
rect 84896 96818 84948 96824
rect 84436 96740 84488 96746
rect 84436 96682 84488 96688
rect 83792 96604 83844 96610
rect 83792 96546 83844 96552
rect 82688 96536 82740 96542
rect 82688 96478 82740 96484
rect 82700 93756 82728 96478
rect 83804 93756 83832 96546
rect 84908 93756 84936 96818
rect 85828 93770 85856 104026
rect 85920 97154 85948 104094
rect 88312 103177 88340 105687
rect 88404 103721 88432 106231
rect 88496 104265 88524 106775
rect 88588 105489 88616 107999
rect 123180 107801 123208 109518
rect 123272 109025 123300 110742
rect 123350 110719 123406 110728
rect 124284 109569 124312 110962
rect 124364 109796 124416 109802
rect 124364 109738 124416 109744
rect 124270 109560 124326 109569
rect 124270 109495 124326 109504
rect 123258 109016 123314 109025
rect 123258 108951 123314 108960
rect 123444 108776 123496 108782
rect 123444 108718 123496 108724
rect 123258 108472 123314 108481
rect 123258 108407 123314 108416
rect 122982 107792 123038 107801
rect 123166 107792 123222 107801
rect 123038 107750 123116 107778
rect 122982 107727 123038 107736
rect 123088 107642 123116 107750
rect 123166 107727 123222 107736
rect 123088 107614 123208 107642
rect 121694 107248 121750 107257
rect 121694 107183 121750 107192
rect 121708 106878 121736 107183
rect 121696 106872 121748 106878
rect 121696 106814 121748 106820
rect 123074 106840 123130 106849
rect 123074 106775 123130 106784
rect 121694 106160 121750 106169
rect 121694 106095 121750 106104
rect 121708 105926 121736 106095
rect 121696 105920 121748 105926
rect 121696 105862 121748 105868
rect 121694 105752 121750 105761
rect 121694 105687 121750 105696
rect 121708 105654 121736 105687
rect 121696 105648 121748 105654
rect 121696 105590 121748 105596
rect 88574 105480 88630 105489
rect 88574 105415 88630 105424
rect 88666 105208 88722 105217
rect 88666 105143 88722 105152
rect 88574 104528 88630 104537
rect 88574 104463 88630 104472
rect 88482 104256 88538 104265
rect 88482 104191 88538 104200
rect 88588 104090 88616 104463
rect 88680 104158 88708 105143
rect 123088 104809 123116 106775
rect 123180 106033 123208 107614
rect 123272 106577 123300 108407
rect 123456 106713 123484 108718
rect 124376 108209 124404 109738
rect 124362 108200 124418 108209
rect 124362 108135 124418 108144
rect 124272 106872 124324 106878
rect 124272 106814 124324 106820
rect 123442 106704 123498 106713
rect 123442 106639 123498 106648
rect 123258 106568 123314 106577
rect 123258 106503 123314 106512
rect 123166 106024 123222 106033
rect 123166 105959 123222 105968
rect 124180 105648 124232 105654
rect 124180 105590 124232 105596
rect 121786 104800 121842 104809
rect 121786 104735 121842 104744
rect 123074 104800 123130 104809
rect 123074 104735 123130 104744
rect 91060 104696 91112 104702
rect 91060 104638 91112 104644
rect 88668 104152 88720 104158
rect 88668 104094 88720 104100
rect 88576 104084 88628 104090
rect 88576 104026 88628 104032
rect 88482 103984 88538 103993
rect 88482 103919 88538 103928
rect 88390 103712 88446 103721
rect 88390 103647 88446 103656
rect 88496 103562 88524 103919
rect 88404 103534 88524 103562
rect 88298 103168 88354 103177
rect 88298 103103 88354 103112
rect 85908 97148 85960 97154
rect 85908 97090 85960 97096
rect 87104 97148 87156 97154
rect 87104 97090 87156 97096
rect 85828 93742 86026 93770
rect 87116 93756 87144 97090
rect 88404 96882 88432 103534
rect 88482 103440 88538 103449
rect 88482 103375 88538 103384
rect 88392 96876 88444 96882
rect 88392 96818 88444 96824
rect 88208 96740 88260 96746
rect 88208 96682 88260 96688
rect 88220 93756 88248 96682
rect 88496 96610 88524 103375
rect 89678 102760 89734 102769
rect 89678 102695 89734 102704
rect 88666 102216 88722 102225
rect 88666 102151 88722 102160
rect 88574 101672 88630 101681
rect 88574 101607 88630 101616
rect 88588 101370 88616 101607
rect 88680 101438 88708 102151
rect 88668 101432 88720 101438
rect 88668 101374 88720 101380
rect 88576 101364 88628 101370
rect 88576 101306 88628 101312
rect 88574 100584 88630 100593
rect 88574 100519 88630 100528
rect 88484 96604 88536 96610
rect 88484 96546 88536 96552
rect 88588 96474 88616 100519
rect 89692 96542 89720 102695
rect 89680 96536 89732 96542
rect 89680 96478 89732 96484
rect 88576 96468 88628 96474
rect 88576 96410 88628 96416
rect 91072 92326 91100 104638
rect 121694 104392 121750 104401
rect 121694 104327 121750 104336
rect 121708 104090 121736 104327
rect 121800 104158 121828 104735
rect 121788 104152 121840 104158
rect 121788 104094 121840 104100
rect 121696 104084 121748 104090
rect 121696 104026 121748 104032
rect 121878 103712 121934 103721
rect 121878 103647 121934 103656
rect 121786 103304 121842 103313
rect 121786 103239 121842 103248
rect 121694 102896 121750 102905
rect 121694 102831 121696 102840
rect 121748 102831 121750 102840
rect 121696 102802 121748 102808
rect 121800 102798 121828 103239
rect 121788 102792 121840 102798
rect 121788 102734 121840 102740
rect 121892 102730 121920 103647
rect 124192 103585 124220 105590
rect 124284 105353 124312 106814
rect 124364 105920 124416 105926
rect 124364 105862 124416 105868
rect 124270 105344 124326 105353
rect 124270 105279 124326 105288
rect 124376 103993 124404 105862
rect 124362 103984 124418 103993
rect 124362 103919 124418 103928
rect 124178 103576 124234 103585
rect 124178 103511 124234 103520
rect 124548 102860 124600 102866
rect 124548 102802 124600 102808
rect 121880 102724 121932 102730
rect 121880 102666 121932 102672
rect 123074 101944 123130 101953
rect 123074 101879 123130 101888
rect 116360 101092 116412 101098
rect 116360 101034 116412 101040
rect 91348 100950 92098 100978
rect 92268 100950 92558 100978
rect 92820 100950 93110 100978
rect 93280 100950 93662 100978
rect 94108 100950 94214 100978
rect 94384 100950 94766 100978
rect 94936 100950 95318 100978
rect 95488 100950 95870 100978
rect 96040 100950 96422 100978
rect 97144 100950 97526 100978
rect 97972 100950 98078 100978
rect 98984 100950 99182 100978
rect 99628 100950 99734 100978
rect 99904 100950 100286 100978
rect 100456 100950 100838 100978
rect 101008 100950 101390 100978
rect 101560 100950 101942 100978
rect 102388 100950 102494 100978
rect 102664 100950 103046 100978
rect 103216 100950 103598 100978
rect 103952 100950 104150 100978
rect 104320 100950 104702 100978
rect 105148 100950 105254 100978
rect 105424 100950 105806 100978
rect 105976 100950 106266 100978
rect 106528 100950 106818 100978
rect 107080 100950 107370 100978
rect 108184 100950 108474 100978
rect 108736 100950 109026 100978
rect 109288 100950 109578 100978
rect 109840 100950 110130 100978
rect 110944 100950 111234 100978
rect 111496 100950 111786 100978
rect 112048 100950 112338 100978
rect 112600 100950 112890 100978
rect 113704 100950 113994 100978
rect 114256 100950 114546 100978
rect 114808 100950 115098 100978
rect 115360 100950 115650 100978
rect 91060 92320 91112 92326
rect 91060 92262 91112 92268
rect 18104 90212 18156 90218
rect 18104 90154 18156 90160
rect 22336 90212 22388 90218
rect 22336 90154 22388 90160
rect 22348 89849 22376 90154
rect 22334 89840 22390 89849
rect 22334 89775 22390 89784
rect 45058 89840 45114 89849
rect 45058 89775 45114 89784
rect 15436 82324 15488 82330
rect 15436 82266 15488 82272
rect 15448 75054 15476 82266
rect 22336 81984 22388 81990
rect 22336 81926 22388 81932
rect 22348 81825 22376 81926
rect 22334 81816 22390 81825
rect 22334 81751 22390 81760
rect 45072 75054 45100 89775
rect 91348 84681 91376 100950
rect 92268 98258 92296 100950
rect 91440 98230 92296 98258
rect 91440 85905 91468 98230
rect 92164 98168 92216 98174
rect 92164 98110 92216 98116
rect 91704 94088 91756 94094
rect 91704 94030 91756 94036
rect 91716 93249 91744 94030
rect 91702 93240 91758 93249
rect 91702 93175 91758 93184
rect 91796 91708 91848 91714
rect 91796 91650 91848 91656
rect 91520 91368 91572 91374
rect 91520 91310 91572 91316
rect 91532 90801 91560 91310
rect 91518 90792 91574 90801
rect 91518 90727 91574 90736
rect 91426 85896 91482 85905
rect 91426 85831 91482 85840
rect 91334 84672 91390 84681
rect 91334 84607 91390 84616
rect 91808 83457 91836 91650
rect 92176 89577 92204 98110
rect 92348 98100 92400 98106
rect 92348 98042 92400 98048
rect 92360 95538 92388 98042
rect 92440 97216 92492 97222
rect 92440 97158 92492 97164
rect 92268 95510 92388 95538
rect 92268 92025 92296 95510
rect 92254 92016 92310 92025
rect 92254 91951 92310 91960
rect 92162 89568 92218 89577
rect 92162 89503 92218 89512
rect 92256 88920 92308 88926
rect 92256 88862 92308 88868
rect 92164 87560 92216 87566
rect 92164 87502 92216 87508
rect 91794 83448 91850 83457
rect 91794 83383 91850 83392
rect 92176 81145 92204 87502
rect 92268 82233 92296 88862
rect 92452 88353 92480 97158
rect 92438 88344 92494 88353
rect 92438 88279 92494 88288
rect 92820 87129 92848 100950
rect 93280 97222 93308 100950
rect 93360 98304 93412 98310
rect 93360 98246 93412 98252
rect 93268 97216 93320 97222
rect 93268 97158 93320 97164
rect 93372 91374 93400 98246
rect 94108 98174 94136 100950
rect 94384 98310 94412 100950
rect 94372 98304 94424 98310
rect 94372 98246 94424 98252
rect 94096 98168 94148 98174
rect 94096 98110 94148 98116
rect 94936 98106 94964 100950
rect 94924 98100 94976 98106
rect 94924 98042 94976 98048
rect 95488 94094 95516 100950
rect 96040 100706 96068 100950
rect 96974 100814 97080 100842
rect 95948 100678 96068 100706
rect 95948 100146 95976 100678
rect 95936 100140 95988 100146
rect 95936 100082 95988 100088
rect 95948 99942 95976 100082
rect 97052 99942 97080 100814
rect 95936 99936 95988 99942
rect 95936 99878 95988 99884
rect 97040 99936 97092 99942
rect 97040 99878 97092 99884
rect 97144 98514 97172 100950
rect 97132 98508 97184 98514
rect 97132 98450 97184 98456
rect 95476 94088 95528 94094
rect 95476 94030 95528 94036
rect 97972 93634 98000 100950
rect 98630 100814 98736 100842
rect 98708 93634 98736 100814
rect 98984 93770 99012 100950
rect 99628 95810 99656 100950
rect 99536 95782 99656 95810
rect 99536 93770 99564 95782
rect 99904 93770 99932 100950
rect 100456 95998 100484 100950
rect 100260 95992 100312 95998
rect 100260 95934 100312 95940
rect 100444 95992 100496 95998
rect 100444 95934 100496 95940
rect 100272 93770 100300 95934
rect 101008 95810 101036 100950
rect 101456 95924 101508 95930
rect 101456 95866 101508 95872
rect 100732 95782 101036 95810
rect 100732 93770 100760 95782
rect 100996 95720 101048 95726
rect 100996 95662 101048 95668
rect 98860 93742 99012 93770
rect 99320 93742 99564 93770
rect 99688 93742 99932 93770
rect 100056 93742 100300 93770
rect 100516 93742 100760 93770
rect 97972 93606 98124 93634
rect 98492 93606 98736 93634
rect 101008 93498 101036 95662
rect 101468 93770 101496 95866
rect 101560 95862 101588 100950
rect 102284 96060 102336 96066
rect 102284 96002 102336 96008
rect 101916 95992 101968 95998
rect 101916 95934 101968 95940
rect 101548 95856 101600 95862
rect 101548 95798 101600 95804
rect 101928 93770 101956 95934
rect 102296 93770 102324 96002
rect 102388 95930 102416 100950
rect 102664 95998 102692 100950
rect 103216 96066 103244 100950
rect 103756 97284 103808 97290
rect 103756 97226 103808 97232
rect 103480 97148 103532 97154
rect 103480 97090 103532 97096
rect 103204 96060 103256 96066
rect 103204 96002 103256 96008
rect 102652 95992 102704 95998
rect 102652 95934 102704 95940
rect 103112 95992 103164 95998
rect 103112 95934 103164 95940
rect 102376 95924 102428 95930
rect 102376 95866 102428 95872
rect 102744 95924 102796 95930
rect 102744 95866 102796 95872
rect 102756 93770 102784 95866
rect 103124 93770 103152 95934
rect 103492 93770 103520 97090
rect 103768 95810 103796 97226
rect 103952 95930 103980 100950
rect 104320 95998 104348 100950
rect 105148 97222 105176 100950
rect 105228 97352 105280 97358
rect 105228 97294 105280 97300
rect 105136 97216 105188 97222
rect 105136 97158 105188 97164
rect 104676 97148 104728 97154
rect 104676 97090 104728 97096
rect 104308 95992 104360 95998
rect 104308 95934 104360 95940
rect 103940 95924 103992 95930
rect 103940 95866 103992 95872
rect 103676 95782 103796 95810
rect 104308 95856 104360 95862
rect 104308 95798 104360 95804
rect 103676 94042 103704 95782
rect 101252 93742 101496 93770
rect 101712 93742 101956 93770
rect 102080 93742 102324 93770
rect 102448 93742 102784 93770
rect 102908 93742 103152 93770
rect 103276 93742 103520 93770
rect 103630 94014 103704 94042
rect 103630 93756 103658 94014
rect 104320 93770 104348 95798
rect 104688 93770 104716 97090
rect 105240 95946 105268 97294
rect 105424 97290 105452 100950
rect 105412 97284 105464 97290
rect 105412 97226 105464 97232
rect 105872 97148 105924 97154
rect 105872 97090 105924 97096
rect 105504 97080 105556 97086
rect 105504 97022 105556 97028
rect 105056 95918 105268 95946
rect 105056 93770 105084 95918
rect 105516 93770 105544 97022
rect 105884 93770 105912 97090
rect 105976 95862 106004 100950
rect 106528 97222 106556 100950
rect 107080 97358 107108 100950
rect 107922 100814 108028 100842
rect 107068 97352 107120 97358
rect 107068 97294 107120 97300
rect 106608 97284 106660 97290
rect 106608 97226 106660 97232
rect 106516 97216 106568 97222
rect 106516 97158 106568 97164
rect 105964 95856 106016 95862
rect 106620 95810 106648 97226
rect 107160 97148 107212 97154
rect 107160 97090 107212 97096
rect 105964 95798 106016 95804
rect 106344 95782 106648 95810
rect 106700 95856 106752 95862
rect 106700 95798 106752 95804
rect 106344 93770 106372 95782
rect 106712 93770 106740 95798
rect 107172 93770 107200 97090
rect 108000 97086 108028 100814
rect 108184 97222 108212 100950
rect 108736 97290 108764 100950
rect 108724 97284 108776 97290
rect 108724 97226 108776 97232
rect 108172 97216 108224 97222
rect 109288 97170 109316 100950
rect 109840 97222 109868 100950
rect 110682 100814 110788 100842
rect 108172 97158 108224 97164
rect 108356 97148 108408 97154
rect 108356 97090 108408 97096
rect 109196 97142 109316 97170
rect 109828 97216 109880 97222
rect 109828 97158 109880 97164
rect 107988 97080 108040 97086
rect 107988 97022 108040 97028
rect 107528 97012 107580 97018
rect 107528 96954 107580 96960
rect 107540 93770 107568 96954
rect 107804 96944 107856 96950
rect 107804 96886 107856 96892
rect 107816 93770 107844 96886
rect 108368 93770 108396 97090
rect 108724 96808 108776 96814
rect 108724 96750 108776 96756
rect 108736 93770 108764 96750
rect 109000 96740 109052 96746
rect 109000 96682 109052 96688
rect 109012 93770 109040 96682
rect 109196 95862 109224 97142
rect 110760 97018 110788 100814
rect 110748 97012 110800 97018
rect 110748 96954 110800 96960
rect 110944 96950 110972 100950
rect 111496 97222 111524 100950
rect 111484 97216 111536 97222
rect 111484 97158 111536 97164
rect 110932 96944 110984 96950
rect 110932 96886 110984 96892
rect 112048 96814 112076 100950
rect 112036 96808 112088 96814
rect 112036 96750 112088 96756
rect 112600 96746 112628 100950
rect 113442 100814 113548 100842
rect 112588 96740 112640 96746
rect 112588 96682 112640 96688
rect 113520 96542 113548 100814
rect 109552 96536 109604 96542
rect 109552 96478 109604 96484
rect 113508 96536 113560 96542
rect 113508 96478 113560 96484
rect 109184 95856 109236 95862
rect 109184 95798 109236 95804
rect 109564 93770 109592 96478
rect 113704 96474 113732 100950
rect 109920 96468 109972 96474
rect 109920 96410 109972 96416
rect 113692 96468 113744 96474
rect 113692 96410 113744 96416
rect 113968 96468 114020 96474
rect 113968 96410 114020 96416
rect 109932 93770 109960 96410
rect 110564 96400 110616 96406
rect 110564 96342 110616 96348
rect 110288 96332 110340 96338
rect 110288 96274 110340 96280
rect 110300 93770 110328 96274
rect 110576 93770 110604 96342
rect 111116 96264 111168 96270
rect 111116 96206 111168 96212
rect 111128 93770 111156 96206
rect 111484 96196 111536 96202
rect 111484 96138 111536 96144
rect 111496 93770 111524 96138
rect 111944 96128 111996 96134
rect 111944 96070 111996 96076
rect 111956 93770 111984 96070
rect 112680 96060 112732 96066
rect 112680 96002 112732 96008
rect 112312 95924 112364 95930
rect 112312 95866 112364 95872
rect 112324 93770 112352 95866
rect 112692 93770 112720 96002
rect 113140 95992 113192 95998
rect 113140 95934 113192 95940
rect 113152 93770 113180 95934
rect 113232 95856 113284 95862
rect 113232 95798 113284 95804
rect 113244 94042 113272 95798
rect 113244 94014 113318 94042
rect 104104 93742 104348 93770
rect 104472 93742 104716 93770
rect 104840 93742 105084 93770
rect 105300 93742 105544 93770
rect 105668 93742 105912 93770
rect 106128 93742 106372 93770
rect 106496 93742 106740 93770
rect 106864 93742 107200 93770
rect 107324 93742 107568 93770
rect 107692 93742 107844 93770
rect 108060 93742 108396 93770
rect 108520 93742 108764 93770
rect 108888 93742 109040 93770
rect 109256 93742 109592 93770
rect 109716 93742 109960 93770
rect 110084 93742 110328 93770
rect 110452 93742 110604 93770
rect 110912 93742 111156 93770
rect 111280 93742 111524 93770
rect 111648 93742 111984 93770
rect 112108 93742 112352 93770
rect 112476 93742 112720 93770
rect 112844 93742 113180 93770
rect 113290 93756 113318 94014
rect 113980 93770 114008 96410
rect 114256 96338 114284 100950
rect 114808 96406 114836 100950
rect 114796 96400 114848 96406
rect 114796 96342 114848 96348
rect 114244 96332 114296 96338
rect 114244 96274 114296 96280
rect 115360 96270 115388 100950
rect 116202 100814 116308 100842
rect 115348 96264 115400 96270
rect 115348 96206 115400 96212
rect 116280 96202 116308 100814
rect 116372 100729 116400 101034
rect 116464 100950 116754 100978
rect 117016 100950 117306 100978
rect 117568 100950 117858 100978
rect 118120 100950 118410 100978
rect 119224 100950 119514 100978
rect 116358 100720 116414 100729
rect 116358 100655 116414 100664
rect 116372 100146 116400 100655
rect 116360 100140 116412 100146
rect 116360 100082 116412 100088
rect 116268 96196 116320 96202
rect 116268 96138 116320 96144
rect 116464 96134 116492 100950
rect 116452 96128 116504 96134
rect 116452 96070 116504 96076
rect 117016 95930 117044 100950
rect 117568 96066 117596 100950
rect 117556 96060 117608 96066
rect 117556 96002 117608 96008
rect 118120 95998 118148 100950
rect 118962 100814 119068 100842
rect 119040 97306 119068 100814
rect 118856 97278 119068 97306
rect 118108 95992 118160 95998
rect 118108 95934 118160 95940
rect 117004 95924 117056 95930
rect 117004 95866 117056 95872
rect 118856 95862 118884 97278
rect 119224 96474 119252 100950
rect 122154 100584 122210 100593
rect 122154 100519 122210 100528
rect 119212 96468 119264 96474
rect 119212 96410 119264 96416
rect 118844 95856 118896 95862
rect 118844 95798 118896 95804
rect 113672 93742 114008 93770
rect 122168 93770 122196 100519
rect 123088 97154 123116 101879
rect 123258 101400 123314 101409
rect 123258 101335 123314 101344
rect 123076 97148 123128 97154
rect 123076 97090 123128 97096
rect 123272 93770 123300 101335
rect 124456 97148 124508 97154
rect 124456 97090 124508 97096
rect 124468 93770 124496 97090
rect 124560 93906 124588 102802
rect 125756 96474 125784 135902
rect 138268 135902 138604 135930
rect 145168 135902 145228 135930
rect 151608 135902 151944 135930
rect 138268 134214 138296 135902
rect 145168 134418 145196 135902
rect 145156 134412 145208 134418
rect 145156 134354 145208 134360
rect 138256 134208 138308 134214
rect 138256 134150 138308 134156
rect 151608 133602 151636 135902
rect 149664 133596 149716 133602
rect 149664 133538 149716 133544
rect 151596 133596 151648 133602
rect 151596 133538 151648 133544
rect 149676 126818 149704 133538
rect 163108 129946 163136 136423
rect 163752 130474 163780 144855
rect 163830 143696 163886 143705
rect 163830 143631 163886 143640
rect 163740 130468 163792 130474
rect 163740 130410 163792 130416
rect 163844 130406 163872 143631
rect 167064 142889 167092 148498
rect 167156 144793 167184 149722
rect 167236 149644 167288 149650
rect 167236 149586 167288 149592
rect 167248 146833 167276 149586
rect 167340 148873 167368 151490
rect 167326 148864 167382 148873
rect 167326 148799 167382 148808
rect 167880 146856 167932 146862
rect 167234 146824 167290 146833
rect 167880 146798 167932 146804
rect 167234 146759 167290 146768
rect 167142 144784 167198 144793
rect 167142 144719 167198 144728
rect 167050 142880 167106 142889
rect 167050 142815 167106 142824
rect 164382 142472 164438 142481
rect 164382 142407 164438 142416
rect 164396 141626 164424 142407
rect 164384 141620 164436 141626
rect 164384 141562 164436 141568
rect 167052 141620 167104 141626
rect 167052 141562 167104 141568
rect 164290 141248 164346 141257
rect 164290 141183 164346 141192
rect 164304 140062 164332 141183
rect 164292 140056 164344 140062
rect 166408 140056 166460 140062
rect 164292 139998 164344 140004
rect 164382 140024 164438 140033
rect 166408 139998 166460 140004
rect 164382 139959 164384 139968
rect 164436 139959 164438 139968
rect 165856 139988 165908 139994
rect 164384 139930 164436 139936
rect 165856 139930 165908 139936
rect 163922 138800 163978 138809
rect 163922 138735 163978 138744
rect 163832 130400 163884 130406
rect 163832 130342 163884 130348
rect 163936 130338 163964 138735
rect 164750 137576 164806 137585
rect 164750 137511 164806 137520
rect 163924 130332 163976 130338
rect 163924 130274 163976 130280
rect 163108 129918 163596 129946
rect 163568 128858 163596 129918
rect 163568 128830 163872 128858
rect 163844 128722 163872 128830
rect 163844 128694 164226 128722
rect 164764 128708 164792 137511
rect 165304 130332 165356 130338
rect 165304 130274 165356 130280
rect 165316 128708 165344 130274
rect 165868 128708 165896 139930
rect 166420 128708 166448 139998
rect 167064 128708 167092 141562
rect 167892 140849 167920 146798
rect 167972 145496 168024 145502
rect 167972 145438 168024 145444
rect 167878 140840 167934 140849
rect 167878 140775 167934 140784
rect 167984 138809 168012 145438
rect 192088 139246 192116 185519
rect 188028 139240 188080 139246
rect 188026 139208 188028 139217
rect 192076 139240 192128 139246
rect 188080 139208 188082 139217
rect 192076 139182 192128 139188
rect 193456 139240 193508 139246
rect 193456 139182 193508 139188
rect 188026 139143 188082 139152
rect 167970 138800 168026 138809
rect 167970 138735 168026 138744
rect 168522 136216 168578 136225
rect 168522 136151 168578 136160
rect 168536 130950 168564 136151
rect 169260 133936 169312 133942
rect 169260 133878 169312 133884
rect 168708 133800 168760 133806
rect 168708 133742 168760 133748
rect 168524 130944 168576 130950
rect 168524 130886 168576 130892
rect 168156 130468 168208 130474
rect 168156 130410 168208 130416
rect 167604 130400 167656 130406
rect 167604 130342 167656 130348
rect 167616 128708 167644 130342
rect 168168 128708 168196 130410
rect 168720 128708 168748 133742
rect 169272 128708 169300 133878
rect 169904 133868 169956 133874
rect 169904 133810 169956 133816
rect 169916 128708 169944 133810
rect 170100 133806 170128 135916
rect 170468 133942 170496 135916
rect 170456 133936 170508 133942
rect 170456 133878 170508 133884
rect 170836 133874 170864 135916
rect 170824 133868 170876 133874
rect 170824 133810 170876 133816
rect 171296 133806 171324 135916
rect 171388 135902 171678 135930
rect 170088 133800 170140 133806
rect 170088 133742 170140 133748
rect 170456 133800 170508 133806
rect 170456 133742 170508 133748
rect 171284 133800 171336 133806
rect 171284 133742 171336 133748
rect 170468 128708 170496 133742
rect 171388 133074 171416 135902
rect 171296 133046 171416 133074
rect 171296 128722 171324 133046
rect 172032 128722 172060 135916
rect 172492 128722 172520 135916
rect 172860 128722 172888 135916
rect 171034 128694 171324 128722
rect 171586 128694 172060 128722
rect 172138 128694 172520 128722
rect 172782 128694 172888 128722
rect 173228 128722 173256 135916
rect 173688 128722 173716 135916
rect 174056 133788 174084 135916
rect 174438 135902 174544 135930
rect 174056 133760 174452 133788
rect 173228 128694 173334 128722
rect 173688 128694 173886 128722
rect 174424 128708 174452 133760
rect 174516 128722 174544 135902
rect 174884 133738 174912 135916
rect 175252 133806 175280 135916
rect 175620 133874 175648 135916
rect 175608 133868 175660 133874
rect 175608 133810 175660 133816
rect 175240 133800 175292 133806
rect 175240 133742 175292 133748
rect 174872 133732 174924 133738
rect 174872 133674 174924 133680
rect 175608 133732 175660 133738
rect 175608 133674 175660 133680
rect 174516 128694 174990 128722
rect 175620 128708 175648 133674
rect 176080 133330 176108 135916
rect 176448 133806 176476 135916
rect 176712 133868 176764 133874
rect 176712 133810 176764 133816
rect 176160 133800 176212 133806
rect 176160 133742 176212 133748
rect 176436 133800 176488 133806
rect 176436 133742 176488 133748
rect 176068 133324 176120 133330
rect 176068 133266 176120 133272
rect 176172 128708 176200 133742
rect 176724 128708 176752 133810
rect 176816 133738 176844 135916
rect 177276 133874 177304 135916
rect 177264 133868 177316 133874
rect 177264 133810 177316 133816
rect 176804 133732 176856 133738
rect 176804 133674 176856 133680
rect 177644 133534 177672 135916
rect 177816 133800 177868 133806
rect 177816 133742 177868 133748
rect 177632 133528 177684 133534
rect 177632 133470 177684 133476
rect 177264 133324 177316 133330
rect 177264 133266 177316 133272
rect 177276 128708 177304 133266
rect 177828 128708 177856 133742
rect 178104 133330 178132 135916
rect 178472 133942 178500 135916
rect 178460 133936 178512 133942
rect 178460 133878 178512 133884
rect 178460 133732 178512 133738
rect 178460 133674 178512 133680
rect 178092 133324 178144 133330
rect 178092 133266 178144 133272
rect 178472 128708 178500 133674
rect 178840 133194 178868 135916
rect 179012 133868 179064 133874
rect 179012 133810 179064 133816
rect 178828 133188 178880 133194
rect 178828 133130 178880 133136
rect 179024 128708 179052 133810
rect 179300 133262 179328 135916
rect 179564 133528 179616 133534
rect 179564 133470 179616 133476
rect 179288 133256 179340 133262
rect 179288 133198 179340 133204
rect 179576 128708 179604 133470
rect 179668 133058 179696 135916
rect 180036 133398 180064 135916
rect 180024 133392 180076 133398
rect 180024 133334 180076 133340
rect 180116 133324 180168 133330
rect 180116 133266 180168 133272
rect 179656 133052 179708 133058
rect 179656 132994 179708 133000
rect 180128 128708 180156 133266
rect 180496 133126 180524 135916
rect 180668 133936 180720 133942
rect 180668 133878 180720 133884
rect 180484 133120 180536 133126
rect 180484 133062 180536 133068
rect 180680 128708 180708 133878
rect 180864 133534 180892 135916
rect 181232 133942 181260 135916
rect 181220 133936 181272 133942
rect 181220 133878 181272 133884
rect 181692 133670 181720 135916
rect 181680 133664 181732 133670
rect 181680 133606 181732 133612
rect 180852 133528 180904 133534
rect 180852 133470 180904 133476
rect 182060 133330 182088 135916
rect 182428 134078 182456 135916
rect 182416 134072 182468 134078
rect 182416 134014 182468 134020
rect 182888 134010 182916 135916
rect 182876 134004 182928 134010
rect 182876 133946 182928 133952
rect 182508 133528 182560 133534
rect 182508 133470 182560 133476
rect 182048 133324 182100 133330
rect 182048 133266 182100 133272
rect 181864 133256 181916 133262
rect 181864 133198 181916 133204
rect 181312 133188 181364 133194
rect 181312 133130 181364 133136
rect 181324 128708 181352 133130
rect 181876 128708 181904 133198
rect 182416 133052 182468 133058
rect 182416 132994 182468 133000
rect 182428 128708 182456 132994
rect 182520 130338 182548 133470
rect 183256 133466 183284 135916
rect 183624 133806 183652 135916
rect 183612 133800 183664 133806
rect 183612 133742 183664 133748
rect 184084 133738 184112 135916
rect 184452 133874 184480 135916
rect 184716 133936 184768 133942
rect 184716 133878 184768 133884
rect 184440 133868 184492 133874
rect 184440 133810 184492 133816
rect 184072 133732 184124 133738
rect 184072 133674 184124 133680
rect 183244 133460 183296 133466
rect 183244 133402 183296 133408
rect 182968 133392 183020 133398
rect 182968 133334 183020 133340
rect 182508 130332 182560 130338
rect 182508 130274 182560 130280
rect 182980 128708 183008 133334
rect 183520 133120 183572 133126
rect 183520 133062 183572 133068
rect 183532 128708 183560 133062
rect 184164 130332 184216 130338
rect 184164 130274 184216 130280
rect 184176 128708 184204 130274
rect 184728 128708 184756 133878
rect 184820 133602 184848 135916
rect 185084 133664 185136 133670
rect 185084 133606 185136 133612
rect 184808 133596 184860 133602
rect 184808 133538 184860 133544
rect 184808 133324 184860 133330
rect 184808 133266 184860 133272
rect 184820 130338 184848 133266
rect 185096 130354 185124 133606
rect 185280 133262 185308 135916
rect 185544 133800 185596 133806
rect 185544 133742 185596 133748
rect 185268 133256 185320 133262
rect 185268 133198 185320 133204
rect 185556 132938 185584 133742
rect 185648 133058 185676 135916
rect 186372 134072 186424 134078
rect 186372 134014 186424 134020
rect 185728 133460 185780 133466
rect 185728 133402 185780 133408
rect 185636 133052 185688 133058
rect 185636 132994 185688 133000
rect 185556 132910 185676 132938
rect 185648 130610 185676 132910
rect 185636 130604 185688 130610
rect 185636 130546 185688 130552
rect 185740 130542 185768 133402
rect 185728 130536 185780 130542
rect 185728 130478 185780 130484
rect 184808 130332 184860 130338
rect 185096 130326 185216 130354
rect 184808 130274 184860 130280
rect 185188 128722 185216 130326
rect 185820 130332 185872 130338
rect 185820 130274 185872 130280
rect 185188 128694 185294 128722
rect 185832 128708 185860 130274
rect 186384 128708 186412 134014
rect 186464 134004 186516 134010
rect 186464 133946 186516 133952
rect 186476 130354 186504 133946
rect 186832 133868 186884 133874
rect 186832 133810 186884 133816
rect 186648 133732 186700 133738
rect 186648 133674 186700 133680
rect 186660 130406 186688 133674
rect 186844 130474 186872 133810
rect 187292 133596 187344 133602
rect 187292 133538 187344 133544
rect 186832 130468 186884 130474
rect 186832 130410 186884 130416
rect 186648 130400 186700 130406
rect 186476 130326 186596 130354
rect 186648 130342 186700 130348
rect 187304 130338 187332 133538
rect 190420 133256 190472 133262
rect 190420 133198 190472 133204
rect 188120 130604 188172 130610
rect 188120 130546 188172 130552
rect 187568 130536 187620 130542
rect 187568 130478 187620 130484
rect 186568 128858 186596 130326
rect 187292 130332 187344 130338
rect 187292 130274 187344 130280
rect 186568 128830 186688 128858
rect 186660 128722 186688 128830
rect 186660 128694 187042 128722
rect 187580 128708 187608 130478
rect 188132 128708 188160 130546
rect 189224 130468 189276 130474
rect 189224 130410 189276 130416
rect 188672 130400 188724 130406
rect 188672 130342 188724 130348
rect 188684 128708 188712 130342
rect 189236 128708 189264 130410
rect 189868 130332 189920 130338
rect 189868 130274 189920 130280
rect 189880 128708 189908 130274
rect 190432 128708 190460 133198
rect 190972 133052 191024 133058
rect 190972 132994 191024 133000
rect 190984 128708 191012 132994
rect 191524 130944 191576 130950
rect 191524 130886 191576 130892
rect 191536 128708 191564 130886
rect 160334 128192 160390 128201
rect 160334 128127 160390 128136
rect 160150 127648 160206 127657
rect 160150 127583 160206 127592
rect 149414 126790 149704 126818
rect 160058 126560 160114 126569
rect 160058 126495 160114 126504
rect 160072 124665 160100 126495
rect 160164 125889 160192 127583
rect 160242 126424 160298 126433
rect 160348 126410 160376 128127
rect 160426 126968 160482 126977
rect 160426 126903 160482 126912
rect 160298 126382 160376 126410
rect 160242 126359 160298 126368
rect 160242 126152 160298 126161
rect 160242 126087 160298 126096
rect 160150 125880 160206 125889
rect 160150 125815 160206 125824
rect 160256 125322 160284 126087
rect 160164 125294 160284 125322
rect 160058 124656 160114 124665
rect 160058 124591 160114 124600
rect 160164 124121 160192 125294
rect 160242 125200 160298 125209
rect 160440 125186 160468 126903
rect 160298 125158 160468 125186
rect 160518 125200 160574 125209
rect 160242 125135 160298 125144
rect 160518 125135 160574 125144
rect 160242 124928 160298 124937
rect 160242 124863 160298 124872
rect 160150 124112 160206 124121
rect 160150 124047 160206 124056
rect 160058 123568 160114 123577
rect 160256 123554 160284 124863
rect 160532 124234 160560 125135
rect 160058 123503 160114 123512
rect 160164 123526 160284 123554
rect 160348 124206 160560 124234
rect 160072 121673 160100 123503
rect 160164 122897 160192 123526
rect 160242 123432 160298 123441
rect 160348 123418 160376 124206
rect 160426 124112 160482 124121
rect 160426 124047 160482 124056
rect 160298 123390 160376 123418
rect 160242 123367 160298 123376
rect 160440 123010 160468 124047
rect 160256 122982 160468 123010
rect 160150 122888 160206 122897
rect 160150 122823 160206 122832
rect 160256 122761 160284 122982
rect 160426 122888 160482 122897
rect 160426 122823 160482 122832
rect 160242 122752 160298 122761
rect 160242 122687 160298 122696
rect 160242 122344 160298 122353
rect 160242 122279 160298 122288
rect 160150 122072 160206 122081
rect 160150 122007 160206 122016
rect 160058 121664 160114 121673
rect 160058 121599 160114 121608
rect 160164 121378 160192 122007
rect 160072 121350 160192 121378
rect 159966 121256 160022 121265
rect 159966 121191 160022 121200
rect 159874 119352 159930 119361
rect 159874 119287 159930 119296
rect 159888 116913 159916 119287
rect 159980 119225 160008 121191
rect 160072 119905 160100 121350
rect 160256 121242 160284 122279
rect 160164 121214 160284 121242
rect 160164 120449 160192 121214
rect 160242 121120 160298 121129
rect 160242 121055 160298 121064
rect 160256 120970 160284 121055
rect 160440 120970 160468 122823
rect 160256 120942 160468 120970
rect 160242 120712 160298 120721
rect 160242 120647 160298 120656
rect 160150 120440 160206 120449
rect 160150 120375 160206 120384
rect 160058 119896 160114 119905
rect 160058 119831 160114 119840
rect 160150 119488 160206 119497
rect 160150 119423 160206 119432
rect 159966 119216 160022 119225
rect 159966 119151 160022 119160
rect 160058 118264 160114 118273
rect 160058 118199 160114 118208
rect 159874 116904 159930 116913
rect 159874 116839 159930 116848
rect 160072 116233 160100 118199
rect 160164 117457 160192 119423
rect 160256 118681 160284 120647
rect 160334 120032 160390 120041
rect 160334 119967 160390 119976
rect 160242 118672 160298 118681
rect 160242 118607 160298 118616
rect 160242 118128 160298 118137
rect 160348 118114 160376 119967
rect 160298 118086 160376 118114
rect 160242 118063 160298 118072
rect 160242 117992 160298 118001
rect 160242 117927 160298 117936
rect 160150 117448 160206 117457
rect 160150 117383 160206 117392
rect 160256 116618 160284 117927
rect 160426 117040 160482 117049
rect 160426 116975 160482 116984
rect 160164 116590 160284 116618
rect 160058 116224 160114 116233
rect 160058 116159 160114 116168
rect 160164 115689 160192 116590
rect 160242 116496 160298 116505
rect 160242 116431 160298 116440
rect 160150 115680 160206 115689
rect 160150 115615 160206 115624
rect 160058 115408 160114 115417
rect 160058 115343 160114 115352
rect 159048 115168 159100 115174
rect 159048 115110 159100 115116
rect 159060 112697 159088 115110
rect 160072 113241 160100 115343
rect 160256 114465 160284 116431
rect 160334 115952 160390 115961
rect 160334 115887 160390 115896
rect 160242 114456 160298 114465
rect 160242 114391 160298 114400
rect 160242 114320 160298 114329
rect 160348 114306 160376 115887
rect 160440 115145 160468 116975
rect 160612 115168 160664 115174
rect 160426 115136 160482 115145
rect 160426 115071 160482 115080
rect 160610 115136 160612 115145
rect 160664 115136 160666 115145
rect 160610 115071 160666 115080
rect 160298 114278 160376 114306
rect 160242 114255 160298 114264
rect 160242 114184 160298 114193
rect 160242 114119 160298 114128
rect 160150 113776 160206 113785
rect 160150 113711 160206 113720
rect 160058 113232 160114 113241
rect 160058 113167 160114 113176
rect 159966 112960 160022 112969
rect 159966 112895 160022 112904
rect 159046 112688 159102 112697
rect 159046 112623 159102 112632
rect 159874 111056 159930 111065
rect 159874 110991 159930 111000
rect 159888 108481 159916 110991
rect 159980 110929 160008 112895
rect 160058 112416 160114 112425
rect 160058 112351 160114 112360
rect 159966 110920 160022 110929
rect 159966 110855 160022 110864
rect 160072 110249 160100 112351
rect 160164 111473 160192 113711
rect 160256 112153 160284 114119
rect 160242 112144 160298 112153
rect 160242 112079 160298 112088
rect 160334 111872 160390 111881
rect 160334 111807 160390 111816
rect 160150 111464 160206 111473
rect 160150 111399 160206 111408
rect 160242 111192 160298 111201
rect 160242 111127 160298 111136
rect 160058 110240 160114 110249
rect 160058 110175 160114 110184
rect 160150 110104 160206 110113
rect 160150 110039 160206 110048
rect 159966 109832 160022 109841
rect 159966 109767 160022 109776
rect 159874 108472 159930 108481
rect 159874 108407 159930 108416
rect 159980 107257 160008 109767
rect 160058 108880 160114 108889
rect 160058 108815 160114 108824
rect 159966 107248 160022 107257
rect 159966 107183 160022 107192
rect 159874 106840 159930 106849
rect 159874 106775 159930 106784
rect 159888 104265 159916 106775
rect 160072 106713 160100 108815
rect 160164 107937 160192 110039
rect 160256 109161 160284 111127
rect 160348 109705 160376 111807
rect 160334 109696 160390 109705
rect 160334 109631 160390 109640
rect 160242 109152 160298 109161
rect 160242 109087 160298 109096
rect 160242 108336 160298 108345
rect 160242 108271 160298 108280
rect 160150 107928 160206 107937
rect 160150 107863 160206 107872
rect 160150 107112 160206 107121
rect 160150 107047 160206 107056
rect 160058 106704 160114 106713
rect 160058 106639 160114 106648
rect 160058 106024 160114 106033
rect 160058 105959 160114 105968
rect 159966 105616 160022 105625
rect 159966 105551 160022 105560
rect 159874 104256 159930 104265
rect 159874 104191 159930 104200
rect 126940 104152 126992 104158
rect 126940 104094 126992 104100
rect 125928 102792 125980 102798
rect 125928 102734 125980 102740
rect 125744 96468 125796 96474
rect 125744 96410 125796 96416
rect 125940 95402 125968 102734
rect 126952 97086 126980 104094
rect 127032 104084 127084 104090
rect 127032 104026 127084 104032
rect 157576 104084 157628 104090
rect 157576 104026 157628 104032
rect 126940 97080 126992 97086
rect 126940 97022 126992 97028
rect 127044 96882 127072 104026
rect 127124 102792 127176 102798
rect 127124 102734 127176 102740
rect 127136 97154 127164 102734
rect 127596 101098 127624 102868
rect 128976 101302 129004 102868
rect 128964 101296 129016 101302
rect 128964 101238 129016 101244
rect 127584 101092 127636 101098
rect 127584 101034 127636 101040
rect 127596 100622 127624 101034
rect 127584 100616 127636 100622
rect 127584 100558 127636 100564
rect 130448 99942 130476 102868
rect 131828 99942 131856 102868
rect 133300 99942 133328 102868
rect 134680 99942 134708 102868
rect 136048 100004 136100 100010
rect 136048 99946 136100 99952
rect 130436 99936 130488 99942
rect 130436 99878 130488 99884
rect 131264 99936 131316 99942
rect 131264 99878 131316 99884
rect 131816 99936 131868 99942
rect 131816 99878 131868 99884
rect 132552 99936 132604 99942
rect 132552 99878 132604 99884
rect 133288 99936 133340 99942
rect 133288 99878 133340 99884
rect 133840 99936 133892 99942
rect 133840 99878 133892 99884
rect 134668 99936 134720 99942
rect 134668 99878 134720 99884
rect 134944 99936 134996 99942
rect 134944 99878 134996 99884
rect 127124 97148 127176 97154
rect 127124 97090 127176 97096
rect 127676 97148 127728 97154
rect 127676 97090 127728 97096
rect 127032 96876 127084 96882
rect 127032 96818 127084 96824
rect 125940 95374 126336 95402
rect 124560 93878 125508 93906
rect 125480 93770 125508 93878
rect 122168 93742 122504 93770
rect 123272 93742 123608 93770
rect 124468 93742 124712 93770
rect 125480 93742 125816 93770
rect 126308 93634 126336 95374
rect 127688 93770 127716 97090
rect 129976 97080 130028 97086
rect 129976 97022 130028 97028
rect 128780 96876 128832 96882
rect 128780 96818 128832 96824
rect 128792 93770 128820 96818
rect 129988 93770 130016 97022
rect 131276 93770 131304 99878
rect 132564 93770 132592 99878
rect 133852 93770 133880 99878
rect 134956 93770 134984 99878
rect 136060 93770 136088 99946
rect 136152 99942 136180 102868
rect 137532 100010 137560 102868
rect 137520 100004 137572 100010
rect 137520 99946 137572 99952
rect 138164 100004 138216 100010
rect 138164 99946 138216 99952
rect 136140 99936 136192 99942
rect 136140 99878 136192 99884
rect 137244 99936 137296 99942
rect 137244 99878 137296 99884
rect 137256 93770 137284 99878
rect 138176 93770 138204 99946
rect 139004 99942 139032 102868
rect 140384 100010 140412 102868
rect 141660 100072 141712 100078
rect 141660 100014 141712 100020
rect 140372 100004 140424 100010
rect 140372 99946 140424 99952
rect 140556 100004 140608 100010
rect 140556 99946 140608 99952
rect 138992 99936 139044 99942
rect 138992 99878 139044 99884
rect 139452 99936 139504 99942
rect 139452 99878 139504 99884
rect 139464 93770 139492 99878
rect 140568 93770 140596 99946
rect 141672 93770 141700 100014
rect 141856 99942 141884 102868
rect 143236 100010 143264 102868
rect 144708 100078 144736 102868
rect 145984 100208 146036 100214
rect 145984 100150 146036 100156
rect 144972 100140 145024 100146
rect 144972 100082 145024 100088
rect 144696 100072 144748 100078
rect 144696 100014 144748 100020
rect 143224 100004 143276 100010
rect 143224 99946 143276 99952
rect 143684 100004 143736 100010
rect 143684 99946 143736 99952
rect 141844 99936 141896 99942
rect 141844 99878 141896 99884
rect 142764 99936 142816 99942
rect 142764 99878 142816 99884
rect 142776 93770 142804 99878
rect 143696 93770 143724 99946
rect 144984 93770 145012 100082
rect 145996 93770 146024 100150
rect 146088 99942 146116 102868
rect 147560 100010 147588 102868
rect 148940 100146 148968 102868
rect 150412 100214 150440 102868
rect 150400 100208 150452 100214
rect 150400 100150 150452 100156
rect 148928 100140 148980 100146
rect 148928 100082 148980 100088
rect 148284 100072 148336 100078
rect 148284 100014 148336 100020
rect 147548 100004 147600 100010
rect 147548 99946 147600 99952
rect 146076 99936 146128 99942
rect 146076 99878 146128 99884
rect 147180 99936 147232 99942
rect 147180 99878 147232 99884
rect 147192 93770 147220 99878
rect 148296 93770 148324 100014
rect 151792 99942 151820 102868
rect 152792 101432 152844 101438
rect 152792 101374 152844 101380
rect 151780 99936 151832 99942
rect 151780 99878 151832 99884
rect 148836 96468 148888 96474
rect 148836 96410 148888 96416
rect 151688 96468 151740 96474
rect 151688 96410 151740 96416
rect 127688 93742 128024 93770
rect 128792 93742 129128 93770
rect 129988 93742 130232 93770
rect 131276 93742 131336 93770
rect 132440 93742 132592 93770
rect 133544 93742 133880 93770
rect 134648 93742 134984 93770
rect 135844 93742 136088 93770
rect 136948 93742 137284 93770
rect 138052 93742 138204 93770
rect 139156 93742 139492 93770
rect 140260 93742 140596 93770
rect 141364 93742 141700 93770
rect 142468 93742 142804 93770
rect 143572 93742 143724 93770
rect 144676 93742 145012 93770
rect 145780 93742 146024 93770
rect 146884 93742 147220 93770
rect 147988 93742 148324 93770
rect 148848 93770 148876 96410
rect 151700 93770 151728 96410
rect 152804 93770 152832 101374
rect 153264 100078 153292 102868
rect 153896 101364 153948 101370
rect 153896 101306 153948 101312
rect 153252 100072 153304 100078
rect 153252 100014 153304 100020
rect 153908 93770 153936 101306
rect 154644 99942 154672 102868
rect 154632 99936 154684 99942
rect 154632 99878 154684 99884
rect 154632 97148 154684 97154
rect 154632 97090 154684 97096
rect 148848 93742 149184 93770
rect 151392 93742 151728 93770
rect 152496 93742 152832 93770
rect 153600 93742 153936 93770
rect 154644 93634 154672 97090
rect 156104 96332 156156 96338
rect 156104 96274 156156 96280
rect 156116 93770 156144 96274
rect 157208 96264 157260 96270
rect 157208 96206 157260 96212
rect 157220 93770 157248 96206
rect 155808 93742 156144 93770
rect 156912 93742 157248 93770
rect 157588 93770 157616 104026
rect 159980 103177 160008 105551
rect 160072 103993 160100 105959
rect 160164 104945 160192 107047
rect 160256 106169 160284 108271
rect 160334 107792 160390 107801
rect 160334 107727 160390 107736
rect 160242 106160 160298 106169
rect 160242 106095 160298 106104
rect 160242 105480 160298 105489
rect 160348 105466 160376 107727
rect 193468 106169 193496 139182
rect 193546 123568 193602 123577
rect 193546 123503 193602 123512
rect 193454 106160 193510 106169
rect 193454 106095 193510 106104
rect 160298 105438 160376 105466
rect 160242 105415 160298 105424
rect 160150 104936 160206 104945
rect 160150 104871 160206 104880
rect 161530 104800 161586 104809
rect 161530 104735 161586 104744
rect 160334 104256 160390 104265
rect 160334 104191 160390 104200
rect 160348 104090 160376 104191
rect 160336 104084 160388 104090
rect 160336 104026 160388 104032
rect 160058 103984 160114 103993
rect 160058 103919 160114 103928
rect 160150 103712 160206 103721
rect 160150 103647 160206 103656
rect 159966 103168 160022 103177
rect 159966 103103 160022 103112
rect 160164 96270 160192 103647
rect 160242 103032 160298 103041
rect 160242 102967 160298 102976
rect 160256 96338 160284 102967
rect 160518 102760 160574 102769
rect 160518 102695 160574 102704
rect 160334 101944 160390 101953
rect 160334 101879 160390 101888
rect 160348 101370 160376 101879
rect 160426 101536 160482 101545
rect 160426 101471 160482 101480
rect 160440 101438 160468 101471
rect 160428 101432 160480 101438
rect 160428 101374 160480 101380
rect 160336 101364 160388 101370
rect 160336 101306 160388 101312
rect 160334 100584 160390 100593
rect 160334 100519 160390 100528
rect 160348 96474 160376 100519
rect 160532 97154 160560 102695
rect 160980 99936 161032 99942
rect 160980 99878 161032 99884
rect 160520 97148 160572 97154
rect 160520 97090 160572 97096
rect 160336 96468 160388 96474
rect 160336 96410 160388 96416
rect 160244 96332 160296 96338
rect 160244 96274 160296 96280
rect 160152 96264 160204 96270
rect 160152 96206 160204 96212
rect 159416 95992 159468 95998
rect 159416 95934 159468 95940
rect 159428 93770 159456 95934
rect 157588 93742 158016 93770
rect 159120 93742 159456 93770
rect 160992 93770 161020 99878
rect 161544 95998 161572 104735
rect 170482 100950 170956 100978
rect 171586 100950 171876 100978
rect 172138 100950 172520 100978
rect 163108 100814 164226 100842
rect 164580 100814 164778 100842
rect 161532 95992 161584 95998
rect 161532 95934 161584 95940
rect 160992 93742 161328 93770
rect 126308 93606 126920 93634
rect 154644 93606 154704 93634
rect 100884 93470 101036 93498
rect 95290 92560 95346 92569
rect 95290 92495 95346 92504
rect 95304 91714 95332 92495
rect 118936 92320 118988 92326
rect 118936 92262 118988 92268
rect 95292 91708 95344 91714
rect 95292 91650 95344 91656
rect 93360 91368 93412 91374
rect 93360 91310 93412 91316
rect 95382 90248 95438 90257
rect 95382 90183 95438 90192
rect 95396 88926 95424 90183
rect 95384 88920 95436 88926
rect 95384 88862 95436 88868
rect 95382 87936 95438 87945
rect 95382 87871 95438 87880
rect 95396 87566 95424 87871
rect 95384 87560 95436 87566
rect 95384 87502 95436 87508
rect 118948 87265 118976 92262
rect 118934 87256 118990 87265
rect 118934 87191 118990 87200
rect 92806 87120 92862 87129
rect 92806 87055 92862 87064
rect 94278 85488 94334 85497
rect 94278 85423 94334 85432
rect 92254 82224 92310 82233
rect 92254 82159 92310 82168
rect 92162 81136 92218 81145
rect 92162 81071 92218 81080
rect 94292 80562 94320 85423
rect 163108 84681 163136 100814
rect 163832 97352 163884 97358
rect 163832 97294 163884 97300
rect 163740 97284 163792 97290
rect 163740 97226 163792 97232
rect 163556 91164 163608 91170
rect 163556 91106 163608 91112
rect 163568 90801 163596 91106
rect 163554 90792 163610 90801
rect 163554 90727 163610 90736
rect 163464 88784 163516 88790
rect 163464 88726 163516 88732
rect 163476 88353 163504 88726
rect 163462 88344 163518 88353
rect 163462 88279 163518 88288
rect 163752 87129 163780 97226
rect 163844 92025 163872 97294
rect 164108 94360 164160 94366
rect 164108 94302 164160 94308
rect 164120 93249 164148 94302
rect 164106 93240 164162 93249
rect 164106 93175 164162 93184
rect 163830 92016 163886 92025
rect 163830 91951 163886 91960
rect 163832 90144 163884 90150
rect 163832 90086 163884 90092
rect 163844 89577 163872 90086
rect 163830 89568 163886 89577
rect 163830 89503 163886 89512
rect 163738 87120 163794 87129
rect 163738 87055 163794 87064
rect 164580 85905 164608 100814
rect 165316 97290 165344 100828
rect 165304 97284 165356 97290
rect 165304 97226 165356 97232
rect 165868 97222 165896 100828
rect 166052 100814 166434 100842
rect 166696 100814 167078 100842
rect 165120 97216 165172 97222
rect 165120 97158 165172 97164
rect 165856 97216 165908 97222
rect 165856 97158 165908 97164
rect 165132 88790 165160 97158
rect 165948 96944 166000 96950
rect 165948 96886 166000 96892
rect 165960 91170 165988 96886
rect 165948 91164 166000 91170
rect 165948 91106 166000 91112
rect 166052 90150 166080 100814
rect 166696 96950 166724 100814
rect 167616 97358 167644 100828
rect 167604 97352 167656 97358
rect 167604 97294 167656 97300
rect 166684 96944 166736 96950
rect 166684 96886 166736 96892
rect 168168 94366 168196 100828
rect 168524 97828 168576 97834
rect 168524 97770 168576 97776
rect 168156 94360 168208 94366
rect 168156 94302 168208 94308
rect 168536 92841 168564 97770
rect 168720 97222 168748 100828
rect 169272 97358 169300 100828
rect 169260 97352 169312 97358
rect 169260 97294 169312 97300
rect 169916 97290 169944 100828
rect 170456 97352 170508 97358
rect 170456 97294 170508 97300
rect 169904 97284 169956 97290
rect 169904 97226 169956 97232
rect 168708 97216 168760 97222
rect 168708 97158 168760 97164
rect 170088 97216 170140 97222
rect 170088 97158 170140 97164
rect 170100 93756 170128 97158
rect 170468 93756 170496 97294
rect 170824 97284 170876 97290
rect 170824 97226 170876 97232
rect 170836 93756 170864 97226
rect 170928 93770 170956 100950
rect 171020 98174 171048 100828
rect 171008 98168 171060 98174
rect 171008 98110 171060 98116
rect 171652 98168 171704 98174
rect 171652 98110 171704 98116
rect 170928 93742 171310 93770
rect 171664 93756 171692 98110
rect 171848 93770 171876 100950
rect 171848 93742 172046 93770
rect 172492 93756 172520 100950
rect 172768 93770 172796 100828
rect 173320 93770 173348 100828
rect 173872 93770 173900 100828
rect 174148 100814 174438 100842
rect 174700 100814 174990 100842
rect 175528 100814 175634 100842
rect 174148 97034 174176 100814
rect 172768 93742 172874 93770
rect 173242 93742 173348 93770
rect 173702 93742 173900 93770
rect 174056 97006 174176 97034
rect 174056 93756 174084 97006
rect 174700 93770 174728 100814
rect 175528 96898 175556 100814
rect 176068 97080 176120 97086
rect 176068 97022 176120 97028
rect 175160 96870 175556 96898
rect 175160 93770 175188 96870
rect 175240 96808 175292 96814
rect 175240 96750 175292 96756
rect 174438 93742 174728 93770
rect 174898 93742 175188 93770
rect 175252 93756 175280 96750
rect 175608 96672 175660 96678
rect 175608 96614 175660 96620
rect 175620 93756 175648 96614
rect 176080 93756 176108 97022
rect 176172 96814 176200 100828
rect 176436 97148 176488 97154
rect 176436 97090 176488 97096
rect 176160 96808 176212 96814
rect 176160 96750 176212 96756
rect 176448 93756 176476 97090
rect 176724 96678 176752 100828
rect 176896 97216 176948 97222
rect 176896 97158 176948 97164
rect 176908 97034 176936 97158
rect 177276 97086 177304 100828
rect 177828 97154 177856 100828
rect 178472 97222 178500 100828
rect 178460 97216 178512 97222
rect 178460 97158 178512 97164
rect 177816 97148 177868 97154
rect 177816 97090 177868 97096
rect 178092 97148 178144 97154
rect 178092 97090 178144 97096
rect 176816 97006 176936 97034
rect 177264 97080 177316 97086
rect 177264 97022 177316 97028
rect 177632 97080 177684 97086
rect 177632 97022 177684 97028
rect 176712 96672 176764 96678
rect 176712 96614 176764 96620
rect 176816 93756 176844 97006
rect 177264 96944 177316 96950
rect 177264 96886 177316 96892
rect 177276 93756 177304 96886
rect 177644 93756 177672 97022
rect 178104 93756 178132 97090
rect 178460 97012 178512 97018
rect 178460 96954 178512 96960
rect 178472 93756 178500 96954
rect 179024 96950 179052 100828
rect 179576 97086 179604 100828
rect 179748 97692 179800 97698
rect 179748 97634 179800 97640
rect 179656 97148 179708 97154
rect 179656 97090 179708 97096
rect 179564 97080 179616 97086
rect 179564 97022 179616 97028
rect 179012 96944 179064 96950
rect 179012 96886 179064 96892
rect 178828 95924 178880 95930
rect 178828 95866 178880 95872
rect 178840 93756 178868 95866
rect 179288 95856 179340 95862
rect 179288 95798 179340 95804
rect 179300 93756 179328 95798
rect 179668 93756 179696 97090
rect 179760 95862 179788 97634
rect 180128 97222 180156 100828
rect 180116 97216 180168 97222
rect 180116 97158 180168 97164
rect 180024 97080 180076 97086
rect 180024 97022 180076 97028
rect 179748 95856 179800 95862
rect 179748 95798 179800 95804
rect 180036 93756 180064 97022
rect 180680 97018 180708 100828
rect 181048 100814 181338 100842
rect 181048 97170 181076 100814
rect 181876 97698 181904 100828
rect 182232 98168 182284 98174
rect 182232 98110 182284 98116
rect 181864 97692 181916 97698
rect 181864 97634 181916 97640
rect 181588 97556 181640 97562
rect 181588 97498 181640 97504
rect 180956 97142 181076 97170
rect 181600 97154 181628 97498
rect 181588 97148 181640 97154
rect 180668 97012 180720 97018
rect 180668 96954 180720 96960
rect 180484 96808 180536 96814
rect 180484 96750 180536 96756
rect 180496 93756 180524 96750
rect 180852 96604 180904 96610
rect 180852 96546 180904 96552
rect 180864 93756 180892 96546
rect 180956 95930 180984 97142
rect 181588 97090 181640 97096
rect 181220 97012 181272 97018
rect 181220 96954 181272 96960
rect 180944 95924 180996 95930
rect 180944 95866 180996 95872
rect 181232 93756 181260 96954
rect 182048 96944 182100 96950
rect 182048 96886 182100 96892
rect 181680 96740 181732 96746
rect 181680 96682 181732 96688
rect 181692 93756 181720 96682
rect 182060 93756 182088 96886
rect 182244 96814 182272 98110
rect 182428 97562 182456 100828
rect 182416 97556 182468 97562
rect 182416 97498 182468 97504
rect 182980 97222 183008 100828
rect 183532 98174 183560 100828
rect 183520 98168 183572 98174
rect 183520 98110 183572 98116
rect 182968 97216 183020 97222
rect 182968 97158 183020 97164
rect 184072 97012 184124 97018
rect 184072 96954 184124 96960
rect 182232 96808 182284 96814
rect 182232 96750 182284 96756
rect 182876 96808 182928 96814
rect 182876 96750 182928 96756
rect 182416 96536 182468 96542
rect 182416 96478 182468 96484
rect 182428 93756 182456 96478
rect 182888 93756 182916 96750
rect 183612 95992 183664 95998
rect 183612 95934 183664 95940
rect 183244 95924 183296 95930
rect 183244 95866 183296 95872
rect 183256 93756 183284 95866
rect 183624 93756 183652 95934
rect 184084 93756 184112 96954
rect 184176 96610 184204 100828
rect 184440 97284 184492 97290
rect 184440 97226 184492 97232
rect 184164 96604 184216 96610
rect 184164 96546 184216 96552
rect 184452 96542 184480 97226
rect 184728 97222 184756 100828
rect 185188 100814 185294 100842
rect 184716 97216 184768 97222
rect 184716 97158 184768 97164
rect 184808 97148 184860 97154
rect 184808 97090 184860 97096
rect 184440 96536 184492 96542
rect 184440 96478 184492 96484
rect 184440 96128 184492 96134
rect 184440 96070 184492 96076
rect 184452 93756 184480 96070
rect 184820 93756 184848 97090
rect 185188 96746 185216 100814
rect 185636 97080 185688 97086
rect 185636 97022 185688 97028
rect 185268 96876 185320 96882
rect 185268 96818 185320 96824
rect 185176 96740 185228 96746
rect 185176 96682 185228 96688
rect 185280 93756 185308 96818
rect 185648 93756 185676 97022
rect 185832 96950 185860 100828
rect 186384 97290 186412 100828
rect 186372 97284 186424 97290
rect 186372 97226 186424 97232
rect 185820 96944 185872 96950
rect 185820 96886 185872 96892
rect 187028 96814 187056 100828
rect 187016 96808 187068 96814
rect 187016 96750 187068 96756
rect 187580 95930 187608 100828
rect 188132 95998 188160 100828
rect 188684 97018 188712 100828
rect 188672 97012 188724 97018
rect 188672 96954 188724 96960
rect 189236 96134 189264 100828
rect 189880 97154 189908 100828
rect 189868 97148 189920 97154
rect 189868 97090 189920 97096
rect 190432 96882 190460 100828
rect 190604 100616 190656 100622
rect 190604 100558 190656 100564
rect 190420 96876 190472 96882
rect 190420 96818 190472 96824
rect 189224 96128 189276 96134
rect 189224 96070 189276 96076
rect 188120 95992 188172 95998
rect 188120 95934 188172 95940
rect 187568 95924 187620 95930
rect 187568 95866 187620 95872
rect 168522 92832 168578 92841
rect 168522 92767 168578 92776
rect 188120 91640 188172 91646
rect 188120 91582 188172 91588
rect 188132 90529 188160 91582
rect 188118 90520 188174 90529
rect 188118 90455 188174 90464
rect 188580 90280 188632 90286
rect 188580 90222 188632 90228
rect 166040 90144 166092 90150
rect 166040 90086 166092 90092
rect 165120 88784 165172 88790
rect 165120 88726 165172 88732
rect 167326 88072 167382 88081
rect 167326 88007 167382 88016
rect 164566 85896 164622 85905
rect 164566 85831 164622 85840
rect 167234 84808 167290 84817
rect 167234 84743 167290 84752
rect 163094 84672 163150 84681
rect 163094 84607 163150 84616
rect 163924 84364 163976 84370
rect 163924 84306 163976 84312
rect 116542 83856 116598 83865
rect 116542 83791 116598 83800
rect 116556 83622 116584 83791
rect 116544 83616 116596 83622
rect 116544 83558 116596 83564
rect 119580 83616 119632 83622
rect 119580 83558 119632 83564
rect 95290 83176 95346 83185
rect 95290 83111 95346 83120
rect 91796 80556 91848 80562
rect 91796 80498 91848 80504
rect 94280 80556 94332 80562
rect 94280 80498 94332 80504
rect 91808 79921 91836 80498
rect 91794 79912 91850 79921
rect 91794 79847 91850 79856
rect 95304 78862 95332 83111
rect 95382 80864 95438 80873
rect 95382 80799 95438 80808
rect 91428 78856 91480 78862
rect 91428 78798 91480 78804
rect 95292 78856 95344 78862
rect 95292 78798 95344 78804
rect 91440 78697 91468 78798
rect 91426 78688 91482 78697
rect 91426 78623 91482 78632
rect 94922 78416 94978 78425
rect 94922 78351 94978 78360
rect 91704 77496 91756 77502
rect 91702 77464 91704 77473
rect 91756 77464 91758 77473
rect 91702 77399 91758 77408
rect 94936 76278 94964 78351
rect 95396 77502 95424 80799
rect 95384 77496 95436 77502
rect 95384 77438 95436 77444
rect 91704 76272 91756 76278
rect 91702 76240 91704 76249
rect 94924 76272 94976 76278
rect 91756 76240 91758 76249
rect 94924 76214 94976 76220
rect 91702 76175 91758 76184
rect 15436 75048 15488 75054
rect 15436 74990 15488 74996
rect 22336 75048 22388 75054
rect 22336 74990 22388 74996
rect 45060 75048 45112 75054
rect 45060 74990 45112 74996
rect 47820 75048 47872 75054
rect 47820 74990 47872 74996
rect 22348 73801 22376 74990
rect 47832 73937 47860 74990
rect 119592 73937 119620 83558
rect 163936 83457 163964 84306
rect 163922 83448 163978 83457
rect 163922 83383 163978 83392
rect 163924 82732 163976 82738
rect 163924 82674 163976 82680
rect 163936 82233 163964 82674
rect 163922 82224 163978 82233
rect 163922 82159 163978 82168
rect 167248 81990 167276 84743
rect 167340 84370 167368 88007
rect 167878 86168 167934 86177
rect 167878 86103 167934 86112
rect 167328 84364 167380 84370
rect 167328 84306 167380 84312
rect 167892 82738 167920 86103
rect 188120 84704 188172 84710
rect 188120 84646 188172 84652
rect 188132 83865 188160 84646
rect 188118 83856 188174 83865
rect 188118 83791 188174 83800
rect 167880 82732 167932 82738
rect 167880 82674 167932 82680
rect 167326 82088 167382 82097
rect 167326 82023 167382 82032
rect 163556 81984 163608 81990
rect 163556 81926 163608 81932
rect 167236 81984 167288 81990
rect 167236 81926 167288 81932
rect 163568 81145 163596 81926
rect 163554 81136 163610 81145
rect 163554 81071 163610 81080
rect 167234 80864 167290 80873
rect 167234 80799 167290 80808
rect 164108 80488 164160 80494
rect 164108 80430 164160 80436
rect 164120 79921 164148 80430
rect 164106 79912 164162 79921
rect 164106 79847 164162 79856
rect 167248 78998 167276 80799
rect 167340 80494 167368 82023
rect 167328 80488 167380 80494
rect 167328 80430 167380 80436
rect 164384 78992 164436 78998
rect 164384 78934 164436 78940
rect 167236 78992 167288 78998
rect 167236 78934 167288 78940
rect 164396 78697 164424 78934
rect 164382 78688 164438 78697
rect 164382 78623 164438 78632
rect 167234 78144 167290 78153
rect 167234 78079 167290 78088
rect 167248 77910 167276 78079
rect 167236 77904 167288 77910
rect 167236 77846 167288 77852
rect 164108 77836 164160 77842
rect 164108 77778 164160 77784
rect 164120 77473 164148 77778
rect 164106 77464 164162 77473
rect 164106 77399 164162 77408
rect 188592 77201 188620 90222
rect 188578 77192 188634 77201
rect 188578 77127 188634 77136
rect 167234 76512 167290 76521
rect 167234 76447 167236 76456
rect 167288 76447 167290 76456
rect 167236 76418 167288 76424
rect 163740 76408 163792 76414
rect 163740 76350 163792 76356
rect 163752 76249 163780 76350
rect 163738 76240 163794 76249
rect 163738 76175 163794 76184
rect 164106 75016 164162 75025
rect 164106 74951 164108 74960
rect 164160 74951 164162 74960
rect 167236 74980 167288 74986
rect 164108 74922 164160 74928
rect 167236 74922 167288 74928
rect 167248 74889 167276 74922
rect 167234 74880 167290 74889
rect 167234 74815 167290 74824
rect 47818 73928 47874 73937
rect 47818 73863 47874 73872
rect 119578 73928 119634 73937
rect 119578 73863 119634 73872
rect 22334 73792 22390 73801
rect 22334 73727 22390 73736
rect 164382 73792 164438 73801
rect 164382 73727 164384 73736
rect 164436 73727 164438 73736
rect 167144 73756 167196 73762
rect 164384 73698 164436 73704
rect 167144 73698 167196 73704
rect 167156 72849 167184 73698
rect 167142 72840 167198 72849
rect 167142 72775 167198 72784
rect 91702 72568 91758 72577
rect 164382 72568 164438 72577
rect 91702 72503 91704 72512
rect 91756 72503 91758 72512
rect 95384 72532 95436 72538
rect 91704 72474 91756 72480
rect 164382 72503 164384 72512
rect 95384 72474 95436 72480
rect 164436 72503 164438 72512
rect 167236 72532 167288 72538
rect 164384 72474 164436 72480
rect 167236 72474 167288 72480
rect 95396 71489 95424 72474
rect 95382 71480 95438 71489
rect 95382 71415 95438 71424
rect 91702 71344 91758 71353
rect 164382 71344 164438 71353
rect 91702 71279 91704 71288
rect 91756 71279 91758 71288
rect 95384 71308 95436 71314
rect 91704 71250 91756 71256
rect 164382 71279 164438 71288
rect 95384 71250 95436 71256
rect 91426 70120 91482 70129
rect 91426 70055 91482 70064
rect 91440 69614 91468 70055
rect 91428 69608 91480 69614
rect 91428 69550 91480 69556
rect 94004 69608 94056 69614
rect 94004 69550 94056 69556
rect 91426 68896 91482 68905
rect 91426 68831 91482 68840
rect 91440 68730 91468 68831
rect 91428 68724 91480 68730
rect 91428 68666 91480 68672
rect 93912 68724 93964 68730
rect 93912 68666 93964 68672
rect 91518 67808 91574 67817
rect 91518 67743 91574 67752
rect 91532 66826 91560 67743
rect 91520 66820 91572 66826
rect 91520 66762 91572 66768
rect 93636 66820 93688 66826
rect 93636 66762 93688 66768
rect 92530 66584 92586 66593
rect 92530 66519 92586 66528
rect 22702 65768 22758 65777
rect 22702 65703 22758 65712
rect 44414 65768 44470 65777
rect 44414 65703 44470 65712
rect 22716 62610 22744 65703
rect 44428 65466 44456 65703
rect 44416 65460 44468 65466
rect 44416 65402 44468 65408
rect 47176 65460 47228 65466
rect 47176 65402 47228 65408
rect 22704 62604 22756 62610
rect 22704 62546 22756 62552
rect 47188 60609 47216 65402
rect 92346 65360 92402 65369
rect 92346 65295 92402 65304
rect 91426 61688 91482 61697
rect 91426 61623 91482 61632
rect 91440 61318 91468 61623
rect 91428 61312 91480 61318
rect 91428 61254 91480 61260
rect 47174 60600 47230 60609
rect 47174 60535 47230 60544
rect 47542 60600 47598 60609
rect 47542 60535 47598 60544
rect 44414 57880 44470 57889
rect 44414 57815 44470 57824
rect 26120 50302 26148 53908
rect 26488 50302 26516 53908
rect 26580 53894 26870 53922
rect 26108 50296 26160 50302
rect 26108 50238 26160 50244
rect 26200 50296 26252 50302
rect 26200 50238 26252 50244
rect 26476 50296 26528 50302
rect 26476 50238 26528 50244
rect 20864 50228 20916 50234
rect 20864 50170 20916 50176
rect 25648 50228 25700 50234
rect 25648 50170 25700 50176
rect 20220 49548 20272 49554
rect 20220 49490 20272 49496
rect 20232 46428 20260 49490
rect 20876 46428 20904 50170
rect 22888 50160 22940 50166
rect 22888 50102 22940 50108
rect 21508 49004 21560 49010
rect 21508 48946 21560 48952
rect 21520 46428 21548 48946
rect 22244 48936 22296 48942
rect 22244 48878 22296 48884
rect 22256 46428 22284 48878
rect 22900 46428 22928 50102
rect 24268 50024 24320 50030
rect 24268 49966 24320 49972
rect 23624 49956 23676 49962
rect 23624 49898 23676 49904
rect 23636 46428 23664 49898
rect 24280 46428 24308 49966
rect 24912 49684 24964 49690
rect 24912 49626 24964 49632
rect 24924 46428 24952 49626
rect 25660 46428 25688 50170
rect 26212 49010 26240 50238
rect 26580 50148 26608 53894
rect 27316 50166 27344 53908
rect 26396 50120 26608 50148
rect 27304 50160 27356 50166
rect 26292 49752 26344 49758
rect 26292 49694 26344 49700
rect 26200 49004 26252 49010
rect 26200 48946 26252 48952
rect 26304 46428 26332 49694
rect 26396 48942 26424 50120
rect 27304 50102 27356 50108
rect 27028 50092 27080 50098
rect 27028 50034 27080 50040
rect 26384 48936 26436 48942
rect 26384 48878 26436 48884
rect 27040 46428 27068 50034
rect 27684 49962 27712 53908
rect 27856 50364 27908 50370
rect 27856 50306 27908 50312
rect 27672 49956 27724 49962
rect 27672 49898 27724 49904
rect 27868 48890 27896 50306
rect 28052 50030 28080 53908
rect 28040 50024 28092 50030
rect 28040 49966 28092 49972
rect 28316 50024 28368 50030
rect 28316 49966 28368 49972
rect 27776 48862 27896 48890
rect 27776 46442 27804 48862
rect 27698 46414 27804 46442
rect 28328 46428 28356 49966
rect 28512 49690 28540 53908
rect 28880 50302 28908 53908
rect 28868 50296 28920 50302
rect 28868 50238 28920 50244
rect 29052 50228 29104 50234
rect 29052 50170 29104 50176
rect 28500 49684 28552 49690
rect 28500 49626 28552 49632
rect 29064 46428 29092 50170
rect 29248 49758 29276 53908
rect 29432 53894 29722 53922
rect 29432 50098 29460 53894
rect 30076 50370 30104 53908
rect 30168 53894 30458 53922
rect 30064 50364 30116 50370
rect 30064 50306 30116 50312
rect 29420 50092 29472 50098
rect 29420 50034 29472 50040
rect 30168 50030 30196 53894
rect 30904 50302 30932 53908
rect 30892 50296 30944 50302
rect 30892 50238 30944 50244
rect 30432 50092 30484 50098
rect 30432 50034 30484 50040
rect 30156 50024 30208 50030
rect 30156 49966 30208 49972
rect 29696 49956 29748 49962
rect 29696 49898 29748 49904
rect 29236 49752 29288 49758
rect 29236 49694 29288 49700
rect 29708 46428 29736 49898
rect 30444 46428 30472 50034
rect 31076 50024 31128 50030
rect 31076 49966 31128 49972
rect 31088 46428 31116 49966
rect 31272 49962 31300 53908
rect 31640 50098 31668 53908
rect 31628 50092 31680 50098
rect 31628 50034 31680 50040
rect 32100 50030 32128 53908
rect 32192 53894 32482 53922
rect 32088 50024 32140 50030
rect 32088 49966 32140 49972
rect 31260 49956 31312 49962
rect 31260 49898 31312 49904
rect 32192 49026 32220 53894
rect 31916 48998 32220 49026
rect 31916 46442 31944 48998
rect 32836 46442 32864 53908
rect 33296 46442 33324 53908
rect 31838 46414 31944 46442
rect 32482 46414 32864 46442
rect 33126 46414 33324 46442
rect 33664 46442 33692 53908
rect 34138 53894 34336 53922
rect 34506 53894 34704 53922
rect 34874 53894 35256 53922
rect 34308 46442 34336 53894
rect 34676 50250 34704 53894
rect 34676 50222 34888 50250
rect 34860 46442 34888 50222
rect 35228 46816 35256 53894
rect 35320 50710 35348 53908
rect 35702 53894 35992 53922
rect 35308 50704 35360 50710
rect 35308 50646 35360 50652
rect 35964 50658 35992 53894
rect 36056 50778 36084 53908
rect 36516 50846 36544 53908
rect 36504 50840 36556 50846
rect 36504 50782 36556 50788
rect 36044 50772 36096 50778
rect 36044 50714 36096 50720
rect 36504 50704 36556 50710
rect 35964 50630 36176 50658
rect 36504 50646 36556 50652
rect 36148 50302 36176 50630
rect 36136 50296 36188 50302
rect 36136 50238 36188 50244
rect 35228 46788 35440 46816
rect 35412 46442 35440 46788
rect 33664 46414 33862 46442
rect 34308 46414 34506 46442
rect 34860 46414 35242 46442
rect 35412 46414 35886 46442
rect 36516 46428 36544 50646
rect 36884 50370 36912 53908
rect 37266 53894 37372 53922
rect 36872 50364 36924 50370
rect 36872 50306 36924 50312
rect 37344 50302 37372 53894
rect 37424 50772 37476 50778
rect 37424 50714 37476 50720
rect 37240 50296 37292 50302
rect 37240 50238 37292 50244
rect 37332 50296 37384 50302
rect 37332 50238 37384 50244
rect 37252 46428 37280 50238
rect 37436 50114 37464 50714
rect 37712 50438 37740 53908
rect 38080 50506 38108 53908
rect 38462 53894 38844 53922
rect 38620 50840 38672 50846
rect 38620 50782 38672 50788
rect 38068 50500 38120 50506
rect 38068 50442 38120 50448
rect 37700 50432 37752 50438
rect 37700 50374 37752 50380
rect 37436 50086 37556 50114
rect 37528 46442 37556 50086
rect 37528 46414 37910 46442
rect 38632 46428 38660 50782
rect 38816 50250 38844 53894
rect 38908 50574 38936 53908
rect 39276 50642 39304 53908
rect 39264 50636 39316 50642
rect 39264 50578 39316 50584
rect 38896 50568 38948 50574
rect 38896 50510 38948 50516
rect 39644 50302 39672 53908
rect 39724 50500 39776 50506
rect 39724 50442 39776 50448
rect 39632 50296 39684 50302
rect 38816 50222 38936 50250
rect 39632 50238 39684 50244
rect 38908 49894 38936 50222
rect 39264 50228 39316 50234
rect 39264 50170 39316 50176
rect 38896 49888 38948 49894
rect 38896 49830 38948 49836
rect 39276 46428 39304 50170
rect 39736 49690 39764 50442
rect 40104 50370 40132 53908
rect 40184 50432 40236 50438
rect 40184 50374 40236 50380
rect 40092 50364 40144 50370
rect 40092 50306 40144 50312
rect 40000 50160 40052 50166
rect 40000 50102 40052 50108
rect 39724 49684 39776 49690
rect 39724 49626 39776 49632
rect 40012 46428 40040 50102
rect 40196 48890 40224 50374
rect 40472 50302 40500 53908
rect 40840 51050 40868 53908
rect 40828 51044 40880 51050
rect 40828 50986 40880 50992
rect 40828 50568 40880 50574
rect 40828 50510 40880 50516
rect 40460 50296 40512 50302
rect 40460 50238 40512 50244
rect 40840 50030 40868 50510
rect 41300 50302 41328 53908
rect 41380 50636 41432 50642
rect 41380 50578 41432 50584
rect 41288 50296 41340 50302
rect 41288 50238 41340 50244
rect 40828 50024 40880 50030
rect 40828 49966 40880 49972
rect 41392 49962 41420 50578
rect 41668 50438 41696 53908
rect 42944 51044 42996 51050
rect 42944 50986 42996 50992
rect 41656 50432 41708 50438
rect 41656 50374 41708 50380
rect 42956 50030 42984 50986
rect 44048 50432 44100 50438
rect 44048 50374 44100 50380
rect 43772 50092 43824 50098
rect 43772 50034 43824 50040
rect 42668 50024 42720 50030
rect 42668 49966 42720 49972
rect 42944 50024 42996 50030
rect 42944 49966 42996 49972
rect 41380 49956 41432 49962
rect 41380 49898 41432 49904
rect 42024 49888 42076 49894
rect 42024 49830 42076 49836
rect 41288 49684 41340 49690
rect 41288 49626 41340 49632
rect 40196 48862 40316 48890
rect 40288 46442 40316 48862
rect 40288 46414 40670 46442
rect 41300 46428 41328 49626
rect 42036 46428 42064 49830
rect 42680 46428 42708 49966
rect 43404 49956 43456 49962
rect 43404 49898 43456 49904
rect 43416 46428 43444 49898
rect 43784 46442 43812 50034
rect 44060 49826 44088 50374
rect 44048 49820 44100 49826
rect 44048 49762 44100 49768
rect 44428 49554 44456 57815
rect 44692 50364 44744 50370
rect 44692 50306 44744 50312
rect 44416 49548 44468 49554
rect 44416 49490 44468 49496
rect 43784 46414 44074 46442
rect 44704 46428 44732 50306
rect 46808 50228 46860 50234
rect 46808 50170 46860 50176
rect 45428 50160 45480 50166
rect 45428 50102 45480 50108
rect 45440 46428 45468 50102
rect 46072 50024 46124 50030
rect 46072 49966 46124 49972
rect 46084 46428 46112 49966
rect 46820 46428 46848 50170
rect 47452 49820 47504 49826
rect 47452 49762 47504 49768
rect 47464 46428 47492 49762
rect 47556 46873 47584 60535
rect 91518 59240 91574 59249
rect 91518 59175 91574 59184
rect 91532 58598 91560 59175
rect 91520 58592 91572 58598
rect 91520 58534 91572 58540
rect 92360 58530 92388 65295
rect 92544 59754 92572 66519
rect 92622 64136 92678 64145
rect 92622 64071 92624 64080
rect 92676 64071 92678 64080
rect 93544 64100 93596 64106
rect 92624 64042 92676 64048
rect 93544 64042 93596 64048
rect 93358 62912 93414 62921
rect 93358 62847 93414 62856
rect 92532 59748 92584 59754
rect 92532 59690 92584 59696
rect 92348 58524 92400 58530
rect 92348 58466 92400 58472
rect 92898 58016 92954 58025
rect 92898 57951 92954 57960
rect 91426 56792 91482 56801
rect 91426 56727 91482 56736
rect 91334 54480 91390 54489
rect 91334 54415 91390 54424
rect 53260 51497 53288 53908
rect 53246 51488 53302 51497
rect 53246 51423 53302 51432
rect 66600 51390 66628 53908
rect 73224 51458 73252 53908
rect 82134 51624 82190 51633
rect 82134 51559 82136 51568
rect 82188 51559 82190 51568
rect 83606 51624 83662 51633
rect 83606 51559 83662 51568
rect 84344 51588 84396 51594
rect 82136 51530 82188 51536
rect 72016 51452 72068 51458
rect 72016 51394 72068 51400
rect 73212 51452 73264 51458
rect 73212 51394 73264 51400
rect 66588 51384 66640 51390
rect 66588 51326 66640 51332
rect 64564 50976 64616 50982
rect 64564 50918 64616 50924
rect 47542 46864 47598 46873
rect 47542 46799 47598 46808
rect 50764 46556 50816 46562
rect 50764 46498 50816 46504
rect 61620 46556 61672 46562
rect 61620 46498 61672 46504
rect 50672 46284 50724 46290
rect 50672 46226 50724 46232
rect 50578 46184 50634 46193
rect 50578 46119 50634 46128
rect 49934 45232 49990 45241
rect 49934 45167 49990 45176
rect 49948 44833 49976 45167
rect 49934 44824 49990 44833
rect 49934 44759 49990 44768
rect 14700 40572 14752 40578
rect 14700 40514 14752 40520
rect 18012 40572 18064 40578
rect 18012 40514 18064 40520
rect 13318 40472 13374 40481
rect 13318 40407 13374 40416
rect 18024 40209 18052 40514
rect 18010 40200 18066 40209
rect 18010 40135 18066 40144
rect 50486 34216 50542 34225
rect 50486 34151 50542 34160
rect 50500 33817 50528 34151
rect 50486 33808 50542 33817
rect 50486 33743 50542 33752
rect 50486 32720 50542 32729
rect 50486 32655 50542 32664
rect 50500 32321 50528 32655
rect 50486 32312 50542 32321
rect 50486 32247 50542 32256
rect 18102 25512 18158 25521
rect 18102 25447 18158 25456
rect 13134 19392 13190 19401
rect 13134 19327 13190 19336
rect 13148 19158 13176 19327
rect 13136 19152 13188 19158
rect 13136 19094 13188 19100
rect 18116 18478 18144 25447
rect 50592 24682 50620 46119
rect 50408 24654 50620 24682
rect 18104 18472 18156 18478
rect 18104 18414 18156 18420
rect 50408 18410 50436 24654
rect 50580 24524 50632 24530
rect 50580 24466 50632 24472
rect 50592 19809 50620 24466
rect 50578 19800 50634 19809
rect 50578 19735 50634 19744
rect 50684 19265 50712 46226
rect 50776 21169 50804 46498
rect 51040 46488 51092 46494
rect 51040 46430 51092 46436
rect 50948 46352 51000 46358
rect 50948 46294 51000 46300
rect 50856 46216 50908 46222
rect 50856 46158 50908 46164
rect 50868 24530 50896 46158
rect 50856 24524 50908 24530
rect 50856 24466 50908 24472
rect 50960 24410 50988 46294
rect 50868 24382 50988 24410
rect 50762 21160 50818 21169
rect 50762 21095 50818 21104
rect 50868 20489 50896 24382
rect 51052 24274 51080 46430
rect 51132 46420 51184 46426
rect 51132 46362 51184 46368
rect 60056 46420 60108 46426
rect 60056 46362 60108 46368
rect 50960 24246 51080 24274
rect 50960 21849 50988 24246
rect 51038 24152 51094 24161
rect 51038 24087 51040 24096
rect 51092 24087 51094 24096
rect 51040 24058 51092 24064
rect 50946 21840 51002 21849
rect 50946 21775 51002 21784
rect 51144 21033 51172 46362
rect 58584 46352 58636 46358
rect 58584 46294 58636 46300
rect 55640 46284 55692 46290
rect 55640 46226 55692 46232
rect 54076 46148 54128 46154
rect 54076 46090 54128 46096
rect 51314 44960 51370 44969
rect 51314 44895 51370 44904
rect 51328 44289 51356 44895
rect 51314 44280 51370 44289
rect 51314 44215 51370 44224
rect 51222 44144 51278 44153
rect 51278 44102 51356 44130
rect 51222 44079 51278 44088
rect 51328 43337 51356 44102
rect 51314 43328 51370 43337
rect 51314 43263 51370 43272
rect 51222 42104 51278 42113
rect 51278 42062 51356 42090
rect 51222 42039 51278 42048
rect 51328 41297 51356 42062
rect 51314 41288 51370 41297
rect 51314 41223 51370 41232
rect 51222 41152 51278 41161
rect 51278 41110 51356 41138
rect 51222 41087 51278 41096
rect 51328 40481 51356 41110
rect 51314 40472 51370 40481
rect 51314 40407 51370 40416
rect 51222 39928 51278 39937
rect 51278 39886 51356 39914
rect 51222 39863 51278 39872
rect 51328 39121 51356 39886
rect 51314 39112 51370 39121
rect 51314 39047 51370 39056
rect 51222 38024 51278 38033
rect 51278 37982 51356 38010
rect 51222 37959 51278 37968
rect 51328 37081 51356 37982
rect 51314 37072 51370 37081
rect 51314 37007 51370 37016
rect 51222 36936 51278 36945
rect 51278 36894 51448 36922
rect 51222 36871 51278 36880
rect 51222 36664 51278 36673
rect 51278 36622 51356 36650
rect 51222 36599 51278 36608
rect 51328 35993 51356 36622
rect 51420 36401 51448 36894
rect 51406 36392 51462 36401
rect 51406 36327 51462 36336
rect 51314 35984 51370 35993
rect 51314 35919 51370 35928
rect 51222 34488 51278 34497
rect 51278 34446 51448 34474
rect 51222 34423 51278 34432
rect 51222 34080 51278 34089
rect 51278 34038 51356 34066
rect 51222 34015 51278 34024
rect 51328 33001 51356 34038
rect 51420 33658 51448 34446
rect 51498 33672 51554 33681
rect 51420 33630 51498 33658
rect 51498 33607 51554 33616
rect 51314 32992 51370 33001
rect 51314 32927 51370 32936
rect 51222 32448 51278 32457
rect 51278 32406 51356 32434
rect 51222 32383 51278 32392
rect 51328 31777 51356 32406
rect 51314 31768 51370 31777
rect 51314 31703 51370 31712
rect 51222 31632 51278 31641
rect 51278 31590 51356 31618
rect 51222 31567 51278 31576
rect 51328 30825 51356 31590
rect 51314 30816 51370 30825
rect 51314 30751 51370 30760
rect 51222 30408 51278 30417
rect 51278 30366 51356 30394
rect 51222 30343 51278 30352
rect 51328 29465 51356 30366
rect 51314 29456 51370 29465
rect 51314 29391 51370 29400
rect 51222 28640 51278 28649
rect 51278 28598 51448 28626
rect 51222 28575 51278 28584
rect 51222 28368 51278 28377
rect 51278 28326 51356 28354
rect 51222 28303 51278 28312
rect 51328 27561 51356 28326
rect 51420 28105 51448 28598
rect 51406 28096 51462 28105
rect 51406 28031 51462 28040
rect 51314 27552 51370 27561
rect 51314 27487 51370 27496
rect 51222 27416 51278 27425
rect 51278 27374 51356 27402
rect 51222 27351 51278 27360
rect 51328 26745 51356 27374
rect 51314 26736 51370 26745
rect 51314 26671 51370 26680
rect 51406 26192 51462 26201
rect 51406 26127 51462 26136
rect 51314 25648 51370 25657
rect 51314 25583 51370 25592
rect 51222 25512 51278 25521
rect 51222 25447 51278 25456
rect 51236 24954 51264 25447
rect 51328 25113 51356 25583
rect 51420 25521 51448 26127
rect 51406 25512 51462 25521
rect 51406 25447 51462 25456
rect 51314 25104 51370 25113
rect 51314 25039 51370 25048
rect 51236 24926 51356 24954
rect 51328 24569 51356 24926
rect 51314 24560 51370 24569
rect 51314 24495 51370 24504
rect 51316 24116 51368 24122
rect 51316 24058 51368 24064
rect 51328 23345 51356 24058
rect 51314 23336 51370 23345
rect 51314 23271 51370 23280
rect 51222 23200 51278 23209
rect 51278 23158 51356 23186
rect 51222 23135 51278 23144
rect 51328 22506 51356 23158
rect 51498 22520 51554 22529
rect 51328 22478 51498 22506
rect 51498 22455 51554 22464
rect 54088 22234 54116 46090
rect 55652 44796 55680 46226
rect 57112 46216 57164 46222
rect 57112 46158 57164 46164
rect 57124 44796 57152 46158
rect 58596 44796 58624 46294
rect 60068 44796 60096 46362
rect 61632 44796 61660 46498
rect 63092 46488 63144 46494
rect 63092 46430 63144 46436
rect 63104 44796 63132 46430
rect 64576 44796 64604 50918
rect 66600 50273 66628 51326
rect 72028 50914 72056 51394
rect 82148 51322 82176 51530
rect 83620 51458 83648 51559
rect 84344 51530 84396 51536
rect 84356 51458 84384 51530
rect 83608 51452 83660 51458
rect 83608 51394 83660 51400
rect 84344 51452 84396 51458
rect 84344 51394 84396 51400
rect 82136 51316 82188 51322
rect 82136 51258 82188 51264
rect 86564 50982 86592 53908
rect 86552 50976 86604 50982
rect 86552 50918 86604 50924
rect 72016 50908 72068 50914
rect 72016 50850 72068 50856
rect 66586 50264 66642 50273
rect 66586 50199 66642 50208
rect 91348 46850 91376 54415
rect 91440 49282 91468 56727
rect 92622 55568 92678 55577
rect 92678 55526 92756 55554
rect 92622 55503 92678 55512
rect 91428 49276 91480 49282
rect 91428 49218 91480 49224
rect 91348 46822 91744 46850
rect 91716 46714 91744 46822
rect 91716 46686 92190 46714
rect 92728 46700 92756 55526
rect 92912 49434 92940 57951
rect 93372 50098 93400 62847
rect 93452 61312 93504 61318
rect 93452 61254 93504 61260
rect 93464 50166 93492 61254
rect 93556 55033 93584 64042
rect 93648 61425 93676 66762
rect 93924 64145 93952 68666
rect 94016 65505 94044 69550
rect 95396 69041 95424 71250
rect 164396 71178 164424 71279
rect 164384 71172 164436 71178
rect 164384 71114 164436 71120
rect 167248 70809 167276 72474
rect 167328 71172 167380 71178
rect 167328 71114 167380 71120
rect 167234 70800 167290 70809
rect 167234 70735 167290 70744
rect 163554 70120 163610 70129
rect 163554 70055 163610 70064
rect 163568 69954 163596 70055
rect 163556 69948 163608 69954
rect 163556 69890 163608 69896
rect 167236 69948 167288 69954
rect 167236 69890 167288 69896
rect 95382 69032 95438 69041
rect 95382 68967 95438 68976
rect 163738 68896 163794 68905
rect 163738 68831 163794 68840
rect 163752 68254 163780 68831
rect 163740 68248 163792 68254
rect 163740 68190 163792 68196
rect 164382 67808 164438 67817
rect 164382 67743 164438 67752
rect 164396 66826 164424 67743
rect 167248 66865 167276 69890
rect 167340 68769 167368 71114
rect 167326 68760 167382 68769
rect 167326 68695 167382 68704
rect 167328 68248 167380 68254
rect 167328 68190 167380 68196
rect 167234 66856 167290 66865
rect 164384 66820 164436 66826
rect 167234 66791 167290 66800
rect 164384 66762 164436 66768
rect 95382 66720 95438 66729
rect 95382 66655 95438 66664
rect 95396 65505 95424 66655
rect 164382 66584 164438 66593
rect 164382 66519 164438 66528
rect 94002 65496 94058 65505
rect 94002 65431 94058 65440
rect 95382 65496 95438 65505
rect 164396 65466 164424 66519
rect 95382 65431 95438 65440
rect 164384 65460 164436 65466
rect 164384 65402 164436 65408
rect 167144 65460 167196 65466
rect 167144 65402 167196 65408
rect 164382 65360 164438 65369
rect 164382 65295 164438 65304
rect 164396 64514 164424 65295
rect 164384 64508 164436 64514
rect 164384 64450 164436 64456
rect 167052 64508 167104 64514
rect 167052 64450 167104 64456
rect 93910 64136 93966 64145
rect 93910 64071 93966 64080
rect 164382 64136 164438 64145
rect 164382 64071 164384 64080
rect 164436 64071 164438 64080
rect 166500 64100 166552 64106
rect 164384 64042 164436 64048
rect 166500 64042 166552 64048
rect 117462 63184 117518 63193
rect 117462 63119 117518 63128
rect 117476 62678 117504 63119
rect 163738 62912 163794 62921
rect 163738 62847 163794 62856
rect 117464 62672 117516 62678
rect 117464 62614 117516 62620
rect 119488 62672 119540 62678
rect 119488 62614 119540 62620
rect 93634 61416 93690 61425
rect 93634 61351 93690 61360
rect 119500 60609 119528 62614
rect 119486 60600 119542 60609
rect 119486 60535 119542 60544
rect 94646 60464 94702 60473
rect 94646 60399 94702 60408
rect 94096 59748 94148 59754
rect 94096 59690 94148 59696
rect 94108 59657 94136 59690
rect 94094 59648 94150 59657
rect 94094 59583 94150 59592
rect 93636 58592 93688 58598
rect 93636 58534 93688 58540
rect 93542 55024 93598 55033
rect 93542 54959 93598 54968
rect 93648 50234 93676 58534
rect 93636 50228 93688 50234
rect 93636 50170 93688 50176
rect 94372 50228 94424 50234
rect 94372 50170 94424 50176
rect 93452 50160 93504 50166
rect 93452 50102 93504 50108
rect 93360 50092 93412 50098
rect 93360 50034 93412 50040
rect 92912 49406 93492 49434
rect 92900 49276 92952 49282
rect 92900 49218 92952 49224
rect 92912 46714 92940 49218
rect 93464 46714 93492 49406
rect 92912 46686 93294 46714
rect 93464 46686 93846 46714
rect 94384 46700 94412 50170
rect 94660 46714 94688 60399
rect 95200 58524 95252 58530
rect 95200 58466 95252 58472
rect 95212 57345 95240 58466
rect 95198 57336 95254 57345
rect 95198 57271 95254 57280
rect 163094 54480 163150 54489
rect 163094 54415 163150 54424
rect 97788 53894 98124 53922
rect 98340 53894 98492 53922
rect 98616 53894 98860 53922
rect 98984 53894 99320 53922
rect 97684 50228 97736 50234
rect 97684 50170 97736 50176
rect 95476 50160 95528 50166
rect 95476 50102 95528 50108
rect 97132 50160 97184 50166
rect 97132 50102 97184 50108
rect 94660 46686 94950 46714
rect 95488 46700 95516 50102
rect 96028 50092 96080 50098
rect 96028 50034 96080 50040
rect 96040 46700 96068 50034
rect 96580 49140 96632 49146
rect 96580 49082 96632 49088
rect 96592 46700 96620 49082
rect 97144 46700 97172 50102
rect 97696 46700 97724 50170
rect 97788 49146 97816 53894
rect 98236 51520 98288 51526
rect 98236 51462 98288 51468
rect 97776 49140 97828 49146
rect 97776 49082 97828 49088
rect 98248 46700 98276 51462
rect 98340 50166 98368 53894
rect 98616 50234 98644 53894
rect 98984 51526 99012 53894
rect 99674 53650 99702 53908
rect 99812 53894 100056 53922
rect 100272 53894 100516 53922
rect 100732 53894 100884 53922
rect 101100 53894 101252 53922
rect 99674 53622 99748 53650
rect 98972 51520 99024 51526
rect 98972 51462 99024 51468
rect 98604 50228 98656 50234
rect 98604 50170 98656 50176
rect 99720 50166 99748 53622
rect 98328 50160 98380 50166
rect 98328 50102 98380 50108
rect 98788 50160 98840 50166
rect 98788 50102 98840 50108
rect 99708 50160 99760 50166
rect 99708 50102 99760 50108
rect 98800 46700 98828 50102
rect 99812 49842 99840 53894
rect 99444 49814 99840 49842
rect 99444 46700 99472 49814
rect 100272 46714 100300 53894
rect 100732 46714 100760 53894
rect 100010 46686 100300 46714
rect 100562 46686 100760 46714
rect 101100 46700 101128 53894
rect 101698 53650 101726 53908
rect 102080 53894 102232 53922
rect 102448 53894 102784 53922
rect 102908 53894 103152 53922
rect 103276 53894 103428 53922
rect 103644 53894 103980 53922
rect 104104 53894 104348 53922
rect 104472 53894 104716 53922
rect 104840 53894 105084 53922
rect 105300 53894 105544 53922
rect 105668 53894 106004 53922
rect 106128 53894 106372 53922
rect 106496 53894 106648 53922
rect 106864 53894 107200 53922
rect 107324 53894 107568 53922
rect 107692 53894 107844 53922
rect 108060 53894 108396 53922
rect 108520 53894 108764 53922
rect 108888 53894 109132 53922
rect 109256 53894 109592 53922
rect 109716 53894 109960 53922
rect 110084 53894 110328 53922
rect 110452 53894 110604 53922
rect 110912 53894 111156 53922
rect 111280 53894 111524 53922
rect 111648 53894 111984 53922
rect 112108 53894 112352 53922
rect 112476 53894 112720 53922
rect 112844 53894 113180 53922
rect 113304 53894 113548 53922
rect 113672 53894 114008 53922
rect 101652 53622 101726 53650
rect 101652 46700 101680 53622
rect 102204 46700 102232 53894
rect 102756 46700 102784 53894
rect 103124 46714 103152 53894
rect 103400 51526 103428 53894
rect 103388 51520 103440 51526
rect 103388 51462 103440 51468
rect 103848 51520 103900 51526
rect 103848 51462 103900 51468
rect 103124 46686 103322 46714
rect 103860 46700 103888 51462
rect 103952 47786 103980 53894
rect 104320 52018 104348 53894
rect 104320 51990 104624 52018
rect 103940 47780 103992 47786
rect 103940 47722 103992 47728
rect 104400 47780 104452 47786
rect 104400 47722 104452 47728
rect 104412 46700 104440 47722
rect 104596 46714 104624 51990
rect 104688 50846 104716 53894
rect 105056 51526 105084 53894
rect 105044 51520 105096 51526
rect 105044 51462 105096 51468
rect 105516 51458 105544 53894
rect 105504 51452 105556 51458
rect 105504 51394 105556 51400
rect 105976 51390 106004 53894
rect 106344 51526 106372 53894
rect 106148 51520 106200 51526
rect 106148 51462 106200 51468
rect 106332 51520 106384 51526
rect 106332 51462 106384 51468
rect 105964 51384 106016 51390
rect 105964 51326 106016 51332
rect 104676 50840 104728 50846
rect 104676 50782 104728 50788
rect 105504 50840 105556 50846
rect 105504 50782 105556 50788
rect 104596 46686 104978 46714
rect 105516 46700 105544 50782
rect 106160 46700 106188 51462
rect 106620 51322 106648 53894
rect 107172 51458 107200 53894
rect 106700 51452 106752 51458
rect 106700 51394 106752 51400
rect 107160 51452 107212 51458
rect 107160 51394 107212 51400
rect 106608 51316 106660 51322
rect 106608 51258 106660 51264
rect 106712 46700 106740 51394
rect 107252 51384 107304 51390
rect 107252 51326 107304 51332
rect 107264 46700 107292 51326
rect 107540 50302 107568 53894
rect 107816 51610 107844 53894
rect 107816 51582 107936 51610
rect 107804 51520 107856 51526
rect 107804 51462 107856 51468
rect 107528 50296 107580 50302
rect 107528 50238 107580 50244
rect 107816 46700 107844 51462
rect 107908 50166 107936 51582
rect 108368 50370 108396 53894
rect 108448 51316 108500 51322
rect 108448 51258 108500 51264
rect 108356 50364 108408 50370
rect 108356 50306 108408 50312
rect 108460 50250 108488 51258
rect 108736 50302 108764 53894
rect 108908 51452 108960 51458
rect 108908 51394 108960 51400
rect 108368 50222 108488 50250
rect 108724 50296 108776 50302
rect 108724 50238 108776 50244
rect 107896 50160 107948 50166
rect 107896 50102 107948 50108
rect 108368 46700 108396 50222
rect 108920 46700 108948 51394
rect 109104 50386 109132 53894
rect 109564 51050 109592 53894
rect 109552 51044 109604 51050
rect 109552 50986 109604 50992
rect 109932 50438 109960 53894
rect 110300 51458 110328 53894
rect 110576 51610 110604 53894
rect 110576 51582 110696 51610
rect 110288 51452 110340 51458
rect 110288 51394 110340 51400
rect 109920 50432 109972 50438
rect 109104 50358 109316 50386
rect 109920 50374 109972 50380
rect 109288 50098 109316 50358
rect 110564 50364 110616 50370
rect 110564 50306 110616 50312
rect 109460 50228 109512 50234
rect 109460 50170 109512 50176
rect 109276 50092 109328 50098
rect 109276 50034 109328 50040
rect 109472 46700 109500 50170
rect 110012 50160 110064 50166
rect 110012 50102 110064 50108
rect 110024 46700 110052 50102
rect 110576 46700 110604 50306
rect 110668 50166 110696 51582
rect 111128 50506 111156 53894
rect 111496 51526 111524 53894
rect 111484 51520 111536 51526
rect 111484 51462 111536 51468
rect 111760 51452 111812 51458
rect 111760 51394 111812 51400
rect 111116 50500 111168 50506
rect 111116 50442 111168 50448
rect 111116 50228 111168 50234
rect 111116 50170 111168 50176
rect 110656 50160 110708 50166
rect 110656 50102 110708 50108
rect 111128 46700 111156 50170
rect 111668 50092 111720 50098
rect 111668 50034 111720 50040
rect 111680 46700 111708 50034
rect 111772 49418 111800 51394
rect 111852 51044 111904 51050
rect 111852 50986 111904 50992
rect 111760 49412 111812 49418
rect 111760 49354 111812 49360
rect 111864 49026 111892 50986
rect 111956 50302 111984 53894
rect 112324 51050 112352 53894
rect 112404 51520 112456 51526
rect 112404 51462 112456 51468
rect 112312 51044 112364 51050
rect 112312 50986 112364 50992
rect 111944 50296 111996 50302
rect 111944 50238 111996 50244
rect 112416 49826 112444 51462
rect 112692 51458 112720 53894
rect 113152 51526 113180 53894
rect 113140 51520 113192 51526
rect 113140 51462 113192 51468
rect 112680 51452 112732 51458
rect 112680 51394 112732 51400
rect 112680 50500 112732 50506
rect 112680 50442 112732 50448
rect 112692 50030 112720 50442
rect 112772 50228 112824 50234
rect 112772 50170 112824 50176
rect 112680 50024 112732 50030
rect 112680 49966 112732 49972
rect 112404 49820 112456 49826
rect 112404 49762 112456 49768
rect 111864 48998 112076 49026
rect 112048 46714 112076 48998
rect 112048 46686 112246 46714
rect 112784 46700 112812 50170
rect 113520 49622 113548 53894
rect 113980 50302 114008 53894
rect 138360 53894 138604 53922
rect 145168 53894 145228 53922
rect 151608 53894 151944 53922
rect 114612 51520 114664 51526
rect 114612 51462 114664 51468
rect 114428 51044 114480 51050
rect 114428 50986 114480 50992
rect 113968 50296 114020 50302
rect 113968 50238 114020 50244
rect 113968 50160 114020 50166
rect 113968 50102 114020 50108
rect 113508 49616 113560 49622
rect 113508 49558 113560 49564
rect 113416 49412 113468 49418
rect 113416 49354 113468 49360
rect 113428 46700 113456 49354
rect 113980 46700 114008 50102
rect 114440 49010 114468 50986
rect 114520 50024 114572 50030
rect 114520 49966 114572 49972
rect 114428 49004 114480 49010
rect 114428 48946 114480 48952
rect 114532 46700 114560 49966
rect 114624 49146 114652 51462
rect 114704 51452 114756 51458
rect 114704 51394 114756 51400
rect 114716 49554 114744 51394
rect 138360 51322 138388 53894
rect 145168 51594 145196 53894
rect 145156 51588 145208 51594
rect 145156 51530 145208 51536
rect 138348 51316 138400 51322
rect 138348 51258 138400 51264
rect 151608 50914 151636 53894
rect 138164 50908 138216 50914
rect 138164 50850 138216 50856
rect 151596 50908 151648 50914
rect 151596 50850 151648 50856
rect 115624 50228 115676 50234
rect 115624 50170 115676 50176
rect 118384 50228 118436 50234
rect 118384 50170 118436 50176
rect 115072 49820 115124 49826
rect 115072 49762 115124 49768
rect 114704 49548 114756 49554
rect 114704 49490 114756 49496
rect 114612 49140 114664 49146
rect 114612 49082 114664 49088
rect 115084 46700 115112 49762
rect 115636 46700 115664 50170
rect 117832 49616 117884 49622
rect 117832 49558 117884 49564
rect 116728 49548 116780 49554
rect 116728 49490 116780 49496
rect 116176 49004 116228 49010
rect 116176 48946 116228 48952
rect 116188 46700 116216 48946
rect 116740 46700 116768 49490
rect 117280 49140 117332 49146
rect 117280 49082 117332 49088
rect 117292 46700 117320 49082
rect 117844 46700 117872 49558
rect 118396 46700 118424 50170
rect 119408 46958 119712 46986
rect 119408 46714 119436 46958
rect 118962 46686 119436 46714
rect 75050 46592 75106 46601
rect 75050 46527 75106 46536
rect 73578 46456 73634 46465
rect 73578 46391 73634 46400
rect 72106 46320 72162 46329
rect 72106 46255 72162 46264
rect 70634 46184 70690 46193
rect 67600 46148 67652 46154
rect 70634 46119 70690 46128
rect 67600 46090 67652 46096
rect 67612 44796 67640 46090
rect 70648 44796 70676 46119
rect 72120 44796 72148 46255
rect 73592 44796 73620 46391
rect 75064 44796 75092 46527
rect 76616 46352 76668 46358
rect 76616 46294 76668 46300
rect 87840 46352 87892 46358
rect 87840 46294 87892 46300
rect 76628 44796 76656 46294
rect 81124 46284 81176 46290
rect 81124 46226 81176 46232
rect 78088 46216 78140 46222
rect 78088 46158 78140 46164
rect 78100 44796 78128 46158
rect 79560 46148 79612 46154
rect 79560 46090 79612 46096
rect 79572 44796 79600 46090
rect 81136 44796 81164 46226
rect 86460 46216 86512 46222
rect 86460 46158 86512 46164
rect 85080 46148 85132 46154
rect 85080 46090 85132 46096
rect 68794 44688 68850 44697
rect 82870 44688 82926 44697
rect 68850 44646 69098 44674
rect 82622 44646 82870 44674
rect 68794 44623 68850 44632
rect 82870 44623 82926 44632
rect 84094 44510 84384 44538
rect 84356 44454 84384 44510
rect 84344 44448 84396 44454
rect 84344 44390 84396 44396
rect 54088 22206 55036 22234
rect 51222 21976 51278 21985
rect 51278 21934 51356 21962
rect 51222 21911 51278 21920
rect 51328 21169 51356 21934
rect 55008 21282 55036 22206
rect 55008 21254 55390 21282
rect 85092 21266 85120 46090
rect 85172 44448 85224 44454
rect 85172 44390 85224 44396
rect 85184 22626 85212 44390
rect 85172 22620 85224 22626
rect 85172 22562 85224 22568
rect 85080 21260 85132 21266
rect 85080 21202 85132 21208
rect 51314 21160 51370 21169
rect 51314 21095 51370 21104
rect 51130 21024 51186 21033
rect 58766 21024 58822 21033
rect 58426 20982 58766 21010
rect 51130 20959 51186 20968
rect 58766 20959 58822 20968
rect 60790 20888 60846 20897
rect 50854 20480 50910 20489
rect 50854 20415 50910 20424
rect 50670 19256 50726 19265
rect 50670 19191 50726 19200
rect 50396 18404 50448 18410
rect 50396 18346 50448 18352
rect 55088 18336 55140 18342
rect 55088 18278 55140 18284
rect 39080 18268 39132 18274
rect 39080 18210 39132 18216
rect 33744 18064 33796 18070
rect 33744 18006 33796 18012
rect 28408 17996 28460 18002
rect 28408 17938 28460 17944
rect 17736 17928 17788 17934
rect 17736 17870 17788 17876
rect 12492 17792 12544 17798
rect 12492 17734 12544 17740
rect 12504 9304 12532 17734
rect 17748 9304 17776 17870
rect 23072 17860 23124 17866
rect 23072 17802 23124 17808
rect 23084 9304 23112 17802
rect 28420 9304 28448 17938
rect 33756 9304 33784 18006
rect 39092 9304 39120 18210
rect 49752 18200 49804 18206
rect 49752 18142 49804 18148
rect 44416 18132 44468 18138
rect 44416 18074 44468 18080
rect 44428 9304 44456 18074
rect 49764 9304 49792 18142
rect 55100 9304 55128 18278
rect 56388 18041 56416 20860
rect 56374 18032 56430 18041
rect 56374 17967 56430 17976
rect 57400 17905 57428 20860
rect 59438 20846 59544 20874
rect 60542 20846 60790 20874
rect 59516 20761 59544 20846
rect 60790 20823 60846 20832
rect 59502 20752 59558 20761
rect 59502 20687 59558 20696
rect 57386 17896 57442 17905
rect 57386 17831 57442 17840
rect 60424 17724 60476 17730
rect 60424 17666 60476 17672
rect 60436 9304 60464 17666
rect 61540 17118 61568 20860
rect 62552 18478 62580 20860
rect 62540 18472 62592 18478
rect 62540 18414 62592 18420
rect 63564 18410 63592 20860
rect 63552 18404 63604 18410
rect 63552 18346 63604 18352
rect 65680 18070 65708 20860
rect 66494 19256 66550 19265
rect 66494 19191 66550 19200
rect 66508 19158 66536 19191
rect 66496 19152 66548 19158
rect 66496 19094 66548 19100
rect 66692 18274 66720 20860
rect 66680 18268 66732 18274
rect 66680 18210 66732 18216
rect 65668 18064 65720 18070
rect 65668 18006 65720 18012
rect 67704 18002 67732 20860
rect 67692 17996 67744 18002
rect 67692 17938 67744 17944
rect 68808 17934 68836 20860
rect 68796 17928 68848 17934
rect 68796 17870 68848 17876
rect 69820 17798 69848 20860
rect 69992 18472 70044 18478
rect 69992 18414 70044 18420
rect 69808 17792 69860 17798
rect 69808 17734 69860 17740
rect 61528 17112 61580 17118
rect 61528 17054 61580 17060
rect 70004 11746 70032 18414
rect 70832 17866 70860 20860
rect 71096 18268 71148 18274
rect 71096 18210 71148 18216
rect 70820 17860 70872 17866
rect 70820 17802 70872 17808
rect 65760 11740 65812 11746
rect 65760 11682 65812 11688
rect 69992 11740 70044 11746
rect 69992 11682 70044 11688
rect 65772 9304 65800 11682
rect 71108 9304 71136 18210
rect 71844 17662 71872 20860
rect 72948 18274 72976 20860
rect 73960 18478 73988 20860
rect 73948 18472 74000 18478
rect 73948 18414 74000 18420
rect 72936 18268 72988 18274
rect 72936 18210 72988 18216
rect 74972 17730 75000 20860
rect 75984 18342 76012 20860
rect 75972 18336 76024 18342
rect 75972 18278 76024 18284
rect 77088 18206 77116 20860
rect 77076 18200 77128 18206
rect 77076 18142 77128 18148
rect 78100 18138 78128 20860
rect 78928 20846 79126 20874
rect 78088 18132 78140 18138
rect 78088 18074 78140 18080
rect 74960 17724 75012 17730
rect 74960 17666 75012 17672
rect 71832 17656 71884 17662
rect 71832 17598 71884 17604
rect 78928 12290 78956 20846
rect 80124 17526 80152 20860
rect 80296 18200 80348 18206
rect 80296 18142 80348 18148
rect 79192 17520 79244 17526
rect 79192 17462 79244 17468
rect 80112 17520 80164 17526
rect 80112 17462 80164 17468
rect 79204 12358 79232 17462
rect 79192 12352 79244 12358
rect 79192 12294 79244 12300
rect 78916 12284 78968 12290
rect 78916 12226 78968 12232
rect 80308 12154 80336 18142
rect 81228 17798 81256 20860
rect 81768 18336 81820 18342
rect 81768 18278 81820 18284
rect 81216 17792 81268 17798
rect 81216 17734 81268 17740
rect 76432 12148 76484 12154
rect 76432 12090 76484 12096
rect 80296 12148 80348 12154
rect 80296 12090 80348 12096
rect 76444 9304 76472 12090
rect 81780 9304 81808 18278
rect 82240 18274 82268 20860
rect 83252 18342 83280 20860
rect 83240 18336 83292 18342
rect 83240 18278 83292 18284
rect 82228 18268 82280 18274
rect 82228 18210 82280 18216
rect 84264 18206 84292 20860
rect 86472 19838 86500 46158
rect 86460 19832 86512 19838
rect 86460 19774 86512 19780
rect 87852 19537 87880 46294
rect 87932 46284 87984 46290
rect 87932 46226 87984 46232
rect 87944 24138 87972 46226
rect 88390 46184 88446 46193
rect 88390 46119 88446 46128
rect 88114 44960 88170 44969
rect 88114 44895 88170 44904
rect 88128 43201 88156 44895
rect 88404 44425 88432 46119
rect 88574 45504 88630 45513
rect 88574 45439 88630 45448
rect 88482 44824 88538 44833
rect 88482 44759 88538 44768
rect 88390 44416 88446 44425
rect 88390 44351 88446 44360
rect 88496 43994 88524 44759
rect 88312 43966 88524 43994
rect 88114 43192 88170 43201
rect 88114 43127 88170 43136
rect 88312 42657 88340 43966
rect 88482 43872 88538 43881
rect 88588 43858 88616 45439
rect 88538 43830 88616 43858
rect 88482 43807 88538 43816
rect 88574 43736 88630 43745
rect 88574 43671 88630 43680
rect 88390 43464 88446 43473
rect 88390 43399 88446 43408
rect 88298 42648 88354 42657
rect 88298 42583 88354 42592
rect 88298 42240 88354 42249
rect 88298 42175 88354 42184
rect 88312 40209 88340 42175
rect 88404 41433 88432 43399
rect 88482 42104 88538 42113
rect 88588 42090 88616 43671
rect 88666 42512 88722 42521
rect 88666 42447 88722 42456
rect 88538 42062 88616 42090
rect 88482 42039 88538 42048
rect 88390 41424 88446 41433
rect 88390 41359 88446 41368
rect 88482 40880 88538 40889
rect 88680 40866 88708 42447
rect 88758 41288 88814 41297
rect 88758 41223 88814 41232
rect 88538 40838 88708 40866
rect 88482 40815 88538 40824
rect 88390 40608 88446 40617
rect 88390 40543 88446 40552
rect 88298 40200 88354 40209
rect 88298 40135 88354 40144
rect 88404 39121 88432 40543
rect 88772 40186 88800 41223
rect 88496 40158 88800 40186
rect 88496 39665 88524 40158
rect 88574 40064 88630 40073
rect 88574 39999 88630 40008
rect 88482 39656 88538 39665
rect 88482 39591 88538 39600
rect 88390 39112 88446 39121
rect 88390 39047 88446 39056
rect 88482 38432 88538 38441
rect 88588 38418 88616 39999
rect 88666 39384 88722 39393
rect 88666 39319 88722 39328
rect 88538 38390 88616 38418
rect 88482 38367 88538 38376
rect 88482 38296 88538 38305
rect 88680 38282 88708 39319
rect 88758 38840 88814 38849
rect 88758 38775 88814 38784
rect 88538 38254 88708 38282
rect 88482 38231 88538 38240
rect 88574 38160 88630 38169
rect 88574 38095 88630 38104
rect 88482 37888 88538 37897
rect 88482 37823 88538 37832
rect 88208 37376 88260 37382
rect 88208 37318 88260 37324
rect 88220 37217 88248 37318
rect 88206 37208 88262 37217
rect 88206 37143 88262 37152
rect 88390 36528 88446 36537
rect 88390 36463 88446 36472
rect 88298 35304 88354 35313
rect 88298 35239 88354 35248
rect 88312 33681 88340 35239
rect 88404 34905 88432 36463
rect 88496 36129 88524 37823
rect 88588 36673 88616 38095
rect 88772 37382 88800 38775
rect 88760 37376 88812 37382
rect 88760 37318 88812 37324
rect 88666 36936 88722 36945
rect 88666 36871 88722 36880
rect 88574 36664 88630 36673
rect 88574 36599 88630 36608
rect 88482 36120 88538 36129
rect 88482 36055 88538 36064
rect 88680 35834 88708 36871
rect 88496 35806 88708 35834
rect 88496 35449 88524 35806
rect 88666 35712 88722 35721
rect 88666 35647 88722 35656
rect 88482 35440 88538 35449
rect 88482 35375 88538 35384
rect 88390 34896 88446 34905
rect 88390 34831 88446 34840
rect 88574 34488 88630 34497
rect 88574 34423 88630 34432
rect 88588 34066 88616 34423
rect 88680 34225 88708 35647
rect 88666 34216 88722 34225
rect 88666 34151 88722 34160
rect 88496 34038 88616 34066
rect 88390 33808 88446 33817
rect 88390 33743 88446 33752
rect 88298 33672 88354 33681
rect 88298 33607 88354 33616
rect 88404 31913 88432 33743
rect 88496 33137 88524 34038
rect 88574 33944 88630 33953
rect 88574 33879 88630 33888
rect 88482 33128 88538 33137
rect 88482 33063 88538 33072
rect 88482 32448 88538 32457
rect 88588 32434 88616 33879
rect 88666 32720 88722 32729
rect 88666 32655 88722 32664
rect 88538 32406 88616 32434
rect 88482 32383 88538 32392
rect 88482 32312 88538 32321
rect 88482 32247 88538 32256
rect 88390 31904 88446 31913
rect 88390 31839 88446 31848
rect 88390 30952 88446 30961
rect 88390 30887 88446 30896
rect 88404 29465 88432 30887
rect 88496 30689 88524 32247
rect 88574 31496 88630 31505
rect 88574 31431 88630 31440
rect 88482 30680 88538 30689
rect 88482 30615 88538 30624
rect 88482 30136 88538 30145
rect 88588 30122 88616 31431
rect 88680 31233 88708 32655
rect 88666 31224 88722 31233
rect 88666 31159 88722 31168
rect 88666 30272 88722 30281
rect 88666 30207 88722 30216
rect 88538 30094 88616 30122
rect 88482 30071 88538 30080
rect 88574 29728 88630 29737
rect 88574 29663 88630 29672
rect 88390 29456 88446 29465
rect 88390 29391 88446 29400
rect 88588 29034 88616 29663
rect 88404 29006 88616 29034
rect 88404 28785 88432 29006
rect 88482 28912 88538 28921
rect 88680 28898 88708 30207
rect 88758 29048 88814 29057
rect 88758 28983 88814 28992
rect 88538 28870 88708 28898
rect 88482 28847 88538 28856
rect 88390 28776 88446 28785
rect 88390 28711 88446 28720
rect 88574 28504 88630 28513
rect 88574 28439 88630 28448
rect 88390 28232 88446 28241
rect 88390 28167 88446 28176
rect 88300 27720 88352 27726
rect 88298 27688 88300 27697
rect 88352 27688 88354 27697
rect 88298 27623 88354 27632
rect 88298 26872 88354 26881
rect 88298 26807 88354 26816
rect 88312 25249 88340 26807
rect 88404 26473 88432 28167
rect 88588 27402 88616 28439
rect 88772 27726 88800 28983
rect 88760 27720 88812 27726
rect 88760 27662 88812 27668
rect 88496 27374 88616 27402
rect 88496 27153 88524 27374
rect 88574 27280 88630 27289
rect 88574 27215 88630 27224
rect 88482 27144 88538 27153
rect 88482 27079 88538 27088
rect 88390 26464 88446 26473
rect 88390 26399 88446 26408
rect 88482 25920 88538 25929
rect 88588 25906 88616 27215
rect 88666 26056 88722 26065
rect 88666 25991 88722 26000
rect 88538 25878 88616 25906
rect 88482 25855 88538 25864
rect 88574 25648 88630 25657
rect 88574 25583 88630 25592
rect 88298 25240 88354 25249
rect 88588 25226 88616 25583
rect 88298 25175 88354 25184
rect 88404 25198 88616 25226
rect 88404 24161 88432 25198
rect 88482 25104 88538 25113
rect 88680 25090 88708 25991
rect 88538 25062 88708 25090
rect 88482 25039 88538 25048
rect 88574 24832 88630 24841
rect 88574 24767 88630 24776
rect 88390 24152 88446 24161
rect 87944 24110 88064 24138
rect 87930 24016 87986 24025
rect 87930 23951 87986 23960
rect 87944 22937 87972 23951
rect 87930 22928 87986 22937
rect 87930 22863 87986 22872
rect 88036 21033 88064 24110
rect 88390 24087 88446 24096
rect 88482 23472 88538 23481
rect 88588 23458 88616 24767
rect 88666 23608 88722 23617
rect 88666 23543 88722 23552
rect 88538 23430 88616 23458
rect 88482 23407 88538 23416
rect 88574 22928 88630 22937
rect 88574 22863 88630 22872
rect 88482 22656 88538 22665
rect 88482 22591 88538 22600
rect 88496 21169 88524 22591
rect 88588 21713 88616 22863
rect 88680 22257 88708 23543
rect 88760 22620 88812 22626
rect 88760 22562 88812 22568
rect 88772 22529 88800 22562
rect 88758 22520 88814 22529
rect 88758 22455 88814 22464
rect 88666 22248 88722 22257
rect 88666 22183 88722 22192
rect 88574 21704 88630 21713
rect 88574 21639 88630 21648
rect 88576 21260 88628 21266
rect 88576 21202 88628 21208
rect 88482 21160 88538 21169
rect 88482 21095 88538 21104
rect 88022 21024 88078 21033
rect 88022 20959 88078 20968
rect 88588 20761 88616 21202
rect 88574 20752 88630 20761
rect 88574 20687 88630 20696
rect 88576 19832 88628 19838
rect 88574 19800 88576 19809
rect 88628 19800 88630 19809
rect 88574 19735 88630 19744
rect 87838 19528 87894 19537
rect 87838 19463 87894 19472
rect 94660 18410 94688 18956
rect 100180 18410 100208 18956
rect 94648 18404 94700 18410
rect 94648 18346 94700 18352
rect 95384 18404 95436 18410
rect 95384 18346 95436 18352
rect 100168 18404 100220 18410
rect 100168 18346 100220 18352
rect 84344 18268 84396 18274
rect 84344 18210 84396 18216
rect 84252 18200 84304 18206
rect 84252 18142 84304 18148
rect 84356 12902 84384 18210
rect 92440 17792 92492 17798
rect 92440 17734 92492 17740
rect 84344 12896 84396 12902
rect 84344 12838 84396 12844
rect 87104 12896 87156 12902
rect 87104 12838 87156 12844
rect 87116 9304 87144 12838
rect 92452 9304 92480 17734
rect 95396 17050 95424 18346
rect 105792 17118 105820 18956
rect 113784 17860 113836 17866
rect 113784 17802 113836 17808
rect 108448 17792 108500 17798
rect 108448 17734 108500 17740
rect 105780 17112 105832 17118
rect 105780 17054 105832 17060
rect 95384 17044 95436 17050
rect 95384 16986 95436 16992
rect 97776 12352 97828 12358
rect 97776 12294 97828 12300
rect 97788 9304 97816 12294
rect 103112 12284 103164 12290
rect 103112 12226 103164 12232
rect 103124 9304 103152 12226
rect 108460 9304 108488 17734
rect 113796 9304 113824 17802
rect 117016 17118 117044 18956
rect 119684 18478 119712 46958
rect 122800 46556 122852 46562
rect 122800 46498 122852 46504
rect 129148 46556 129200 46562
rect 129148 46498 129200 46504
rect 122340 46488 122392 46494
rect 122340 46430 122392 46436
rect 121694 45096 121750 45105
rect 121694 45031 121750 45040
rect 121708 44930 121736 45031
rect 121696 44924 121748 44930
rect 121696 44866 121748 44872
rect 121694 44824 121750 44833
rect 121694 44759 121696 44768
rect 121748 44759 121750 44768
rect 121696 44730 121748 44736
rect 121694 43464 121750 43473
rect 121694 43399 121696 43408
rect 121748 43399 121750 43408
rect 121696 43370 121748 43376
rect 121694 42240 121750 42249
rect 121694 42175 121750 42184
rect 121708 42074 121736 42175
rect 121696 42068 121748 42074
rect 121696 42010 121748 42016
rect 121694 40880 121750 40889
rect 121694 40815 121750 40824
rect 121708 40714 121736 40815
rect 121696 40708 121748 40714
rect 121696 40650 121748 40656
rect 121786 38840 121842 38849
rect 121786 38775 121842 38784
rect 121800 38470 121828 38775
rect 121788 38464 121840 38470
rect 121694 38432 121750 38441
rect 121788 38406 121840 38412
rect 121694 38367 121750 38376
rect 121708 38266 121736 38367
rect 121696 38260 121748 38266
rect 121696 38202 121748 38208
rect 121694 37888 121750 37897
rect 121694 37823 121696 37832
rect 121748 37823 121750 37832
rect 121696 37794 121748 37800
rect 121694 35304 121750 35313
rect 121694 35239 121750 35248
rect 121708 35138 121736 35239
rect 121696 35132 121748 35138
rect 121696 35074 121748 35080
rect 121694 34488 121750 34497
rect 121694 34423 121750 34432
rect 121708 34050 121736 34423
rect 121696 34044 121748 34050
rect 121696 33986 121748 33992
rect 121694 33808 121750 33817
rect 121694 33743 121696 33752
rect 121748 33743 121750 33752
rect 121696 33714 121748 33720
rect 121694 32448 121750 32457
rect 121694 32383 121696 32392
rect 121748 32383 121750 32392
rect 121696 32354 121748 32360
rect 121694 31224 121750 31233
rect 121694 31159 121750 31168
rect 121708 31058 121736 31159
rect 121696 31052 121748 31058
rect 121696 30994 121748 31000
rect 121694 29184 121750 29193
rect 121694 29119 121750 29128
rect 121708 28882 121736 29119
rect 121696 28876 121748 28882
rect 121696 28818 121748 28824
rect 121694 28640 121750 28649
rect 121694 28575 121750 28584
rect 121708 28542 121736 28575
rect 121696 28536 121748 28542
rect 121696 28478 121748 28484
rect 121694 28232 121750 28241
rect 121694 28167 121696 28176
rect 121748 28167 121750 28176
rect 121696 28138 121748 28144
rect 121694 24832 121750 24841
rect 121694 24767 121750 24776
rect 121708 24258 121736 24767
rect 121696 24252 121748 24258
rect 121696 24194 121748 24200
rect 122352 19537 122380 46430
rect 122432 46420 122484 46426
rect 122432 46362 122484 46368
rect 122444 20761 122472 46362
rect 122524 46352 122576 46358
rect 122524 46294 122576 46300
rect 122536 39914 122564 46294
rect 122708 46216 122760 46222
rect 122708 46158 122760 46164
rect 122536 39886 122656 39914
rect 122524 39212 122576 39218
rect 122524 39154 122576 39160
rect 122430 20752 122486 20761
rect 122430 20687 122486 20696
rect 122536 19809 122564 39154
rect 122628 21169 122656 39886
rect 122720 21985 122748 46158
rect 122812 39218 122840 46498
rect 127676 46488 127728 46494
rect 127676 46430 127728 46436
rect 126480 46284 126532 46290
rect 126480 46226 126532 46232
rect 122982 46184 123038 46193
rect 122892 46148 122944 46154
rect 123038 46142 123208 46170
rect 122982 46119 123038 46128
rect 122892 46090 122944 46096
rect 122800 39212 122852 39218
rect 122800 39154 122852 39160
rect 122904 22529 122932 46090
rect 122982 45504 123038 45513
rect 123038 45462 123116 45490
rect 122982 45439 123038 45448
rect 123088 44289 123116 45462
rect 123180 44425 123208 46142
rect 123536 44924 123588 44930
rect 123536 44866 123588 44872
rect 123352 44788 123404 44794
rect 123352 44730 123404 44736
rect 123166 44416 123222 44425
rect 123166 44351 123222 44360
rect 123074 44280 123130 44289
rect 123074 44215 123130 44224
rect 122982 43736 123038 43745
rect 122982 43671 123038 43680
rect 122996 43450 123024 43671
rect 122996 43422 123116 43450
rect 122982 42512 123038 42521
rect 122982 42447 123038 42456
rect 122996 42226 123024 42447
rect 123088 42385 123116 43422
rect 123364 43065 123392 44730
rect 123548 43201 123576 44866
rect 124364 43428 124416 43434
rect 124364 43370 124416 43376
rect 123534 43192 123590 43201
rect 123534 43127 123590 43136
rect 123350 43056 123406 43065
rect 123350 42991 123406 43000
rect 123074 42376 123130 42385
rect 123074 42311 123130 42320
rect 122996 42198 123208 42226
rect 123180 41297 123208 42198
rect 124272 42068 124324 42074
rect 124272 42010 124324 42016
rect 122982 41288 123038 41297
rect 123166 41288 123222 41297
rect 123038 41246 123116 41274
rect 122982 41223 123038 41232
rect 123088 39937 123116 41246
rect 123166 41223 123222 41232
rect 124284 40481 124312 42010
rect 124376 41977 124404 43370
rect 124362 41968 124418 41977
rect 124362 41903 124418 41912
rect 124364 40708 124416 40714
rect 124364 40650 124416 40656
rect 124270 40472 124326 40481
rect 124270 40407 124326 40416
rect 123166 40064 123222 40073
rect 123166 39999 123222 40008
rect 123074 39928 123130 39937
rect 123074 39863 123130 39872
rect 122982 39384 123038 39393
rect 123038 39342 123116 39370
rect 122982 39319 123038 39328
rect 123088 38305 123116 39342
rect 123180 38985 123208 39999
rect 124376 39121 124404 40650
rect 124362 39112 124418 39121
rect 124362 39047 124418 39056
rect 123166 38976 123222 38985
rect 123166 38911 123222 38920
rect 123904 38464 123956 38470
rect 123904 38406 123956 38412
rect 123074 38296 123130 38305
rect 123074 38231 123130 38240
rect 123444 38260 123496 38266
rect 123444 38202 123496 38208
rect 123456 37081 123484 38202
rect 123916 37761 123944 38406
rect 124364 37852 124416 37858
rect 124364 37794 124416 37800
rect 123902 37752 123958 37761
rect 123902 37687 123958 37696
rect 123442 37072 123498 37081
rect 123442 37007 123498 37016
rect 122982 36936 123038 36945
rect 123038 36894 123116 36922
rect 122982 36871 123038 36880
rect 123088 35993 123116 36894
rect 123258 36528 123314 36537
rect 123258 36463 123314 36472
rect 123074 35984 123130 35993
rect 123074 35919 123130 35928
rect 122982 35712 123038 35721
rect 122982 35647 123038 35656
rect 122996 35154 123024 35647
rect 122996 35126 123208 35154
rect 123180 34633 123208 35126
rect 123272 34905 123300 36463
rect 124376 36401 124404 37794
rect 124362 36392 124418 36401
rect 124362 36327 124418 36336
rect 123628 35132 123680 35138
rect 123628 35074 123680 35080
rect 123258 34896 123314 34905
rect 123258 34831 123314 34840
rect 123166 34624 123222 34633
rect 123166 34559 123222 34568
rect 122982 33944 123038 33953
rect 123038 33902 123116 33930
rect 122982 33879 123038 33888
rect 123088 33001 123116 33902
rect 123640 33681 123668 35074
rect 124364 34044 124416 34050
rect 124364 33986 124416 33992
rect 124272 33772 124324 33778
rect 124272 33714 124324 33720
rect 123626 33672 123682 33681
rect 123626 33607 123682 33616
rect 123074 32992 123130 33001
rect 123074 32927 123130 32936
rect 122982 32856 123038 32865
rect 122982 32791 123038 32800
rect 122996 32434 123024 32791
rect 122996 32406 123116 32434
rect 123088 31777 123116 32406
rect 123996 32412 124048 32418
rect 123996 32354 124048 32360
rect 123074 31768 123130 31777
rect 123074 31703 123130 31712
rect 122982 31496 123038 31505
rect 123038 31454 123116 31482
rect 122982 31431 123038 31440
rect 123088 30553 123116 31454
rect 124008 30689 124036 32354
rect 124284 32185 124312 33714
rect 124376 33545 124404 33986
rect 124362 33536 124418 33545
rect 124362 33471 124418 33480
rect 124270 32176 124326 32185
rect 124270 32111 124326 32120
rect 124364 31052 124416 31058
rect 124364 30994 124416 31000
rect 123994 30680 124050 30689
rect 123994 30615 124050 30624
rect 123074 30544 123130 30553
rect 123074 30479 123130 30488
rect 123166 30272 123222 30281
rect 123166 30207 123222 30216
rect 122982 29728 123038 29737
rect 123038 29686 123116 29714
rect 122982 29663 123038 29672
rect 123088 28785 123116 29686
rect 123180 29329 123208 30207
rect 124376 29465 124404 30994
rect 124362 29456 124418 29465
rect 124362 29391 124418 29400
rect 123166 29320 123222 29329
rect 123166 29255 123222 29264
rect 123536 28876 123588 28882
rect 123536 28818 123588 28824
rect 123074 28776 123130 28785
rect 123074 28711 123130 28720
rect 123548 28105 123576 28818
rect 124364 28536 124416 28542
rect 124364 28478 124416 28484
rect 124088 28196 124140 28202
rect 124088 28138 124140 28144
rect 123534 28096 123590 28105
rect 123534 28031 123590 28040
rect 122982 27280 123038 27289
rect 123038 27238 123116 27266
rect 122982 27215 123038 27224
rect 123088 26337 123116 27238
rect 123258 26872 123314 26881
rect 123258 26807 123314 26816
rect 123074 26328 123130 26337
rect 123074 26263 123130 26272
rect 123166 26056 123222 26065
rect 123166 25991 123222 26000
rect 122982 25512 123038 25521
rect 123038 25470 123116 25498
rect 122982 25447 123038 25456
rect 123088 24569 123116 25470
rect 123180 25113 123208 25991
rect 123272 25249 123300 26807
rect 124100 26745 124128 28138
rect 124376 27561 124404 28478
rect 124362 27552 124418 27561
rect 124362 27487 124418 27496
rect 124086 26736 124142 26745
rect 124086 26671 124142 26680
rect 123258 25240 123314 25249
rect 123258 25175 123314 25184
rect 123166 25104 123222 25113
rect 123166 25039 123222 25048
rect 123074 24560 123130 24569
rect 123074 24495 123130 24504
rect 123444 24252 123496 24258
rect 123444 24194 123496 24200
rect 122982 24152 123038 24161
rect 123038 24110 123116 24138
rect 122982 24087 123038 24096
rect 123088 23345 123116 24110
rect 123456 23889 123484 24194
rect 123442 23880 123498 23889
rect 123442 23815 123498 23824
rect 123258 23608 123314 23617
rect 123258 23543 123314 23552
rect 123074 23336 123130 23345
rect 123074 23271 123130 23280
rect 122982 23064 123038 23073
rect 122982 22999 123038 23008
rect 122996 22642 123024 22999
rect 123166 22656 123222 22665
rect 122996 22614 123116 22642
rect 122890 22520 122946 22529
rect 122890 22455 122946 22464
rect 123088 22121 123116 22614
rect 123166 22591 123222 22600
rect 123074 22112 123130 22121
rect 123074 22047 123130 22056
rect 122706 21976 122762 21985
rect 122706 21911 122762 21920
rect 123180 21169 123208 22591
rect 123272 22529 123300 23543
rect 123258 22520 123314 22529
rect 123258 22455 123314 22464
rect 122614 21160 122670 21169
rect 122614 21095 122670 21104
rect 123166 21160 123222 21169
rect 123166 21095 123222 21104
rect 122522 19800 122578 19809
rect 122522 19735 122578 19744
rect 122338 19528 122394 19537
rect 122338 19463 122394 19472
rect 119672 18472 119724 18478
rect 119672 18414 119724 18420
rect 124456 17996 124508 18002
rect 124456 17938 124508 17944
rect 119120 17928 119172 17934
rect 119120 17870 119172 17876
rect 117004 17112 117056 17118
rect 117004 17054 117056 17060
rect 119132 9304 119160 17870
rect 124468 9304 124496 17938
rect 126492 17118 126520 46226
rect 127688 44796 127716 46430
rect 129160 44796 129188 46498
rect 130620 46420 130672 46426
rect 130620 46362 130672 46368
rect 130632 44796 130660 46362
rect 132092 46352 132144 46358
rect 132092 46294 132144 46300
rect 132104 44796 132132 46294
rect 136600 46284 136652 46290
rect 136600 46226 136652 46232
rect 133656 46216 133708 46222
rect 133656 46158 133708 46164
rect 133668 44796 133696 46158
rect 135128 46148 135180 46154
rect 135128 46090 135180 46096
rect 135140 44796 135168 46090
rect 136612 44796 136640 46226
rect 138176 44796 138204 50850
rect 163108 46850 163136 54415
rect 163752 49758 163780 62847
rect 163830 61688 163886 61697
rect 163830 61623 163886 61632
rect 163844 50166 163872 61623
rect 165118 60464 165174 60473
rect 165118 60399 165174 60408
rect 164382 59240 164438 59249
rect 164382 59175 164438 59184
rect 164396 58598 164424 59175
rect 164384 58592 164436 58598
rect 164384 58534 164436 58540
rect 164382 58016 164438 58025
rect 164382 57951 164438 57960
rect 164396 57170 164424 57951
rect 164384 57164 164436 57170
rect 164384 57106 164436 57112
rect 165026 56792 165082 56801
rect 165026 56727 165082 56736
rect 164566 55568 164622 55577
rect 164566 55503 164622 55512
rect 163832 50160 163884 50166
rect 163832 50102 163884 50108
rect 163740 49752 163792 49758
rect 163740 49694 163792 49700
rect 163108 46822 163872 46850
rect 142670 46728 142726 46737
rect 163844 46714 163872 46822
rect 164580 46714 164608 55503
rect 165040 46714 165068 56727
rect 165132 50234 165160 60399
rect 166040 58592 166092 58598
rect 166040 58534 166092 58540
rect 165948 57164 166000 57170
rect 165948 57106 166000 57112
rect 165120 50228 165172 50234
rect 165120 50170 165172 50176
rect 165960 46714 165988 57106
rect 163844 46686 164226 46714
rect 164580 46686 164778 46714
rect 165040 46686 165330 46714
rect 165882 46686 165988 46714
rect 166052 46714 166080 58534
rect 166512 56801 166540 64042
rect 167064 58841 167092 64450
rect 167156 60881 167184 65402
rect 167340 64825 167368 68190
rect 190616 67506 190644 100558
rect 190984 97086 191012 100828
rect 191536 97834 191564 100828
rect 193468 100622 193496 106095
rect 193560 101302 193588 123503
rect 193548 101296 193600 101302
rect 193548 101238 193600 101244
rect 193456 100616 193508 100622
rect 193456 100558 193508 100564
rect 191524 97828 191576 97834
rect 191524 97770 191576 97776
rect 190972 97080 191024 97086
rect 190972 97022 191024 97028
rect 189960 67500 190012 67506
rect 189960 67442 190012 67448
rect 190604 67500 190656 67506
rect 190604 67442 190656 67448
rect 167880 66820 167932 66826
rect 167880 66762 167932 66768
rect 167326 64816 167382 64825
rect 167326 64751 167382 64760
rect 167892 62785 167920 66762
rect 167878 62776 167934 62785
rect 167878 62711 167934 62720
rect 167142 60872 167198 60881
rect 167142 60807 167198 60816
rect 167050 58832 167106 58841
rect 167050 58767 167106 58776
rect 189972 57986 190000 67442
rect 187936 57980 187988 57986
rect 187936 57922 187988 57928
rect 189960 57980 190012 57986
rect 189960 57922 190012 57928
rect 187948 57209 187976 57922
rect 187934 57200 187990 57209
rect 187934 57135 187990 57144
rect 166498 56792 166554 56801
rect 166498 56727 166554 56736
rect 168522 54480 168578 54489
rect 168522 54415 168578 54424
rect 167052 50228 167104 50234
rect 167052 50170 167104 50176
rect 166052 46686 166434 46714
rect 167064 46700 167092 50170
rect 167604 50160 167656 50166
rect 167604 50102 167656 50108
rect 167616 46700 167644 50102
rect 168156 49752 168208 49758
rect 168156 49694 168208 49700
rect 168168 46700 168196 49694
rect 168536 49554 168564 54415
rect 169904 50228 169956 50234
rect 169904 50170 169956 50176
rect 168708 50160 168760 50166
rect 168708 50102 168760 50108
rect 168524 49548 168576 49554
rect 168524 49490 168576 49496
rect 168720 46700 168748 50102
rect 169260 50092 169312 50098
rect 169260 50034 169312 50040
rect 169272 46700 169300 50034
rect 169916 46700 169944 50170
rect 170100 50166 170128 53908
rect 170088 50160 170140 50166
rect 170088 50102 170140 50108
rect 170468 50098 170496 53908
rect 170836 50234 170864 53908
rect 170928 53894 171310 53922
rect 170824 50228 170876 50234
rect 170824 50170 170876 50176
rect 170456 50092 170508 50098
rect 170456 50034 170508 50040
rect 170928 46714 170956 53894
rect 171664 50234 171692 53908
rect 171756 53894 172046 53922
rect 171008 50228 171060 50234
rect 171008 50170 171060 50176
rect 171652 50228 171704 50234
rect 171652 50170 171704 50176
rect 170482 46686 170956 46714
rect 171020 46700 171048 50170
rect 171756 46714 171784 53894
rect 172492 46714 172520 53908
rect 172860 46714 172888 53908
rect 171586 46686 171784 46714
rect 172138 46686 172520 46714
rect 172782 46686 172888 46714
rect 173228 46714 173256 53908
rect 173688 46714 173716 53908
rect 173964 53894 174070 53922
rect 174438 53894 174728 53922
rect 173964 51594 173992 53894
rect 173952 51588 174004 51594
rect 173952 51530 174004 51536
rect 174136 51588 174188 51594
rect 174136 51530 174188 51536
rect 174148 46714 174176 51530
rect 174700 46714 174728 53894
rect 174884 51526 174912 53908
rect 175252 51594 175280 53908
rect 175240 51588 175292 51594
rect 175240 51530 175292 51536
rect 174872 51520 174924 51526
rect 174872 51462 174924 51468
rect 175516 51520 175568 51526
rect 175516 51462 175568 51468
rect 175528 46714 175556 51462
rect 175620 50778 175648 53908
rect 175608 50772 175660 50778
rect 175608 50714 175660 50720
rect 176080 50370 176108 53908
rect 176160 51588 176212 51594
rect 176160 51530 176212 51536
rect 176068 50364 176120 50370
rect 176068 50306 176120 50312
rect 173228 46686 173334 46714
rect 173688 46686 173886 46714
rect 174148 46686 174438 46714
rect 174700 46686 174990 46714
rect 175528 46686 175634 46714
rect 176172 46700 176200 51530
rect 176448 50438 176476 53908
rect 176712 50772 176764 50778
rect 176712 50714 176764 50720
rect 176436 50432 176488 50438
rect 176436 50374 176488 50380
rect 176724 46700 176752 50714
rect 176816 50302 176844 53908
rect 177276 50506 177304 53908
rect 177264 50500 177316 50506
rect 177264 50442 177316 50448
rect 177644 50370 177672 53908
rect 178118 53894 178224 53922
rect 177816 50432 177868 50438
rect 177816 50374 177868 50380
rect 177264 50364 177316 50370
rect 177264 50306 177316 50312
rect 177632 50364 177684 50370
rect 177632 50306 177684 50312
rect 176804 50296 176856 50302
rect 176804 50238 176856 50244
rect 177276 46700 177304 50306
rect 177828 46700 177856 50374
rect 178196 50250 178224 53894
rect 178472 50438 178500 53908
rect 178840 50642 178868 53908
rect 179314 53894 179512 53922
rect 178828 50636 178880 50642
rect 178828 50578 178880 50584
rect 179012 50500 179064 50506
rect 179012 50442 179064 50448
rect 178460 50432 178512 50438
rect 178460 50374 178512 50380
rect 178196 50222 178316 50250
rect 178288 50166 178316 50222
rect 178460 50228 178512 50234
rect 178460 50170 178512 50176
rect 178276 50160 178328 50166
rect 178276 50102 178328 50108
rect 178472 46700 178500 50170
rect 179024 46700 179052 50442
rect 179484 50302 179512 53894
rect 179668 50574 179696 53908
rect 180036 50710 180064 53908
rect 180024 50704 180076 50710
rect 180024 50646 180076 50652
rect 179656 50568 179708 50574
rect 179656 50510 179708 50516
rect 180496 50370 180524 53908
rect 180878 53894 180984 53922
rect 180956 50794 180984 53894
rect 180956 50766 181168 50794
rect 180944 50636 180996 50642
rect 180944 50578 180996 50584
rect 180668 50432 180720 50438
rect 180668 50374 180720 50380
rect 179564 50364 179616 50370
rect 179564 50306 179616 50312
rect 180484 50364 180536 50370
rect 180484 50306 180536 50312
rect 179472 50296 179524 50302
rect 179472 50238 179524 50244
rect 179576 46700 179604 50306
rect 180116 50160 180168 50166
rect 180116 50102 180168 50108
rect 180128 46700 180156 50102
rect 180680 46700 180708 50374
rect 180956 50352 180984 50578
rect 180956 50324 181076 50352
rect 181048 46714 181076 50324
rect 181140 50030 181168 50766
rect 181232 50302 181260 53908
rect 181692 50506 181720 53908
rect 182074 53894 182364 53922
rect 182048 50704 182100 50710
rect 182048 50646 182100 50652
rect 182336 50658 182364 53894
rect 182428 50778 182456 53908
rect 182416 50772 182468 50778
rect 182416 50714 182468 50720
rect 181680 50500 181732 50506
rect 181680 50442 181732 50448
rect 181220 50296 181272 50302
rect 181220 50238 181272 50244
rect 181864 50228 181916 50234
rect 181864 50170 181916 50176
rect 181128 50024 181180 50030
rect 181128 49966 181180 49972
rect 181048 46686 181338 46714
rect 181876 46700 181904 50170
rect 182060 49010 182088 50646
rect 182336 50630 182548 50658
rect 182324 50568 182376 50574
rect 182324 50510 182376 50516
rect 182336 50114 182364 50510
rect 182336 50086 182456 50114
rect 182048 49004 182100 49010
rect 182048 48946 182100 48952
rect 182428 46700 182456 50086
rect 182520 49894 182548 50630
rect 182888 50438 182916 53908
rect 182876 50432 182928 50438
rect 182876 50374 182928 50380
rect 183256 50302 183284 53908
rect 183624 50574 183652 53908
rect 184084 50642 184112 53908
rect 184072 50636 184124 50642
rect 184072 50578 184124 50584
rect 183612 50568 183664 50574
rect 183612 50510 183664 50516
rect 184452 50506 184480 53908
rect 183428 50500 183480 50506
rect 183428 50442 183480 50448
rect 184440 50500 184492 50506
rect 184440 50442 184492 50448
rect 183244 50296 183296 50302
rect 183244 50238 183296 50244
rect 183440 49962 183468 50442
rect 184820 50370 184848 53908
rect 184992 50772 185044 50778
rect 184992 50714 185044 50720
rect 184900 50432 184952 50438
rect 184900 50374 184952 50380
rect 184808 50364 184860 50370
rect 184808 50306 184860 50312
rect 183520 50228 183572 50234
rect 183520 50170 183572 50176
rect 183428 49956 183480 49962
rect 183428 49898 183480 49904
rect 182508 49888 182560 49894
rect 182508 49830 182560 49836
rect 182968 49004 183020 49010
rect 182968 48946 183020 48952
rect 182980 46700 183008 48946
rect 183532 46700 183560 50170
rect 184716 50160 184768 50166
rect 184716 50102 184768 50108
rect 184164 50024 184216 50030
rect 184164 49966 184216 49972
rect 184176 46700 184204 49966
rect 184728 46700 184756 50102
rect 184912 50098 184940 50374
rect 185004 50166 185032 50714
rect 185280 50438 185308 53908
rect 185268 50432 185320 50438
rect 185268 50374 185320 50380
rect 185648 50302 185676 53908
rect 186280 50636 186332 50642
rect 186280 50578 186332 50584
rect 185636 50296 185688 50302
rect 185636 50238 185688 50244
rect 184992 50160 185044 50166
rect 184992 50102 185044 50108
rect 184900 50092 184952 50098
rect 184900 50034 184952 50040
rect 185268 49956 185320 49962
rect 185268 49898 185320 49904
rect 185280 46700 185308 49898
rect 185820 49888 185872 49894
rect 185820 49830 185872 49836
rect 185832 46700 185860 49830
rect 186292 49690 186320 50578
rect 188120 50568 188172 50574
rect 188120 50510 188172 50516
rect 186464 50500 186516 50506
rect 186464 50442 186516 50448
rect 186372 50160 186424 50166
rect 186372 50102 186424 50108
rect 186280 49684 186332 49690
rect 186280 49626 186332 49632
rect 186384 46700 186412 50102
rect 186476 49826 186504 50442
rect 187752 50432 187804 50438
rect 187752 50374 187804 50380
rect 187568 50228 187620 50234
rect 187568 50170 187620 50176
rect 187016 50092 187068 50098
rect 187016 50034 187068 50040
rect 186464 49820 186516 49826
rect 186464 49762 186516 49768
rect 187028 46700 187056 50034
rect 187580 46700 187608 50170
rect 187764 49962 187792 50374
rect 187752 49956 187804 49962
rect 187752 49898 187804 49904
rect 188132 46700 188160 50510
rect 189868 50364 189920 50370
rect 189868 50306 189920 50312
rect 189224 49820 189276 49826
rect 189224 49762 189276 49768
rect 188672 49684 188724 49690
rect 188672 49626 188724 49632
rect 188684 46700 188712 49626
rect 189236 46700 189264 49762
rect 189880 46700 189908 50306
rect 190972 50024 191024 50030
rect 190972 49966 191024 49972
rect 190420 49956 190472 49962
rect 190420 49898 190472 49904
rect 190432 46700 190460 49898
rect 190984 46700 191012 49966
rect 191524 49548 191576 49554
rect 191524 49490 191576 49496
rect 191536 46700 191564 49490
rect 142670 46663 142726 46672
rect 142684 44796 142712 46663
rect 145614 46592 145670 46601
rect 145614 46527 145670 46536
rect 144142 46320 144198 46329
rect 144142 46255 144198 46264
rect 144156 44796 144184 46255
rect 145628 44796 145656 46527
rect 147086 46456 147142 46465
rect 147086 46391 147142 46400
rect 148652 46420 148704 46426
rect 147100 44796 147128 46391
rect 148652 46362 148704 46368
rect 158220 46420 158272 46426
rect 158220 46362 158272 46368
rect 148664 44796 148692 46362
rect 150124 46352 150176 46358
rect 150124 46294 150176 46300
rect 150136 44796 150164 46294
rect 151596 46284 151648 46290
rect 151596 46226 151648 46232
rect 151608 44796 151636 46226
rect 153160 46148 153212 46154
rect 153160 46090 153212 46096
rect 153172 44796 153200 46090
rect 154658 44794 154764 44810
rect 154658 44788 154776 44794
rect 154658 44782 154724 44788
rect 154724 44730 154776 44736
rect 156840 44788 156892 44794
rect 156840 44730 156892 44736
rect 139726 44688 139782 44697
rect 139662 44646 139726 44674
rect 139726 44623 139782 44632
rect 140922 44688 140978 44697
rect 140978 44646 141134 44674
rect 140922 44623 140978 44632
rect 156130 44510 156512 44538
rect 156484 39762 156512 44510
rect 156472 39756 156524 39762
rect 156472 39698 156524 39704
rect 156852 22558 156880 44730
rect 156932 39756 156984 39762
rect 156932 39698 156984 39704
rect 156944 22626 156972 39698
rect 156932 22620 156984 22626
rect 156932 22562 156984 22568
rect 156840 22552 156892 22558
rect 156840 22494 156892 22500
rect 129698 21024 129754 21033
rect 129450 20982 129698 21010
rect 130710 21024 130766 21033
rect 130462 20982 130710 21010
rect 129698 20959 129754 20968
rect 130710 20959 130766 20968
rect 135862 20888 135918 20897
rect 135614 20860 135862 20874
rect 127412 18313 127440 20860
rect 127398 18304 127454 18313
rect 127398 18239 127454 18248
rect 128424 18041 128452 20860
rect 128410 18032 128466 18041
rect 128410 17967 128466 17976
rect 131460 17905 131488 20860
rect 132564 18177 132592 20860
rect 132550 18168 132606 18177
rect 132550 18103 132606 18112
rect 131446 17896 131502 17905
rect 131446 17831 131502 17840
rect 133576 17118 133604 20860
rect 134588 18410 134616 20860
rect 135600 20846 135862 20860
rect 134576 18404 134628 18410
rect 134576 18346 134628 18352
rect 126480 17112 126532 17118
rect 126480 17054 126532 17060
rect 133564 17112 133616 17118
rect 133564 17054 133616 17060
rect 135600 17050 135628 20846
rect 135862 20823 135918 20832
rect 138268 20846 138742 20874
rect 139754 20846 139860 20874
rect 135588 17044 135640 17050
rect 135588 16986 135640 16992
rect 138268 12358 138296 20846
rect 135128 12352 135180 12358
rect 135128 12294 135180 12300
rect 138256 12352 138308 12358
rect 138256 12294 138308 12300
rect 129792 12284 129844 12290
rect 129792 12226 129844 12232
rect 129804 9304 129832 12226
rect 135140 9304 135168 12294
rect 139832 12290 139860 20846
rect 140844 18002 140872 20860
rect 140832 17996 140884 18002
rect 140832 17938 140884 17944
rect 141856 17934 141884 20860
rect 141844 17928 141896 17934
rect 141844 17870 141896 17876
rect 142868 17866 142896 20860
rect 143776 18336 143828 18342
rect 143776 18278 143828 18284
rect 142856 17860 142908 17866
rect 142856 17802 142908 17808
rect 143788 12562 143816 18278
rect 143880 17798 143908 20860
rect 144984 18342 145012 20860
rect 145996 18342 146024 20860
rect 144972 18336 145024 18342
rect 144972 18278 145024 18284
rect 145156 18336 145208 18342
rect 145156 18278 145208 18284
rect 145984 18336 146036 18342
rect 145984 18278 146036 18284
rect 143868 17792 143920 17798
rect 143868 17734 143920 17740
rect 145168 12698 145196 18278
rect 145800 18064 145852 18070
rect 145800 18006 145852 18012
rect 145156 12692 145208 12698
rect 145156 12634 145208 12640
rect 143776 12556 143828 12562
rect 143776 12498 143828 12504
rect 140464 12352 140516 12358
rect 140464 12294 140516 12300
rect 139820 12284 139872 12290
rect 139820 12226 139872 12232
rect 140476 9304 140504 12294
rect 145812 9304 145840 18006
rect 147008 17798 147036 20860
rect 146996 17792 147048 17798
rect 146996 17734 147048 17740
rect 148020 17186 148048 20860
rect 149124 18070 149152 20860
rect 149112 18064 149164 18070
rect 149112 18006 149164 18012
rect 148008 17180 148060 17186
rect 148008 17122 148060 17128
rect 150136 12358 150164 20860
rect 150584 17180 150636 17186
rect 150584 17122 150636 17128
rect 150124 12352 150176 12358
rect 150124 12294 150176 12300
rect 150596 12154 150624 17122
rect 151148 12290 151176 20860
rect 152160 12358 152188 20860
rect 153264 12426 153292 20860
rect 154276 12494 154304 20860
rect 154816 17792 154868 17798
rect 154816 17734 154868 17740
rect 154828 12970 154856 17734
rect 154816 12964 154868 12970
rect 154816 12906 154868 12912
rect 155288 12630 155316 20860
rect 156300 12766 156328 20860
rect 158232 19838 158260 46362
rect 159600 46352 159652 46358
rect 159600 46294 159652 46300
rect 158312 46148 158364 46154
rect 158312 46090 158364 46096
rect 158324 21266 158352 46090
rect 159048 38600 159100 38606
rect 159048 38542 159100 38548
rect 159060 37897 159088 38542
rect 159046 37888 159102 37897
rect 159046 37823 159102 37832
rect 159048 28196 159100 28202
rect 159048 28138 159100 28144
rect 159060 26473 159088 28138
rect 159046 26464 159102 26473
rect 159046 26399 159102 26408
rect 158956 25204 159008 25210
rect 158956 25146 159008 25152
rect 158968 24161 158996 25146
rect 158954 24152 159010 24161
rect 158954 24087 159010 24096
rect 159048 22688 159100 22694
rect 159048 22630 159100 22636
rect 158312 21260 158364 21266
rect 158312 21202 158364 21208
rect 159060 21169 159088 22630
rect 159046 21160 159102 21169
rect 159046 21095 159102 21104
rect 158220 19832 158272 19838
rect 159612 19809 159640 46294
rect 159692 46284 159744 46290
rect 159692 46226 159744 46232
rect 159704 20761 159732 46226
rect 160242 46184 160298 46193
rect 160242 46119 160298 46128
rect 160150 44960 160206 44969
rect 160150 44895 160206 44904
rect 160058 44824 160114 44833
rect 160058 44759 160114 44768
rect 160072 43706 160100 44759
rect 159784 43700 159836 43706
rect 159784 43642 159836 43648
rect 160060 43700 160112 43706
rect 160060 43642 160112 43648
rect 159796 42657 159824 43642
rect 160164 43586 160192 44895
rect 160256 44425 160284 46119
rect 160334 45504 160390 45513
rect 160334 45439 160390 45448
rect 160242 44416 160298 44425
rect 160242 44351 160298 44360
rect 160242 43872 160298 43881
rect 160348 43858 160376 45439
rect 160298 43830 160376 43858
rect 160242 43807 160298 43816
rect 160334 43736 160390 43745
rect 160334 43671 160390 43680
rect 160072 43558 160192 43586
rect 160072 43201 160100 43558
rect 160150 43464 160206 43473
rect 160150 43399 160206 43408
rect 160058 43192 160114 43201
rect 160058 43127 160114 43136
rect 159782 42648 159838 42657
rect 159782 42583 159838 42592
rect 160058 42240 160114 42249
rect 160058 42175 160114 42184
rect 160072 40209 160100 42175
rect 160164 41433 160192 43399
rect 160348 42634 160376 43671
rect 160256 42606 160376 42634
rect 160256 42113 160284 42606
rect 160334 42512 160390 42521
rect 160334 42447 160390 42456
rect 160242 42104 160298 42113
rect 160242 42039 160298 42048
rect 160150 41424 160206 41433
rect 160150 41359 160206 41368
rect 160242 40880 160298 40889
rect 160348 40866 160376 42447
rect 160426 41288 160482 41297
rect 160426 41223 160482 41232
rect 160298 40838 160376 40866
rect 160242 40815 160298 40824
rect 160242 40608 160298 40617
rect 160242 40543 160298 40552
rect 160058 40200 160114 40209
rect 160058 40135 160114 40144
rect 160256 39121 160284 40543
rect 160334 40064 160390 40073
rect 160334 39999 160390 40008
rect 160242 39112 160298 39121
rect 160242 39047 160298 39056
rect 160242 38432 160298 38441
rect 160348 38418 160376 39999
rect 160440 39665 160468 41223
rect 160426 39656 160482 39665
rect 160426 39591 160482 39600
rect 160518 39384 160574 39393
rect 160518 39319 160574 39328
rect 160426 38840 160482 38849
rect 160426 38775 160482 38784
rect 160298 38390 160376 38418
rect 160242 38367 160298 38376
rect 160334 38296 160390 38305
rect 160334 38231 160390 38240
rect 160150 38024 160206 38033
rect 160150 37959 160206 37968
rect 160164 36129 160192 37959
rect 160348 37058 160376 38231
rect 160440 37897 160468 38775
rect 160532 38606 160560 39319
rect 160520 38600 160572 38606
rect 160520 38542 160572 38548
rect 160426 37888 160482 37897
rect 160426 37823 160482 37832
rect 160256 37030 160376 37058
rect 160256 36673 160284 37030
rect 160334 36936 160390 36945
rect 160334 36871 160390 36880
rect 160242 36664 160298 36673
rect 160242 36599 160298 36608
rect 160242 36528 160298 36537
rect 160242 36463 160298 36472
rect 160150 36120 160206 36129
rect 160150 36055 160206 36064
rect 160058 35168 160114 35177
rect 160058 35103 160114 35112
rect 160072 33681 160100 35103
rect 160256 34905 160284 36463
rect 160348 35449 160376 36871
rect 160426 35712 160482 35721
rect 160426 35647 160482 35656
rect 160334 35440 160390 35449
rect 160334 35375 160390 35384
rect 160242 34896 160298 34905
rect 160242 34831 160298 34840
rect 160334 34488 160390 34497
rect 160334 34423 160390 34432
rect 160150 33808 160206 33817
rect 160150 33743 160206 33752
rect 160058 33672 160114 33681
rect 160058 33607 160114 33616
rect 160058 32312 160114 32321
rect 160058 32247 160114 32256
rect 160072 30689 160100 32247
rect 160164 31913 160192 33743
rect 160242 33128 160298 33137
rect 160348 33114 160376 34423
rect 160440 34225 160468 35647
rect 160426 34216 160482 34225
rect 160426 34151 160482 34160
rect 160426 33944 160482 33953
rect 160426 33879 160482 33888
rect 160298 33086 160376 33114
rect 160242 33063 160298 33072
rect 160242 32448 160298 32457
rect 160440 32434 160468 33879
rect 160518 32720 160574 32729
rect 160518 32655 160574 32664
rect 160298 32406 160468 32434
rect 160242 32383 160298 32392
rect 160150 31904 160206 31913
rect 160150 31839 160206 31848
rect 160532 31618 160560 32655
rect 160256 31590 160560 31618
rect 160256 31233 160284 31590
rect 160334 31496 160390 31505
rect 160334 31431 160390 31440
rect 160242 31224 160298 31233
rect 160242 31159 160298 31168
rect 160150 30952 160206 30961
rect 160150 30887 160206 30896
rect 160058 30680 160114 30689
rect 160058 30615 160114 30624
rect 160164 29465 160192 30887
rect 160242 30136 160298 30145
rect 160348 30122 160376 31431
rect 160426 30272 160482 30281
rect 160426 30207 160482 30216
rect 160298 30094 160376 30122
rect 160242 30071 160298 30080
rect 160334 29728 160390 29737
rect 160334 29663 160390 29672
rect 160150 29456 160206 29465
rect 160150 29391 160206 29400
rect 160348 29170 160376 29663
rect 160164 29142 160376 29170
rect 160164 28241 160192 29142
rect 160440 29034 160468 30207
rect 160256 29006 160468 29034
rect 160518 29048 160574 29057
rect 160256 28921 160284 29006
rect 160518 28983 160574 28992
rect 160242 28912 160298 28921
rect 160242 28847 160298 28856
rect 160334 28504 160390 28513
rect 160334 28439 160390 28448
rect 160150 28232 160206 28241
rect 160150 28167 160206 28176
rect 160348 27402 160376 28439
rect 160532 28241 160560 28983
rect 160518 28232 160574 28241
rect 160518 28167 160574 28176
rect 160702 28232 160758 28241
rect 160702 28167 160704 28176
rect 160756 28167 160758 28176
rect 160704 28138 160756 28144
rect 160256 27374 160376 27402
rect 160256 27153 160284 27374
rect 160334 27280 160390 27289
rect 160334 27215 160390 27224
rect 160242 27144 160298 27153
rect 160242 27079 160298 27088
rect 160150 26872 160206 26881
rect 160150 26807 160206 26816
rect 160164 25249 160192 26807
rect 160242 25920 160298 25929
rect 160348 25906 160376 27215
rect 160426 26056 160482 26065
rect 160426 25991 160482 26000
rect 160298 25878 160376 25906
rect 160242 25855 160298 25864
rect 160334 25512 160390 25521
rect 160334 25447 160390 25456
rect 160150 25240 160206 25249
rect 160348 25210 160376 25447
rect 160150 25175 160206 25184
rect 160336 25204 160388 25210
rect 160336 25146 160388 25152
rect 160242 25104 160298 25113
rect 160440 25090 160468 25991
rect 160298 25062 160468 25090
rect 160242 25039 160298 25048
rect 160334 24832 160390 24841
rect 160334 24767 160390 24776
rect 160242 23472 160298 23481
rect 160348 23458 160376 24767
rect 160426 24288 160482 24297
rect 160426 24223 160482 24232
rect 160298 23430 160376 23458
rect 160242 23407 160298 23416
rect 160242 22928 160298 22937
rect 160440 22914 160468 24223
rect 160518 23608 160574 23617
rect 160518 23543 160574 23552
rect 160298 22886 160468 22914
rect 160242 22863 160298 22872
rect 160532 22665 160560 23543
rect 160610 22928 160666 22937
rect 160610 22863 160666 22872
rect 160518 22656 160574 22665
rect 160428 22620 160480 22626
rect 160518 22591 160574 22600
rect 160428 22562 160480 22568
rect 160440 22529 160468 22562
rect 160520 22552 160572 22558
rect 160426 22520 160482 22529
rect 160520 22494 160572 22500
rect 160426 22455 160482 22464
rect 160532 21985 160560 22494
rect 160518 21976 160574 21985
rect 160518 21911 160574 21920
rect 160624 21826 160652 22863
rect 160704 22688 160756 22694
rect 160702 22656 160704 22665
rect 160756 22656 160758 22665
rect 160702 22591 160758 22600
rect 160256 21798 160652 21826
rect 160256 21713 160284 21798
rect 160242 21704 160298 21713
rect 160242 21639 160298 21648
rect 160336 21260 160388 21266
rect 160336 21202 160388 21208
rect 160348 21169 160376 21202
rect 160334 21160 160390 21169
rect 160334 21095 160390 21104
rect 159690 20752 159746 20761
rect 159690 20687 159746 20696
rect 196872 20625 196900 190998
rect 196964 173042 196992 208911
rect 198238 185448 198294 185457
rect 198238 185383 198294 185392
rect 196952 173036 197004 173042
rect 196952 172978 197004 172984
rect 197596 164808 197648 164814
rect 197596 164750 197648 164756
rect 197608 161929 197636 164750
rect 197594 161920 197650 161929
rect 197594 161855 197650 161864
rect 196950 138392 197006 138401
rect 196950 138327 197006 138336
rect 196964 84710 196992 138327
rect 198252 91646 198280 185383
rect 201274 114728 201330 114737
rect 201274 114663 201330 114672
rect 201288 114601 201316 114663
rect 201274 114592 201330 114601
rect 201274 114527 201330 114536
rect 198240 91640 198292 91646
rect 198240 91582 198292 91588
rect 197594 91200 197650 91209
rect 197594 91135 197650 91144
rect 197608 90286 197636 91135
rect 197596 90280 197648 90286
rect 197596 90222 197648 90228
rect 196952 84704 197004 84710
rect 196952 84646 197004 84652
rect 197594 67672 197650 67681
rect 197594 67607 197650 67616
rect 197608 67506 197636 67607
rect 197596 67500 197648 67506
rect 197596 67442 197648 67448
rect 201274 44144 201330 44153
rect 201274 44079 201330 44088
rect 201288 43881 201316 44079
rect 201274 43872 201330 43881
rect 201274 43807 201330 43816
rect 196858 20616 196914 20625
rect 196858 20551 196914 20560
rect 160336 19832 160388 19838
rect 158220 19774 158272 19780
rect 159598 19800 159654 19809
rect 160336 19774 160388 19780
rect 159598 19735 159654 19744
rect 160348 19537 160376 19774
rect 160334 19528 160390 19537
rect 160334 19463 160390 19472
rect 168536 17050 168564 18956
rect 177828 17089 177856 18956
rect 187120 17118 187148 18956
rect 187108 17112 187160 17118
rect 177814 17080 177870 17089
rect 168524 17044 168576 17050
rect 187108 17054 187160 17060
rect 177814 17015 177870 17024
rect 168524 16986 168576 16992
rect 156472 12964 156524 12970
rect 156472 12906 156524 12912
rect 156288 12760 156340 12766
rect 156288 12702 156340 12708
rect 155276 12624 155328 12630
rect 155276 12566 155328 12572
rect 154264 12488 154316 12494
rect 154264 12430 154316 12436
rect 153252 12420 153304 12426
rect 153252 12362 153304 12368
rect 152148 12352 152200 12358
rect 152148 12294 152200 12300
rect 151136 12284 151188 12290
rect 151136 12226 151188 12232
rect 150584 12148 150636 12154
rect 150584 12090 150636 12096
rect 151136 12148 151188 12154
rect 151136 12090 151188 12096
rect 151148 9304 151176 12090
rect 156484 9304 156512 12906
rect 172480 12760 172532 12766
rect 172480 12702 172532 12708
rect 161808 12692 161860 12698
rect 161808 12634 161860 12640
rect 161820 9304 161848 12634
rect 167144 12556 167196 12562
rect 167144 12498 167196 12504
rect 167156 9304 167184 12498
rect 172492 9304 172520 12702
rect 177816 12624 177868 12630
rect 177816 12566 177868 12572
rect 177828 9304 177856 12566
rect 183152 12488 183204 12494
rect 183152 12430 183204 12436
rect 183164 9304 183192 12430
rect 188488 12420 188540 12426
rect 188488 12362 188540 12368
rect 188500 9304 188528 12362
rect 193824 12352 193876 12358
rect 193824 12294 193876 12300
rect 193836 9304 193864 12294
rect 199160 12284 199212 12290
rect 199160 12226 199212 12232
rect 199172 9304 199200 12226
rect 12490 8824 12546 9304
rect 17734 8824 17790 9304
rect 23070 8824 23126 9304
rect 28406 8824 28462 9304
rect 33742 8824 33798 9304
rect 39078 8824 39134 9304
rect 44414 8824 44470 9304
rect 49750 8824 49806 9304
rect 55086 8824 55142 9304
rect 60422 8824 60478 9304
rect 65758 8824 65814 9304
rect 71094 8824 71150 9304
rect 76430 8824 76486 9304
rect 81766 8824 81822 9304
rect 87102 8824 87158 9304
rect 92438 8824 92494 9304
rect 97774 8824 97830 9304
rect 103110 8824 103166 9304
rect 108446 8824 108502 9304
rect 113782 8824 113838 9304
rect 119118 8824 119174 9304
rect 124454 8824 124510 9304
rect 129790 8824 129846 9304
rect 135126 8824 135182 9304
rect 140462 8824 140518 9304
rect 145798 8824 145854 9304
rect 151134 8824 151190 9304
rect 156470 8824 156526 9304
rect 161806 8824 161862 9304
rect 167142 8824 167198 9304
rect 172478 8824 172534 9304
rect 177814 8824 177870 9304
rect 183150 8824 183206 9304
rect 188486 8824 188542 9304
rect 193822 8824 193878 9304
rect 199158 8824 199214 9304
<< via2 >>
rect 33374 213136 33430 213192
rect 39446 213136 39502 213192
rect 49290 210416 49346 210472
rect 13318 210144 13374 210200
rect 14698 188928 14754 188984
rect 13318 167712 13374 167768
rect 13410 146496 13466 146552
rect 13318 125280 13374 125336
rect 13318 104064 13374 104120
rect 13226 82848 13282 82904
rect 13318 61632 13374 61688
rect 49934 209872 49990 209928
rect 51314 209328 51370 209384
rect 49934 208920 49990 208976
rect 73210 210280 73266 210336
rect 120866 210416 120922 210472
rect 138806 210688 138862 210744
rect 88574 209872 88630 209928
rect 88666 208784 88722 208840
rect 51498 208376 51554 208432
rect 51314 208240 51370 208296
rect 51314 208104 51370 208160
rect 51406 207560 51462 207616
rect 51314 207016 51370 207072
rect 51314 206744 51370 206800
rect 88574 208240 88630 208296
rect 51498 207424 51554 207480
rect 88482 207152 88538 207208
rect 88666 207832 88722 207888
rect 88666 207696 88722 207752
rect 88482 206608 88538 206664
rect 88758 207152 88814 207208
rect 51498 206472 51554 206528
rect 51406 206064 51462 206120
rect 51314 205928 51370 205984
rect 88850 206608 88906 206664
rect 88758 206200 88814 206256
rect 87194 205928 87250 205984
rect 51590 205520 51646 205576
rect 51314 205248 51370 205304
rect 51498 205248 51554 205304
rect 88482 205792 88538 205848
rect 87194 204840 87250 204896
rect 51406 204704 51462 204760
rect 51590 204704 51646 204760
rect 51314 204024 51370 204080
rect 51314 203888 51370 203944
rect 51498 203616 51554 203672
rect 88482 203616 88538 203672
rect 88666 204840 88722 204896
rect 88666 204296 88722 204352
rect 51406 203344 51462 203400
rect 51406 203072 51462 203128
rect 51314 202936 51370 202992
rect 51314 202392 51370 202448
rect 50302 201984 50358 202040
rect 50486 201984 50542 202040
rect 51222 201848 51278 201904
rect 88758 203752 88814 203808
rect 88666 203480 88722 203536
rect 88482 202392 88538 202448
rect 88850 203208 88906 203264
rect 88574 202256 88630 202312
rect 51498 201848 51554 201904
rect 51406 201712 51462 201768
rect 88942 202664 88998 202720
rect 88850 202120 88906 202176
rect 51498 201304 51554 201360
rect 51314 201032 51370 201088
rect 51406 200760 51462 200816
rect 51314 200488 51370 200544
rect 51314 200216 51370 200272
rect 87194 201168 87250 201224
rect 88574 201440 88630 201496
rect 88482 200624 88538 200680
rect 88482 200080 88538 200136
rect 122982 209872 123038 209928
rect 122982 209328 123038 209384
rect 123074 208784 123130 208840
rect 145614 210280 145670 210336
rect 160334 210416 160390 210472
rect 123258 208376 123314 208432
rect 123074 208240 123130 208296
rect 122982 208104 123038 208160
rect 123166 207560 123222 207616
rect 123074 207016 123130 207072
rect 122982 206744 123038 206800
rect 122982 206472 123038 206528
rect 122154 205928 122210 205984
rect 123258 207424 123314 207480
rect 123166 206064 123222 206120
rect 123074 205928 123130 205984
rect 123258 205248 123314 205304
rect 123074 205112 123130 205168
rect 122982 204704 123038 204760
rect 122982 204160 123038 204216
rect 124362 204432 124418 204488
rect 123258 204024 123314 204080
rect 123166 203616 123222 203672
rect 123074 203344 123130 203400
rect 123074 202936 123130 202992
rect 122982 202392 123038 202448
rect 88666 200896 88722 200952
rect 51498 199944 51554 200000
rect 51498 199536 51554 199592
rect 51406 198992 51462 199048
rect 51406 198856 51462 198912
rect 51314 198720 51370 198776
rect 51314 198448 51370 198504
rect 88482 199400 88538 199456
rect 88758 200352 88814 200408
rect 88850 199808 88906 199864
rect 51590 197904 51646 197960
rect 51498 197632 51554 197688
rect 51406 197496 51462 197552
rect 51498 197360 51554 197416
rect 51406 196680 51462 196736
rect 51314 196408 51370 196464
rect 51314 196136 51370 196192
rect 88758 199264 88814 199320
rect 88942 199300 88944 199320
rect 88944 199300 88996 199320
rect 88996 199300 88998 199320
rect 88942 199264 88998 199300
rect 88942 198720 88998 198776
rect 88482 198176 88538 198232
rect 88666 198176 88722 198232
rect 87194 197632 87250 197688
rect 87194 197088 87250 197144
rect 88574 197632 88630 197688
rect 88482 196408 88538 196464
rect 51590 196272 51646 196328
rect 88482 196272 88538 196328
rect 88666 197088 88722 197144
rect 121786 196680 121842 196736
rect 89218 196408 89274 196464
rect 88574 195864 88630 195920
rect 51498 195728 51554 195784
rect 88482 195728 88538 195784
rect 51498 195592 51554 195648
rect 51406 195048 51462 195104
rect 51406 194776 51462 194832
rect 51314 194504 51370 194560
rect 51314 193824 51370 193880
rect 88390 195320 88446 195376
rect 88298 194232 88354 194288
rect 51590 194096 51646 194152
rect 51498 193688 51554 193744
rect 51406 193280 51462 193336
rect 51314 193008 51370 193064
rect 49934 185936 49990 185992
rect 50210 185256 50266 185312
rect 50118 184712 50174 184768
rect 50026 184168 50082 184224
rect 49934 183080 49990 183136
rect 20218 180496 20274 180552
rect 51498 192736 51554 192792
rect 51406 192056 51462 192112
rect 51406 191648 51462 191704
rect 51314 191512 51370 191568
rect 51314 190424 51370 190480
rect 51590 192328 51646 192384
rect 51682 192192 51738 192248
rect 51590 190968 51646 191024
rect 51498 190832 51554 190888
rect 51498 189880 51554 189936
rect 51406 189200 51462 189256
rect 51406 189064 51462 189120
rect 51314 188112 51370 188168
rect 51314 187840 51370 187896
rect 50670 187024 50726 187080
rect 51682 190288 51738 190344
rect 51590 189064 51646 189120
rect 51590 188792 51646 188848
rect 51498 187976 51554 188032
rect 51498 187568 51554 187624
rect 51406 187296 51462 187352
rect 51314 186072 51370 186128
rect 51590 186752 51646 186808
rect 51958 186480 52014 186536
rect 51498 185392 51554 185448
rect 51314 183624 51370 183680
rect 88482 194096 88538 194152
rect 89218 195184 89274 195240
rect 88666 194776 88722 194832
rect 88390 193416 88446 193472
rect 122246 194504 122302 194560
rect 88758 193688 88814 193744
rect 88482 192872 88538 192928
rect 88390 192600 88446 192656
rect 88298 192192 88354 192248
rect 88298 191376 88354 191432
rect 87194 191104 87250 191160
rect 88206 189744 88262 189800
rect 82226 184984 82282 185040
rect 77166 177232 77222 177288
rect 88850 193144 88906 193200
rect 122982 201848 123038 201904
rect 123258 203072 123314 203128
rect 123166 201848 123222 201904
rect 123258 201712 123314 201768
rect 123166 201304 123222 201360
rect 123074 201032 123130 201088
rect 122982 200760 123038 200816
rect 123074 200488 123130 200544
rect 122982 199536 123038 199592
rect 123166 199944 123222 200000
rect 123166 199808 123222 199864
rect 123074 199128 123130 199184
rect 122982 198720 123038 198776
rect 123166 198720 123222 198776
rect 123166 198448 123222 198504
rect 123074 197768 123130 197824
rect 123074 197496 123130 197552
rect 122982 197360 123038 197416
rect 123258 197904 123314 197960
rect 123166 196408 123222 196464
rect 123074 196136 123130 196192
rect 122982 195048 123038 195104
rect 123258 196272 123314 196328
rect 123166 195728 123222 195784
rect 123166 195592 123222 195648
rect 123074 194504 123130 194560
rect 124178 194912 124234 194968
rect 123258 193824 123314 193880
rect 123166 193688 123222 193744
rect 123074 193280 123130 193336
rect 122982 193008 123038 193064
rect 88574 191920 88630 191976
rect 88482 191648 88538 191704
rect 88390 190424 88446 190480
rect 88390 190288 88446 190344
rect 88298 189200 88354 189256
rect 88482 189880 88538 189936
rect 122154 191648 122210 191704
rect 123166 192736 123222 192792
rect 123074 191512 123130 191568
rect 122982 190968 123038 191024
rect 88666 190832 88722 190888
rect 122982 189336 123038 189392
rect 88758 189200 88814 189256
rect 88482 188656 88538 188712
rect 88666 188656 88722 188712
rect 88390 188112 88446 188168
rect 88206 187432 88262 187488
rect 88390 187432 88446 187488
rect 87194 186208 87250 186264
rect 88482 187296 88538 187352
rect 123350 192192 123406 192248
rect 123258 192056 123314 192112
rect 123258 191920 123314 191976
rect 123166 190832 123222 190888
rect 123166 190424 123222 190480
rect 123074 189064 123130 189120
rect 121970 188812 122026 188848
rect 121970 188792 121972 188812
rect 121972 188792 122024 188812
rect 122024 188792 122026 188812
rect 88850 188112 88906 188168
rect 122982 188112 123038 188168
rect 88574 186908 88630 186944
rect 88574 186888 88576 186908
rect 88576 186888 88628 186908
rect 88628 186888 88630 186908
rect 123258 190288 123314 190344
rect 123258 189880 123314 189936
rect 123166 188112 123222 188168
rect 123350 189472 123406 189528
rect 123258 187976 123314 188032
rect 123074 187296 123130 187352
rect 122430 187024 122486 187080
rect 88574 186344 88630 186400
rect 88574 185800 88630 185856
rect 88482 185664 88538 185720
rect 88666 185256 88722 185312
rect 88390 185120 88446 185176
rect 88574 184168 88630 184224
rect 89218 184712 89274 184768
rect 122338 184712 122394 184768
rect 87838 183624 87894 183680
rect 88574 183080 88630 183136
rect 122154 183080 122210 183136
rect 45058 171792 45114 171848
rect 22242 163768 22298 163824
rect 48462 169208 48518 169264
rect 47818 155880 47874 155936
rect 22334 155744 22390 155800
rect 22334 147720 22390 147776
rect 45794 147720 45850 147776
rect 45794 142552 45850 142608
rect 44414 139832 44470 139888
rect 92162 172744 92218 172800
rect 122890 186480 122946 186536
rect 123534 187568 123590 187624
rect 123350 186752 123406 186808
rect 123074 186072 123130 186128
rect 122982 185936 123038 185992
rect 122890 185256 122946 185312
rect 123534 185120 123590 185176
rect 122982 184168 123038 184224
rect 123074 183624 123130 183680
rect 160334 209872 160390 209928
rect 160242 208376 160298 208432
rect 160426 209328 160482 209384
rect 160242 207832 160298 207888
rect 191706 208920 191762 208976
rect 160518 208784 160574 208840
rect 160150 207560 160206 207616
rect 159046 207188 159048 207208
rect 159048 207188 159100 207208
rect 159100 207188 159102 207208
rect 159046 207152 159102 207188
rect 159046 206608 159102 206664
rect 160610 207832 160666 207888
rect 160426 207016 160482 207072
rect 160334 206472 160390 206528
rect 160150 206064 160206 206120
rect 160518 205928 160574 205984
rect 160242 205384 160298 205440
rect 160334 205248 160390 205304
rect 160150 204840 160206 204896
rect 160518 204840 160574 204896
rect 160426 204704 160482 204760
rect 160334 203888 160390 203944
rect 160242 203616 160298 203672
rect 160242 202392 160298 202448
rect 160518 203616 160574 203672
rect 160426 203480 160482 203536
rect 160610 203072 160666 203128
rect 160426 202392 160482 202448
rect 159046 201848 159102 201904
rect 160518 201848 160574 201904
rect 158954 201168 159010 201224
rect 160150 200760 160206 200816
rect 160334 201304 160390 201360
rect 160242 200624 160298 200680
rect 160242 199400 160298 199456
rect 160518 200624 160574 200680
rect 160518 200216 160574 200272
rect 160242 199264 160298 199320
rect 160150 198856 160206 198912
rect 160058 198448 160114 198504
rect 158954 198176 159010 198232
rect 160426 198992 160482 199048
rect 160242 197904 160298 197960
rect 160150 197632 160206 197688
rect 160058 196408 160114 196464
rect 160242 197088 160298 197144
rect 160518 197360 160574 197416
rect 160242 196680 160298 196736
rect 160150 195864 160206 195920
rect 160150 195592 160206 195648
rect 158954 195184 159010 195240
rect 159966 194504 160022 194560
rect 160058 193824 160114 193880
rect 159966 192192 160022 192248
rect 160334 196136 160390 196192
rect 160242 194640 160298 194696
rect 160242 194096 160298 194152
rect 160426 195048 160482 195104
rect 160150 193416 160206 193472
rect 160518 193280 160574 193336
rect 160242 192872 160298 192928
rect 160150 192736 160206 192792
rect 160058 192056 160114 192112
rect 160058 191648 160114 191704
rect 158954 189880 159010 189936
rect 159966 189608 160022 189664
rect 160242 191104 160298 191160
rect 160610 192192 160666 192248
rect 160242 190968 160298 191024
rect 160150 190832 160206 190888
rect 160150 190424 160206 190480
rect 160058 189200 160114 189256
rect 160058 188792 160114 188848
rect 159966 187432 160022 187488
rect 160334 189336 160390 189392
rect 160242 188656 160298 188712
rect 160150 188112 160206 188168
rect 160150 187568 160206 187624
rect 160058 186208 160114 186264
rect 154354 184984 154410 185040
rect 148834 177232 148890 177288
rect 160242 186888 160298 186944
rect 160426 188112 160482 188168
rect 160978 187024 161034 187080
rect 160518 186480 160574 186536
rect 160242 185664 160298 185720
rect 160610 185936 160666 185992
rect 160334 185256 160390 185312
rect 160150 185120 160206 185176
rect 159598 183624 159654 183680
rect 160334 183080 160390 183136
rect 196950 208920 197006 208976
rect 194742 191104 194798 191160
rect 192074 185528 192130 185584
rect 161254 184712 161310 184768
rect 161070 184168 161126 184224
rect 92622 175192 92678 175248
rect 163186 175192 163242 175248
rect 94554 174512 94610 174568
rect 92346 173968 92402 174024
rect 92254 171520 92310 171576
rect 92070 170296 92126 170352
rect 91978 169072 92034 169128
rect 91426 167848 91482 167904
rect 91334 166624 91390 166680
rect 91978 165400 92034 165456
rect 95014 172200 95070 172256
rect 94830 169888 94886 169944
rect 163186 169108 163188 169128
rect 163188 169108 163240 169128
rect 163240 169108 163242 169128
rect 163186 169072 163242 169108
rect 118934 168956 118990 168992
rect 118934 168936 118936 168956
rect 118936 168936 118988 168956
rect 118988 168936 118990 168956
rect 95382 167440 95438 167496
rect 94186 165128 94242 165184
rect 92622 164176 92678 164232
rect 91702 163088 91758 163144
rect 94094 162816 94150 162872
rect 92622 161900 92624 161920
rect 92624 161900 92676 161920
rect 92676 161900 92678 161920
rect 92622 161864 92678 161900
rect 91978 160640 92034 160696
rect 94002 160368 94058 160424
rect 91978 159416 92034 159472
rect 91978 158192 92034 158248
rect 94002 158056 94058 158112
rect 91794 156968 91850 157024
rect 91426 154520 91482 154576
rect 94738 153432 94794 153488
rect 91794 153296 91850 153352
rect 91702 152072 91758 152128
rect 91426 150848 91482 150904
rect 91334 149760 91390 149816
rect 91702 148536 91758 148592
rect 91426 147312 91482 147368
rect 93358 146088 93414 146144
rect 91978 144864 92034 144920
rect 91794 143640 91850 143696
rect 91794 142416 91850 142472
rect 91702 141736 91758 141792
rect 51222 128136 51278 128192
rect 51406 127592 51462 127648
rect 51314 127048 51370 127104
rect 51222 126912 51278 126968
rect 51222 126096 51278 126152
rect 51498 126368 51554 126424
rect 51406 125824 51462 125880
rect 51314 125688 51370 125744
rect 51222 125144 51278 125200
rect 51406 124736 51462 124792
rect 51314 124464 51370 124520
rect 51222 124056 51278 124112
rect 51314 123920 51370 123976
rect 18102 123512 18158 123568
rect 18010 114128 18066 114184
rect 51498 124600 51554 124656
rect 51498 123512 51554 123568
rect 51406 123240 51462 123296
rect 51314 122832 51370 122888
rect 51406 122696 51462 122752
rect 51406 122016 51462 122072
rect 51314 121472 51370 121528
rect 51222 120656 51278 120712
rect 51222 119976 51278 120032
rect 51130 119316 51186 119352
rect 51130 119296 51132 119316
rect 51132 119296 51184 119316
rect 51184 119296 51186 119316
rect 51774 122288 51830 122344
rect 51498 121608 51554 121664
rect 51498 121064 51554 121120
rect 51406 120248 51462 120304
rect 51406 119432 51462 119488
rect 51314 119024 51370 119080
rect 51314 118480 51370 118536
rect 51222 118208 51278 118264
rect 51774 120384 51830 120440
rect 51498 119160 51554 119216
rect 51498 117936 51554 117992
rect 51406 117800 51462 117856
rect 50578 116984 50634 117040
rect 51222 116440 51278 116496
rect 51222 115896 51278 115952
rect 51406 116168 51462 116224
rect 51590 117256 51646 117312
rect 51498 116032 51554 116088
rect 51590 115488 51646 115544
rect 51406 115352 51462 115408
rect 51314 114944 51370 115000
rect 51314 114264 51370 114320
rect 51314 114128 51370 114184
rect 51222 112904 51278 112960
rect 51498 115080 51554 115136
rect 51406 113584 51462 113640
rect 51590 113720 51646 113776
rect 51498 113040 51554 113096
rect 51498 112496 51554 112552
rect 51314 112224 51370 112280
rect 51222 111816 51278 111872
rect 51222 111156 51278 111192
rect 51222 111136 51224 111156
rect 51224 111136 51276 111156
rect 51276 111136 51278 111156
rect 51222 111000 51278 111056
rect 51314 110864 51370 110920
rect 51590 111952 51646 112008
rect 51498 110728 51554 110784
rect 51406 110048 51462 110104
rect 51590 110048 51646 110104
rect 51314 108960 51370 109016
rect 51222 108824 51278 108880
rect 51222 108280 51278 108336
rect 51222 107056 51278 107112
rect 51498 109640 51554 109696
rect 51406 108144 51462 108200
rect 51406 107872 51462 107928
rect 51314 106512 51370 106568
rect 51222 105968 51278 106024
rect 51682 109504 51738 109560
rect 51498 107736 51554 107792
rect 51498 106784 51554 106840
rect 51406 105968 51462 106024
rect 51406 105424 51462 105480
rect 51314 105288 51370 105344
rect 50670 104744 50726 104800
rect 50486 101072 50542 101128
rect 20494 97808 20550 97864
rect 50946 104200 51002 104256
rect 50762 103112 50818 103168
rect 51314 103928 51370 103984
rect 51222 103656 51278 103712
rect 51590 106648 51646 106704
rect 51498 104744 51554 104800
rect 51406 103520 51462 103576
rect 51406 102704 51462 102760
rect 51222 101888 51278 101944
rect 51314 101344 51370 101400
rect 82134 133032 82190 133088
rect 83606 133032 83662 133088
rect 92530 141192 92586 141248
rect 92622 139988 92678 140024
rect 92622 139968 92624 139988
rect 92624 139968 92676 139988
rect 92676 139968 92678 139988
rect 93266 138744 93322 138800
rect 92070 137520 92126 137576
rect 92162 136432 92218 136488
rect 93358 136976 93414 137032
rect 95382 150984 95438 151040
rect 94186 148672 94242 148728
rect 94002 145544 94058 145600
rect 94370 143912 94426 143968
rect 95382 141600 95438 141656
rect 93542 138608 93598 138664
rect 164382 174004 164384 174024
rect 164384 174004 164436 174024
rect 164436 174004 164438 174024
rect 164382 173968 164438 174004
rect 164290 172780 164292 172800
rect 164292 172780 164344 172800
rect 164344 172780 164346 172800
rect 164290 172744 164346 172780
rect 164014 171556 164016 171576
rect 164016 171556 164068 171576
rect 164068 171556 164070 171576
rect 164014 171520 164070 171556
rect 163370 170332 163372 170352
rect 163372 170332 163424 170352
rect 163424 170332 163426 170352
rect 163370 170296 163426 170332
rect 168522 174784 168578 174840
rect 188026 172472 188082 172528
rect 167510 170432 167566 170488
rect 167326 168120 167382 168176
rect 164382 167848 164438 167904
rect 163278 166624 163334 166680
rect 167234 166216 167290 166272
rect 163186 165400 163242 165456
rect 116542 165128 116598 165184
rect 164290 164176 164346 164232
rect 188026 165808 188082 165864
rect 167970 164040 168026 164096
rect 164290 163124 164292 163144
rect 164292 163124 164344 163144
rect 164344 163124 164346 163144
rect 164290 163088 164346 163124
rect 164290 161900 164292 161920
rect 164292 161900 164344 161920
rect 164344 161900 164346 161920
rect 164290 161864 164346 161900
rect 164382 160640 164438 160696
rect 168430 162156 168486 162192
rect 168430 162136 168432 162156
rect 168432 162136 168484 162156
rect 168484 162136 168486 162156
rect 168522 160776 168578 160832
rect 164290 159416 164346 159472
rect 168522 158464 168578 158520
rect 164290 158228 164292 158248
rect 164292 158228 164344 158248
rect 164344 158228 164346 158248
rect 164290 158192 164346 158228
rect 164290 156988 164346 157024
rect 164290 156968 164292 156988
rect 164292 156968 164344 156988
rect 164344 156968 164346 156988
rect 168522 156832 168578 156888
rect 119578 155880 119634 155936
rect 164382 155744 164438 155800
rect 167142 154792 167198 154848
rect 163370 154540 163426 154576
rect 163370 154520 163372 154540
rect 163372 154520 163424 154540
rect 163424 154520 163426 154540
rect 164382 153296 164438 153352
rect 167142 152752 167198 152808
rect 164382 152072 164438 152128
rect 163922 150848 163978 150904
rect 167234 150712 167290 150768
rect 164382 149780 164438 149816
rect 164382 149760 164384 149780
rect 164384 149760 164436 149780
rect 164436 149760 164438 149780
rect 164382 148556 164438 148592
rect 164382 148536 164384 148556
rect 164384 148536 164436 148556
rect 164436 148536 164438 148556
rect 164382 147312 164438 147368
rect 164382 146088 164438 146144
rect 116818 145544 116874 145600
rect 163738 144864 163794 144920
rect 116818 142588 116820 142608
rect 116820 142588 116872 142608
rect 116872 142588 116874 142608
rect 116818 142552 116874 142588
rect 118934 142588 118936 142608
rect 118936 142588 118988 142608
rect 118988 142588 118990 142608
rect 118934 142552 118990 142588
rect 163094 136432 163150 136488
rect 88574 128408 88630 128464
rect 88390 127864 88446 127920
rect 88298 126640 88354 126696
rect 88482 126368 88538 126424
rect 123074 128136 123130 128192
rect 88666 127320 88722 127376
rect 88482 126096 88538 126152
rect 88390 125824 88446 125880
rect 88298 124600 88354 124656
rect 121694 127184 121750 127240
rect 123166 127728 123222 127784
rect 123074 127048 123130 127104
rect 121786 126504 121842 126560
rect 121694 126132 121696 126152
rect 121696 126132 121748 126152
rect 121748 126132 121750 126152
rect 121694 126096 121750 126132
rect 123166 125824 123222 125880
rect 88758 125552 88814 125608
rect 88482 125144 88538 125200
rect 88482 124872 88538 124928
rect 88390 124056 88446 124112
rect 88390 123784 88446 123840
rect 87746 123376 87802 123432
rect 88206 122560 88262 122616
rect 88298 122016 88354 122072
rect 88206 120384 88262 120440
rect 121694 125416 121750 125472
rect 123166 124872 123222 124928
rect 88666 124328 88722 124384
rect 88574 123240 88630 123296
rect 88482 122832 88538 122888
rect 88390 121608 88446 121664
rect 88390 121472 88446 121528
rect 88298 119840 88354 119896
rect 88298 119704 88354 119760
rect 88206 119296 88262 119352
rect 88114 117936 88170 117992
rect 88482 121064 88538 121120
rect 122982 124056 123038 124112
rect 121694 123648 121750 123704
rect 122982 122832 123038 122888
rect 121694 122424 121750 122480
rect 88666 122152 88722 122208
rect 121694 122036 121750 122072
rect 121694 122016 121696 122036
rect 121696 122016 121748 122036
rect 121748 122016 121750 122036
rect 123994 125688 124050 125744
rect 124362 124600 124418 124656
rect 123902 124464 123958 124520
rect 123718 123920 123774 123976
rect 123166 123240 123222 123296
rect 123074 122696 123130 122752
rect 123074 121472 123130 121528
rect 121694 121200 121750 121256
rect 88482 120792 88538 120848
rect 88390 119160 88446 119216
rect 122982 120656 123038 120712
rect 88574 120248 88630 120304
rect 88482 118616 88538 118672
rect 88390 118480 88446 118536
rect 88298 117392 88354 117448
rect 88206 116848 88262 116904
rect 88482 118072 88538 118128
rect 122982 119976 123038 120032
rect 121694 119568 121750 119624
rect 123534 121608 123590 121664
rect 123442 120384 123498 120440
rect 123350 120248 123406 120304
rect 123258 119296 123314 119352
rect 123166 119024 123222 119080
rect 123074 118480 123130 118536
rect 121694 118344 121750 118400
rect 123166 117936 123222 117992
rect 88666 117392 88722 117448
rect 88482 116712 88538 116768
rect 88390 116168 88446 116224
rect 88114 115624 88170 115680
rect 88390 115624 88446 115680
rect 88206 115216 88262 115272
rect 88114 113856 88170 113912
rect 88022 113312 88078 113368
rect 88298 114400 88354 114456
rect 88206 112632 88262 112688
rect 88574 116168 88630 116224
rect 88482 114944 88538 115000
rect 88482 114264 88538 114320
rect 122982 116984 123038 117040
rect 123074 116440 123130 116496
rect 121694 115896 121750 115952
rect 121694 115488 121750 115544
rect 88666 115080 88722 115136
rect 121694 115116 121696 115136
rect 121696 115116 121748 115136
rect 121748 115116 121750 115136
rect 121694 115080 121750 115116
rect 124362 119160 124418 119216
rect 124270 117800 124326 117856
rect 123258 117256 123314 117312
rect 123166 116032 123222 116088
rect 124362 116168 124418 116224
rect 124270 115488 124326 115544
rect 123074 114944 123130 115000
rect 121694 114264 121750 114320
rect 122982 113720 123038 113776
rect 88390 113176 88446 113232
rect 88482 112632 88538 112688
rect 88298 112088 88354 112144
rect 88298 111544 88354 111600
rect 88114 111408 88170 111464
rect 88022 110864 88078 110920
rect 88206 109776 88262 109832
rect 88114 109232 88170 109288
rect 88022 107464 88078 107520
rect 85170 106820 85172 106840
rect 85172 106820 85224 106840
rect 85224 106820 85226 106840
rect 85170 106784 85226 106820
rect 88390 111000 88446 111056
rect 88298 109096 88354 109152
rect 88298 108552 88354 108608
rect 88206 107192 88262 107248
rect 88114 106648 88170 106704
rect 121694 112496 121750 112552
rect 88666 112088 88722 112144
rect 88574 110320 88630 110376
rect 88482 110184 88538 110240
rect 123258 112904 123314 112960
rect 122982 111816 123038 111872
rect 121694 111272 121750 111328
rect 123166 111816 123222 111872
rect 123166 111000 123222 111056
rect 123258 110864 123314 110920
rect 123994 113584 124050 113640
rect 124362 114264 124418 114320
rect 124270 113040 124326 113096
rect 123442 112088 123498 112144
rect 121694 110048 121750 110104
rect 123074 110048 123130 110104
rect 88390 108416 88446 108472
rect 88666 109640 88722 109696
rect 122982 109640 123038 109696
rect 121694 108960 121750 109016
rect 88574 108008 88630 108064
rect 88482 107872 88538 107928
rect 88482 106784 88538 106840
rect 88390 106240 88446 106296
rect 88298 106104 88354 106160
rect 88298 105696 88354 105752
rect 88022 104880 88078 104936
rect 55546 100936 55602 100992
rect 56742 100936 56798 100992
rect 123350 110728 123406 110784
rect 124270 109504 124326 109560
rect 123258 108960 123314 109016
rect 123258 108416 123314 108472
rect 122982 107736 123038 107792
rect 123166 107736 123222 107792
rect 121694 107192 121750 107248
rect 123074 106784 123130 106840
rect 121694 106104 121750 106160
rect 121694 105696 121750 105752
rect 88574 105424 88630 105480
rect 88666 105152 88722 105208
rect 88574 104472 88630 104528
rect 88482 104200 88538 104256
rect 124362 108144 124418 108200
rect 123442 106648 123498 106704
rect 123258 106512 123314 106568
rect 123166 105968 123222 106024
rect 121786 104744 121842 104800
rect 123074 104744 123130 104800
rect 88482 103928 88538 103984
rect 88390 103656 88446 103712
rect 88298 103112 88354 103168
rect 88482 103384 88538 103440
rect 89678 102704 89734 102760
rect 88666 102160 88722 102216
rect 88574 101616 88630 101672
rect 88574 100528 88630 100584
rect 121694 104336 121750 104392
rect 121878 103656 121934 103712
rect 121786 103248 121842 103304
rect 121694 102860 121750 102896
rect 121694 102840 121696 102860
rect 121696 102840 121748 102860
rect 121748 102840 121750 102860
rect 124270 105288 124326 105344
rect 124362 103928 124418 103984
rect 124178 103520 124234 103576
rect 123074 101888 123130 101944
rect 22334 89784 22390 89840
rect 45058 89784 45114 89840
rect 22334 81760 22390 81816
rect 91702 93184 91758 93240
rect 91518 90736 91574 90792
rect 91426 85840 91482 85896
rect 91334 84616 91390 84672
rect 92254 91960 92310 92016
rect 92162 89512 92218 89568
rect 91794 83392 91850 83448
rect 92438 88288 92494 88344
rect 116358 100664 116414 100720
rect 122154 100528 122210 100584
rect 123258 101344 123314 101400
rect 163830 143640 163886 143696
rect 167326 148808 167382 148864
rect 167234 146768 167290 146824
rect 167142 144728 167198 144784
rect 167050 142824 167106 142880
rect 164382 142416 164438 142472
rect 164290 141192 164346 141248
rect 164382 139988 164438 140024
rect 164382 139968 164384 139988
rect 164384 139968 164436 139988
rect 164436 139968 164438 139988
rect 163922 138744 163978 138800
rect 164750 137520 164806 137576
rect 167878 140784 167934 140840
rect 188026 139188 188028 139208
rect 188028 139188 188080 139208
rect 188080 139188 188082 139208
rect 188026 139152 188082 139188
rect 167970 138744 168026 138800
rect 168522 136160 168578 136216
rect 160334 128136 160390 128192
rect 160150 127592 160206 127648
rect 160058 126504 160114 126560
rect 160242 126368 160298 126424
rect 160426 126912 160482 126968
rect 160242 126096 160298 126152
rect 160150 125824 160206 125880
rect 160058 124600 160114 124656
rect 160242 125144 160298 125200
rect 160518 125144 160574 125200
rect 160242 124872 160298 124928
rect 160150 124056 160206 124112
rect 160058 123512 160114 123568
rect 160242 123376 160298 123432
rect 160426 124056 160482 124112
rect 160150 122832 160206 122888
rect 160426 122832 160482 122888
rect 160242 122696 160298 122752
rect 160242 122288 160298 122344
rect 160150 122016 160206 122072
rect 160058 121608 160114 121664
rect 159966 121200 160022 121256
rect 159874 119296 159930 119352
rect 160242 121064 160298 121120
rect 160242 120656 160298 120712
rect 160150 120384 160206 120440
rect 160058 119840 160114 119896
rect 160150 119432 160206 119488
rect 159966 119160 160022 119216
rect 160058 118208 160114 118264
rect 159874 116848 159930 116904
rect 160334 119976 160390 120032
rect 160242 118616 160298 118672
rect 160242 118072 160298 118128
rect 160242 117936 160298 117992
rect 160150 117392 160206 117448
rect 160426 116984 160482 117040
rect 160058 116168 160114 116224
rect 160242 116440 160298 116496
rect 160150 115624 160206 115680
rect 160058 115352 160114 115408
rect 160334 115896 160390 115952
rect 160242 114400 160298 114456
rect 160242 114264 160298 114320
rect 160426 115080 160482 115136
rect 160610 115116 160612 115136
rect 160612 115116 160664 115136
rect 160664 115116 160666 115136
rect 160610 115080 160666 115116
rect 160242 114128 160298 114184
rect 160150 113720 160206 113776
rect 160058 113176 160114 113232
rect 159966 112904 160022 112960
rect 159046 112632 159102 112688
rect 159874 111000 159930 111056
rect 160058 112360 160114 112416
rect 159966 110864 160022 110920
rect 160242 112088 160298 112144
rect 160334 111816 160390 111872
rect 160150 111408 160206 111464
rect 160242 111136 160298 111192
rect 160058 110184 160114 110240
rect 160150 110048 160206 110104
rect 159966 109776 160022 109832
rect 159874 108416 159930 108472
rect 160058 108824 160114 108880
rect 159966 107192 160022 107248
rect 159874 106784 159930 106840
rect 160334 109640 160390 109696
rect 160242 109096 160298 109152
rect 160242 108280 160298 108336
rect 160150 107872 160206 107928
rect 160150 107056 160206 107112
rect 160058 106648 160114 106704
rect 160058 105968 160114 106024
rect 159966 105560 160022 105616
rect 159874 104200 159930 104256
rect 160334 107736 160390 107792
rect 160242 106104 160298 106160
rect 160242 105424 160298 105480
rect 193546 123512 193602 123568
rect 193454 106104 193510 106160
rect 160150 104880 160206 104936
rect 161530 104744 161586 104800
rect 160334 104200 160390 104256
rect 160058 103928 160114 103984
rect 160150 103656 160206 103712
rect 159966 103112 160022 103168
rect 160242 102976 160298 103032
rect 160518 102704 160574 102760
rect 160334 101888 160390 101944
rect 160426 101480 160482 101536
rect 160334 100528 160390 100584
rect 95290 92504 95346 92560
rect 95382 90192 95438 90248
rect 95382 87880 95438 87936
rect 118934 87200 118990 87256
rect 92806 87064 92862 87120
rect 94278 85432 94334 85488
rect 92254 82168 92310 82224
rect 92162 81080 92218 81136
rect 163554 90736 163610 90792
rect 163462 88288 163518 88344
rect 164106 93184 164162 93240
rect 163830 91960 163886 92016
rect 163830 89512 163886 89568
rect 163738 87064 163794 87120
rect 168522 92776 168578 92832
rect 188118 90464 188174 90520
rect 167326 88016 167382 88072
rect 164566 85840 164622 85896
rect 167234 84752 167290 84808
rect 163094 84616 163150 84672
rect 116542 83800 116598 83856
rect 95290 83120 95346 83176
rect 91794 79856 91850 79912
rect 95382 80808 95438 80864
rect 91426 78632 91482 78688
rect 94922 78360 94978 78416
rect 91702 77444 91704 77464
rect 91704 77444 91756 77464
rect 91756 77444 91758 77464
rect 91702 77408 91758 77444
rect 91702 76220 91704 76240
rect 91704 76220 91756 76240
rect 91756 76220 91758 76240
rect 91702 76184 91758 76220
rect 163922 83392 163978 83448
rect 163922 82168 163978 82224
rect 167878 86112 167934 86168
rect 188118 83800 188174 83856
rect 167326 82032 167382 82088
rect 163554 81080 163610 81136
rect 167234 80808 167290 80864
rect 164106 79856 164162 79912
rect 164382 78632 164438 78688
rect 167234 78088 167290 78144
rect 164106 77408 164162 77464
rect 188578 77136 188634 77192
rect 167234 76476 167290 76512
rect 167234 76456 167236 76476
rect 167236 76456 167288 76476
rect 167288 76456 167290 76476
rect 163738 76184 163794 76240
rect 164106 74980 164162 75016
rect 164106 74960 164108 74980
rect 164108 74960 164160 74980
rect 164160 74960 164162 74980
rect 167234 74824 167290 74880
rect 47818 73872 47874 73928
rect 119578 73872 119634 73928
rect 22334 73736 22390 73792
rect 164382 73756 164438 73792
rect 164382 73736 164384 73756
rect 164384 73736 164436 73756
rect 164436 73736 164438 73756
rect 167142 72784 167198 72840
rect 91702 72532 91758 72568
rect 91702 72512 91704 72532
rect 91704 72512 91756 72532
rect 91756 72512 91758 72532
rect 164382 72532 164438 72568
rect 164382 72512 164384 72532
rect 164384 72512 164436 72532
rect 164436 72512 164438 72532
rect 95382 71424 95438 71480
rect 91702 71308 91758 71344
rect 91702 71288 91704 71308
rect 91704 71288 91756 71308
rect 91756 71288 91758 71308
rect 164382 71288 164438 71344
rect 91426 70064 91482 70120
rect 91426 68840 91482 68896
rect 91518 67752 91574 67808
rect 92530 66528 92586 66584
rect 22702 65712 22758 65768
rect 44414 65712 44470 65768
rect 92346 65304 92402 65360
rect 91426 61632 91482 61688
rect 47174 60544 47230 60600
rect 47542 60544 47598 60600
rect 44414 57824 44470 57880
rect 91518 59184 91574 59240
rect 92622 64100 92678 64136
rect 92622 64080 92624 64100
rect 92624 64080 92676 64100
rect 92676 64080 92678 64100
rect 93358 62856 93414 62912
rect 92898 57960 92954 58016
rect 91426 56736 91482 56792
rect 91334 54424 91390 54480
rect 53246 51432 53302 51488
rect 82134 51588 82190 51624
rect 82134 51568 82136 51588
rect 82136 51568 82188 51588
rect 82188 51568 82190 51588
rect 83606 51568 83662 51624
rect 47542 46808 47598 46864
rect 50578 46128 50634 46184
rect 49934 45176 49990 45232
rect 49934 44768 49990 44824
rect 13318 40416 13374 40472
rect 18010 40144 18066 40200
rect 50486 34160 50542 34216
rect 50486 33752 50542 33808
rect 50486 32664 50542 32720
rect 50486 32256 50542 32312
rect 18102 25456 18158 25512
rect 13134 19336 13190 19392
rect 50578 19744 50634 19800
rect 50762 21104 50818 21160
rect 51038 24116 51094 24152
rect 51038 24096 51040 24116
rect 51040 24096 51092 24116
rect 51092 24096 51094 24116
rect 50946 21784 51002 21840
rect 51314 44904 51370 44960
rect 51314 44224 51370 44280
rect 51222 44088 51278 44144
rect 51314 43272 51370 43328
rect 51222 42048 51278 42104
rect 51314 41232 51370 41288
rect 51222 41096 51278 41152
rect 51314 40416 51370 40472
rect 51222 39872 51278 39928
rect 51314 39056 51370 39112
rect 51222 37968 51278 38024
rect 51314 37016 51370 37072
rect 51222 36880 51278 36936
rect 51222 36608 51278 36664
rect 51406 36336 51462 36392
rect 51314 35928 51370 35984
rect 51222 34432 51278 34488
rect 51222 34024 51278 34080
rect 51498 33616 51554 33672
rect 51314 32936 51370 32992
rect 51222 32392 51278 32448
rect 51314 31712 51370 31768
rect 51222 31576 51278 31632
rect 51314 30760 51370 30816
rect 51222 30352 51278 30408
rect 51314 29400 51370 29456
rect 51222 28584 51278 28640
rect 51222 28312 51278 28368
rect 51406 28040 51462 28096
rect 51314 27496 51370 27552
rect 51222 27360 51278 27416
rect 51314 26680 51370 26736
rect 51406 26136 51462 26192
rect 51314 25592 51370 25648
rect 51222 25456 51278 25512
rect 51406 25456 51462 25512
rect 51314 25048 51370 25104
rect 51314 24504 51370 24560
rect 51314 23280 51370 23336
rect 51222 23144 51278 23200
rect 51498 22464 51554 22520
rect 66586 50208 66642 50264
rect 92622 55512 92678 55568
rect 167234 70744 167290 70800
rect 163554 70064 163610 70120
rect 95382 68976 95438 69032
rect 163738 68840 163794 68896
rect 164382 67752 164438 67808
rect 167326 68704 167382 68760
rect 167234 66800 167290 66856
rect 95382 66664 95438 66720
rect 164382 66528 164438 66584
rect 94002 65440 94058 65496
rect 95382 65440 95438 65496
rect 164382 65304 164438 65360
rect 93910 64080 93966 64136
rect 164382 64100 164438 64136
rect 164382 64080 164384 64100
rect 164384 64080 164436 64100
rect 164436 64080 164438 64100
rect 117462 63128 117518 63184
rect 163738 62856 163794 62912
rect 93634 61360 93690 61416
rect 119486 60544 119542 60600
rect 94646 60408 94702 60464
rect 94094 59592 94150 59648
rect 93542 54968 93598 55024
rect 95198 57280 95254 57336
rect 163094 54424 163150 54480
rect 75050 46536 75106 46592
rect 73578 46400 73634 46456
rect 72106 46264 72162 46320
rect 70634 46128 70690 46184
rect 68794 44632 68850 44688
rect 82870 44632 82926 44688
rect 51222 21920 51278 21976
rect 51314 21104 51370 21160
rect 51130 20968 51186 21024
rect 58766 20968 58822 21024
rect 50854 20424 50910 20480
rect 50670 19200 50726 19256
rect 56374 17976 56430 18032
rect 60790 20832 60846 20888
rect 59502 20696 59558 20752
rect 57386 17840 57442 17896
rect 66494 19200 66550 19256
rect 88390 46128 88446 46184
rect 88114 44904 88170 44960
rect 88574 45448 88630 45504
rect 88482 44768 88538 44824
rect 88390 44360 88446 44416
rect 88114 43136 88170 43192
rect 88482 43816 88538 43872
rect 88574 43680 88630 43736
rect 88390 43408 88446 43464
rect 88298 42592 88354 42648
rect 88298 42184 88354 42240
rect 88482 42048 88538 42104
rect 88666 42456 88722 42512
rect 88390 41368 88446 41424
rect 88482 40824 88538 40880
rect 88758 41232 88814 41288
rect 88390 40552 88446 40608
rect 88298 40144 88354 40200
rect 88574 40008 88630 40064
rect 88482 39600 88538 39656
rect 88390 39056 88446 39112
rect 88482 38376 88538 38432
rect 88666 39328 88722 39384
rect 88482 38240 88538 38296
rect 88758 38784 88814 38840
rect 88574 38104 88630 38160
rect 88482 37832 88538 37888
rect 88206 37152 88262 37208
rect 88390 36472 88446 36528
rect 88298 35248 88354 35304
rect 88666 36880 88722 36936
rect 88574 36608 88630 36664
rect 88482 36064 88538 36120
rect 88666 35656 88722 35712
rect 88482 35384 88538 35440
rect 88390 34840 88446 34896
rect 88574 34432 88630 34488
rect 88666 34160 88722 34216
rect 88390 33752 88446 33808
rect 88298 33616 88354 33672
rect 88574 33888 88630 33944
rect 88482 33072 88538 33128
rect 88482 32392 88538 32448
rect 88666 32664 88722 32720
rect 88482 32256 88538 32312
rect 88390 31848 88446 31904
rect 88390 30896 88446 30952
rect 88574 31440 88630 31496
rect 88482 30624 88538 30680
rect 88482 30080 88538 30136
rect 88666 31168 88722 31224
rect 88666 30216 88722 30272
rect 88574 29672 88630 29728
rect 88390 29400 88446 29456
rect 88482 28856 88538 28912
rect 88758 28992 88814 29048
rect 88390 28720 88446 28776
rect 88574 28448 88630 28504
rect 88390 28176 88446 28232
rect 88298 27668 88300 27688
rect 88300 27668 88352 27688
rect 88352 27668 88354 27688
rect 88298 27632 88354 27668
rect 88298 26816 88354 26872
rect 88574 27224 88630 27280
rect 88482 27088 88538 27144
rect 88390 26408 88446 26464
rect 88482 25864 88538 25920
rect 88666 26000 88722 26056
rect 88574 25592 88630 25648
rect 88298 25184 88354 25240
rect 88482 25048 88538 25104
rect 88574 24776 88630 24832
rect 87930 23960 87986 24016
rect 87930 22872 87986 22928
rect 88390 24096 88446 24152
rect 88482 23416 88538 23472
rect 88666 23552 88722 23608
rect 88574 22872 88630 22928
rect 88482 22600 88538 22656
rect 88758 22464 88814 22520
rect 88666 22192 88722 22248
rect 88574 21648 88630 21704
rect 88482 21104 88538 21160
rect 88022 20968 88078 21024
rect 88574 20696 88630 20752
rect 88574 19780 88576 19800
rect 88576 19780 88628 19800
rect 88628 19780 88630 19800
rect 88574 19744 88630 19780
rect 87838 19472 87894 19528
rect 121694 45040 121750 45096
rect 121694 44788 121750 44824
rect 121694 44768 121696 44788
rect 121696 44768 121748 44788
rect 121748 44768 121750 44788
rect 121694 43428 121750 43464
rect 121694 43408 121696 43428
rect 121696 43408 121748 43428
rect 121748 43408 121750 43428
rect 121694 42184 121750 42240
rect 121694 40824 121750 40880
rect 121786 38784 121842 38840
rect 121694 38376 121750 38432
rect 121694 37852 121750 37888
rect 121694 37832 121696 37852
rect 121696 37832 121748 37852
rect 121748 37832 121750 37852
rect 121694 35248 121750 35304
rect 121694 34432 121750 34488
rect 121694 33772 121750 33808
rect 121694 33752 121696 33772
rect 121696 33752 121748 33772
rect 121748 33752 121750 33772
rect 121694 32412 121750 32448
rect 121694 32392 121696 32412
rect 121696 32392 121748 32412
rect 121748 32392 121750 32412
rect 121694 31168 121750 31224
rect 121694 29128 121750 29184
rect 121694 28584 121750 28640
rect 121694 28196 121750 28232
rect 121694 28176 121696 28196
rect 121696 28176 121748 28196
rect 121748 28176 121750 28196
rect 121694 24776 121750 24832
rect 122430 20696 122486 20752
rect 122982 46128 123038 46184
rect 122982 45448 123038 45504
rect 123166 44360 123222 44416
rect 123074 44224 123130 44280
rect 122982 43680 123038 43736
rect 122982 42456 123038 42512
rect 123534 43136 123590 43192
rect 123350 43000 123406 43056
rect 123074 42320 123130 42376
rect 122982 41232 123038 41288
rect 123166 41232 123222 41288
rect 124362 41912 124418 41968
rect 124270 40416 124326 40472
rect 123166 40008 123222 40064
rect 123074 39872 123130 39928
rect 122982 39328 123038 39384
rect 124362 39056 124418 39112
rect 123166 38920 123222 38976
rect 123074 38240 123130 38296
rect 123902 37696 123958 37752
rect 123442 37016 123498 37072
rect 122982 36880 123038 36936
rect 123258 36472 123314 36528
rect 123074 35928 123130 35984
rect 122982 35656 123038 35712
rect 124362 36336 124418 36392
rect 123258 34840 123314 34896
rect 123166 34568 123222 34624
rect 122982 33888 123038 33944
rect 123626 33616 123682 33672
rect 123074 32936 123130 32992
rect 122982 32800 123038 32856
rect 123074 31712 123130 31768
rect 122982 31440 123038 31496
rect 124362 33480 124418 33536
rect 124270 32120 124326 32176
rect 123994 30624 124050 30680
rect 123074 30488 123130 30544
rect 123166 30216 123222 30272
rect 122982 29672 123038 29728
rect 124362 29400 124418 29456
rect 123166 29264 123222 29320
rect 123074 28720 123130 28776
rect 123534 28040 123590 28096
rect 122982 27224 123038 27280
rect 123258 26816 123314 26872
rect 123074 26272 123130 26328
rect 123166 26000 123222 26056
rect 122982 25456 123038 25512
rect 124362 27496 124418 27552
rect 124086 26680 124142 26736
rect 123258 25184 123314 25240
rect 123166 25048 123222 25104
rect 123074 24504 123130 24560
rect 122982 24096 123038 24152
rect 123442 23824 123498 23880
rect 123258 23552 123314 23608
rect 123074 23280 123130 23336
rect 122982 23008 123038 23064
rect 122890 22464 122946 22520
rect 123166 22600 123222 22656
rect 123074 22056 123130 22112
rect 122706 21920 122762 21976
rect 123258 22464 123314 22520
rect 122614 21104 122670 21160
rect 123166 21104 123222 21160
rect 122522 19744 122578 19800
rect 122338 19472 122394 19528
rect 163830 61632 163886 61688
rect 165118 60408 165174 60464
rect 164382 59184 164438 59240
rect 164382 57960 164438 58016
rect 165026 56736 165082 56792
rect 164566 55512 164622 55568
rect 142670 46672 142726 46728
rect 167326 64760 167382 64816
rect 167878 62720 167934 62776
rect 167142 60816 167198 60872
rect 167050 58776 167106 58832
rect 187934 57144 187990 57200
rect 166498 56736 166554 56792
rect 168522 54424 168578 54480
rect 145614 46536 145670 46592
rect 144142 46264 144198 46320
rect 147086 46400 147142 46456
rect 139726 44632 139782 44688
rect 140922 44632 140978 44688
rect 129698 20968 129754 21024
rect 130710 20968 130766 21024
rect 127398 18248 127454 18304
rect 128410 17976 128466 18032
rect 132550 18112 132606 18168
rect 131446 17840 131502 17896
rect 135862 20832 135918 20888
rect 159046 37832 159102 37888
rect 159046 26408 159102 26464
rect 158954 24096 159010 24152
rect 159046 21104 159102 21160
rect 160242 46128 160298 46184
rect 160150 44904 160206 44960
rect 160058 44768 160114 44824
rect 160334 45448 160390 45504
rect 160242 44360 160298 44416
rect 160242 43816 160298 43872
rect 160334 43680 160390 43736
rect 160150 43408 160206 43464
rect 160058 43136 160114 43192
rect 159782 42592 159838 42648
rect 160058 42184 160114 42240
rect 160334 42456 160390 42512
rect 160242 42048 160298 42104
rect 160150 41368 160206 41424
rect 160242 40824 160298 40880
rect 160426 41232 160482 41288
rect 160242 40552 160298 40608
rect 160058 40144 160114 40200
rect 160334 40008 160390 40064
rect 160242 39056 160298 39112
rect 160242 38376 160298 38432
rect 160426 39600 160482 39656
rect 160518 39328 160574 39384
rect 160426 38784 160482 38840
rect 160334 38240 160390 38296
rect 160150 37968 160206 38024
rect 160426 37832 160482 37888
rect 160334 36880 160390 36936
rect 160242 36608 160298 36664
rect 160242 36472 160298 36528
rect 160150 36064 160206 36120
rect 160058 35112 160114 35168
rect 160426 35656 160482 35712
rect 160334 35384 160390 35440
rect 160242 34840 160298 34896
rect 160334 34432 160390 34488
rect 160150 33752 160206 33808
rect 160058 33616 160114 33672
rect 160058 32256 160114 32312
rect 160242 33072 160298 33128
rect 160426 34160 160482 34216
rect 160426 33888 160482 33944
rect 160242 32392 160298 32448
rect 160518 32664 160574 32720
rect 160150 31848 160206 31904
rect 160334 31440 160390 31496
rect 160242 31168 160298 31224
rect 160150 30896 160206 30952
rect 160058 30624 160114 30680
rect 160242 30080 160298 30136
rect 160426 30216 160482 30272
rect 160334 29672 160390 29728
rect 160150 29400 160206 29456
rect 160518 28992 160574 29048
rect 160242 28856 160298 28912
rect 160334 28448 160390 28504
rect 160150 28176 160206 28232
rect 160518 28176 160574 28232
rect 160702 28196 160758 28232
rect 160702 28176 160704 28196
rect 160704 28176 160756 28196
rect 160756 28176 160758 28196
rect 160334 27224 160390 27280
rect 160242 27088 160298 27144
rect 160150 26816 160206 26872
rect 160242 25864 160298 25920
rect 160426 26000 160482 26056
rect 160334 25456 160390 25512
rect 160150 25184 160206 25240
rect 160242 25048 160298 25104
rect 160334 24776 160390 24832
rect 160242 23416 160298 23472
rect 160426 24232 160482 24288
rect 160242 22872 160298 22928
rect 160518 23552 160574 23608
rect 160610 22872 160666 22928
rect 160518 22600 160574 22656
rect 160426 22464 160482 22520
rect 160518 21920 160574 21976
rect 160702 22636 160704 22656
rect 160704 22636 160756 22656
rect 160756 22636 160758 22656
rect 160702 22600 160758 22636
rect 160242 21648 160298 21704
rect 160334 21104 160390 21160
rect 159690 20696 159746 20752
rect 198238 185392 198294 185448
rect 197594 161864 197650 161920
rect 196950 138336 197006 138392
rect 201274 114672 201330 114728
rect 201274 114536 201330 114592
rect 197594 91144 197650 91200
rect 197594 67616 197650 67672
rect 201274 44088 201330 44144
rect 201274 43816 201330 43872
rect 196858 20560 196914 20616
rect 159598 19744 159654 19800
rect 160334 19472 160390 19528
rect 177814 17024 177870 17080
<< metal3 >>
rect 23566 213132 23572 213196
rect 23636 213194 23642 213196
rect 33369 213194 33435 213197
rect 23636 213192 33435 213194
rect 23636 213136 33374 213192
rect 33430 213136 33435 213192
rect 23636 213134 33435 213136
rect 23636 213132 23642 213134
rect 33369 213131 33435 213134
rect 39441 213194 39507 213197
rect 187142 213194 187148 213196
rect 39441 213192 187148 213194
rect 39441 213136 39446 213192
rect 39502 213136 187148 213192
rect 39441 213134 187148 213136
rect 39441 213131 39507 213134
rect 187142 213132 187148 213134
rect 187212 213132 187218 213196
rect 138801 210746 138867 210749
rect 190638 210746 190644 210748
rect 138801 210744 190644 210746
rect 138801 210688 138806 210744
rect 138862 210688 190644 210744
rect 138801 210686 190644 210688
rect 138801 210683 138867 210686
rect 190638 210684 190644 210686
rect 190708 210684 190714 210748
rect 49285 210474 49351 210477
rect 120861 210474 120927 210477
rect 47524 210472 49351 210474
rect 47524 210416 49290 210472
rect 49346 210416 49351 210472
rect 47524 210414 49351 210416
rect 119836 210472 120927 210474
rect 119836 210416 120866 210472
rect 120922 210416 120927 210472
rect 119836 210414 120927 210416
rect 49285 210411 49351 210414
rect 120861 210411 120927 210414
rect 160329 210474 160395 210477
rect 160329 210472 163996 210474
rect 160329 210416 160334 210472
rect 160390 210416 163996 210472
rect 160329 210414 163996 210416
rect 160329 210411 160395 210414
rect 73205 210338 73271 210341
rect 81710 210338 81716 210340
rect 73205 210336 81716 210338
rect 73205 210280 73210 210336
rect 73266 210280 81716 210336
rect 73205 210278 81716 210280
rect 73205 210275 73271 210278
rect 81710 210276 81716 210278
rect 81780 210276 81786 210340
rect 145609 210338 145675 210341
rect 153470 210338 153476 210340
rect 145609 210336 153476 210338
rect 145609 210280 145614 210336
rect 145670 210280 153476 210336
rect 145609 210278 153476 210280
rect 145609 210275 145675 210278
rect 153470 210276 153476 210278
rect 153540 210276 153546 210340
rect 9896 210202 10376 210232
rect 13313 210202 13379 210205
rect 9896 210200 13379 210202
rect 9896 210144 13318 210200
rect 13374 210144 13379 210200
rect 9896 210142 13379 210144
rect 9896 210112 10376 210142
rect 13313 210139 13379 210142
rect 49929 209930 49995 209933
rect 47524 209928 49995 209930
rect 47524 209872 49934 209928
rect 49990 209872 49995 209928
rect 47524 209870 49995 209872
rect 49929 209867 49995 209870
rect 88569 209930 88635 209933
rect 122977 209930 123043 209933
rect 88569 209928 92052 209930
rect 88569 209872 88574 209928
rect 88630 209872 92052 209928
rect 88569 209870 92052 209872
rect 119836 209928 123043 209930
rect 119836 209872 122982 209928
rect 123038 209872 123043 209928
rect 119836 209870 123043 209872
rect 88569 209867 88635 209870
rect 122977 209867 123043 209870
rect 160329 209930 160395 209933
rect 160329 209928 163996 209930
rect 160329 209872 160334 209928
rect 160390 209872 163996 209928
rect 160329 209870 163996 209872
rect 160329 209867 160395 209870
rect 51309 209386 51375 209389
rect 122977 209386 123043 209389
rect 47524 209384 51375 209386
rect 47524 209328 51314 209384
rect 51370 209328 51375 209384
rect 47524 209326 51375 209328
rect 51309 209323 51375 209326
rect 88526 209326 92052 209386
rect 119836 209384 123043 209386
rect 119836 209328 122982 209384
rect 123038 209328 123043 209384
rect 119836 209326 123043 209328
rect 49929 208978 49995 208981
rect 49929 208976 51418 208978
rect 49929 208920 49934 208976
rect 49990 208920 51418 208976
rect 49929 208918 51418 208920
rect 49929 208915 49995 208918
rect 51358 208842 51418 208918
rect 88526 208842 88586 209326
rect 122977 209323 123043 209326
rect 160421 209386 160487 209389
rect 160421 209384 163996 209386
rect 160421 209328 160426 209384
rect 160482 209328 163996 209384
rect 160421 209326 163996 209328
rect 160421 209323 160487 209326
rect 191701 208978 191767 208981
rect 196945 208978 197011 208981
rect 201416 208978 201896 209008
rect 191701 208976 191810 208978
rect 191701 208920 191706 208976
rect 191762 208920 191810 208976
rect 191701 208915 191810 208920
rect 196945 208976 201896 208978
rect 196945 208920 196950 208976
rect 197006 208920 201896 208976
rect 196945 208918 201896 208920
rect 196945 208915 197011 208918
rect 47494 208434 47554 208812
rect 51358 208782 55098 208842
rect 55038 208472 55098 208782
rect 84846 208782 88586 208842
rect 88661 208842 88727 208845
rect 123069 208842 123135 208845
rect 160513 208842 160579 208845
rect 88661 208840 92052 208842
rect 88661 208784 88666 208840
rect 88722 208784 92052 208840
rect 123069 208840 127042 208842
rect 88661 208782 92052 208784
rect 51493 208434 51559 208437
rect 47494 208432 51559 208434
rect 47494 208376 51498 208432
rect 51554 208376 51559 208432
rect 84846 208404 84906 208782
rect 88661 208779 88727 208782
rect 119806 208434 119866 208812
rect 123069 208784 123074 208840
rect 123130 208784 127042 208840
rect 123069 208782 127042 208784
rect 123069 208779 123135 208782
rect 126982 208472 127042 208782
rect 160513 208840 163996 208842
rect 160513 208784 160518 208840
rect 160574 208784 163996 208840
rect 160513 208782 163996 208784
rect 160513 208779 160579 208782
rect 123253 208434 123319 208437
rect 160237 208434 160303 208437
rect 119806 208432 123319 208434
rect 47494 208374 51559 208376
rect 119806 208376 123258 208432
rect 123314 208376 123319 208432
rect 119806 208374 123319 208376
rect 156820 208432 160303 208434
rect 156820 208376 160242 208432
rect 160298 208376 160303 208432
rect 156820 208374 160303 208376
rect 51493 208371 51559 208374
rect 123253 208371 123319 208374
rect 160237 208371 160303 208374
rect 51309 208298 51375 208301
rect 88569 208298 88635 208301
rect 123069 208298 123135 208301
rect 51309 208296 55098 208298
rect 51309 208240 51314 208296
rect 51370 208240 55098 208296
rect 51309 208238 55098 208240
rect 51309 208235 51375 208238
rect 51309 208162 51375 208165
rect 47524 208160 51375 208162
rect 47524 208104 51314 208160
rect 51370 208104 51375 208160
rect 47524 208102 51375 208104
rect 51309 208099 51375 208102
rect 55038 207928 55098 208238
rect 88569 208296 92052 208298
rect 88569 208240 88574 208296
rect 88630 208240 92052 208296
rect 88569 208238 92052 208240
rect 123069 208296 127042 208298
rect 123069 208240 123074 208296
rect 123130 208240 127042 208296
rect 123069 208238 127042 208240
rect 88569 208235 88635 208238
rect 123069 208235 123135 208238
rect 122977 208162 123043 208165
rect 119836 208160 123043 208162
rect 119836 208104 122982 208160
rect 123038 208104 123043 208160
rect 119836 208102 123043 208104
rect 122977 208099 123043 208102
rect 126982 207928 127042 208238
rect 88661 207890 88727 207893
rect 160237 207890 160303 207893
rect 84876 207888 88727 207890
rect 84876 207832 88666 207888
rect 88722 207832 88727 207888
rect 84876 207830 88727 207832
rect 156820 207888 160303 207890
rect 156820 207832 160242 207888
rect 160298 207832 160303 207888
rect 156820 207830 160303 207832
rect 88661 207827 88727 207830
rect 160237 207827 160303 207830
rect 160605 207890 160671 207893
rect 163966 207890 164026 208132
rect 191750 207928 191810 208915
rect 201416 208888 201896 208918
rect 160605 207888 164026 207890
rect 160605 207832 160610 207888
rect 160666 207832 164026 207888
rect 160605 207830 164026 207832
rect 160605 207827 160671 207830
rect 88661 207754 88727 207757
rect 88661 207752 92052 207754
rect 88661 207696 88666 207752
rect 88722 207696 92052 207752
rect 88661 207694 92052 207696
rect 88661 207691 88727 207694
rect 51401 207618 51467 207621
rect 123161 207618 123227 207621
rect 47524 207616 51467 207618
rect 47524 207560 51406 207616
rect 51462 207560 51467 207616
rect 47524 207558 51467 207560
rect 119836 207616 123227 207618
rect 119836 207560 123166 207616
rect 123222 207560 123227 207616
rect 119836 207558 123227 207560
rect 51401 207555 51467 207558
rect 123161 207555 123227 207558
rect 160145 207618 160211 207621
rect 160145 207616 163996 207618
rect 160145 207560 160150 207616
rect 160206 207560 163996 207616
rect 160145 207558 163996 207560
rect 160145 207555 160211 207558
rect 51493 207482 51559 207485
rect 123253 207482 123319 207485
rect 51493 207480 55098 207482
rect 51493 207424 51498 207480
rect 51554 207424 55098 207480
rect 51493 207422 55098 207424
rect 51493 207419 51559 207422
rect 55038 207248 55098 207422
rect 123253 207480 127042 207482
rect 123253 207424 123258 207480
rect 123314 207424 127042 207480
rect 123253 207422 127042 207424
rect 123253 207419 123319 207422
rect 126982 207248 127042 207422
rect 88477 207210 88543 207213
rect 84876 207208 88543 207210
rect 84876 207152 88482 207208
rect 88538 207152 88543 207208
rect 84876 207150 88543 207152
rect 88477 207147 88543 207150
rect 88753 207210 88819 207213
rect 159041 207210 159107 207213
rect 88753 207208 92052 207210
rect 88753 207152 88758 207208
rect 88814 207152 92052 207208
rect 88753 207150 92052 207152
rect 156820 207208 159107 207210
rect 156820 207152 159046 207208
rect 159102 207152 159107 207208
rect 156820 207150 159107 207152
rect 88753 207147 88819 207150
rect 159041 207147 159107 207150
rect 51309 207074 51375 207077
rect 123069 207074 123135 207077
rect 160421 207074 160487 207077
rect 51309 207072 55098 207074
rect 47494 206802 47554 207044
rect 51309 207016 51314 207072
rect 51370 207016 55098 207072
rect 123069 207072 127042 207074
rect 51309 207014 55098 207016
rect 51309 207011 51375 207014
rect 51309 206802 51375 206805
rect 47494 206800 51375 206802
rect 47494 206744 51314 206800
rect 51370 206744 51375 206800
rect 47494 206742 51375 206744
rect 51309 206739 51375 206742
rect 55038 206704 55098 207014
rect 119806 206802 119866 207044
rect 123069 207016 123074 207072
rect 123130 207016 127042 207072
rect 123069 207014 127042 207016
rect 123069 207011 123135 207014
rect 122977 206802 123043 206805
rect 119806 206800 123043 206802
rect 119806 206744 122982 206800
rect 123038 206744 123043 206800
rect 119806 206742 123043 206744
rect 122977 206739 123043 206742
rect 126982 206704 127042 207014
rect 160421 207072 163996 207074
rect 160421 207016 160426 207072
rect 160482 207016 163996 207072
rect 160421 207014 163996 207016
rect 160421 207011 160487 207014
rect 88477 206666 88543 206669
rect 84876 206664 88543 206666
rect 84876 206608 88482 206664
rect 88538 206608 88543 206664
rect 84876 206606 88543 206608
rect 88477 206603 88543 206606
rect 88845 206666 88911 206669
rect 159041 206666 159107 206669
rect 88845 206664 92052 206666
rect 88845 206608 88850 206664
rect 88906 206608 92052 206664
rect 88845 206606 92052 206608
rect 156820 206664 159107 206666
rect 156820 206608 159046 206664
rect 159102 206608 159107 206664
rect 156820 206606 159107 206608
rect 88845 206603 88911 206606
rect 159041 206603 159107 206606
rect 51493 206530 51559 206533
rect 122977 206530 123043 206533
rect 47524 206528 51559 206530
rect 47524 206472 51498 206528
rect 51554 206472 51559 206528
rect 47524 206470 51559 206472
rect 119836 206528 123043 206530
rect 119836 206472 122982 206528
rect 123038 206472 123043 206528
rect 119836 206470 123043 206472
rect 51493 206467 51559 206470
rect 122977 206467 123043 206470
rect 160329 206530 160395 206533
rect 160329 206528 163996 206530
rect 160329 206472 160334 206528
rect 160390 206472 163996 206528
rect 160329 206470 163996 206472
rect 160329 206467 160395 206470
rect 88753 206258 88819 206261
rect 88526 206256 88819 206258
rect 88526 206200 88758 206256
rect 88814 206200 88819 206256
rect 88526 206198 88819 206200
rect 51401 206122 51467 206125
rect 88526 206122 88586 206198
rect 88753 206195 88819 206198
rect 51401 206120 55068 206122
rect 51401 206064 51406 206120
rect 51462 206064 55068 206120
rect 51401 206062 55068 206064
rect 84876 206062 88586 206122
rect 123161 206122 123227 206125
rect 160145 206122 160211 206125
rect 123161 206120 127012 206122
rect 123161 206064 123166 206120
rect 123222 206064 127012 206120
rect 123161 206062 127012 206064
rect 156820 206120 160211 206122
rect 156820 206064 160150 206120
rect 160206 206064 160211 206120
rect 156820 206062 160211 206064
rect 51401 206059 51467 206062
rect 123161 206059 123227 206062
rect 160145 206059 160211 206062
rect 51309 205986 51375 205989
rect 87189 205986 87255 205989
rect 122149 205986 122215 205989
rect 51309 205984 55098 205986
rect 47494 205578 47554 205956
rect 51309 205928 51314 205984
rect 51370 205928 55098 205984
rect 51309 205926 55098 205928
rect 51309 205923 51375 205926
rect 51585 205578 51651 205581
rect 47494 205576 51651 205578
rect 47494 205520 51590 205576
rect 51646 205520 51651 205576
rect 47494 205518 51651 205520
rect 51585 205515 51651 205518
rect 55038 205480 55098 205926
rect 87189 205984 92052 205986
rect 87189 205928 87194 205984
rect 87250 205928 92052 205984
rect 87189 205926 92052 205928
rect 119836 205984 122215 205986
rect 119836 205928 122154 205984
rect 122210 205928 122215 205984
rect 119836 205926 122215 205928
rect 87189 205923 87255 205926
rect 122149 205923 122215 205926
rect 123069 205986 123135 205989
rect 160513 205986 160579 205989
rect 123069 205984 127042 205986
rect 123069 205928 123074 205984
rect 123130 205928 127042 205984
rect 123069 205926 127042 205928
rect 123069 205923 123135 205926
rect 88477 205850 88543 205853
rect 84846 205848 88543 205850
rect 84846 205792 88482 205848
rect 88538 205792 88543 205848
rect 84846 205790 88543 205792
rect 84846 205412 84906 205790
rect 88477 205787 88543 205790
rect 126982 205480 127042 205926
rect 160513 205984 163996 205986
rect 160513 205928 160518 205984
rect 160574 205928 163996 205984
rect 160513 205926 163996 205928
rect 160513 205923 160579 205926
rect 160237 205442 160303 205445
rect 88526 205382 92052 205442
rect 156820 205440 160303 205442
rect 156820 205384 160242 205440
rect 160298 205384 160303 205440
rect 156820 205382 160303 205384
rect 51309 205306 51375 205309
rect 47524 205304 51375 205306
rect 47524 205248 51314 205304
rect 51370 205248 51375 205304
rect 47524 205246 51375 205248
rect 51309 205243 51375 205246
rect 51493 205306 51559 205309
rect 51493 205304 55098 205306
rect 51493 205248 51498 205304
rect 51554 205248 55098 205304
rect 51493 205246 55098 205248
rect 51493 205243 51559 205246
rect 55038 204936 55098 205246
rect 87189 204898 87255 204901
rect 84876 204896 87255 204898
rect 84876 204840 87194 204896
rect 87250 204840 87255 204896
rect 84876 204838 87255 204840
rect 87189 204835 87255 204838
rect 51401 204762 51467 204765
rect 47524 204760 51467 204762
rect 47524 204704 51406 204760
rect 51462 204704 51467 204760
rect 47524 204702 51467 204704
rect 51401 204699 51467 204702
rect 51585 204762 51651 204765
rect 88526 204762 88586 205382
rect 160237 205379 160303 205382
rect 123253 205306 123319 205309
rect 119836 205304 123319 205306
rect 119836 205248 123258 205304
rect 123314 205248 123319 205304
rect 119836 205246 123319 205248
rect 123253 205243 123319 205246
rect 160329 205306 160395 205309
rect 160329 205304 163996 205306
rect 160329 205248 160334 205304
rect 160390 205248 163996 205304
rect 160329 205246 163996 205248
rect 160329 205243 160395 205246
rect 123069 205170 123135 205173
rect 123069 205168 127042 205170
rect 123069 205112 123074 205168
rect 123130 205112 127042 205168
rect 123069 205110 127042 205112
rect 123069 205107 123135 205110
rect 126982 204936 127042 205110
rect 88661 204898 88727 204901
rect 160145 204898 160211 204901
rect 160513 204898 160579 204901
rect 88661 204896 92052 204898
rect 88661 204840 88666 204896
rect 88722 204840 92052 204896
rect 88661 204838 92052 204840
rect 156820 204896 160211 204898
rect 156820 204840 160150 204896
rect 160206 204840 160211 204896
rect 156820 204838 160211 204840
rect 88661 204835 88727 204838
rect 160145 204835 160211 204838
rect 160286 204896 160579 204898
rect 160286 204840 160518 204896
rect 160574 204840 160579 204896
rect 160286 204838 160579 204840
rect 122977 204762 123043 204765
rect 160286 204762 160346 204838
rect 160513 204835 160579 204838
rect 51585 204760 55098 204762
rect 51585 204704 51590 204760
rect 51646 204704 55098 204760
rect 51585 204702 55098 204704
rect 51585 204699 51651 204702
rect 55038 204256 55098 204702
rect 84846 204702 88586 204762
rect 119836 204760 123043 204762
rect 119836 204704 122982 204760
rect 123038 204704 123043 204760
rect 119836 204702 123043 204704
rect 84846 204188 84906 204702
rect 122977 204699 123043 204702
rect 156790 204702 160346 204762
rect 160421 204762 160487 204765
rect 160421 204760 163996 204762
rect 160421 204704 160426 204760
rect 160482 204704 163996 204760
rect 160421 204702 163996 204704
rect 124357 204490 124423 204493
rect 124357 204488 127042 204490
rect 124357 204432 124362 204488
rect 124418 204432 127042 204488
rect 124357 204430 127042 204432
rect 124357 204427 124423 204430
rect 88661 204354 88727 204357
rect 88661 204352 92052 204354
rect 88661 204296 88666 204352
rect 88722 204296 92052 204352
rect 88661 204294 92052 204296
rect 88661 204291 88727 204294
rect 126982 204256 127042 204430
rect 122977 204218 123043 204221
rect 119836 204216 123043 204218
rect 47494 203946 47554 204188
rect 119836 204160 122982 204216
rect 123038 204160 123043 204216
rect 156790 204188 156850 204702
rect 160421 204699 160487 204702
rect 119836 204158 123043 204160
rect 122977 204155 123043 204158
rect 51309 204082 51375 204085
rect 123253 204082 123319 204085
rect 51309 204080 55098 204082
rect 51309 204024 51314 204080
rect 51370 204024 55098 204080
rect 51309 204022 55098 204024
rect 51309 204019 51375 204022
rect 51309 203946 51375 203949
rect 47494 203944 51375 203946
rect 47494 203888 51314 203944
rect 51370 203888 51375 203944
rect 47494 203886 51375 203888
rect 51309 203883 51375 203886
rect 55038 203712 55098 204022
rect 123253 204080 127042 204082
rect 123253 204024 123258 204080
rect 123314 204024 127042 204080
rect 123253 204022 127042 204024
rect 123253 204019 123319 204022
rect 88753 203810 88819 203813
rect 88753 203808 92052 203810
rect 88753 203752 88758 203808
rect 88814 203752 92052 203808
rect 88753 203750 92052 203752
rect 88753 203747 88819 203750
rect 126982 203712 127042 204022
rect 160329 203946 160395 203949
rect 163966 203946 164026 204188
rect 160329 203944 164026 203946
rect 160329 203888 160334 203944
rect 160390 203888 164026 203944
rect 160329 203886 164026 203888
rect 160329 203883 160395 203886
rect 51493 203674 51559 203677
rect 88477 203674 88543 203677
rect 123161 203674 123227 203677
rect 160237 203674 160303 203677
rect 47524 203672 51559 203674
rect 47524 203616 51498 203672
rect 51554 203616 51559 203672
rect 47524 203614 51559 203616
rect 84876 203672 88543 203674
rect 84876 203616 88482 203672
rect 88538 203616 88543 203672
rect 84876 203614 88543 203616
rect 119836 203672 123227 203674
rect 119836 203616 123166 203672
rect 123222 203616 123227 203672
rect 119836 203614 123227 203616
rect 156820 203672 160303 203674
rect 156820 203616 160242 203672
rect 160298 203616 160303 203672
rect 156820 203614 160303 203616
rect 51493 203611 51559 203614
rect 88477 203611 88543 203614
rect 123161 203611 123227 203614
rect 160237 203611 160303 203614
rect 160513 203674 160579 203677
rect 160513 203672 163996 203674
rect 160513 203616 160518 203672
rect 160574 203616 163996 203672
rect 160513 203614 163996 203616
rect 160513 203611 160579 203614
rect 88661 203538 88727 203541
rect 160421 203538 160487 203541
rect 88526 203536 88727 203538
rect 88526 203480 88666 203536
rect 88722 203480 88727 203536
rect 88526 203478 88727 203480
rect 51401 203402 51467 203405
rect 88526 203402 88586 203478
rect 88661 203475 88727 203478
rect 160286 203536 160487 203538
rect 160286 203480 160426 203536
rect 160482 203480 160487 203536
rect 160286 203478 160487 203480
rect 51401 203400 55098 203402
rect 51401 203344 51406 203400
rect 51462 203344 55098 203400
rect 51401 203342 55098 203344
rect 51401 203339 51467 203342
rect 55038 203168 55098 203342
rect 84846 203342 88586 203402
rect 123069 203402 123135 203405
rect 160286 203402 160346 203478
rect 160421 203475 160487 203478
rect 123069 203400 127042 203402
rect 123069 203344 123074 203400
rect 123130 203344 127042 203400
rect 123069 203342 127042 203344
rect 51401 203130 51467 203133
rect 47524 203128 51467 203130
rect 47524 203072 51406 203128
rect 51462 203072 51467 203128
rect 84846 203100 84906 203342
rect 123069 203339 123135 203342
rect 88845 203266 88911 203269
rect 88845 203264 92052 203266
rect 88845 203208 88850 203264
rect 88906 203208 92052 203264
rect 88845 203206 92052 203208
rect 88845 203203 88911 203206
rect 126982 203168 127042 203342
rect 156790 203342 160346 203402
rect 123253 203130 123319 203133
rect 119836 203128 123319 203130
rect 47524 203070 51467 203072
rect 119836 203072 123258 203128
rect 123314 203072 123319 203128
rect 156790 203100 156850 203342
rect 160605 203130 160671 203133
rect 160605 203128 163996 203130
rect 119836 203070 123319 203072
rect 51401 203067 51467 203070
rect 123253 203067 123319 203070
rect 160605 203072 160610 203128
rect 160666 203072 163996 203128
rect 160605 203070 163996 203072
rect 160605 203067 160671 203070
rect 51309 202994 51375 202997
rect 123069 202994 123135 202997
rect 51309 202992 55098 202994
rect 51309 202936 51314 202992
rect 51370 202936 55098 202992
rect 51309 202934 55098 202936
rect 51309 202931 51375 202934
rect 55038 202488 55098 202934
rect 123069 202992 127042 202994
rect 123069 202936 123074 202992
rect 123130 202936 127042 202992
rect 123069 202934 127042 202936
rect 123069 202931 123135 202934
rect 88937 202722 89003 202725
rect 88937 202720 92052 202722
rect 88937 202664 88942 202720
rect 88998 202664 92052 202720
rect 88937 202662 92052 202664
rect 88937 202659 89003 202662
rect 126982 202488 127042 202934
rect 51309 202450 51375 202453
rect 88477 202450 88543 202453
rect 122977 202450 123043 202453
rect 160237 202450 160303 202453
rect 47524 202448 51375 202450
rect 47524 202392 51314 202448
rect 51370 202392 51375 202448
rect 47524 202390 51375 202392
rect 84876 202448 88543 202450
rect 84876 202392 88482 202448
rect 88538 202392 88543 202448
rect 84876 202390 88543 202392
rect 119836 202448 123043 202450
rect 119836 202392 122982 202448
rect 123038 202392 123043 202448
rect 119836 202390 123043 202392
rect 156820 202448 160303 202450
rect 156820 202392 160242 202448
rect 160298 202392 160303 202448
rect 156820 202390 160303 202392
rect 51309 202387 51375 202390
rect 88477 202387 88543 202390
rect 122977 202387 123043 202390
rect 160237 202387 160303 202390
rect 160421 202450 160487 202453
rect 160421 202448 163996 202450
rect 160421 202392 160426 202448
rect 160482 202392 163996 202448
rect 160421 202390 163996 202392
rect 160421 202387 160487 202390
rect 88569 202314 88635 202317
rect 88569 202312 91530 202314
rect 88569 202256 88574 202312
rect 88630 202256 91530 202312
rect 88569 202254 91530 202256
rect 88569 202251 88635 202254
rect 91470 202246 91530 202254
rect 91470 202186 92052 202246
rect 88845 202178 88911 202181
rect 88526 202176 88911 202178
rect 88526 202120 88850 202176
rect 88906 202120 88911 202176
rect 88526 202118 88911 202120
rect 50297 202042 50363 202045
rect 50481 202042 50547 202045
rect 88526 202042 88586 202118
rect 88845 202115 88911 202118
rect 50297 202040 50547 202042
rect 50297 201984 50302 202040
rect 50358 201984 50486 202040
rect 50542 201984 50547 202040
rect 50297 201982 50547 201984
rect 50297 201979 50363 201982
rect 50481 201979 50547 201982
rect 84846 201982 88586 202042
rect 51217 201906 51283 201909
rect 47524 201904 51283 201906
rect 47524 201848 51222 201904
rect 51278 201848 51283 201904
rect 47524 201846 51283 201848
rect 51217 201843 51283 201846
rect 51493 201906 51559 201909
rect 51493 201904 55068 201906
rect 51493 201848 51498 201904
rect 51554 201848 55068 201904
rect 84846 201876 84906 201982
rect 122977 201906 123043 201909
rect 119836 201904 123043 201906
rect 51493 201846 55068 201848
rect 119836 201848 122982 201904
rect 123038 201848 123043 201904
rect 119836 201846 123043 201848
rect 51493 201843 51559 201846
rect 122977 201843 123043 201846
rect 123161 201906 123227 201909
rect 159041 201906 159107 201909
rect 123161 201904 127012 201906
rect 123161 201848 123166 201904
rect 123222 201848 127012 201904
rect 123161 201846 127012 201848
rect 156820 201904 159107 201906
rect 156820 201848 159046 201904
rect 159102 201848 159107 201904
rect 156820 201846 159107 201848
rect 123161 201843 123227 201846
rect 159041 201843 159107 201846
rect 160513 201906 160579 201909
rect 160513 201904 163996 201906
rect 160513 201848 160518 201904
rect 160574 201848 163996 201904
rect 160513 201846 163996 201848
rect 160513 201843 160579 201846
rect 51401 201770 51467 201773
rect 123253 201770 123319 201773
rect 51401 201768 55098 201770
rect 51401 201712 51406 201768
rect 51462 201712 55098 201768
rect 51401 201710 55098 201712
rect 51401 201707 51467 201710
rect 51493 201362 51559 201365
rect 47524 201360 51559 201362
rect 47524 201304 51498 201360
rect 51554 201304 51559 201360
rect 47524 201302 51559 201304
rect 51493 201299 51559 201302
rect 55038 201264 55098 201710
rect 123253 201768 127042 201770
rect 123253 201712 123258 201768
rect 123314 201712 127042 201768
rect 123253 201710 127042 201712
rect 123253 201707 123319 201710
rect 88569 201498 88635 201501
rect 88569 201496 92052 201498
rect 88569 201440 88574 201496
rect 88630 201440 92052 201496
rect 88569 201438 92052 201440
rect 88569 201435 88635 201438
rect 123161 201362 123227 201365
rect 119836 201360 123227 201362
rect 119836 201304 123166 201360
rect 123222 201304 123227 201360
rect 119836 201302 123227 201304
rect 123161 201299 123227 201302
rect 126982 201264 127042 201710
rect 160329 201362 160395 201365
rect 160329 201360 163996 201362
rect 160329 201304 160334 201360
rect 160390 201304 163996 201360
rect 160329 201302 163996 201304
rect 160329 201299 160395 201302
rect 87189 201226 87255 201229
rect 158949 201226 159015 201229
rect 84876 201224 87255 201226
rect 84876 201168 87194 201224
rect 87250 201168 87255 201224
rect 84876 201166 87255 201168
rect 156820 201224 159015 201226
rect 156820 201168 158954 201224
rect 159010 201168 159015 201224
rect 156820 201166 159015 201168
rect 87189 201163 87255 201166
rect 158949 201163 159015 201166
rect 51309 201090 51375 201093
rect 123069 201090 123135 201093
rect 51309 201088 55098 201090
rect 51309 201032 51314 201088
rect 51370 201032 55098 201088
rect 51309 201030 55098 201032
rect 51309 201027 51375 201030
rect 51401 200818 51467 200821
rect 47524 200816 51467 200818
rect 47524 200760 51406 200816
rect 51462 200760 51467 200816
rect 47524 200758 51467 200760
rect 51401 200755 51467 200758
rect 55038 200720 55098 201030
rect 123069 201088 127042 201090
rect 123069 201032 123074 201088
rect 123130 201032 127042 201088
rect 123069 201030 127042 201032
rect 123069 201027 123135 201030
rect 88661 200954 88727 200957
rect 88661 200952 92052 200954
rect 88661 200896 88666 200952
rect 88722 200896 92052 200952
rect 88661 200894 92052 200896
rect 88661 200891 88727 200894
rect 122977 200818 123043 200821
rect 119836 200816 123043 200818
rect 119836 200760 122982 200816
rect 123038 200760 123043 200816
rect 119836 200758 123043 200760
rect 122977 200755 123043 200758
rect 126982 200720 127042 201030
rect 160145 200818 160211 200821
rect 160145 200816 163996 200818
rect 160145 200760 160150 200816
rect 160206 200760 163996 200816
rect 160145 200758 163996 200760
rect 160145 200755 160211 200758
rect 88477 200682 88543 200685
rect 160237 200682 160303 200685
rect 160513 200682 160579 200685
rect 84876 200680 88543 200682
rect 84876 200624 88482 200680
rect 88538 200624 88543 200680
rect 84876 200622 88543 200624
rect 156820 200680 160303 200682
rect 156820 200624 160242 200680
rect 160298 200624 160303 200680
rect 156820 200622 160303 200624
rect 88477 200619 88543 200622
rect 160237 200619 160303 200622
rect 160470 200680 160579 200682
rect 160470 200624 160518 200680
rect 160574 200624 160579 200680
rect 160470 200619 160579 200624
rect 51309 200546 51375 200549
rect 123069 200546 123135 200549
rect 160470 200546 160530 200619
rect 51309 200544 55098 200546
rect 51309 200488 51314 200544
rect 51370 200488 55098 200544
rect 51309 200486 55098 200488
rect 51309 200483 51375 200486
rect 51309 200274 51375 200277
rect 47524 200272 51375 200274
rect 47524 200216 51314 200272
rect 51370 200216 51375 200272
rect 47524 200214 51375 200216
rect 51309 200211 51375 200214
rect 55038 200176 55098 200486
rect 123069 200544 127042 200546
rect 123069 200488 123074 200544
rect 123130 200488 127042 200544
rect 123069 200486 127042 200488
rect 123069 200483 123135 200486
rect 88753 200410 88819 200413
rect 88753 200408 92052 200410
rect 88753 200352 88758 200408
rect 88814 200352 92052 200408
rect 88753 200350 92052 200352
rect 88753 200347 88819 200350
rect 88477 200138 88543 200141
rect 84876 200136 88543 200138
rect 84876 200080 88482 200136
rect 88538 200080 88543 200136
rect 84876 200078 88543 200080
rect 88477 200075 88543 200078
rect 51493 200002 51559 200005
rect 51493 200000 55098 200002
rect 51493 199944 51498 200000
rect 51554 199944 55098 200000
rect 51493 199942 55098 199944
rect 51493 199939 51559 199942
rect 51493 199594 51559 199597
rect 47524 199592 51559 199594
rect 47524 199536 51498 199592
rect 51554 199536 51559 199592
rect 47524 199534 51559 199536
rect 51493 199531 51559 199534
rect 55038 199496 55098 199942
rect 88845 199866 88911 199869
rect 119806 199866 119866 200244
rect 126982 200176 127042 200486
rect 156790 200486 160530 200546
rect 156790 200108 156850 200486
rect 160513 200274 160579 200277
rect 160513 200272 163996 200274
rect 160513 200216 160518 200272
rect 160574 200216 163996 200272
rect 160513 200214 163996 200216
rect 160513 200211 160579 200214
rect 123161 200002 123227 200005
rect 123161 200000 127042 200002
rect 123161 199944 123166 200000
rect 123222 199944 127042 200000
rect 123161 199942 127042 199944
rect 123161 199939 123227 199942
rect 123161 199866 123227 199869
rect 88845 199864 92052 199866
rect 88845 199808 88850 199864
rect 88906 199808 92052 199864
rect 88845 199806 92052 199808
rect 119806 199864 123227 199866
rect 119806 199808 123166 199864
rect 123222 199808 123227 199864
rect 119806 199806 123227 199808
rect 88845 199803 88911 199806
rect 123161 199803 123227 199806
rect 122977 199594 123043 199597
rect 119836 199592 123043 199594
rect 119836 199536 122982 199592
rect 123038 199536 123043 199592
rect 119836 199534 123043 199536
rect 122977 199531 123043 199534
rect 126982 199496 127042 199942
rect 88477 199458 88543 199461
rect 160237 199458 160303 199461
rect 84876 199456 88543 199458
rect 84876 199400 88482 199456
rect 88538 199400 88543 199456
rect 84876 199398 88543 199400
rect 156820 199456 160303 199458
rect 156820 199400 160242 199456
rect 160298 199400 160303 199456
rect 156820 199398 160303 199400
rect 88477 199395 88543 199398
rect 160237 199395 160303 199398
rect 88753 199322 88819 199325
rect 88480 199320 88819 199322
rect 88480 199264 88758 199320
rect 88814 199264 88819 199320
rect 88480 199262 88819 199264
rect 88480 199186 88540 199262
rect 88753 199259 88819 199262
rect 88937 199322 89003 199325
rect 160237 199322 160303 199325
rect 163966 199322 164026 199564
rect 88937 199320 92052 199322
rect 88937 199264 88942 199320
rect 88998 199264 92052 199320
rect 88937 199262 92052 199264
rect 160237 199320 164026 199322
rect 160237 199264 160242 199320
rect 160298 199264 164026 199320
rect 160237 199262 164026 199264
rect 88937 199259 89003 199262
rect 160237 199259 160303 199262
rect 84846 199126 88540 199186
rect 123069 199186 123135 199189
rect 123069 199184 127042 199186
rect 123069 199128 123074 199184
rect 123130 199128 127042 199184
rect 123069 199126 127042 199128
rect 51401 199050 51467 199053
rect 51401 199048 54546 199050
rect 47494 198914 47554 199020
rect 51401 198992 51406 199048
rect 51462 198992 54546 199048
rect 51401 198990 54546 198992
rect 51401 198987 51467 198990
rect 54486 198982 54546 198990
rect 54486 198922 55068 198982
rect 51401 198914 51467 198917
rect 47494 198912 51467 198914
rect 47494 198856 51406 198912
rect 51462 198856 51467 198912
rect 84846 198884 84906 199126
rect 123069 199123 123135 199126
rect 47494 198854 51467 198856
rect 51401 198851 51467 198854
rect 51309 198778 51375 198781
rect 88937 198778 89003 198781
rect 119806 198778 119866 199020
rect 126982 198952 127042 199126
rect 160421 199050 160487 199053
rect 160421 199048 163996 199050
rect 160421 198992 160426 199048
rect 160482 198992 163996 199048
rect 160421 198990 163996 198992
rect 160421 198987 160487 198990
rect 160145 198914 160211 198917
rect 156820 198912 160211 198914
rect 156820 198856 160150 198912
rect 160206 198856 160211 198912
rect 156820 198854 160211 198856
rect 160145 198851 160211 198854
rect 122977 198778 123043 198781
rect 51309 198776 55098 198778
rect 51309 198720 51314 198776
rect 51370 198720 55098 198776
rect 51309 198718 55098 198720
rect 51309 198715 51375 198718
rect 51309 198506 51375 198509
rect 47524 198504 51375 198506
rect 47524 198448 51314 198504
rect 51370 198448 51375 198504
rect 47524 198446 51375 198448
rect 51309 198443 51375 198446
rect 55038 198272 55098 198718
rect 88937 198776 92052 198778
rect 88937 198720 88942 198776
rect 88998 198720 92052 198776
rect 88937 198718 92052 198720
rect 119806 198776 123043 198778
rect 119806 198720 122982 198776
rect 123038 198720 123043 198776
rect 119806 198718 123043 198720
rect 88937 198715 89003 198718
rect 122977 198715 123043 198718
rect 123161 198778 123227 198781
rect 123161 198776 127042 198778
rect 123161 198720 123166 198776
rect 123222 198720 127042 198776
rect 123161 198718 127042 198720
rect 123161 198715 123227 198718
rect 123161 198506 123227 198509
rect 119836 198504 123227 198506
rect 119836 198448 123166 198504
rect 123222 198448 123227 198504
rect 119836 198446 123227 198448
rect 123161 198443 123227 198446
rect 126982 198272 127042 198718
rect 160053 198506 160119 198509
rect 160053 198504 163996 198506
rect 160053 198448 160058 198504
rect 160114 198448 163996 198504
rect 160053 198446 163996 198448
rect 160053 198443 160119 198446
rect 88477 198234 88543 198237
rect 84876 198232 88543 198234
rect 84876 198176 88482 198232
rect 88538 198176 88543 198232
rect 84876 198174 88543 198176
rect 88477 198171 88543 198174
rect 88661 198234 88727 198237
rect 158949 198234 159015 198237
rect 88661 198232 92052 198234
rect 88661 198176 88666 198232
rect 88722 198176 92052 198232
rect 88661 198174 92052 198176
rect 156820 198232 159015 198234
rect 156820 198176 158954 198232
rect 159010 198176 159015 198232
rect 156820 198174 159015 198176
rect 88661 198171 88727 198174
rect 158949 198171 159015 198174
rect 51585 197962 51651 197965
rect 123253 197962 123319 197965
rect 47524 197960 51651 197962
rect 47524 197904 51590 197960
rect 51646 197904 51651 197960
rect 47524 197902 51651 197904
rect 119836 197960 123319 197962
rect 119836 197904 123258 197960
rect 123314 197904 123319 197960
rect 119836 197902 123319 197904
rect 51585 197899 51651 197902
rect 123253 197899 123319 197902
rect 160237 197962 160303 197965
rect 160237 197960 163996 197962
rect 160237 197904 160242 197960
rect 160298 197904 163996 197960
rect 160237 197902 163996 197904
rect 160237 197899 160303 197902
rect 123069 197826 123135 197829
rect 123069 197824 126490 197826
rect 123069 197768 123074 197824
rect 123130 197768 126490 197824
rect 123069 197766 126490 197768
rect 123069 197763 123135 197766
rect 126430 197758 126490 197766
rect 126430 197698 127012 197758
rect 51493 197690 51559 197693
rect 87189 197690 87255 197693
rect 51493 197688 55068 197690
rect 51493 197632 51498 197688
rect 51554 197632 55068 197688
rect 51493 197630 55068 197632
rect 84876 197688 87255 197690
rect 84876 197632 87194 197688
rect 87250 197632 87255 197688
rect 84876 197630 87255 197632
rect 51493 197627 51559 197630
rect 87189 197627 87255 197630
rect 88569 197690 88635 197693
rect 160145 197690 160211 197693
rect 88569 197688 92052 197690
rect 88569 197632 88574 197688
rect 88630 197632 92052 197688
rect 88569 197630 92052 197632
rect 156820 197688 160211 197690
rect 156820 197632 160150 197688
rect 160206 197632 160211 197688
rect 156820 197630 160211 197632
rect 88569 197627 88635 197630
rect 160145 197627 160211 197630
rect 51401 197554 51467 197557
rect 123069 197554 123135 197557
rect 51401 197552 55098 197554
rect 51401 197496 51406 197552
rect 51462 197496 55098 197552
rect 51401 197494 55098 197496
rect 51401 197491 51467 197494
rect 51493 197418 51559 197421
rect 47524 197416 51559 197418
rect 47524 197360 51498 197416
rect 51554 197360 51559 197416
rect 47524 197358 51559 197360
rect 51493 197355 51559 197358
rect 55038 197184 55098 197494
rect 123069 197552 127042 197554
rect 123069 197496 123074 197552
rect 123130 197496 127042 197552
rect 123069 197494 127042 197496
rect 123069 197491 123135 197494
rect 122977 197418 123043 197421
rect 119836 197416 123043 197418
rect 119836 197360 122982 197416
rect 123038 197360 123043 197416
rect 119836 197358 123043 197360
rect 122977 197355 123043 197358
rect 126982 197184 127042 197494
rect 160513 197418 160579 197421
rect 160513 197416 163996 197418
rect 160513 197360 160518 197416
rect 160574 197360 163996 197416
rect 160513 197358 163996 197360
rect 160513 197355 160579 197358
rect 191558 197356 191564 197420
rect 191628 197356 191634 197420
rect 87189 197146 87255 197149
rect 84876 197144 87255 197146
rect 84876 197088 87194 197144
rect 87250 197088 87255 197144
rect 84876 197086 87255 197088
rect 87189 197083 87255 197086
rect 88661 197146 88727 197149
rect 160237 197146 160303 197149
rect 88661 197144 92052 197146
rect 88661 197088 88666 197144
rect 88722 197088 92052 197144
rect 88661 197086 92052 197088
rect 156820 197144 160303 197146
rect 156820 197088 160242 197144
rect 160298 197088 160303 197144
rect 156820 197086 160303 197088
rect 88661 197083 88727 197086
rect 160237 197083 160303 197086
rect 191566 196776 191626 197356
rect 51401 196738 51467 196741
rect 121781 196738 121847 196741
rect 47524 196736 51467 196738
rect 47524 196680 51406 196736
rect 51462 196680 51467 196736
rect 47524 196678 51467 196680
rect 119836 196736 121847 196738
rect 119836 196680 121786 196736
rect 121842 196680 121847 196736
rect 119836 196678 121847 196680
rect 51401 196675 51467 196678
rect 121781 196675 121847 196678
rect 160237 196738 160303 196741
rect 160237 196736 163996 196738
rect 160237 196680 160242 196736
rect 160298 196680 163996 196736
rect 160237 196678 163996 196680
rect 160237 196675 160303 196678
rect 51309 196466 51375 196469
rect 88477 196466 88543 196469
rect 51309 196464 55068 196466
rect 51309 196408 51314 196464
rect 51370 196408 55068 196464
rect 51309 196406 55068 196408
rect 84876 196464 88543 196466
rect 84876 196408 88482 196464
rect 88538 196408 88543 196464
rect 84876 196406 88543 196408
rect 51309 196403 51375 196406
rect 88477 196403 88543 196406
rect 89213 196466 89279 196469
rect 123161 196466 123227 196469
rect 160053 196466 160119 196469
rect 89213 196464 92052 196466
rect 89213 196408 89218 196464
rect 89274 196408 92052 196464
rect 89213 196406 92052 196408
rect 123161 196464 127012 196466
rect 123161 196408 123166 196464
rect 123222 196408 127012 196464
rect 123161 196406 127012 196408
rect 156820 196464 160119 196466
rect 156820 196408 160058 196464
rect 160114 196408 160119 196464
rect 156820 196406 160119 196408
rect 89213 196403 89279 196406
rect 123161 196403 123227 196406
rect 160053 196403 160119 196406
rect 51585 196330 51651 196333
rect 88477 196330 88543 196333
rect 51585 196328 55098 196330
rect 51585 196272 51590 196328
rect 51646 196272 55098 196328
rect 51585 196270 55098 196272
rect 51585 196267 51651 196270
rect 51309 196194 51375 196197
rect 47524 196192 51375 196194
rect 47524 196136 51314 196192
rect 51370 196136 51375 196192
rect 47524 196134 51375 196136
rect 51309 196131 51375 196134
rect 55038 195960 55098 196270
rect 84846 196328 88543 196330
rect 84846 196272 88482 196328
rect 88538 196272 88543 196328
rect 84846 196270 88543 196272
rect 84846 195892 84906 196270
rect 88477 196267 88543 196270
rect 123253 196330 123319 196333
rect 123253 196328 127042 196330
rect 123253 196272 123258 196328
rect 123314 196272 127042 196328
rect 123253 196270 127042 196272
rect 123253 196267 123319 196270
rect 123069 196194 123135 196197
rect 119836 196192 123135 196194
rect 119836 196136 123074 196192
rect 123130 196136 123135 196192
rect 119836 196134 123135 196136
rect 123069 196131 123135 196134
rect 126982 195960 127042 196270
rect 160329 196194 160395 196197
rect 160329 196192 163996 196194
rect 160329 196136 160334 196192
rect 160390 196136 163996 196192
rect 160329 196134 163996 196136
rect 160329 196131 160395 196134
rect 88569 195922 88635 195925
rect 160145 195922 160211 195925
rect 88569 195920 92052 195922
rect 88569 195864 88574 195920
rect 88630 195864 92052 195920
rect 88569 195862 92052 195864
rect 156820 195920 160211 195922
rect 156820 195864 160150 195920
rect 160206 195864 160211 195920
rect 156820 195862 160211 195864
rect 88569 195859 88635 195862
rect 160145 195859 160211 195862
rect 51493 195786 51559 195789
rect 88477 195786 88543 195789
rect 51493 195784 55098 195786
rect 51493 195728 51498 195784
rect 51554 195728 55098 195784
rect 51493 195726 55098 195728
rect 51493 195723 51559 195726
rect 51493 195650 51559 195653
rect 47524 195648 51559 195650
rect 47524 195592 51498 195648
rect 51554 195592 51559 195648
rect 47524 195590 51559 195592
rect 51493 195587 51559 195590
rect 55038 195280 55098 195726
rect 84846 195784 88543 195786
rect 84846 195728 88482 195784
rect 88538 195728 88543 195784
rect 84846 195726 88543 195728
rect 84846 195212 84906 195726
rect 88477 195723 88543 195726
rect 123161 195786 123227 195789
rect 123161 195784 127042 195786
rect 123161 195728 123166 195784
rect 123222 195728 127042 195784
rect 123161 195726 127042 195728
rect 123161 195723 123227 195726
rect 123161 195650 123227 195653
rect 119836 195648 123227 195650
rect 119836 195592 123166 195648
rect 123222 195592 123227 195648
rect 119836 195590 123227 195592
rect 123161 195587 123227 195590
rect 88385 195378 88451 195381
rect 88385 195376 92052 195378
rect 88385 195320 88390 195376
rect 88446 195320 92052 195376
rect 88385 195318 92052 195320
rect 88385 195315 88451 195318
rect 126982 195280 127042 195726
rect 160145 195650 160211 195653
rect 160145 195648 163996 195650
rect 160145 195592 160150 195648
rect 160206 195592 163996 195648
rect 160145 195590 163996 195592
rect 160145 195587 160211 195590
rect 89213 195242 89279 195245
rect 158949 195242 159015 195245
rect 88480 195240 89279 195242
rect 88480 195184 89218 195240
rect 89274 195184 89279 195240
rect 88480 195182 89279 195184
rect 156820 195240 159015 195242
rect 156820 195184 158954 195240
rect 159010 195184 159015 195240
rect 156820 195182 159015 195184
rect 51401 195106 51467 195109
rect 88480 195106 88540 195182
rect 89213 195179 89279 195182
rect 158949 195179 159015 195182
rect 122977 195106 123043 195109
rect 51401 195104 55098 195106
rect 47494 194834 47554 195076
rect 51401 195048 51406 195104
rect 51462 195048 55098 195104
rect 51401 195046 55098 195048
rect 51401 195043 51467 195046
rect 51401 194834 51467 194837
rect 47494 194832 51467 194834
rect 47494 194776 51406 194832
rect 51462 194776 51467 194832
rect 47494 194774 51467 194776
rect 51401 194771 51467 194774
rect 55038 194736 55098 195046
rect 84846 195046 88540 195106
rect 119836 195104 123043 195106
rect 119836 195048 122982 195104
rect 123038 195048 123043 195104
rect 119836 195046 123043 195048
rect 84846 194668 84906 195046
rect 122977 195043 123043 195046
rect 160421 195106 160487 195109
rect 160421 195104 163996 195106
rect 160421 195048 160426 195104
rect 160482 195048 163996 195104
rect 160421 195046 163996 195048
rect 160421 195043 160487 195046
rect 124173 194970 124239 194973
rect 124173 194968 127042 194970
rect 124173 194912 124178 194968
rect 124234 194912 127042 194968
rect 124173 194910 127042 194912
rect 124173 194907 124239 194910
rect 88661 194834 88727 194837
rect 88661 194832 92052 194834
rect 88661 194776 88666 194832
rect 88722 194776 92052 194832
rect 88661 194774 92052 194776
rect 88661 194771 88727 194774
rect 126982 194736 127042 194910
rect 160237 194698 160303 194701
rect 156820 194696 160303 194698
rect 156820 194640 160242 194696
rect 160298 194640 160303 194696
rect 156820 194638 160303 194640
rect 160237 194635 160303 194638
rect 51309 194562 51375 194565
rect 122241 194562 122307 194565
rect 51309 194560 55098 194562
rect 47494 194154 47554 194532
rect 51309 194504 51314 194560
rect 51370 194504 55098 194560
rect 51309 194502 55098 194504
rect 119836 194560 122307 194562
rect 119836 194504 122246 194560
rect 122302 194504 122307 194560
rect 119836 194502 122307 194504
rect 51309 194499 51375 194502
rect 55038 194192 55098 194502
rect 122241 194499 122307 194502
rect 123069 194562 123135 194565
rect 159961 194562 160027 194565
rect 123069 194560 127042 194562
rect 123069 194504 123074 194560
rect 123130 194504 127042 194560
rect 123069 194502 127042 194504
rect 123069 194499 123135 194502
rect 88293 194290 88359 194293
rect 88293 194288 92052 194290
rect 88293 194232 88298 194288
rect 88354 194232 92052 194288
rect 88293 194230 92052 194232
rect 88293 194227 88359 194230
rect 126982 194192 127042 194502
rect 159961 194560 163996 194562
rect 159961 194504 159966 194560
rect 160022 194504 163996 194560
rect 159961 194502 163996 194504
rect 159961 194499 160027 194502
rect 51585 194154 51651 194157
rect 88477 194154 88543 194157
rect 160237 194154 160303 194157
rect 47494 194152 51651 194154
rect 47494 194096 51590 194152
rect 51646 194096 51651 194152
rect 47494 194094 51651 194096
rect 84876 194152 88543 194154
rect 84876 194096 88482 194152
rect 88538 194096 88543 194152
rect 84876 194094 88543 194096
rect 156820 194152 160303 194154
rect 156820 194096 160242 194152
rect 160298 194096 160303 194152
rect 156820 194094 160303 194096
rect 51585 194091 51651 194094
rect 88477 194091 88543 194094
rect 160237 194091 160303 194094
rect 51309 193882 51375 193885
rect 123253 193882 123319 193885
rect 47524 193880 51375 193882
rect 47524 193824 51314 193880
rect 51370 193824 51375 193880
rect 47524 193822 51375 193824
rect 119836 193880 123319 193882
rect 119836 193824 123258 193880
rect 123314 193824 123319 193880
rect 119836 193822 123319 193824
rect 51309 193819 51375 193822
rect 123253 193819 123319 193822
rect 160053 193882 160119 193885
rect 160053 193880 163996 193882
rect 160053 193824 160058 193880
rect 160114 193824 163996 193880
rect 160053 193822 163996 193824
rect 160053 193819 160119 193822
rect 51493 193746 51559 193749
rect 88753 193746 88819 193749
rect 123161 193746 123227 193749
rect 51493 193744 55098 193746
rect 51493 193688 51498 193744
rect 51554 193688 55098 193744
rect 51493 193686 55098 193688
rect 51493 193683 51559 193686
rect 55038 193512 55098 193686
rect 88753 193744 92052 193746
rect 88753 193688 88758 193744
rect 88814 193688 92052 193744
rect 88753 193686 92052 193688
rect 123161 193744 127042 193746
rect 123161 193688 123166 193744
rect 123222 193688 127042 193744
rect 123161 193686 127042 193688
rect 88753 193683 88819 193686
rect 123161 193683 123227 193686
rect 126982 193512 127042 193686
rect 88385 193474 88451 193477
rect 160145 193474 160211 193477
rect 84876 193472 88451 193474
rect 84876 193416 88390 193472
rect 88446 193416 88451 193472
rect 84876 193414 88451 193416
rect 156820 193472 160211 193474
rect 156820 193416 160150 193472
rect 160206 193416 160211 193472
rect 156820 193414 160211 193416
rect 88385 193411 88451 193414
rect 160145 193411 160211 193414
rect 51401 193338 51467 193341
rect 123069 193338 123135 193341
rect 160513 193338 160579 193341
rect 51401 193336 55098 193338
rect 47494 193066 47554 193308
rect 51401 193280 51406 193336
rect 51462 193280 55098 193336
rect 123069 193336 127042 193338
rect 51401 193278 55098 193280
rect 51401 193275 51467 193278
rect 51309 193066 51375 193069
rect 47494 193064 51375 193066
rect 47494 193008 51314 193064
rect 51370 193008 51375 193064
rect 47494 193006 51375 193008
rect 51309 193003 51375 193006
rect 55038 192968 55098 193278
rect 88845 193202 88911 193205
rect 88845 193200 92052 193202
rect 88845 193144 88850 193200
rect 88906 193144 92052 193200
rect 88845 193142 92052 193144
rect 88845 193139 88911 193142
rect 119806 193066 119866 193308
rect 123069 193280 123074 193336
rect 123130 193280 127042 193336
rect 123069 193278 127042 193280
rect 123069 193275 123135 193278
rect 122977 193066 123043 193069
rect 119806 193064 123043 193066
rect 119806 193008 122982 193064
rect 123038 193008 123043 193064
rect 119806 193006 123043 193008
rect 122977 193003 123043 193006
rect 126982 192968 127042 193278
rect 160513 193336 163996 193338
rect 160513 193280 160518 193336
rect 160574 193280 163996 193336
rect 160513 193278 163996 193280
rect 160513 193275 160579 193278
rect 88477 192930 88543 192933
rect 160237 192930 160303 192933
rect 84876 192928 88543 192930
rect 84876 192872 88482 192928
rect 88538 192872 88543 192928
rect 84876 192870 88543 192872
rect 156820 192928 160303 192930
rect 156820 192872 160242 192928
rect 160298 192872 160303 192928
rect 156820 192870 160303 192872
rect 88477 192867 88543 192870
rect 160237 192867 160303 192870
rect 51493 192794 51559 192797
rect 123161 192794 123227 192797
rect 47524 192792 51559 192794
rect 47524 192736 51498 192792
rect 51554 192736 51559 192792
rect 47524 192734 51559 192736
rect 119836 192792 123227 192794
rect 119836 192736 123166 192792
rect 123222 192736 123227 192792
rect 119836 192734 123227 192736
rect 51493 192731 51559 192734
rect 123161 192731 123227 192734
rect 160145 192794 160211 192797
rect 160145 192792 163996 192794
rect 160145 192736 160150 192792
rect 160206 192736 163996 192792
rect 160145 192734 163996 192736
rect 160145 192731 160211 192734
rect 88385 192658 88451 192661
rect 88385 192656 92052 192658
rect 88385 192600 88390 192656
rect 88446 192600 92052 192656
rect 88385 192598 92052 192600
rect 88385 192595 88451 192598
rect 51585 192386 51651 192389
rect 51585 192384 51970 192386
rect 51585 192328 51590 192384
rect 51646 192328 51970 192384
rect 51585 192326 51970 192328
rect 51585 192323 51651 192326
rect 51677 192250 51743 192253
rect 47524 192248 51743 192250
rect 47524 192192 51682 192248
rect 51738 192192 51743 192248
rect 47524 192190 51743 192192
rect 51910 192250 51970 192326
rect 88293 192250 88359 192253
rect 51910 192190 55068 192250
rect 84876 192248 88359 192250
rect 84876 192192 88298 192248
rect 88354 192192 88359 192248
rect 123345 192250 123411 192253
rect 159961 192250 160027 192253
rect 123345 192248 127012 192250
rect 84876 192190 88359 192192
rect 51677 192187 51743 192190
rect 88293 192187 88359 192190
rect 51401 192114 51467 192117
rect 51401 192112 55098 192114
rect 51401 192056 51406 192112
rect 51462 192056 55098 192112
rect 51401 192054 55098 192056
rect 51401 192051 51467 192054
rect 55038 191744 55098 192054
rect 88569 191978 88635 191981
rect 119806 191978 119866 192220
rect 123345 192192 123350 192248
rect 123406 192192 127012 192248
rect 123345 192190 127012 192192
rect 156820 192248 160027 192250
rect 156820 192192 159966 192248
rect 160022 192192 160027 192248
rect 156820 192190 160027 192192
rect 123345 192187 123411 192190
rect 159961 192187 160027 192190
rect 160605 192250 160671 192253
rect 160605 192248 163996 192250
rect 160605 192192 160610 192248
rect 160666 192192 163996 192248
rect 160605 192190 163996 192192
rect 160605 192187 160671 192190
rect 123253 192114 123319 192117
rect 160053 192114 160119 192117
rect 123253 192112 127042 192114
rect 123253 192056 123258 192112
rect 123314 192056 127042 192112
rect 123253 192054 127042 192056
rect 123253 192051 123319 192054
rect 123253 191978 123319 191981
rect 88569 191976 92052 191978
rect 88569 191920 88574 191976
rect 88630 191920 92052 191976
rect 88569 191918 92052 191920
rect 119806 191976 123319 191978
rect 119806 191920 123258 191976
rect 123314 191920 123319 191976
rect 119806 191918 123319 191920
rect 88569 191915 88635 191918
rect 123253 191915 123319 191918
rect 126982 191744 127042 192054
rect 156790 192112 160119 192114
rect 156790 192056 160058 192112
rect 160114 192056 160119 192112
rect 156790 192054 160119 192056
rect 51401 191706 51467 191709
rect 88477 191706 88543 191709
rect 122149 191706 122215 191709
rect 47524 191704 51467 191706
rect 47524 191648 51406 191704
rect 51462 191648 51467 191704
rect 47524 191646 51467 191648
rect 84876 191704 88543 191706
rect 84876 191648 88482 191704
rect 88538 191648 88543 191704
rect 84876 191646 88543 191648
rect 119836 191704 122215 191706
rect 119836 191648 122154 191704
rect 122210 191648 122215 191704
rect 156790 191676 156850 192054
rect 160053 192051 160119 192054
rect 160053 191706 160119 191709
rect 160053 191704 163996 191706
rect 119836 191646 122215 191648
rect 51401 191643 51467 191646
rect 88477 191643 88543 191646
rect 122149 191643 122215 191646
rect 160053 191648 160058 191704
rect 160114 191648 163996 191704
rect 160053 191646 163996 191648
rect 160053 191643 160119 191646
rect 51309 191570 51375 191573
rect 123069 191570 123135 191573
rect 51309 191568 55098 191570
rect 51309 191512 51314 191568
rect 51370 191512 55098 191568
rect 51309 191510 55098 191512
rect 51309 191507 51375 191510
rect 55038 191200 55098 191510
rect 123069 191568 127042 191570
rect 123069 191512 123074 191568
rect 123130 191512 127042 191568
rect 123069 191510 127042 191512
rect 123069 191507 123135 191510
rect 88293 191434 88359 191437
rect 88293 191432 92052 191434
rect 88293 191376 88298 191432
rect 88354 191376 92052 191432
rect 88293 191374 92052 191376
rect 88293 191371 88359 191374
rect 126982 191200 127042 191510
rect 87189 191162 87255 191165
rect 160237 191162 160303 191165
rect 194737 191162 194803 191165
rect 84876 191160 87255 191162
rect 84876 191104 87194 191160
rect 87250 191104 87255 191160
rect 84876 191102 87255 191104
rect 156820 191160 160303 191162
rect 156820 191104 160242 191160
rect 160298 191104 160303 191160
rect 156820 191102 160303 191104
rect 191780 191160 194803 191162
rect 191780 191104 194742 191160
rect 194798 191104 194803 191160
rect 191780 191102 194803 191104
rect 87189 191099 87255 191102
rect 160237 191099 160303 191102
rect 194737 191099 194803 191102
rect 51585 191026 51651 191029
rect 122977 191026 123043 191029
rect 47524 191024 51651 191026
rect 47524 190968 51590 191024
rect 51646 190968 51651 191024
rect 47524 190966 51651 190968
rect 119836 191024 123043 191026
rect 119836 190968 122982 191024
rect 123038 190968 123043 191024
rect 119836 190966 123043 190968
rect 51585 190963 51651 190966
rect 122977 190963 123043 190966
rect 160237 191026 160303 191029
rect 160237 191024 163996 191026
rect 160237 190968 160242 191024
rect 160298 190968 163996 191024
rect 160237 190966 163996 190968
rect 160237 190963 160303 190966
rect 51493 190890 51559 190893
rect 88661 190890 88727 190893
rect 123161 190890 123227 190893
rect 160145 190890 160211 190893
rect 51493 190888 55098 190890
rect 51493 190832 51498 190888
rect 51554 190832 55098 190888
rect 51493 190830 55098 190832
rect 51493 190827 51559 190830
rect 55038 190520 55098 190830
rect 88661 190888 92052 190890
rect 88661 190832 88666 190888
rect 88722 190832 92052 190888
rect 88661 190830 92052 190832
rect 123161 190888 127042 190890
rect 123161 190832 123166 190888
rect 123222 190832 127042 190888
rect 123161 190830 127042 190832
rect 88661 190827 88727 190830
rect 123161 190827 123227 190830
rect 126982 190520 127042 190830
rect 156790 190888 160211 190890
rect 156790 190832 160150 190888
rect 160206 190832 160211 190888
rect 156790 190830 160211 190832
rect 51309 190482 51375 190485
rect 88385 190482 88451 190485
rect 123161 190482 123227 190485
rect 47524 190480 51375 190482
rect 47524 190424 51314 190480
rect 51370 190424 51375 190480
rect 47524 190422 51375 190424
rect 84876 190480 88451 190482
rect 84876 190424 88390 190480
rect 88446 190424 88451 190480
rect 84876 190422 88451 190424
rect 119836 190480 123227 190482
rect 119836 190424 123166 190480
rect 123222 190424 123227 190480
rect 156790 190452 156850 190830
rect 160145 190827 160211 190830
rect 160145 190482 160211 190485
rect 160145 190480 163996 190482
rect 119836 190422 123227 190424
rect 51309 190419 51375 190422
rect 88385 190419 88451 190422
rect 123161 190419 123227 190422
rect 160145 190424 160150 190480
rect 160206 190424 163996 190480
rect 160145 190422 163996 190424
rect 160145 190419 160211 190422
rect 51677 190346 51743 190349
rect 88385 190346 88451 190349
rect 123253 190346 123319 190349
rect 51677 190344 55098 190346
rect 51677 190288 51682 190344
rect 51738 190288 55098 190344
rect 51677 190286 55098 190288
rect 51677 190283 51743 190286
rect 55038 189976 55098 190286
rect 88385 190344 92052 190346
rect 88385 190288 88390 190344
rect 88446 190288 92052 190344
rect 88385 190286 92052 190288
rect 123253 190344 127042 190346
rect 123253 190288 123258 190344
rect 123314 190288 127042 190344
rect 123253 190286 127042 190288
rect 88385 190283 88451 190286
rect 123253 190283 123319 190286
rect 126982 189976 127042 190286
rect 51493 189938 51559 189941
rect 88477 189938 88543 189941
rect 123253 189938 123319 189941
rect 158949 189938 159015 189941
rect 47524 189936 51559 189938
rect 47524 189880 51498 189936
rect 51554 189880 51559 189936
rect 47524 189878 51559 189880
rect 84876 189936 88543 189938
rect 84876 189880 88482 189936
rect 88538 189880 88543 189936
rect 84876 189878 88543 189880
rect 119836 189936 123319 189938
rect 119836 189880 123258 189936
rect 123314 189880 123319 189936
rect 119836 189878 123319 189880
rect 156820 189936 159015 189938
rect 156820 189880 158954 189936
rect 159010 189880 159015 189936
rect 156820 189878 159015 189880
rect 51493 189875 51559 189878
rect 88477 189875 88543 189878
rect 123253 189875 123319 189878
rect 158949 189875 159015 189878
rect 88201 189802 88267 189805
rect 88201 189800 92052 189802
rect 88201 189744 88206 189800
rect 88262 189744 92052 189800
rect 88201 189742 92052 189744
rect 88201 189739 88267 189742
rect 159961 189666 160027 189669
rect 163966 189666 164026 189908
rect 159961 189664 164026 189666
rect 159961 189608 159966 189664
rect 160022 189608 164026 189664
rect 159961 189606 164026 189608
rect 159961 189603 160027 189606
rect 123345 189530 123411 189533
rect 123345 189528 127042 189530
rect 123345 189472 123350 189528
rect 123406 189472 127042 189528
rect 123345 189470 127042 189472
rect 123345 189467 123411 189470
rect 122977 189394 123043 189397
rect 119836 189392 123043 189394
rect 47494 189122 47554 189364
rect 119836 189336 122982 189392
rect 123038 189336 123043 189392
rect 119836 189334 123043 189336
rect 122977 189331 123043 189334
rect 126982 189296 127042 189470
rect 160329 189394 160395 189397
rect 160329 189392 163996 189394
rect 160329 189336 160334 189392
rect 160390 189336 163996 189392
rect 160329 189334 163996 189336
rect 160329 189331 160395 189334
rect 51401 189258 51467 189261
rect 88293 189258 88359 189261
rect 51401 189256 55068 189258
rect 51401 189200 51406 189256
rect 51462 189200 55068 189256
rect 51401 189198 55068 189200
rect 84876 189256 88359 189258
rect 84876 189200 88298 189256
rect 88354 189200 88359 189256
rect 84876 189198 88359 189200
rect 51401 189195 51467 189198
rect 88293 189195 88359 189198
rect 88753 189258 88819 189261
rect 160053 189258 160119 189261
rect 88753 189256 92052 189258
rect 88753 189200 88758 189256
rect 88814 189200 92052 189256
rect 88753 189198 92052 189200
rect 156820 189256 160119 189258
rect 156820 189200 160058 189256
rect 160114 189200 160119 189256
rect 156820 189198 160119 189200
rect 88753 189195 88819 189198
rect 160053 189195 160119 189198
rect 51401 189122 51467 189125
rect 47494 189120 51467 189122
rect 47494 189064 51406 189120
rect 51462 189064 51467 189120
rect 47494 189062 51467 189064
rect 51401 189059 51467 189062
rect 51585 189122 51651 189125
rect 123069 189122 123135 189125
rect 51585 189120 55098 189122
rect 51585 189064 51590 189120
rect 51646 189064 55098 189120
rect 51585 189062 55098 189064
rect 51585 189059 51651 189062
rect 9896 188986 10376 189016
rect 14693 188986 14759 188989
rect 9896 188984 14759 188986
rect 9896 188928 14698 188984
rect 14754 188928 14759 188984
rect 9896 188926 14759 188928
rect 9896 188896 10376 188926
rect 14693 188923 14759 188926
rect 51585 188850 51651 188853
rect 47524 188848 51651 188850
rect 47524 188792 51590 188848
rect 51646 188792 51651 188848
rect 47524 188790 51651 188792
rect 51585 188787 51651 188790
rect 55038 188752 55098 189062
rect 123069 189120 127042 189122
rect 123069 189064 123074 189120
rect 123130 189064 127042 189120
rect 123069 189062 127042 189064
rect 123069 189059 123135 189062
rect 121965 188850 122031 188853
rect 119836 188848 122031 188850
rect 119836 188792 121970 188848
rect 122026 188792 122031 188848
rect 119836 188790 122031 188792
rect 121965 188787 122031 188790
rect 126982 188752 127042 189062
rect 160053 188850 160119 188853
rect 160053 188848 163996 188850
rect 160053 188792 160058 188848
rect 160114 188792 163996 188848
rect 160053 188790 163996 188792
rect 160053 188787 160119 188790
rect 88477 188714 88543 188717
rect 84876 188712 88543 188714
rect 84876 188656 88482 188712
rect 88538 188656 88543 188712
rect 84876 188654 88543 188656
rect 88477 188651 88543 188654
rect 88661 188714 88727 188717
rect 160237 188714 160303 188717
rect 88661 188712 92052 188714
rect 88661 188656 88666 188712
rect 88722 188656 92052 188712
rect 88661 188654 92052 188656
rect 156820 188712 160303 188714
rect 156820 188656 160242 188712
rect 160298 188656 160303 188712
rect 156820 188654 160303 188656
rect 88661 188651 88727 188654
rect 160237 188651 160303 188654
rect 51309 188170 51375 188173
rect 88385 188170 88451 188173
rect 51309 188168 55068 188170
rect 47494 187898 47554 188140
rect 51309 188112 51314 188168
rect 51370 188112 55068 188168
rect 51309 188110 55068 188112
rect 84876 188168 88451 188170
rect 84876 188112 88390 188168
rect 88446 188112 88451 188168
rect 84876 188110 88451 188112
rect 51309 188107 51375 188110
rect 88385 188107 88451 188110
rect 88845 188170 88911 188173
rect 122977 188170 123043 188173
rect 88845 188168 92052 188170
rect 88845 188112 88850 188168
rect 88906 188112 92052 188168
rect 88845 188110 92052 188112
rect 119836 188168 123043 188170
rect 119836 188112 122982 188168
rect 123038 188112 123043 188168
rect 119836 188110 123043 188112
rect 88845 188107 88911 188110
rect 122977 188107 123043 188110
rect 123161 188170 123227 188173
rect 160145 188170 160211 188173
rect 123161 188168 127012 188170
rect 123161 188112 123166 188168
rect 123222 188112 127012 188168
rect 123161 188110 127012 188112
rect 156820 188168 160211 188170
rect 156820 188112 160150 188168
rect 160206 188112 160211 188168
rect 156820 188110 160211 188112
rect 123161 188107 123227 188110
rect 160145 188107 160211 188110
rect 160421 188170 160487 188173
rect 160421 188168 163996 188170
rect 160421 188112 160426 188168
rect 160482 188112 163996 188168
rect 160421 188110 163996 188112
rect 160421 188107 160487 188110
rect 51493 188034 51559 188037
rect 123253 188034 123319 188037
rect 51493 188032 55098 188034
rect 51493 187976 51498 188032
rect 51554 187976 55098 188032
rect 51493 187974 55098 187976
rect 51493 187971 51559 187974
rect 51309 187898 51375 187901
rect 47494 187896 51375 187898
rect 47494 187840 51314 187896
rect 51370 187840 51375 187896
rect 47494 187838 51375 187840
rect 51309 187835 51375 187838
rect 51493 187626 51559 187629
rect 47524 187624 51559 187626
rect 47524 187568 51498 187624
rect 51554 187568 51559 187624
rect 47524 187566 51559 187568
rect 51493 187563 51559 187566
rect 55038 187528 55098 187974
rect 123253 188032 127042 188034
rect 123253 187976 123258 188032
rect 123314 187976 127042 188032
rect 123253 187974 127042 187976
rect 123253 187971 123319 187974
rect 123529 187626 123595 187629
rect 119836 187624 123595 187626
rect 119836 187568 123534 187624
rect 123590 187568 123595 187624
rect 119836 187566 123595 187568
rect 123529 187563 123595 187566
rect 126982 187528 127042 187974
rect 160145 187626 160211 187629
rect 160145 187624 163996 187626
rect 160145 187568 160150 187624
rect 160206 187568 163996 187624
rect 160145 187566 163996 187568
rect 160145 187563 160211 187566
rect 88201 187490 88267 187493
rect 84876 187488 88267 187490
rect 84876 187432 88206 187488
rect 88262 187432 88267 187488
rect 84876 187430 88267 187432
rect 88201 187427 88267 187430
rect 88385 187490 88451 187493
rect 159961 187490 160027 187493
rect 88385 187488 92052 187490
rect 88385 187432 88390 187488
rect 88446 187432 92052 187488
rect 88385 187430 92052 187432
rect 156820 187488 160027 187490
rect 156820 187432 159966 187488
rect 160022 187432 160027 187488
rect 156820 187430 160027 187432
rect 88385 187427 88451 187430
rect 159961 187427 160027 187430
rect 51401 187354 51467 187357
rect 88477 187354 88543 187357
rect 51401 187352 55098 187354
rect 51401 187296 51406 187352
rect 51462 187296 55098 187352
rect 51401 187294 55098 187296
rect 51401 187291 51467 187294
rect 50665 187082 50731 187085
rect 47524 187080 50731 187082
rect 47524 187024 50670 187080
rect 50726 187024 50731 187080
rect 47524 187022 50731 187024
rect 50665 187019 50731 187022
rect 55038 186984 55098 187294
rect 84846 187352 88543 187354
rect 84846 187296 88482 187352
rect 88538 187296 88543 187352
rect 84846 187294 88543 187296
rect 84846 186916 84906 187294
rect 88477 187291 88543 187294
rect 123069 187354 123135 187357
rect 123069 187352 127042 187354
rect 123069 187296 123074 187352
rect 123130 187296 127042 187352
rect 123069 187294 127042 187296
rect 123069 187291 123135 187294
rect 122425 187082 122491 187085
rect 119836 187080 122491 187082
rect 119836 187024 122430 187080
rect 122486 187024 122491 187080
rect 119836 187022 122491 187024
rect 122425 187019 122491 187022
rect 126982 186984 127042 187294
rect 160973 187082 161039 187085
rect 160973 187080 163996 187082
rect 160973 187024 160978 187080
rect 161034 187024 163996 187080
rect 160973 187022 163996 187024
rect 160973 187019 161039 187022
rect 88569 186946 88635 186949
rect 160237 186946 160303 186949
rect 88569 186944 92052 186946
rect 88569 186888 88574 186944
rect 88630 186888 92052 186944
rect 88569 186886 92052 186888
rect 156820 186944 160303 186946
rect 156820 186888 160242 186944
rect 160298 186888 160303 186944
rect 156820 186886 160303 186888
rect 88569 186883 88635 186886
rect 160237 186883 160303 186886
rect 51585 186810 51651 186813
rect 123345 186810 123411 186813
rect 51585 186808 55098 186810
rect 51585 186752 51590 186808
rect 51646 186752 55098 186808
rect 51585 186750 55098 186752
rect 51585 186747 51651 186750
rect 51953 186538 52019 186541
rect 47524 186536 52019 186538
rect 47524 186480 51958 186536
rect 52014 186480 52019 186536
rect 47524 186478 52019 186480
rect 51953 186475 52019 186478
rect 55038 186304 55098 186750
rect 123345 186808 127042 186810
rect 123345 186752 123350 186808
rect 123406 186752 127042 186808
rect 123345 186750 127042 186752
rect 123345 186747 123411 186750
rect 122885 186538 122951 186541
rect 119836 186536 122951 186538
rect 119836 186480 122890 186536
rect 122946 186480 122951 186536
rect 119836 186478 122951 186480
rect 122885 186475 122951 186478
rect 88569 186402 88635 186405
rect 88569 186400 92052 186402
rect 88569 186344 88574 186400
rect 88630 186344 92052 186400
rect 88569 186342 92052 186344
rect 88569 186339 88635 186342
rect 126982 186304 127042 186750
rect 160513 186538 160579 186541
rect 160513 186536 163996 186538
rect 160513 186480 160518 186536
rect 160574 186480 163996 186536
rect 160513 186478 163996 186480
rect 160513 186475 160579 186478
rect 87189 186266 87255 186269
rect 160053 186266 160119 186269
rect 84876 186264 87255 186266
rect 84876 186208 87194 186264
rect 87250 186208 87255 186264
rect 84876 186206 87255 186208
rect 156820 186264 160119 186266
rect 156820 186208 160058 186264
rect 160114 186208 160119 186264
rect 156820 186206 160119 186208
rect 87189 186203 87255 186206
rect 160053 186203 160119 186206
rect 51309 186130 51375 186133
rect 123069 186130 123135 186133
rect 51309 186128 55098 186130
rect 51309 186072 51314 186128
rect 51370 186072 55098 186128
rect 51309 186070 55098 186072
rect 51309 186067 51375 186070
rect 49929 185994 49995 185997
rect 47524 185992 49995 185994
rect 47524 185936 49934 185992
rect 49990 185936 49995 185992
rect 47524 185934 49995 185936
rect 49929 185931 49995 185934
rect 55038 185760 55098 186070
rect 123069 186128 127042 186130
rect 123069 186072 123074 186128
rect 123130 186072 127042 186128
rect 123069 186070 127042 186072
rect 123069 186067 123135 186070
rect 122977 185994 123043 185997
rect 119836 185992 123043 185994
rect 119836 185936 122982 185992
rect 123038 185936 123043 185992
rect 119836 185934 123043 185936
rect 122977 185931 123043 185934
rect 88569 185858 88635 185861
rect 88569 185856 92052 185858
rect 88569 185800 88574 185856
rect 88630 185800 92052 185856
rect 88569 185798 92052 185800
rect 88569 185795 88635 185798
rect 126982 185760 127042 186070
rect 160605 185994 160671 185997
rect 160605 185992 163996 185994
rect 160605 185936 160610 185992
rect 160666 185936 163996 185992
rect 160605 185934 163996 185936
rect 160605 185931 160671 185934
rect 88477 185722 88543 185725
rect 160237 185722 160303 185725
rect 84876 185720 88543 185722
rect 84876 185664 88482 185720
rect 88538 185664 88543 185720
rect 84876 185662 88543 185664
rect 156820 185720 160303 185722
rect 156820 185664 160242 185720
rect 160298 185664 160303 185720
rect 156820 185662 160303 185664
rect 88477 185659 88543 185662
rect 160237 185659 160303 185662
rect 192069 185586 192135 185589
rect 191780 185584 192135 185586
rect 191780 185528 192074 185584
rect 192130 185528 192135 185584
rect 191780 185526 192135 185528
rect 192069 185523 192135 185526
rect 51493 185450 51559 185453
rect 198233 185450 198299 185453
rect 201416 185450 201896 185480
rect 51493 185448 55098 185450
rect 51493 185392 51498 185448
rect 51554 185392 55098 185448
rect 51493 185390 55098 185392
rect 51493 185387 51559 185390
rect 50205 185314 50271 185317
rect 47524 185312 50271 185314
rect 47524 185256 50210 185312
rect 50266 185256 50271 185312
rect 47524 185254 50271 185256
rect 50205 185251 50271 185254
rect 55038 185216 55098 185390
rect 198233 185448 201896 185450
rect 198233 185392 198238 185448
rect 198294 185392 201896 185448
rect 198233 185390 201896 185392
rect 198233 185387 198299 185390
rect 201416 185360 201896 185390
rect 88661 185314 88727 185317
rect 122885 185314 122951 185317
rect 88661 185312 92052 185314
rect 88661 185256 88666 185312
rect 88722 185256 92052 185312
rect 88661 185254 92052 185256
rect 119836 185312 122951 185314
rect 119836 185256 122890 185312
rect 122946 185256 122951 185312
rect 119836 185254 122951 185256
rect 88661 185251 88727 185254
rect 122885 185251 122951 185254
rect 160329 185314 160395 185317
rect 160329 185312 163996 185314
rect 160329 185256 160334 185312
rect 160390 185256 163996 185312
rect 160329 185254 163996 185256
rect 160329 185251 160395 185254
rect 88385 185178 88451 185181
rect 84876 185176 88451 185178
rect 84876 185120 88390 185176
rect 88446 185120 88451 185176
rect 84876 185118 88451 185120
rect 88385 185115 88451 185118
rect 123529 185178 123595 185181
rect 160145 185178 160211 185181
rect 123529 185176 127012 185178
rect 123529 185120 123534 185176
rect 123590 185120 127012 185176
rect 123529 185118 127012 185120
rect 156820 185176 160211 185178
rect 156820 185120 160150 185176
rect 160206 185120 160211 185176
rect 156820 185118 160211 185120
rect 123529 185115 123595 185118
rect 160145 185115 160211 185118
rect 81710 184980 81716 185044
rect 81780 185042 81786 185044
rect 82221 185042 82287 185045
rect 81780 185040 82287 185042
rect 81780 184984 82226 185040
rect 82282 184984 82287 185040
rect 81780 184982 82287 184984
rect 81780 184980 81786 184982
rect 82221 184979 82287 184982
rect 153470 184980 153476 185044
rect 153540 185042 153546 185044
rect 154349 185042 154415 185045
rect 153540 185040 154415 185042
rect 153540 184984 154354 185040
rect 154410 184984 154415 185040
rect 153540 184982 154415 184984
rect 153540 184980 153546 184982
rect 154349 184979 154415 184982
rect 50113 184770 50179 184773
rect 47524 184768 50179 184770
rect 47524 184712 50118 184768
rect 50174 184712 50179 184768
rect 47524 184710 50179 184712
rect 50113 184707 50179 184710
rect 89213 184770 89279 184773
rect 122333 184770 122399 184773
rect 89213 184768 92052 184770
rect 89213 184712 89218 184768
rect 89274 184712 92052 184768
rect 89213 184710 92052 184712
rect 119836 184768 122399 184770
rect 119836 184712 122338 184768
rect 122394 184712 122399 184768
rect 119836 184710 122399 184712
rect 89213 184707 89279 184710
rect 122333 184707 122399 184710
rect 161249 184770 161315 184773
rect 161249 184768 163996 184770
rect 161249 184712 161254 184768
rect 161310 184712 163996 184768
rect 161249 184710 163996 184712
rect 161249 184707 161315 184710
rect 50021 184226 50087 184229
rect 47524 184224 50087 184226
rect 47524 184168 50026 184224
rect 50082 184168 50087 184224
rect 47524 184166 50087 184168
rect 50021 184163 50087 184166
rect 88569 184226 88635 184229
rect 122977 184226 123043 184229
rect 88569 184224 92052 184226
rect 88569 184168 88574 184224
rect 88630 184168 92052 184224
rect 88569 184166 92052 184168
rect 119836 184224 123043 184226
rect 119836 184168 122982 184224
rect 123038 184168 123043 184224
rect 119836 184166 123043 184168
rect 88569 184163 88635 184166
rect 122977 184163 123043 184166
rect 161065 184226 161131 184229
rect 161065 184224 163996 184226
rect 161065 184168 161070 184224
rect 161126 184168 163996 184224
rect 161065 184166 163996 184168
rect 161065 184163 161131 184166
rect 51309 183682 51375 183685
rect 47524 183680 51375 183682
rect 47524 183624 51314 183680
rect 51370 183624 51375 183680
rect 47524 183622 51375 183624
rect 51309 183619 51375 183622
rect 87833 183682 87899 183685
rect 123069 183682 123135 183685
rect 87833 183680 92052 183682
rect 87833 183624 87838 183680
rect 87894 183624 92052 183680
rect 87833 183622 92052 183624
rect 119836 183680 123135 183682
rect 119836 183624 123074 183680
rect 123130 183624 123135 183680
rect 119836 183622 123135 183624
rect 87833 183619 87899 183622
rect 123069 183619 123135 183622
rect 159593 183682 159659 183685
rect 159593 183680 163996 183682
rect 159593 183624 159598 183680
rect 159654 183624 163996 183680
rect 159593 183622 163996 183624
rect 159593 183619 159659 183622
rect 49929 183138 49995 183141
rect 47524 183136 49995 183138
rect 47524 183080 49934 183136
rect 49990 183080 49995 183136
rect 47524 183078 49995 183080
rect 49929 183075 49995 183078
rect 88569 183138 88635 183141
rect 122149 183138 122215 183141
rect 88569 183136 92052 183138
rect 88569 183080 88574 183136
rect 88630 183080 92052 183136
rect 88569 183078 92052 183080
rect 119836 183136 122215 183138
rect 119836 183080 122154 183136
rect 122210 183080 122215 183136
rect 119836 183078 122215 183080
rect 88569 183075 88635 183078
rect 122149 183075 122215 183078
rect 160329 183138 160395 183141
rect 160329 183136 163996 183138
rect 160329 183080 160334 183136
rect 160390 183080 163996 183136
rect 160329 183078 163996 183080
rect 160329 183075 160395 183078
rect 20213 180554 20279 180557
rect 40310 180554 40316 180556
rect 20213 180552 40316 180554
rect 20213 180496 20218 180552
rect 20274 180496 40316 180552
rect 20213 180494 40316 180496
rect 20213 180491 20279 180494
rect 40310 180492 40316 180494
rect 40380 180492 40386 180556
rect 77161 177290 77227 177293
rect 89070 177290 89076 177292
rect 77161 177288 89076 177290
rect 77161 177232 77166 177288
rect 77222 177232 89076 177288
rect 77161 177230 89076 177232
rect 77161 177227 77227 177230
rect 89070 177228 89076 177230
rect 89140 177228 89146 177292
rect 138750 177228 138756 177292
rect 138820 177290 138826 177292
rect 148829 177290 148895 177293
rect 138820 177288 148895 177290
rect 138820 177232 148834 177288
rect 148890 177232 148895 177288
rect 138820 177230 148895 177232
rect 138820 177228 138826 177230
rect 148829 177227 148895 177230
rect 92617 175250 92683 175253
rect 163181 175250 163247 175253
rect 89844 175248 92683 175250
rect 89844 175192 92622 175248
rect 92678 175192 92683 175248
rect 89844 175190 92683 175192
rect 161788 175248 163247 175250
rect 161788 175192 163186 175248
rect 163242 175192 163247 175248
rect 161788 175190 163247 175192
rect 92617 175187 92683 175190
rect 163181 175187 163247 175190
rect 168517 174842 168583 174845
rect 168517 174840 170068 174842
rect 168517 174784 168522 174840
rect 168578 174784 170068 174840
rect 168517 174782 170068 174784
rect 168517 174779 168583 174782
rect 94549 174570 94615 174573
rect 94549 174568 97940 174570
rect 94549 174512 94554 174568
rect 94610 174512 97940 174568
rect 94549 174510 97940 174512
rect 94549 174507 94615 174510
rect 92341 174026 92407 174029
rect 164377 174026 164443 174029
rect 89844 174024 92407 174026
rect 89844 173968 92346 174024
rect 92402 173968 92407 174024
rect 89844 173966 92407 173968
rect 161788 174024 164443 174026
rect 161788 173968 164382 174024
rect 164438 173968 164443 174024
rect 161788 173966 164443 173968
rect 92341 173963 92407 173966
rect 164377 173963 164443 173966
rect 92157 172802 92223 172805
rect 164285 172802 164351 172805
rect 89844 172800 92223 172802
rect 89844 172744 92162 172800
rect 92218 172744 92223 172800
rect 89844 172742 92223 172744
rect 161788 172800 164351 172802
rect 161788 172744 164290 172800
rect 164346 172744 164351 172800
rect 161788 172742 164351 172744
rect 92157 172739 92223 172742
rect 164285 172739 164351 172742
rect 95009 172258 95075 172261
rect 95009 172256 97940 172258
rect 95009 172200 95014 172256
rect 95070 172200 97940 172256
rect 95009 172198 97940 172200
rect 95009 172195 95075 172198
rect 168374 172060 168380 172124
rect 168444 172122 168450 172124
rect 170038 172122 170098 172704
rect 188021 172530 188087 172533
rect 185892 172528 188087 172530
rect 185892 172472 188026 172528
rect 188082 172472 188087 172528
rect 185892 172470 188087 172472
rect 188021 172467 188087 172470
rect 168444 172062 170098 172122
rect 168444 172060 168450 172062
rect 23566 171788 23572 171852
rect 23636 171850 23642 171852
rect 45053 171850 45119 171853
rect 23636 171790 25996 171850
rect 41820 171848 45119 171850
rect 41820 171792 45058 171848
rect 45114 171792 45119 171848
rect 41820 171790 45119 171792
rect 23636 171788 23642 171790
rect 45053 171787 45119 171790
rect 92249 171578 92315 171581
rect 164009 171578 164075 171581
rect 89844 171576 92315 171578
rect 89844 171520 92254 171576
rect 92310 171520 92315 171576
rect 89844 171518 92315 171520
rect 161788 171576 164075 171578
rect 161788 171520 164014 171576
rect 164070 171520 164075 171576
rect 161788 171518 164075 171520
rect 92249 171515 92315 171518
rect 164009 171515 164075 171518
rect 167505 170490 167571 170493
rect 170038 170490 170098 170664
rect 167505 170488 170098 170490
rect 167505 170432 167510 170488
rect 167566 170432 170098 170488
rect 167505 170430 170098 170432
rect 167505 170427 167571 170430
rect 92065 170354 92131 170357
rect 163365 170354 163431 170357
rect 89844 170352 92131 170354
rect 89844 170296 92070 170352
rect 92126 170296 92131 170352
rect 89844 170294 92131 170296
rect 161788 170352 163431 170354
rect 161788 170296 163370 170352
rect 163426 170296 163431 170352
rect 161788 170294 163431 170296
rect 92065 170291 92131 170294
rect 163365 170291 163431 170294
rect 94825 169946 94891 169949
rect 94825 169944 97940 169946
rect 94825 169888 94830 169944
rect 94886 169888 97940 169944
rect 94825 169886 97940 169888
rect 94825 169883 94891 169886
rect 48457 169266 48523 169269
rect 48457 169264 49916 169266
rect 48457 169208 48462 169264
rect 48518 169208 49916 169264
rect 48457 169206 49916 169208
rect 48457 169203 48523 169206
rect 91973 169130 92039 169133
rect 89844 169128 92039 169130
rect 89844 169072 91978 169128
rect 92034 169072 92039 169128
rect 89844 169070 92039 169072
rect 91973 169067 92039 169070
rect 118929 168994 118995 168997
rect 122014 168994 122074 169168
rect 163181 169130 163247 169133
rect 161788 169128 163247 169130
rect 161788 169072 163186 169128
rect 163242 169072 163247 169128
rect 161788 169070 163247 169072
rect 163181 169067 163247 169070
rect 118929 168992 122074 168994
rect 118929 168936 118934 168992
rect 118990 168936 122074 168992
rect 118929 168934 122074 168936
rect 118929 168931 118995 168934
rect 167321 168178 167387 168181
rect 170038 168178 170098 168760
rect 167321 168176 170098 168178
rect 167321 168120 167326 168176
rect 167382 168120 170098 168176
rect 167321 168118 170098 168120
rect 167321 168115 167387 168118
rect 91421 167906 91487 167909
rect 164377 167906 164443 167909
rect 89844 167904 91487 167906
rect 89844 167848 91426 167904
rect 91482 167848 91487 167904
rect 89844 167846 91487 167848
rect 161788 167904 164443 167906
rect 161788 167848 164382 167904
rect 164438 167848 164443 167904
rect 161788 167846 164443 167848
rect 91421 167843 91487 167846
rect 164377 167843 164443 167846
rect 9896 167770 10376 167800
rect 13313 167770 13379 167773
rect 9896 167768 13379 167770
rect 9896 167712 13318 167768
rect 13374 167712 13379 167768
rect 9896 167710 13379 167712
rect 9896 167680 10376 167710
rect 13313 167707 13379 167710
rect 95377 167498 95443 167501
rect 95377 167496 97940 167498
rect 95377 167440 95382 167496
rect 95438 167440 97940 167496
rect 95377 167438 97940 167440
rect 95377 167435 95443 167438
rect 91329 166682 91395 166685
rect 163273 166682 163339 166685
rect 89844 166680 91395 166682
rect 89844 166624 91334 166680
rect 91390 166624 91395 166680
rect 89844 166622 91395 166624
rect 161788 166680 163339 166682
rect 161788 166624 163278 166680
rect 163334 166624 163339 166680
rect 161788 166622 163339 166624
rect 91329 166619 91395 166622
rect 163273 166619 163339 166622
rect 167229 166274 167295 166277
rect 170038 166274 170098 166720
rect 167229 166272 170098 166274
rect 167229 166216 167234 166272
rect 167290 166216 170098 166272
rect 167229 166214 170098 166216
rect 167229 166211 167295 166214
rect 188021 165866 188087 165869
rect 185892 165864 188087 165866
rect 185892 165808 188026 165864
rect 188082 165808 188087 165864
rect 185892 165806 188087 165808
rect 188021 165803 188087 165806
rect 91973 165458 92039 165461
rect 89844 165456 92039 165458
rect 89844 165400 91978 165456
rect 92034 165400 92039 165456
rect 89844 165398 92039 165400
rect 91973 165395 92039 165398
rect 94181 165186 94247 165189
rect 113734 165186 113794 165768
rect 163181 165458 163247 165461
rect 161788 165456 163247 165458
rect 161788 165400 163186 165456
rect 163242 165400 163247 165456
rect 161788 165398 163247 165400
rect 163181 165395 163247 165398
rect 116537 165186 116603 165189
rect 94181 165184 97940 165186
rect 94181 165128 94186 165184
rect 94242 165128 97940 165184
rect 94181 165126 97940 165128
rect 113734 165184 116603 165186
rect 113734 165128 116542 165184
rect 116598 165128 116603 165184
rect 113734 165126 116603 165128
rect 94181 165123 94247 165126
rect 116537 165123 116603 165126
rect 41598 164172 41604 164236
rect 41668 164172 41674 164236
rect 92617 164234 92683 164237
rect 164285 164234 164351 164237
rect 89844 164232 92683 164234
rect 89844 164176 92622 164232
rect 92678 164176 92683 164232
rect 89844 164174 92683 164176
rect 161788 164232 164351 164234
rect 161788 164176 164290 164232
rect 164346 164176 164351 164232
rect 161788 164174 164351 164176
rect 22237 163826 22303 163829
rect 22237 163824 25996 163826
rect 22237 163768 22242 163824
rect 22298 163768 25996 163824
rect 41606 163796 41666 164172
rect 92617 164171 92683 164174
rect 164285 164171 164351 164174
rect 167965 164098 168031 164101
rect 170038 164098 170098 164680
rect 167965 164096 170098 164098
rect 167965 164040 167970 164096
rect 168026 164040 170098 164096
rect 167965 164038 170098 164040
rect 167965 164035 168031 164038
rect 22237 163766 25996 163768
rect 22237 163763 22303 163766
rect 91697 163146 91763 163149
rect 164285 163146 164351 163149
rect 89844 163144 91763 163146
rect 89844 163088 91702 163144
rect 91758 163088 91763 163144
rect 89844 163086 91763 163088
rect 161788 163144 164351 163146
rect 161788 163088 164290 163144
rect 164346 163088 164351 163144
rect 161788 163086 164351 163088
rect 91697 163083 91763 163086
rect 164285 163083 164351 163086
rect 94089 162874 94155 162877
rect 94089 162872 97940 162874
rect 94089 162816 94094 162872
rect 94150 162816 97940 162872
rect 94089 162814 97940 162816
rect 94089 162811 94155 162814
rect 168425 162194 168491 162197
rect 170038 162194 170098 162776
rect 168425 162192 170098 162194
rect 168425 162136 168430 162192
rect 168486 162136 170098 162192
rect 168425 162134 170098 162136
rect 168425 162131 168491 162134
rect 92617 161922 92683 161925
rect 164285 161922 164351 161925
rect 89844 161920 92683 161922
rect 89844 161864 92622 161920
rect 92678 161864 92683 161920
rect 89844 161862 92683 161864
rect 161788 161920 164351 161922
rect 161788 161864 164290 161920
rect 164346 161864 164351 161920
rect 161788 161862 164351 161864
rect 92617 161859 92683 161862
rect 164285 161859 164351 161862
rect 197589 161922 197655 161925
rect 201416 161922 201896 161952
rect 197589 161920 201896 161922
rect 197589 161864 197594 161920
rect 197650 161864 201896 161920
rect 197589 161862 201896 161864
rect 197589 161859 197655 161862
rect 201416 161832 201896 161862
rect 168517 160834 168583 160837
rect 168517 160832 170068 160834
rect 168517 160776 168522 160832
rect 168578 160776 170068 160832
rect 168517 160774 170068 160776
rect 168517 160771 168583 160774
rect 91973 160698 92039 160701
rect 164377 160698 164443 160701
rect 89844 160696 92039 160698
rect 89844 160640 91978 160696
rect 92034 160640 92039 160696
rect 89844 160638 92039 160640
rect 161788 160696 164443 160698
rect 161788 160640 164382 160696
rect 164438 160640 164443 160696
rect 161788 160638 164443 160640
rect 91973 160635 92039 160638
rect 164377 160635 164443 160638
rect 93997 160426 94063 160429
rect 93997 160424 97940 160426
rect 93997 160368 94002 160424
rect 94058 160368 97940 160424
rect 93997 160366 97940 160368
rect 93997 160363 94063 160366
rect 91973 159474 92039 159477
rect 164285 159474 164351 159477
rect 89844 159472 92039 159474
rect 89844 159416 91978 159472
rect 92034 159416 92039 159472
rect 89844 159414 92039 159416
rect 161788 159472 164351 159474
rect 161788 159416 164290 159472
rect 164346 159416 164351 159472
rect 161788 159414 164351 159416
rect 91973 159411 92039 159414
rect 164285 159411 164351 159414
rect 191190 159202 191196 159204
rect 185892 159142 191196 159202
rect 191190 159140 191196 159142
rect 191260 159140 191266 159204
rect 168517 158522 168583 158525
rect 170038 158522 170098 158696
rect 168517 158520 170098 158522
rect 168517 158464 168522 158520
rect 168578 158464 170098 158520
rect 168517 158462 170098 158464
rect 168517 158459 168583 158462
rect 91973 158250 92039 158253
rect 164285 158250 164351 158253
rect 89844 158248 92039 158250
rect 89844 158192 91978 158248
rect 92034 158192 92039 158248
rect 89844 158190 92039 158192
rect 161788 158248 164351 158250
rect 161788 158192 164290 158248
rect 164346 158192 164351 158248
rect 161788 158190 164351 158192
rect 91973 158187 92039 158190
rect 164285 158187 164351 158190
rect 93997 158114 94063 158117
rect 93997 158112 97940 158114
rect 93997 158056 94002 158112
rect 94058 158056 97940 158112
rect 93997 158054 97940 158056
rect 93997 158051 94063 158054
rect 91789 157026 91855 157029
rect 164285 157026 164351 157029
rect 89844 157024 91855 157026
rect 89844 156968 91794 157024
rect 91850 156968 91855 157024
rect 89844 156966 91855 156968
rect 161788 157024 164351 157026
rect 161788 156968 164290 157024
rect 164346 156968 164351 157024
rect 161788 156966 164351 156968
rect 91789 156963 91855 156966
rect 164285 156963 164351 156966
rect 168517 156890 168583 156893
rect 168517 156888 170068 156890
rect 168517 156832 168522 156888
rect 168578 156832 170068 156888
rect 168517 156830 170068 156832
rect 168517 156827 168583 156830
rect 47813 155938 47879 155941
rect 119573 155938 119639 155941
rect 47813 155936 49916 155938
rect 47813 155880 47818 155936
rect 47874 155880 49916 155936
rect 47813 155878 49916 155880
rect 119573 155936 122044 155938
rect 119573 155880 119578 155936
rect 119634 155880 122044 155936
rect 119573 155878 122044 155880
rect 47813 155875 47879 155878
rect 119573 155875 119639 155878
rect 22329 155802 22395 155805
rect 44358 155802 44364 155804
rect 22329 155800 25996 155802
rect 22329 155744 22334 155800
rect 22390 155744 25996 155800
rect 22329 155742 25996 155744
rect 41820 155742 44364 155802
rect 22329 155739 22395 155742
rect 44358 155740 44364 155742
rect 44428 155740 44434 155804
rect 164377 155802 164443 155805
rect 161788 155800 164443 155802
rect 89814 155258 89874 155772
rect 97910 155258 97970 155772
rect 161788 155744 164382 155800
rect 164438 155744 164443 155800
rect 161788 155742 164443 155744
rect 164377 155739 164443 155742
rect 89814 155198 97970 155258
rect 167137 154850 167203 154853
rect 167137 154848 170068 154850
rect 167137 154792 167142 154848
rect 167198 154792 170068 154848
rect 167137 154790 170068 154792
rect 167137 154787 167203 154790
rect 91421 154578 91487 154581
rect 163365 154578 163431 154581
rect 89844 154576 91487 154578
rect 89844 154520 91426 154576
rect 91482 154520 91487 154576
rect 89844 154518 91487 154520
rect 161788 154576 163431 154578
rect 161788 154520 163370 154576
rect 163426 154520 163431 154576
rect 161788 154518 163431 154520
rect 91421 154515 91487 154518
rect 163365 154515 163431 154518
rect 94733 153490 94799 153493
rect 94733 153488 97940 153490
rect 94733 153432 94738 153488
rect 94794 153432 97940 153488
rect 94733 153430 97940 153432
rect 94733 153427 94799 153430
rect 91789 153354 91855 153357
rect 164377 153354 164443 153357
rect 89844 153352 91855 153354
rect 89844 153296 91794 153352
rect 91850 153296 91855 153352
rect 89844 153294 91855 153296
rect 161788 153352 164443 153354
rect 161788 153296 164382 153352
rect 164438 153296 164443 153352
rect 161788 153294 164443 153296
rect 91789 153291 91855 153294
rect 164377 153291 164443 153294
rect 167137 152810 167203 152813
rect 167137 152808 170068 152810
rect 167137 152752 167142 152808
rect 167198 152752 170068 152808
rect 167137 152750 170068 152752
rect 167137 152747 167203 152750
rect 186038 152538 186044 152540
rect 185892 152478 186044 152538
rect 186038 152476 186044 152478
rect 186108 152476 186114 152540
rect 91697 152130 91763 152133
rect 164377 152130 164443 152133
rect 89844 152128 91763 152130
rect 89844 152072 91702 152128
rect 91758 152072 91763 152128
rect 89844 152070 91763 152072
rect 161788 152128 164443 152130
rect 161788 152072 164382 152128
rect 164438 152072 164443 152128
rect 161788 152070 164443 152072
rect 91697 152067 91763 152070
rect 164377 152067 164443 152070
rect 95377 151042 95443 151045
rect 95377 151040 97940 151042
rect 95377 150984 95382 151040
rect 95438 150984 97940 151040
rect 95377 150982 97940 150984
rect 95377 150979 95443 150982
rect 91421 150906 91487 150909
rect 163917 150906 163983 150909
rect 89844 150904 91487 150906
rect 89844 150848 91426 150904
rect 91482 150848 91487 150904
rect 89844 150846 91487 150848
rect 161788 150904 163983 150906
rect 161788 150848 163922 150904
rect 163978 150848 163983 150904
rect 161788 150846 163983 150848
rect 91421 150843 91487 150846
rect 163917 150843 163983 150846
rect 167229 150770 167295 150773
rect 167229 150768 170068 150770
rect 167229 150712 167234 150768
rect 167290 150712 170068 150768
rect 167229 150710 170068 150712
rect 167229 150707 167295 150710
rect 91329 149818 91395 149821
rect 164377 149818 164443 149821
rect 89844 149816 91395 149818
rect 89844 149760 91334 149816
rect 91390 149760 91395 149816
rect 89844 149758 91395 149760
rect 161788 149816 164443 149818
rect 161788 149760 164382 149816
rect 164438 149760 164443 149816
rect 161788 149758 164443 149760
rect 91329 149755 91395 149758
rect 164377 149755 164443 149758
rect 167321 148866 167387 148869
rect 167321 148864 170068 148866
rect 167321 148808 167326 148864
rect 167382 148808 170068 148864
rect 167321 148806 170068 148808
rect 167321 148803 167387 148806
rect 94181 148730 94247 148733
rect 94181 148728 97940 148730
rect 94181 148672 94186 148728
rect 94242 148672 97940 148728
rect 94181 148670 97940 148672
rect 94181 148667 94247 148670
rect 91697 148594 91763 148597
rect 164377 148594 164443 148597
rect 89844 148592 91763 148594
rect 89844 148536 91702 148592
rect 91758 148536 91763 148592
rect 89844 148534 91763 148536
rect 161788 148592 164443 148594
rect 161788 148536 164382 148592
rect 164438 148536 164443 148592
rect 161788 148534 164443 148536
rect 91697 148531 91763 148534
rect 164377 148531 164443 148534
rect 22329 147778 22395 147781
rect 45789 147778 45855 147781
rect 22329 147776 25996 147778
rect 22329 147720 22334 147776
rect 22390 147720 25996 147776
rect 22329 147718 25996 147720
rect 41820 147776 45855 147778
rect 41820 147720 45794 147776
rect 45850 147720 45855 147776
rect 41820 147718 45855 147720
rect 22329 147715 22395 147718
rect 45789 147715 45855 147718
rect 91421 147370 91487 147373
rect 164377 147370 164443 147373
rect 89844 147368 91487 147370
rect 89844 147312 91426 147368
rect 91482 147312 91487 147368
rect 89844 147310 91487 147312
rect 161788 147368 164443 147370
rect 161788 147312 164382 147368
rect 164438 147312 164443 147368
rect 161788 147310 164443 147312
rect 91421 147307 91487 147310
rect 164377 147307 164443 147310
rect 167229 146826 167295 146829
rect 167229 146824 170068 146826
rect 167229 146768 167234 146824
rect 167290 146768 170068 146824
rect 167229 146766 170068 146768
rect 167229 146763 167295 146766
rect 9896 146554 10376 146584
rect 13405 146554 13471 146557
rect 9896 146552 13471 146554
rect 9896 146496 13410 146552
rect 13466 146496 13471 146552
rect 9896 146494 13471 146496
rect 9896 146464 10376 146494
rect 13405 146491 13471 146494
rect 93353 146146 93419 146149
rect 89844 146144 93419 146146
rect 89844 146088 93358 146144
rect 93414 146088 93419 146144
rect 89844 146086 93419 146088
rect 93353 146083 93419 146086
rect 93997 145602 94063 145605
rect 97910 145602 97970 146388
rect 164377 146146 164443 146149
rect 161788 146144 164443 146146
rect 161788 146088 164382 146144
rect 164438 146088 164443 146144
rect 161788 146086 164443 146088
rect 164377 146083 164443 146086
rect 190638 145874 190644 145876
rect 185892 145814 190644 145874
rect 190638 145812 190644 145814
rect 190708 145812 190714 145876
rect 93997 145600 97970 145602
rect 93997 145544 94002 145600
rect 94058 145544 97970 145600
rect 93997 145542 97970 145544
rect 113734 145602 113794 145776
rect 116813 145602 116879 145605
rect 113734 145600 116879 145602
rect 113734 145544 116818 145600
rect 116874 145544 116879 145600
rect 113734 145542 116879 145544
rect 93997 145539 94063 145542
rect 116813 145539 116879 145542
rect 91973 144922 92039 144925
rect 163733 144922 163799 144925
rect 89844 144920 92039 144922
rect 89844 144864 91978 144920
rect 92034 144864 92039 144920
rect 89844 144862 92039 144864
rect 161788 144920 163799 144922
rect 161788 144864 163738 144920
rect 163794 144864 163799 144920
rect 161788 144862 163799 144864
rect 91973 144859 92039 144862
rect 163733 144859 163799 144862
rect 167137 144786 167203 144789
rect 167137 144784 170068 144786
rect 167137 144728 167142 144784
rect 167198 144728 170068 144784
rect 167137 144726 170068 144728
rect 167137 144723 167203 144726
rect 94365 143970 94431 143973
rect 94365 143968 97940 143970
rect 94365 143912 94370 143968
rect 94426 143912 97940 143968
rect 94365 143910 97940 143912
rect 94365 143907 94431 143910
rect 91789 143698 91855 143701
rect 163825 143698 163891 143701
rect 89844 143696 91855 143698
rect 89844 143640 91794 143696
rect 91850 143640 91855 143696
rect 89844 143638 91855 143640
rect 161788 143696 163891 143698
rect 161788 143640 163830 143696
rect 163886 143640 163891 143696
rect 161788 143638 163891 143640
rect 91789 143635 91855 143638
rect 163825 143635 163891 143638
rect 167045 142882 167111 142885
rect 167045 142880 170068 142882
rect 167045 142824 167050 142880
rect 167106 142824 170068 142880
rect 167045 142822 170068 142824
rect 167045 142819 167111 142822
rect 45789 142610 45855 142613
rect 116813 142612 116879 142613
rect 46382 142610 46388 142612
rect 45789 142608 46388 142610
rect 45789 142552 45794 142608
rect 45850 142552 46388 142608
rect 45789 142550 46388 142552
rect 45789 142547 45855 142550
rect 46382 142548 46388 142550
rect 46452 142610 46458 142612
rect 46452 142550 49916 142610
rect 116813 142608 116860 142612
rect 116924 142610 116930 142612
rect 118929 142610 118995 142613
rect 116813 142552 116818 142608
rect 46452 142548 46458 142550
rect 116813 142548 116860 142552
rect 116924 142550 116970 142610
rect 118929 142608 122044 142610
rect 118929 142552 118934 142608
rect 118990 142552 122044 142608
rect 118929 142550 122044 142552
rect 116924 142548 116930 142550
rect 116813 142547 116879 142548
rect 118929 142547 118995 142550
rect 91789 142474 91855 142477
rect 164377 142474 164443 142477
rect 89844 142472 91855 142474
rect 89844 142416 91794 142472
rect 91850 142416 91855 142472
rect 89844 142414 91855 142416
rect 161788 142472 164443 142474
rect 161788 142416 164382 142472
rect 164438 142416 164443 142472
rect 161788 142414 164443 142416
rect 91789 142411 91855 142414
rect 164377 142411 164443 142414
rect 89622 141732 89628 141796
rect 89692 141794 89698 141796
rect 91697 141794 91763 141797
rect 89692 141792 91763 141794
rect 89692 141736 91702 141792
rect 91758 141736 91763 141792
rect 89692 141734 91763 141736
rect 89692 141732 89698 141734
rect 91697 141731 91763 141734
rect 95377 141658 95443 141661
rect 95377 141656 97940 141658
rect 95377 141600 95382 141656
rect 95438 141600 97940 141656
rect 95377 141598 97940 141600
rect 95377 141595 95443 141598
rect 92525 141250 92591 141253
rect 164285 141250 164351 141253
rect 89844 141248 92591 141250
rect 89844 141192 92530 141248
rect 92586 141192 92591 141248
rect 89844 141190 92591 141192
rect 161788 141248 164351 141250
rect 161788 141192 164290 141248
rect 164346 141192 164351 141248
rect 161788 141190 164351 141192
rect 92525 141187 92591 141190
rect 164285 141187 164351 141190
rect 167873 140842 167939 140845
rect 167873 140840 170068 140842
rect 167873 140784 167878 140840
rect 167934 140784 170068 140840
rect 167873 140782 170068 140784
rect 167873 140779 167939 140782
rect 26142 140372 26148 140436
rect 26212 140372 26218 140436
rect 26150 139860 26210 140372
rect 92617 140026 92683 140029
rect 164377 140026 164443 140029
rect 89844 140024 92683 140026
rect 89844 139968 92622 140024
rect 92678 139968 92683 140024
rect 89844 139966 92683 139968
rect 161788 140024 164443 140026
rect 161788 139968 164382 140024
rect 164438 139968 164443 140024
rect 161788 139966 164443 139968
rect 92617 139963 92683 139966
rect 164377 139963 164443 139966
rect 44409 139890 44475 139893
rect 41820 139888 44475 139890
rect 41820 139832 44414 139888
rect 44470 139832 44475 139888
rect 41820 139830 44475 139832
rect 44409 139827 44475 139830
rect 93261 138802 93327 138805
rect 89844 138800 93327 138802
rect 89844 138744 93266 138800
rect 93322 138744 93327 138800
rect 89844 138742 93327 138744
rect 93261 138739 93327 138742
rect 93537 138666 93603 138669
rect 97910 138666 97970 139316
rect 188021 139210 188087 139213
rect 185892 139208 188087 139210
rect 185892 139152 188026 139208
rect 188082 139152 188087 139208
rect 185892 139150 188087 139152
rect 188021 139147 188087 139150
rect 163917 138802 163983 138805
rect 161788 138800 163983 138802
rect 161788 138744 163922 138800
rect 163978 138744 163983 138800
rect 161788 138742 163983 138744
rect 163917 138739 163983 138742
rect 167965 138802 168031 138805
rect 167965 138800 170068 138802
rect 167965 138744 167970 138800
rect 168026 138744 170068 138800
rect 167965 138742 170068 138744
rect 167965 138739 168031 138742
rect 93537 138664 97970 138666
rect 93537 138608 93542 138664
rect 93598 138608 97970 138664
rect 93537 138606 97970 138608
rect 93537 138603 93603 138606
rect 196945 138394 197011 138397
rect 201416 138394 201896 138424
rect 196945 138392 201896 138394
rect 196945 138336 196950 138392
rect 197006 138336 201896 138392
rect 196945 138334 201896 138336
rect 196945 138331 197011 138334
rect 201416 138304 201896 138334
rect 92065 137578 92131 137581
rect 164745 137578 164811 137581
rect 89844 137576 92131 137578
rect 89844 137520 92070 137576
rect 92126 137520 92131 137576
rect 89844 137518 92131 137520
rect 161788 137576 164811 137578
rect 161788 137520 164750 137576
rect 164806 137520 164811 137576
rect 161788 137518 164811 137520
rect 92065 137515 92131 137518
rect 164745 137515 164811 137518
rect 93353 137034 93419 137037
rect 93353 137032 97940 137034
rect 93353 136976 93358 137032
rect 93414 136976 97940 137032
rect 93353 136974 97940 136976
rect 93353 136971 93419 136974
rect 92157 136490 92223 136493
rect 163089 136490 163155 136493
rect 89844 136488 92223 136490
rect 89844 136432 92162 136488
rect 92218 136432 92223 136488
rect 89844 136430 92223 136432
rect 161788 136488 163155 136490
rect 161788 136432 163094 136488
rect 163150 136432 163155 136488
rect 161788 136430 163155 136432
rect 92157 136427 92223 136430
rect 163089 136427 163155 136430
rect 168517 136218 168583 136221
rect 170038 136218 170098 136800
rect 168517 136216 170098 136218
rect 168517 136160 168522 136216
rect 168578 136160 170098 136216
rect 168517 136158 170098 136160
rect 168517 136155 168583 136158
rect 82129 133090 82195 133093
rect 83601 133092 83667 133093
rect 82262 133090 82268 133092
rect 82129 133088 82268 133090
rect 82129 133032 82134 133088
rect 82190 133032 82268 133088
rect 82129 133030 82268 133032
rect 82129 133027 82195 133030
rect 82262 133028 82268 133030
rect 82332 133028 82338 133092
rect 83550 133090 83556 133092
rect 83510 133030 83556 133090
rect 83620 133088 83667 133092
rect 83662 133032 83667 133088
rect 83550 133028 83556 133030
rect 83620 133028 83667 133032
rect 83601 133027 83667 133028
rect 47862 128194 47922 128504
rect 91470 128470 92052 128530
rect 88569 128466 88635 128469
rect 91470 128466 91530 128470
rect 88569 128464 91530 128466
rect 88569 128408 88574 128464
rect 88630 128408 91530 128464
rect 88569 128406 91530 128408
rect 88569 128403 88635 128406
rect 51217 128194 51283 128197
rect 47862 128192 51283 128194
rect 47862 128136 51222 128192
rect 51278 128136 51283 128192
rect 47862 128134 51283 128136
rect 119806 128194 119866 128504
rect 123069 128194 123135 128197
rect 119806 128192 123135 128194
rect 119806 128136 123074 128192
rect 123130 128136 123135 128192
rect 119806 128134 123135 128136
rect 51217 128131 51283 128134
rect 123069 128131 123135 128134
rect 160329 128194 160395 128197
rect 163966 128194 164026 128504
rect 160329 128192 164026 128194
rect 160329 128136 160334 128192
rect 160390 128136 164026 128192
rect 160329 128134 164026 128136
rect 160329 128131 160395 128134
rect 47862 127650 47922 127960
rect 91470 127926 92052 127986
rect 88385 127922 88451 127925
rect 91470 127922 91530 127926
rect 88385 127920 91530 127922
rect 88385 127864 88390 127920
rect 88446 127864 91530 127920
rect 88385 127862 91530 127864
rect 88385 127859 88451 127862
rect 119806 127786 119866 127960
rect 123161 127786 123227 127789
rect 119806 127784 123227 127786
rect 119806 127728 123166 127784
rect 123222 127728 123227 127784
rect 119806 127726 123227 127728
rect 123161 127723 123227 127726
rect 51401 127650 51467 127653
rect 47862 127648 51467 127650
rect 47862 127592 51406 127648
rect 51462 127592 51467 127648
rect 47862 127590 51467 127592
rect 51401 127587 51467 127590
rect 160145 127650 160211 127653
rect 163966 127650 164026 127960
rect 160145 127648 164026 127650
rect 160145 127592 160150 127648
rect 160206 127592 164026 127648
rect 160145 127590 164026 127592
rect 160145 127587 160211 127590
rect 47862 126970 47922 127416
rect 91470 127382 92052 127442
rect 88661 127378 88727 127381
rect 91470 127378 91530 127382
rect 88661 127376 91530 127378
rect 88661 127320 88666 127376
rect 88722 127320 91530 127376
rect 88661 127318 91530 127320
rect 88661 127315 88727 127318
rect 119806 127242 119866 127416
rect 121689 127242 121755 127245
rect 119806 127240 121755 127242
rect 119806 127184 121694 127240
rect 121750 127184 121755 127240
rect 119806 127182 121755 127184
rect 121689 127179 121755 127182
rect 51309 127106 51375 127109
rect 123069 127106 123135 127109
rect 51309 127104 55098 127106
rect 51309 127048 51314 127104
rect 51370 127048 55098 127104
rect 51309 127046 55098 127048
rect 51309 127043 51375 127046
rect 51217 126970 51283 126973
rect 47862 126968 51283 126970
rect 47862 126912 51222 126968
rect 51278 126912 51283 126968
rect 47862 126910 51283 126912
rect 51217 126907 51283 126910
rect 47862 126426 47922 126736
rect 55038 126464 55098 127046
rect 123069 127104 127042 127106
rect 123069 127048 123074 127104
rect 123130 127048 127042 127104
rect 123069 127046 127042 127048
rect 123069 127043 123135 127046
rect 91470 126702 92052 126762
rect 88293 126698 88359 126701
rect 91470 126698 91530 126702
rect 88293 126696 91530 126698
rect 88293 126640 88298 126696
rect 88354 126640 91530 126696
rect 88293 126638 91530 126640
rect 88293 126635 88359 126638
rect 119806 126562 119866 126736
rect 121781 126562 121847 126565
rect 119806 126560 121847 126562
rect 119806 126504 121786 126560
rect 121842 126504 121847 126560
rect 119806 126502 121847 126504
rect 121781 126499 121847 126502
rect 126982 126464 127042 127046
rect 160421 126970 160487 126973
rect 163966 126970 164026 127416
rect 160421 126968 164026 126970
rect 160421 126912 160426 126968
rect 160482 126912 164026 126968
rect 160421 126910 164026 126912
rect 160421 126907 160487 126910
rect 160053 126562 160119 126565
rect 163966 126562 164026 126736
rect 160053 126560 164026 126562
rect 160053 126504 160058 126560
rect 160114 126504 164026 126560
rect 160053 126502 164026 126504
rect 160053 126499 160119 126502
rect 51493 126426 51559 126429
rect 88477 126426 88543 126429
rect 160237 126426 160303 126429
rect 47862 126424 51559 126426
rect 47862 126368 51498 126424
rect 51554 126368 51559 126424
rect 47862 126366 51559 126368
rect 84876 126424 88543 126426
rect 84876 126368 88482 126424
rect 88538 126368 88543 126424
rect 84876 126366 88543 126368
rect 156820 126424 160303 126426
rect 156820 126368 160242 126424
rect 160298 126368 160303 126424
rect 156820 126366 160303 126368
rect 51493 126363 51559 126366
rect 88477 126363 88543 126366
rect 160237 126363 160303 126366
rect 47862 126154 47922 126192
rect 91470 126158 92052 126218
rect 51217 126154 51283 126157
rect 47862 126152 51283 126154
rect 47862 126096 51222 126152
rect 51278 126096 51283 126152
rect 47862 126094 51283 126096
rect 51217 126091 51283 126094
rect 88477 126154 88543 126157
rect 91470 126154 91530 126158
rect 88477 126152 91530 126154
rect 88477 126096 88482 126152
rect 88538 126096 91530 126152
rect 88477 126094 91530 126096
rect 119806 126154 119866 126192
rect 121689 126154 121755 126157
rect 119806 126152 121755 126154
rect 119806 126096 121694 126152
rect 121750 126096 121755 126152
rect 119806 126094 121755 126096
rect 88477 126091 88543 126094
rect 121689 126091 121755 126094
rect 160237 126154 160303 126157
rect 163966 126154 164026 126192
rect 160237 126152 164026 126154
rect 160237 126096 160242 126152
rect 160298 126096 164026 126152
rect 160237 126094 164026 126096
rect 160237 126091 160303 126094
rect 51401 125882 51467 125885
rect 88385 125882 88451 125885
rect 51401 125880 55068 125882
rect 51401 125824 51406 125880
rect 51462 125824 55068 125880
rect 51401 125822 55068 125824
rect 84876 125880 88451 125882
rect 84876 125824 88390 125880
rect 88446 125824 88451 125880
rect 84876 125822 88451 125824
rect 51401 125819 51467 125822
rect 88385 125819 88451 125822
rect 123161 125882 123227 125885
rect 160145 125882 160211 125885
rect 123161 125880 127012 125882
rect 123161 125824 123166 125880
rect 123222 125824 127012 125880
rect 123161 125822 127012 125824
rect 156820 125880 160211 125882
rect 156820 125824 160150 125880
rect 160206 125824 160211 125880
rect 156820 125822 160211 125824
rect 123161 125819 123227 125822
rect 160145 125819 160211 125822
rect 51309 125746 51375 125749
rect 123989 125746 124055 125749
rect 51309 125744 55098 125746
rect 51309 125688 51314 125744
rect 51370 125688 55098 125744
rect 51309 125686 55098 125688
rect 51309 125683 51375 125686
rect 9896 125338 10376 125368
rect 13313 125338 13379 125341
rect 9896 125336 13379 125338
rect 9896 125280 13318 125336
rect 13374 125280 13379 125336
rect 9896 125278 13379 125280
rect 9896 125248 10376 125278
rect 13313 125275 13379 125278
rect 47862 125202 47922 125648
rect 55038 125240 55098 125686
rect 123989 125744 127042 125746
rect 123989 125688 123994 125744
rect 124050 125688 127042 125744
rect 123989 125686 127042 125688
rect 123989 125683 124055 125686
rect 91470 125614 92052 125674
rect 88753 125610 88819 125613
rect 91470 125610 91530 125614
rect 88753 125608 91530 125610
rect 88753 125552 88758 125608
rect 88814 125552 91530 125608
rect 88753 125550 91530 125552
rect 88753 125547 88819 125550
rect 119806 125474 119866 125648
rect 121689 125474 121755 125477
rect 119806 125472 121755 125474
rect 119806 125416 121694 125472
rect 121750 125416 121755 125472
rect 119806 125414 121755 125416
rect 121689 125411 121755 125414
rect 126982 125240 127042 125686
rect 51217 125202 51283 125205
rect 88477 125202 88543 125205
rect 160237 125202 160303 125205
rect 47862 125200 51283 125202
rect 47862 125144 51222 125200
rect 51278 125144 51283 125200
rect 47862 125142 51283 125144
rect 84876 125200 88543 125202
rect 84876 125144 88482 125200
rect 88538 125144 88543 125200
rect 84876 125142 88543 125144
rect 156820 125200 160303 125202
rect 156820 125144 160242 125200
rect 160298 125144 160303 125200
rect 156820 125142 160303 125144
rect 51217 125139 51283 125142
rect 88477 125139 88543 125142
rect 160237 125139 160303 125142
rect 160513 125202 160579 125205
rect 163966 125202 164026 125648
rect 160513 125200 164026 125202
rect 160513 125144 160518 125200
rect 160574 125144 164026 125200
rect 160513 125142 164026 125144
rect 160513 125139 160579 125142
rect 47862 124794 47922 124968
rect 91470 124934 92052 124994
rect 88477 124930 88543 124933
rect 91470 124930 91530 124934
rect 88477 124928 91530 124930
rect 88477 124872 88482 124928
rect 88538 124872 91530 124928
rect 88477 124870 91530 124872
rect 119806 124930 119866 124968
rect 123161 124930 123227 124933
rect 119806 124928 123227 124930
rect 119806 124872 123166 124928
rect 123222 124872 123227 124928
rect 119806 124870 123227 124872
rect 88477 124867 88543 124870
rect 123161 124867 123227 124870
rect 160237 124930 160303 124933
rect 163966 124930 164026 124968
rect 160237 124928 164026 124930
rect 160237 124872 160242 124928
rect 160298 124872 164026 124928
rect 160237 124870 164026 124872
rect 160237 124867 160303 124870
rect 51401 124794 51467 124797
rect 47862 124792 51467 124794
rect 47862 124736 51406 124792
rect 51462 124736 51467 124792
rect 47862 124734 51467 124736
rect 51401 124731 51467 124734
rect 51493 124658 51559 124661
rect 88293 124658 88359 124661
rect 51493 124656 55068 124658
rect 51493 124600 51498 124656
rect 51554 124600 55068 124656
rect 51493 124598 55068 124600
rect 84876 124656 88359 124658
rect 84876 124600 88298 124656
rect 88354 124600 88359 124656
rect 84876 124598 88359 124600
rect 51493 124595 51559 124598
rect 88293 124595 88359 124598
rect 124357 124658 124423 124661
rect 160053 124658 160119 124661
rect 124357 124656 127012 124658
rect 124357 124600 124362 124656
rect 124418 124600 127012 124656
rect 124357 124598 127012 124600
rect 156820 124656 160119 124658
rect 156820 124600 160058 124656
rect 160114 124600 160119 124656
rect 156820 124598 160119 124600
rect 124357 124595 124423 124598
rect 160053 124595 160119 124598
rect 51309 124522 51375 124525
rect 123897 124522 123963 124525
rect 51309 124520 55098 124522
rect 51309 124464 51314 124520
rect 51370 124464 55098 124520
rect 51309 124462 55098 124464
rect 51309 124459 51375 124462
rect 18097 123570 18163 123573
rect 19894 123570 19954 124152
rect 47862 124114 47922 124424
rect 55038 124152 55098 124462
rect 123897 124520 127042 124522
rect 123897 124464 123902 124520
rect 123958 124464 127042 124520
rect 123897 124462 127042 124464
rect 123897 124459 123963 124462
rect 91470 124390 92052 124450
rect 88661 124386 88727 124389
rect 91470 124386 91530 124390
rect 88661 124384 91530 124386
rect 88661 124328 88666 124384
rect 88722 124328 91530 124384
rect 88661 124326 91530 124328
rect 88661 124323 88727 124326
rect 51217 124114 51283 124117
rect 88385 124114 88451 124117
rect 47862 124112 51283 124114
rect 47862 124056 51222 124112
rect 51278 124056 51283 124112
rect 47862 124054 51283 124056
rect 84876 124112 88451 124114
rect 84876 124056 88390 124112
rect 88446 124056 88451 124112
rect 84876 124054 88451 124056
rect 119806 124114 119866 124424
rect 126982 124152 127042 124462
rect 122977 124114 123043 124117
rect 160145 124114 160211 124117
rect 119806 124112 123043 124114
rect 119806 124056 122982 124112
rect 123038 124056 123043 124112
rect 119806 124054 123043 124056
rect 156820 124112 160211 124114
rect 156820 124056 160150 124112
rect 160206 124056 160211 124112
rect 156820 124054 160211 124056
rect 51217 124051 51283 124054
rect 88385 124051 88451 124054
rect 122977 124051 123043 124054
rect 160145 124051 160211 124054
rect 160421 124114 160487 124117
rect 163966 124114 164026 124424
rect 160421 124112 164026 124114
rect 160421 124056 160426 124112
rect 160482 124056 164026 124112
rect 160421 124054 164026 124056
rect 160421 124051 160487 124054
rect 51309 123978 51375 123981
rect 123713 123978 123779 123981
rect 51309 123976 55098 123978
rect 51309 123920 51314 123976
rect 51370 123920 55098 123976
rect 51309 123918 55098 123920
rect 51309 123915 51375 123918
rect 18097 123568 19954 123570
rect 18097 123512 18102 123568
rect 18158 123512 19954 123568
rect 18097 123510 19954 123512
rect 47862 123570 47922 123880
rect 51493 123570 51559 123573
rect 47862 123568 51559 123570
rect 47862 123512 51498 123568
rect 51554 123512 51559 123568
rect 47862 123510 51559 123512
rect 18097 123507 18163 123510
rect 51493 123507 51559 123510
rect 55038 123472 55098 123918
rect 123713 123976 127042 123978
rect 123713 123920 123718 123976
rect 123774 123920 127042 123976
rect 123713 123918 127042 123920
rect 123713 123915 123779 123918
rect 91470 123846 92052 123906
rect 88385 123842 88451 123845
rect 91470 123842 91530 123846
rect 88385 123840 91530 123842
rect 88385 123784 88390 123840
rect 88446 123784 91530 123840
rect 88385 123782 91530 123784
rect 88385 123779 88451 123782
rect 119806 123706 119866 123880
rect 121689 123706 121755 123709
rect 119806 123704 121755 123706
rect 119806 123648 121694 123704
rect 121750 123648 121755 123704
rect 119806 123646 121755 123648
rect 121689 123643 121755 123646
rect 126982 123472 127042 123918
rect 160053 123570 160119 123573
rect 163966 123570 164026 123880
rect 160053 123568 164026 123570
rect 160053 123512 160058 123568
rect 160114 123512 164026 123568
rect 160053 123510 164026 123512
rect 191750 123570 191810 124148
rect 193541 123570 193607 123573
rect 191750 123568 193607 123570
rect 191750 123512 193546 123568
rect 193602 123512 193607 123568
rect 191750 123510 193607 123512
rect 160053 123507 160119 123510
rect 193541 123507 193607 123510
rect 87741 123434 87807 123437
rect 160237 123434 160303 123437
rect 84876 123432 87807 123434
rect 84876 123376 87746 123432
rect 87802 123376 87807 123432
rect 84876 123374 87807 123376
rect 156820 123432 160303 123434
rect 156820 123376 160242 123432
rect 160298 123376 160303 123432
rect 156820 123374 160303 123376
rect 87741 123371 87807 123374
rect 160237 123371 160303 123374
rect 47862 122890 47922 123336
rect 91470 123302 92052 123362
rect 51401 123298 51467 123301
rect 88569 123298 88635 123301
rect 91470 123298 91530 123302
rect 51401 123296 55098 123298
rect 51401 123240 51406 123296
rect 51462 123240 55098 123296
rect 51401 123238 55098 123240
rect 51401 123235 51467 123238
rect 55038 122928 55098 123238
rect 88569 123296 91530 123298
rect 88569 123240 88574 123296
rect 88630 123240 91530 123296
rect 88569 123238 91530 123240
rect 88569 123235 88635 123238
rect 51309 122890 51375 122893
rect 88477 122890 88543 122893
rect 47862 122888 51375 122890
rect 47862 122832 51314 122888
rect 51370 122832 51375 122888
rect 47862 122830 51375 122832
rect 84876 122888 88543 122890
rect 84876 122832 88482 122888
rect 88538 122832 88543 122888
rect 84876 122830 88543 122832
rect 119806 122890 119866 123336
rect 123161 123298 123227 123301
rect 123161 123296 127042 123298
rect 123161 123240 123166 123296
rect 123222 123240 127042 123296
rect 123161 123238 127042 123240
rect 123161 123235 123227 123238
rect 126982 122928 127042 123238
rect 122977 122890 123043 122893
rect 160145 122890 160211 122893
rect 119806 122888 123043 122890
rect 119806 122832 122982 122888
rect 123038 122832 123043 122888
rect 119806 122830 123043 122832
rect 156820 122888 160211 122890
rect 156820 122832 160150 122888
rect 160206 122832 160211 122888
rect 156820 122830 160211 122832
rect 51309 122827 51375 122830
rect 88477 122827 88543 122830
rect 122977 122827 123043 122830
rect 160145 122827 160211 122830
rect 160421 122890 160487 122893
rect 163966 122890 164026 123336
rect 160421 122888 164026 122890
rect 160421 122832 160426 122888
rect 160482 122832 164026 122888
rect 160421 122830 164026 122832
rect 160421 122827 160487 122830
rect 51401 122754 51467 122757
rect 123069 122754 123135 122757
rect 160237 122754 160303 122757
rect 51401 122752 55098 122754
rect 51401 122696 51406 122752
rect 51462 122696 55098 122752
rect 51401 122694 55098 122696
rect 51401 122691 51467 122694
rect 47862 122346 47922 122656
rect 51769 122346 51835 122349
rect 47862 122344 51835 122346
rect 47862 122288 51774 122344
rect 51830 122288 51835 122344
rect 47862 122286 51835 122288
rect 51769 122283 51835 122286
rect 55038 122248 55098 122694
rect 123069 122752 127042 122754
rect 123069 122696 123074 122752
rect 123130 122696 127042 122752
rect 123069 122694 127042 122696
rect 123069 122691 123135 122694
rect 91470 122622 92052 122682
rect 88201 122618 88267 122621
rect 91470 122618 91530 122622
rect 88201 122616 91530 122618
rect 88201 122560 88206 122616
rect 88262 122560 91530 122616
rect 88201 122558 91530 122560
rect 88201 122555 88267 122558
rect 119806 122482 119866 122656
rect 121689 122482 121755 122485
rect 119806 122480 121755 122482
rect 119806 122424 121694 122480
rect 121750 122424 121755 122480
rect 119806 122422 121755 122424
rect 121689 122419 121755 122422
rect 126982 122248 127042 122694
rect 156790 122752 160303 122754
rect 156790 122696 160242 122752
rect 160298 122696 160303 122752
rect 156790 122694 160303 122696
rect 88661 122210 88727 122213
rect 84876 122208 88727 122210
rect 84876 122152 88666 122208
rect 88722 122152 88727 122208
rect 156790 122180 156850 122694
rect 160237 122691 160303 122694
rect 160237 122346 160303 122349
rect 163966 122346 164026 122656
rect 160237 122344 164026 122346
rect 160237 122288 160242 122344
rect 160298 122288 164026 122344
rect 160237 122286 164026 122288
rect 160237 122283 160303 122286
rect 84876 122150 88727 122152
rect 88661 122147 88727 122150
rect 47862 122074 47922 122112
rect 91470 122078 92052 122138
rect 51401 122074 51467 122077
rect 47862 122072 51467 122074
rect 47862 122016 51406 122072
rect 51462 122016 51467 122072
rect 47862 122014 51467 122016
rect 51401 122011 51467 122014
rect 88293 122074 88359 122077
rect 91470 122074 91530 122078
rect 88293 122072 91530 122074
rect 88293 122016 88298 122072
rect 88354 122016 91530 122072
rect 88293 122014 91530 122016
rect 119806 122074 119866 122112
rect 121689 122074 121755 122077
rect 119806 122072 121755 122074
rect 119806 122016 121694 122072
rect 121750 122016 121755 122072
rect 119806 122014 121755 122016
rect 88293 122011 88359 122014
rect 121689 122011 121755 122014
rect 160145 122074 160211 122077
rect 163966 122074 164026 122112
rect 160145 122072 164026 122074
rect 160145 122016 160150 122072
rect 160206 122016 164026 122072
rect 160145 122014 164026 122016
rect 160145 122011 160211 122014
rect 51493 121666 51559 121669
rect 88385 121666 88451 121669
rect 51493 121664 55068 121666
rect 51493 121608 51498 121664
rect 51554 121608 55068 121664
rect 51493 121606 55068 121608
rect 84876 121664 88451 121666
rect 84876 121608 88390 121664
rect 88446 121608 88451 121664
rect 84876 121606 88451 121608
rect 51493 121603 51559 121606
rect 88385 121603 88451 121606
rect 123529 121666 123595 121669
rect 160053 121666 160119 121669
rect 123529 121664 127012 121666
rect 123529 121608 123534 121664
rect 123590 121608 127012 121664
rect 123529 121606 127012 121608
rect 156820 121664 160119 121666
rect 156820 121608 160058 121664
rect 160114 121608 160119 121664
rect 156820 121606 160119 121608
rect 123529 121603 123595 121606
rect 160053 121603 160119 121606
rect 47862 121122 47922 121568
rect 91470 121534 92052 121594
rect 51309 121530 51375 121533
rect 88385 121530 88451 121533
rect 91470 121530 91530 121534
rect 51309 121528 55098 121530
rect 51309 121472 51314 121528
rect 51370 121472 55098 121528
rect 51309 121470 55098 121472
rect 51309 121467 51375 121470
rect 55038 121160 55098 121470
rect 88385 121528 91530 121530
rect 88385 121472 88390 121528
rect 88446 121472 91530 121528
rect 88385 121470 91530 121472
rect 88385 121467 88451 121470
rect 119806 121258 119866 121568
rect 123069 121530 123135 121533
rect 123069 121528 127042 121530
rect 123069 121472 123074 121528
rect 123130 121472 127042 121528
rect 123069 121470 127042 121472
rect 123069 121467 123135 121470
rect 121689 121258 121755 121261
rect 119806 121256 121755 121258
rect 119806 121200 121694 121256
rect 121750 121200 121755 121256
rect 119806 121198 121755 121200
rect 121689 121195 121755 121198
rect 126982 121160 127042 121470
rect 159961 121258 160027 121261
rect 163966 121258 164026 121568
rect 159961 121256 164026 121258
rect 159961 121200 159966 121256
rect 160022 121200 164026 121256
rect 159961 121198 164026 121200
rect 159961 121195 160027 121198
rect 51493 121122 51559 121125
rect 88477 121122 88543 121125
rect 160237 121122 160303 121125
rect 47862 121120 51559 121122
rect 47862 121064 51498 121120
rect 51554 121064 51559 121120
rect 47862 121062 51559 121064
rect 84876 121120 88543 121122
rect 84876 121064 88482 121120
rect 88538 121064 88543 121120
rect 84876 121062 88543 121064
rect 156820 121120 160303 121122
rect 156820 121064 160242 121120
rect 160298 121064 160303 121120
rect 156820 121062 160303 121064
rect 51493 121059 51559 121062
rect 88477 121059 88543 121062
rect 160237 121059 160303 121062
rect 47862 120714 47922 120888
rect 91470 120854 92052 120914
rect 88477 120850 88543 120853
rect 91470 120850 91530 120854
rect 88477 120848 91530 120850
rect 88477 120792 88482 120848
rect 88538 120792 91530 120848
rect 88477 120790 91530 120792
rect 88477 120787 88543 120790
rect 51217 120714 51283 120717
rect 47862 120712 51283 120714
rect 47862 120656 51222 120712
rect 51278 120656 51283 120712
rect 47862 120654 51283 120656
rect 119806 120714 119866 120888
rect 122977 120714 123043 120717
rect 119806 120712 123043 120714
rect 119806 120656 122982 120712
rect 123038 120656 123043 120712
rect 119806 120654 123043 120656
rect 51217 120651 51283 120654
rect 122977 120651 123043 120654
rect 160237 120714 160303 120717
rect 163966 120714 164026 120888
rect 160237 120712 164026 120714
rect 160237 120656 160242 120712
rect 160298 120656 164026 120712
rect 160237 120654 164026 120656
rect 160237 120651 160303 120654
rect 51769 120442 51835 120445
rect 88201 120442 88267 120445
rect 51769 120440 55068 120442
rect 51769 120384 51774 120440
rect 51830 120384 55068 120440
rect 51769 120382 55068 120384
rect 84876 120440 88267 120442
rect 84876 120384 88206 120440
rect 88262 120384 88267 120440
rect 84876 120382 88267 120384
rect 51769 120379 51835 120382
rect 88201 120379 88267 120382
rect 123437 120442 123503 120445
rect 160145 120442 160211 120445
rect 123437 120440 127012 120442
rect 123437 120384 123442 120440
rect 123498 120384 127012 120440
rect 123437 120382 127012 120384
rect 156820 120440 160211 120442
rect 156820 120384 160150 120440
rect 160206 120384 160211 120440
rect 156820 120382 160211 120384
rect 123437 120379 123503 120382
rect 160145 120379 160211 120382
rect 47862 120034 47922 120344
rect 91470 120310 92052 120370
rect 51401 120306 51467 120309
rect 88569 120306 88635 120309
rect 91470 120306 91530 120310
rect 51401 120304 55098 120306
rect 51401 120248 51406 120304
rect 51462 120248 55098 120304
rect 51401 120246 55098 120248
rect 51401 120243 51467 120246
rect 51217 120034 51283 120037
rect 47862 120032 51283 120034
rect 47862 119976 51222 120032
rect 51278 119976 51283 120032
rect 47862 119974 51283 119976
rect 51217 119971 51283 119974
rect 55038 119936 55098 120246
rect 88569 120304 91530 120306
rect 88569 120248 88574 120304
rect 88630 120248 91530 120304
rect 88569 120246 91530 120248
rect 88569 120243 88635 120246
rect 119806 120034 119866 120344
rect 123345 120306 123411 120309
rect 123345 120304 127042 120306
rect 123345 120248 123350 120304
rect 123406 120248 127042 120304
rect 123345 120246 127042 120248
rect 123345 120243 123411 120246
rect 122977 120034 123043 120037
rect 119806 120032 123043 120034
rect 119806 119976 122982 120032
rect 123038 119976 123043 120032
rect 119806 119974 123043 119976
rect 122977 119971 123043 119974
rect 126982 119936 127042 120246
rect 160329 120034 160395 120037
rect 163966 120034 164026 120344
rect 160329 120032 164026 120034
rect 160329 119976 160334 120032
rect 160390 119976 164026 120032
rect 160329 119974 164026 119976
rect 160329 119971 160395 119974
rect 88293 119898 88359 119901
rect 160053 119898 160119 119901
rect 84876 119896 88359 119898
rect 84876 119840 88298 119896
rect 88354 119840 88359 119896
rect 84876 119838 88359 119840
rect 156820 119896 160119 119898
rect 156820 119840 160058 119896
rect 160114 119840 160119 119896
rect 156820 119838 160119 119840
rect 88293 119835 88359 119838
rect 160053 119835 160119 119838
rect 47862 119490 47922 119800
rect 91470 119766 92052 119826
rect 88293 119762 88359 119765
rect 91470 119762 91530 119766
rect 88293 119760 91530 119762
rect 88293 119704 88298 119760
rect 88354 119704 91530 119760
rect 88293 119702 91530 119704
rect 88293 119699 88359 119702
rect 119806 119626 119866 119800
rect 121689 119626 121755 119629
rect 119806 119624 121755 119626
rect 119806 119568 121694 119624
rect 121750 119568 121755 119624
rect 119806 119566 121755 119568
rect 121689 119563 121755 119566
rect 51401 119490 51467 119493
rect 47862 119488 51467 119490
rect 47862 119432 51406 119488
rect 51462 119432 51467 119488
rect 47862 119430 51467 119432
rect 51401 119427 51467 119430
rect 160145 119490 160211 119493
rect 163966 119490 164026 119800
rect 160145 119488 164026 119490
rect 160145 119432 160150 119488
rect 160206 119432 164026 119488
rect 160145 119430 164026 119432
rect 160145 119427 160211 119430
rect 51125 119354 51191 119357
rect 47862 119352 51191 119354
rect 47862 119296 51130 119352
rect 51186 119296 51191 119352
rect 47862 119294 51191 119296
rect 47862 119256 47922 119294
rect 51125 119291 51191 119294
rect 88201 119354 88267 119357
rect 123253 119354 123319 119357
rect 88201 119352 91530 119354
rect 88201 119296 88206 119352
rect 88262 119296 91530 119352
rect 88201 119294 91530 119296
rect 88201 119291 88267 119294
rect 91470 119286 91530 119294
rect 119806 119352 123319 119354
rect 119806 119296 123258 119352
rect 123314 119296 123319 119352
rect 119806 119294 123319 119296
rect 91470 119226 92052 119286
rect 119806 119256 119866 119294
rect 123253 119291 123319 119294
rect 159869 119354 159935 119357
rect 159869 119352 164026 119354
rect 159869 119296 159874 119352
rect 159930 119296 164026 119352
rect 159869 119294 164026 119296
rect 159869 119291 159935 119294
rect 163966 119256 164026 119294
rect 51493 119218 51559 119221
rect 88385 119218 88451 119221
rect 51493 119216 55068 119218
rect 51493 119160 51498 119216
rect 51554 119160 55068 119216
rect 51493 119158 55068 119160
rect 84876 119216 88451 119218
rect 84876 119160 88390 119216
rect 88446 119160 88451 119216
rect 84876 119158 88451 119160
rect 51493 119155 51559 119158
rect 88385 119155 88451 119158
rect 124357 119218 124423 119221
rect 159961 119218 160027 119221
rect 124357 119216 127012 119218
rect 124357 119160 124362 119216
rect 124418 119160 127012 119216
rect 124357 119158 127012 119160
rect 156820 119216 160027 119218
rect 156820 119160 159966 119216
rect 160022 119160 160027 119216
rect 156820 119158 160027 119160
rect 124357 119155 124423 119158
rect 159961 119155 160027 119158
rect 51309 119082 51375 119085
rect 123161 119082 123227 119085
rect 51309 119080 55098 119082
rect 51309 119024 51314 119080
rect 51370 119024 55098 119080
rect 51309 119022 55098 119024
rect 51309 119019 51375 119022
rect 55038 118712 55098 119022
rect 123161 119080 127042 119082
rect 123161 119024 123166 119080
rect 123222 119024 127042 119080
rect 123161 119022 127042 119024
rect 123161 119019 123227 119022
rect 126982 118712 127042 119022
rect 88477 118674 88543 118677
rect 160237 118674 160303 118677
rect 84876 118672 88543 118674
rect 84876 118616 88482 118672
rect 88538 118616 88543 118672
rect 84876 118614 88543 118616
rect 156820 118672 160303 118674
rect 156820 118616 160242 118672
rect 160298 118616 160303 118672
rect 156820 118614 160303 118616
rect 88477 118611 88543 118614
rect 160237 118611 160303 118614
rect 47862 118266 47922 118576
rect 91470 118542 92052 118602
rect 51309 118538 51375 118541
rect 88385 118538 88451 118541
rect 91470 118538 91530 118542
rect 51309 118536 55098 118538
rect 51309 118480 51314 118536
rect 51370 118480 55098 118536
rect 51309 118478 55098 118480
rect 51309 118475 51375 118478
rect 51217 118266 51283 118269
rect 47862 118264 51283 118266
rect 47862 118208 51222 118264
rect 51278 118208 51283 118264
rect 47862 118206 51283 118208
rect 51217 118203 51283 118206
rect 55038 118168 55098 118478
rect 88385 118536 91530 118538
rect 88385 118480 88390 118536
rect 88446 118480 91530 118536
rect 88385 118478 91530 118480
rect 88385 118475 88451 118478
rect 119806 118402 119866 118576
rect 123069 118538 123135 118541
rect 123069 118536 127042 118538
rect 123069 118480 123074 118536
rect 123130 118480 127042 118536
rect 123069 118478 127042 118480
rect 123069 118475 123135 118478
rect 121689 118402 121755 118405
rect 119806 118400 121755 118402
rect 119806 118344 121694 118400
rect 121750 118344 121755 118400
rect 119806 118342 121755 118344
rect 121689 118339 121755 118342
rect 126982 118168 127042 118478
rect 160053 118266 160119 118269
rect 163966 118266 164026 118576
rect 160053 118264 164026 118266
rect 160053 118208 160058 118264
rect 160114 118208 164026 118264
rect 160053 118206 164026 118208
rect 160053 118203 160119 118206
rect 88477 118130 88543 118133
rect 160237 118130 160303 118133
rect 84876 118128 88543 118130
rect 84876 118072 88482 118128
rect 88538 118072 88543 118128
rect 84876 118070 88543 118072
rect 156820 118128 160303 118130
rect 156820 118072 160242 118128
rect 160298 118072 160303 118128
rect 156820 118070 160303 118072
rect 88477 118067 88543 118070
rect 160237 118067 160303 118070
rect 47862 117994 47922 118032
rect 91470 117998 92052 118058
rect 51493 117994 51559 117997
rect 47862 117992 51559 117994
rect 47862 117936 51498 117992
rect 51554 117936 51559 117992
rect 47862 117934 51559 117936
rect 51493 117931 51559 117934
rect 88109 117994 88175 117997
rect 91470 117994 91530 117998
rect 88109 117992 91530 117994
rect 88109 117936 88114 117992
rect 88170 117936 91530 117992
rect 88109 117934 91530 117936
rect 119806 117994 119866 118032
rect 123161 117994 123227 117997
rect 119806 117992 123227 117994
rect 119806 117936 123166 117992
rect 123222 117936 123227 117992
rect 119806 117934 123227 117936
rect 88109 117931 88175 117934
rect 123161 117931 123227 117934
rect 160237 117994 160303 117997
rect 163966 117994 164026 118032
rect 160237 117992 164026 117994
rect 160237 117936 160242 117992
rect 160298 117936 164026 117992
rect 160237 117934 164026 117936
rect 160237 117931 160303 117934
rect 51401 117858 51467 117861
rect 124265 117858 124331 117861
rect 51401 117856 55098 117858
rect 51401 117800 51406 117856
rect 51462 117800 55098 117856
rect 51401 117798 55098 117800
rect 51401 117795 51467 117798
rect 55038 117488 55098 117798
rect 124265 117856 127042 117858
rect 124265 117800 124270 117856
rect 124326 117800 127042 117856
rect 124265 117798 127042 117800
rect 124265 117795 124331 117798
rect 47862 117042 47922 117488
rect 91470 117454 92052 117514
rect 126982 117488 127042 117798
rect 88293 117450 88359 117453
rect 84876 117448 88359 117450
rect 84876 117392 88298 117448
rect 88354 117392 88359 117448
rect 84876 117390 88359 117392
rect 88293 117387 88359 117390
rect 88661 117450 88727 117453
rect 91470 117450 91530 117454
rect 88661 117448 91530 117450
rect 88661 117392 88666 117448
rect 88722 117392 91530 117448
rect 88661 117390 91530 117392
rect 88661 117387 88727 117390
rect 51585 117314 51651 117317
rect 51585 117312 55098 117314
rect 51585 117256 51590 117312
rect 51646 117256 55098 117312
rect 51585 117254 55098 117256
rect 51585 117251 51651 117254
rect 50573 117042 50639 117045
rect 47862 117040 50639 117042
rect 47862 116984 50578 117040
rect 50634 116984 50639 117040
rect 47862 116982 50639 116984
rect 50573 116979 50639 116982
rect 55038 116944 55098 117254
rect 119806 117042 119866 117488
rect 160145 117450 160211 117453
rect 156820 117448 160211 117450
rect 156820 117392 160150 117448
rect 160206 117392 160211 117448
rect 156820 117390 160211 117392
rect 160145 117387 160211 117390
rect 123253 117314 123319 117317
rect 123253 117312 127042 117314
rect 123253 117256 123258 117312
rect 123314 117256 127042 117312
rect 123253 117254 127042 117256
rect 123253 117251 123319 117254
rect 122977 117042 123043 117045
rect 119806 117040 123043 117042
rect 119806 116984 122982 117040
rect 123038 116984 123043 117040
rect 119806 116982 123043 116984
rect 122977 116979 123043 116982
rect 126982 116944 127042 117254
rect 160421 117042 160487 117045
rect 163966 117042 164026 117488
rect 160421 117040 164026 117042
rect 160421 116984 160426 117040
rect 160482 116984 164026 117040
rect 160421 116982 164026 116984
rect 160421 116979 160487 116982
rect 88201 116906 88267 116909
rect 159869 116906 159935 116909
rect 84876 116904 88267 116906
rect 84876 116848 88206 116904
rect 88262 116848 88267 116904
rect 84876 116846 88267 116848
rect 156820 116904 159935 116906
rect 156820 116848 159874 116904
rect 159930 116848 159935 116904
rect 156820 116846 159935 116848
rect 88201 116843 88267 116846
rect 159869 116843 159935 116846
rect 47862 116498 47922 116808
rect 91470 116774 92052 116834
rect 88477 116770 88543 116773
rect 91470 116770 91530 116774
rect 88477 116768 91530 116770
rect 88477 116712 88482 116768
rect 88538 116712 91530 116768
rect 88477 116710 91530 116712
rect 88477 116707 88543 116710
rect 51217 116498 51283 116501
rect 47862 116496 51283 116498
rect 47862 116440 51222 116496
rect 51278 116440 51283 116496
rect 47862 116438 51283 116440
rect 119806 116498 119866 116808
rect 123069 116498 123135 116501
rect 119806 116496 123135 116498
rect 119806 116440 123074 116496
rect 123130 116440 123135 116496
rect 119806 116438 123135 116440
rect 51217 116435 51283 116438
rect 123069 116435 123135 116438
rect 160237 116498 160303 116501
rect 163966 116498 164026 116808
rect 160237 116496 164026 116498
rect 160237 116440 160242 116496
rect 160298 116440 164026 116496
rect 160237 116438 164026 116440
rect 160237 116435 160303 116438
rect 47862 115954 47922 116264
rect 91470 116230 92052 116290
rect 51401 116226 51467 116229
rect 88385 116226 88451 116229
rect 51401 116224 55068 116226
rect 51401 116168 51406 116224
rect 51462 116168 55068 116224
rect 51401 116166 55068 116168
rect 84876 116224 88451 116226
rect 84876 116168 88390 116224
rect 88446 116168 88451 116224
rect 84876 116166 88451 116168
rect 51401 116163 51467 116166
rect 88385 116163 88451 116166
rect 88569 116226 88635 116229
rect 91470 116226 91530 116230
rect 88569 116224 91530 116226
rect 88569 116168 88574 116224
rect 88630 116168 91530 116224
rect 88569 116166 91530 116168
rect 88569 116163 88635 116166
rect 51493 116090 51559 116093
rect 51493 116088 55098 116090
rect 51493 116032 51498 116088
rect 51554 116032 55098 116088
rect 51493 116030 55098 116032
rect 51493 116027 51559 116030
rect 51217 115954 51283 115957
rect 47862 115952 51283 115954
rect 47862 115896 51222 115952
rect 51278 115896 51283 115952
rect 47862 115894 51283 115896
rect 51217 115891 51283 115894
rect 55038 115720 55098 116030
rect 119806 115954 119866 116264
rect 124357 116226 124423 116229
rect 160053 116226 160119 116229
rect 124357 116224 127012 116226
rect 124357 116168 124362 116224
rect 124418 116168 127012 116224
rect 124357 116166 127012 116168
rect 156820 116224 160119 116226
rect 156820 116168 160058 116224
rect 160114 116168 160119 116224
rect 156820 116166 160119 116168
rect 124357 116163 124423 116166
rect 160053 116163 160119 116166
rect 123161 116090 123227 116093
rect 123161 116088 127042 116090
rect 123161 116032 123166 116088
rect 123222 116032 127042 116088
rect 123161 116030 127042 116032
rect 123161 116027 123227 116030
rect 121689 115954 121755 115957
rect 119806 115952 121755 115954
rect 119806 115896 121694 115952
rect 121750 115896 121755 115952
rect 119806 115894 121755 115896
rect 121689 115891 121755 115894
rect 47862 115410 47922 115720
rect 91470 115686 92052 115746
rect 126982 115720 127042 116030
rect 160329 115954 160395 115957
rect 163966 115954 164026 116264
rect 160329 115952 164026 115954
rect 160329 115896 160334 115952
rect 160390 115896 164026 115952
rect 160329 115894 164026 115896
rect 160329 115891 160395 115894
rect 88109 115682 88175 115685
rect 84876 115680 88175 115682
rect 84876 115624 88114 115680
rect 88170 115624 88175 115680
rect 84876 115622 88175 115624
rect 88109 115619 88175 115622
rect 88385 115682 88451 115685
rect 91470 115682 91530 115686
rect 88385 115680 91530 115682
rect 88385 115624 88390 115680
rect 88446 115624 91530 115680
rect 88385 115622 91530 115624
rect 88385 115619 88451 115622
rect 51585 115546 51651 115549
rect 119806 115546 119866 115720
rect 160145 115682 160211 115685
rect 156820 115680 160211 115682
rect 156820 115624 160150 115680
rect 160206 115624 160211 115680
rect 156820 115622 160211 115624
rect 160145 115619 160211 115622
rect 121689 115546 121755 115549
rect 51585 115544 55098 115546
rect 51585 115488 51590 115544
rect 51646 115488 55098 115544
rect 51585 115486 55098 115488
rect 119806 115544 121755 115546
rect 119806 115488 121694 115544
rect 121750 115488 121755 115544
rect 119806 115486 121755 115488
rect 51585 115483 51651 115486
rect 51401 115410 51467 115413
rect 47862 115408 51467 115410
rect 47862 115352 51406 115408
rect 51462 115352 51467 115408
rect 47862 115350 51467 115352
rect 51401 115347 51467 115350
rect 55038 115176 55098 115486
rect 121689 115483 121755 115486
rect 124265 115546 124331 115549
rect 124265 115544 127042 115546
rect 124265 115488 124270 115544
rect 124326 115488 127042 115544
rect 124265 115486 127042 115488
rect 124265 115483 124331 115486
rect 88201 115274 88267 115277
rect 88201 115272 91530 115274
rect 88201 115216 88206 115272
rect 88262 115216 91530 115272
rect 88201 115214 91530 115216
rect 88201 115211 88267 115214
rect 91470 115206 91530 115214
rect 47862 115138 47922 115176
rect 91470 115146 92052 115206
rect 126982 115176 127042 115486
rect 160053 115410 160119 115413
rect 163966 115410 164026 115720
rect 160053 115408 164026 115410
rect 160053 115352 160058 115408
rect 160114 115352 164026 115408
rect 160053 115350 164026 115352
rect 160053 115347 160119 115350
rect 51493 115138 51559 115141
rect 88661 115138 88727 115141
rect 47862 115136 51559 115138
rect 47862 115080 51498 115136
rect 51554 115080 51559 115136
rect 47862 115078 51559 115080
rect 84876 115136 88727 115138
rect 84876 115080 88666 115136
rect 88722 115080 88727 115136
rect 84876 115078 88727 115080
rect 119806 115138 119866 115176
rect 121689 115138 121755 115141
rect 160421 115138 160487 115141
rect 119806 115136 121755 115138
rect 119806 115080 121694 115136
rect 121750 115080 121755 115136
rect 119806 115078 121755 115080
rect 156820 115136 160487 115138
rect 156820 115080 160426 115136
rect 160482 115080 160487 115136
rect 156820 115078 160487 115080
rect 51493 115075 51559 115078
rect 88661 115075 88727 115078
rect 121689 115075 121755 115078
rect 160421 115075 160487 115078
rect 160605 115138 160671 115141
rect 163966 115138 164026 115176
rect 160605 115136 164026 115138
rect 160605 115080 160610 115136
rect 160666 115080 164026 115136
rect 160605 115078 164026 115080
rect 160605 115075 160671 115078
rect 51309 115002 51375 115005
rect 88477 115002 88543 115005
rect 51309 115000 55098 115002
rect 51309 114944 51314 115000
rect 51370 114944 55098 115000
rect 51309 114942 55098 114944
rect 51309 114939 51375 114942
rect 18005 114186 18071 114189
rect 19894 114186 19954 114768
rect 55038 114496 55098 114942
rect 84846 115000 88543 115002
rect 84846 114944 88482 115000
rect 88538 114944 88543 115000
rect 84846 114942 88543 114944
rect 18005 114184 19954 114186
rect 18005 114128 18010 114184
rect 18066 114128 19954 114184
rect 18005 114126 19954 114128
rect 47862 114186 47922 114496
rect 84846 114428 84906 114942
rect 88477 114939 88543 114942
rect 123069 115002 123135 115005
rect 123069 115000 127042 115002
rect 123069 114944 123074 115000
rect 123130 114944 127042 115000
rect 123069 114942 127042 114944
rect 123069 114939 123135 114942
rect 91470 114462 92052 114522
rect 126982 114496 127042 114942
rect 191558 114940 191564 115004
rect 191628 114940 191634 115004
rect 191566 114768 191626 114940
rect 201269 114730 201335 114733
rect 201416 114730 201896 114760
rect 201269 114728 201896 114730
rect 201269 114672 201274 114728
rect 201330 114672 201896 114728
rect 201269 114670 201896 114672
rect 201269 114667 201335 114670
rect 201416 114640 201896 114670
rect 191742 114532 191748 114596
rect 191812 114594 191818 114596
rect 201269 114594 201335 114597
rect 191812 114592 201335 114594
rect 191812 114536 201274 114592
rect 201330 114536 201335 114592
rect 191812 114534 201335 114536
rect 191812 114532 191818 114534
rect 201269 114531 201335 114534
rect 88293 114458 88359 114461
rect 91470 114458 91530 114462
rect 88293 114456 91530 114458
rect 88293 114400 88298 114456
rect 88354 114400 91530 114456
rect 88293 114398 91530 114400
rect 88293 114395 88359 114398
rect 51309 114322 51375 114325
rect 88477 114322 88543 114325
rect 51309 114320 55098 114322
rect 51309 114264 51314 114320
rect 51370 114264 55098 114320
rect 51309 114262 55098 114264
rect 51309 114259 51375 114262
rect 51309 114186 51375 114189
rect 47862 114184 51375 114186
rect 47862 114128 51314 114184
rect 51370 114128 51375 114184
rect 47862 114126 51375 114128
rect 18005 114123 18071 114126
rect 51309 114123 51375 114126
rect 55038 113952 55098 114262
rect 84846 114320 88543 114322
rect 84846 114264 88482 114320
rect 88538 114264 88543 114320
rect 84846 114262 88543 114264
rect 119806 114322 119866 114496
rect 160237 114458 160303 114461
rect 156820 114456 160303 114458
rect 156820 114400 160242 114456
rect 160298 114400 160303 114456
rect 156820 114398 160303 114400
rect 160237 114395 160303 114398
rect 121689 114322 121755 114325
rect 119806 114320 121755 114322
rect 119806 114264 121694 114320
rect 121750 114264 121755 114320
rect 119806 114262 121755 114264
rect 47862 113778 47922 113952
rect 84846 113884 84906 114262
rect 88477 114259 88543 114262
rect 121689 114259 121755 114262
rect 124357 114322 124423 114325
rect 160237 114322 160303 114325
rect 124357 114320 127042 114322
rect 124357 114264 124362 114320
rect 124418 114264 127042 114320
rect 124357 114262 127042 114264
rect 124357 114259 124423 114262
rect 91470 113918 92052 113978
rect 126982 113952 127042 114262
rect 156790 114320 160303 114322
rect 156790 114264 160242 114320
rect 160298 114264 160303 114320
rect 156790 114262 160303 114264
rect 88109 113914 88175 113917
rect 91470 113914 91530 113918
rect 88109 113912 91530 113914
rect 88109 113856 88114 113912
rect 88170 113856 91530 113912
rect 88109 113854 91530 113856
rect 88109 113851 88175 113854
rect 51585 113778 51651 113781
rect 47862 113776 51651 113778
rect 47862 113720 51590 113776
rect 51646 113720 51651 113776
rect 47862 113718 51651 113720
rect 119806 113778 119866 113952
rect 156790 113884 156850 114262
rect 160237 114259 160303 114262
rect 160237 114186 160303 114189
rect 163966 114186 164026 114496
rect 160237 114184 164026 114186
rect 160237 114128 160242 114184
rect 160298 114128 164026 114184
rect 160237 114126 164026 114128
rect 160237 114123 160303 114126
rect 122977 113778 123043 113781
rect 119806 113776 123043 113778
rect 119806 113720 122982 113776
rect 123038 113720 123043 113776
rect 119806 113718 123043 113720
rect 51585 113715 51651 113718
rect 122977 113715 123043 113718
rect 160145 113778 160211 113781
rect 163966 113778 164026 113952
rect 160145 113776 164026 113778
rect 160145 113720 160150 113776
rect 160206 113720 164026 113776
rect 160145 113718 164026 113720
rect 160145 113715 160211 113718
rect 51401 113642 51467 113645
rect 123989 113642 124055 113645
rect 51401 113640 55098 113642
rect 51401 113584 51406 113640
rect 51462 113584 55098 113640
rect 51401 113582 55098 113584
rect 51401 113579 51467 113582
rect 47862 112962 47922 113408
rect 55038 113272 55098 113582
rect 123989 113640 127042 113642
rect 123989 113584 123994 113640
rect 124050 113584 127042 113640
rect 123989 113582 127042 113584
rect 123989 113579 124055 113582
rect 91470 113374 92052 113434
rect 88017 113370 88083 113373
rect 91470 113370 91530 113374
rect 88017 113368 91530 113370
rect 88017 113312 88022 113368
rect 88078 113312 91530 113368
rect 88017 113310 91530 113312
rect 88017 113307 88083 113310
rect 88385 113234 88451 113237
rect 84876 113232 88451 113234
rect 84876 113176 88390 113232
rect 88446 113176 88451 113232
rect 84876 113174 88451 113176
rect 88385 113171 88451 113174
rect 51493 113098 51559 113101
rect 51493 113096 55098 113098
rect 51493 113040 51498 113096
rect 51554 113040 55098 113096
rect 51493 113038 55098 113040
rect 51493 113035 51559 113038
rect 51217 112962 51283 112965
rect 47862 112960 51283 112962
rect 47862 112904 51222 112960
rect 51278 112904 51283 112960
rect 47862 112902 51283 112904
rect 51217 112899 51283 112902
rect 55038 112728 55098 113038
rect 119806 112962 119866 113408
rect 126982 113272 127042 113582
rect 160053 113234 160119 113237
rect 156820 113232 160119 113234
rect 156820 113176 160058 113232
rect 160114 113176 160119 113232
rect 156820 113174 160119 113176
rect 160053 113171 160119 113174
rect 124265 113098 124331 113101
rect 124265 113096 127042 113098
rect 124265 113040 124270 113096
rect 124326 113040 127042 113096
rect 124265 113038 127042 113040
rect 124265 113035 124331 113038
rect 123253 112962 123319 112965
rect 119806 112960 123319 112962
rect 119806 112904 123258 112960
rect 123314 112904 123319 112960
rect 119806 112902 123319 112904
rect 123253 112899 123319 112902
rect 47862 112554 47922 112728
rect 91470 112694 92052 112754
rect 126982 112728 127042 113038
rect 159961 112962 160027 112965
rect 163966 112962 164026 113408
rect 159961 112960 164026 112962
rect 159961 112904 159966 112960
rect 160022 112904 164026 112960
rect 159961 112902 164026 112904
rect 159961 112899 160027 112902
rect 88201 112690 88267 112693
rect 84876 112688 88267 112690
rect 84876 112632 88206 112688
rect 88262 112632 88267 112688
rect 84876 112630 88267 112632
rect 88201 112627 88267 112630
rect 88477 112690 88543 112693
rect 91470 112690 91530 112694
rect 88477 112688 91530 112690
rect 88477 112632 88482 112688
rect 88538 112632 91530 112688
rect 88477 112630 91530 112632
rect 88477 112627 88543 112630
rect 51493 112554 51559 112557
rect 47862 112552 51559 112554
rect 47862 112496 51498 112552
rect 51554 112496 51559 112552
rect 47862 112494 51559 112496
rect 119806 112554 119866 112728
rect 159041 112690 159107 112693
rect 156820 112688 159107 112690
rect 156820 112632 159046 112688
rect 159102 112632 159107 112688
rect 156820 112630 159107 112632
rect 159041 112627 159107 112630
rect 121689 112554 121755 112557
rect 119806 112552 121755 112554
rect 119806 112496 121694 112552
rect 121750 112496 121755 112552
rect 119806 112494 121755 112496
rect 51493 112491 51559 112494
rect 121689 112491 121755 112494
rect 160053 112418 160119 112421
rect 163966 112418 164026 112728
rect 160053 112416 164026 112418
rect 160053 112360 160058 112416
rect 160114 112360 164026 112416
rect 160053 112358 164026 112360
rect 160053 112355 160119 112358
rect 51309 112282 51375 112285
rect 51309 112280 54546 112282
rect 51309 112224 51314 112280
rect 51370 112224 54546 112280
rect 51309 112222 54546 112224
rect 51309 112219 51375 112222
rect 54486 112214 54546 112222
rect 47862 111874 47922 112184
rect 54486 112154 55068 112214
rect 91470 112150 92052 112210
rect 88293 112146 88359 112149
rect 84876 112144 88359 112146
rect 84876 112088 88298 112144
rect 88354 112088 88359 112144
rect 84876 112086 88359 112088
rect 88293 112083 88359 112086
rect 88661 112146 88727 112149
rect 91470 112146 91530 112150
rect 88661 112144 91530 112146
rect 88661 112088 88666 112144
rect 88722 112088 91530 112144
rect 88661 112086 91530 112088
rect 88661 112083 88727 112086
rect 51585 112010 51651 112013
rect 51585 112008 55098 112010
rect 51585 111952 51590 112008
rect 51646 111952 55098 112008
rect 51585 111950 55098 111952
rect 51585 111947 51651 111950
rect 51217 111874 51283 111877
rect 47862 111872 51283 111874
rect 47862 111816 51222 111872
rect 51278 111816 51283 111872
rect 47862 111814 51283 111816
rect 51217 111811 51283 111814
rect 47862 111194 47922 111640
rect 55038 111504 55098 111950
rect 119806 111874 119866 112184
rect 123437 112146 123503 112149
rect 160237 112146 160303 112149
rect 123437 112144 127012 112146
rect 123437 112088 123442 112144
rect 123498 112088 127012 112144
rect 123437 112086 127012 112088
rect 156820 112144 160303 112146
rect 156820 112088 160242 112144
rect 160298 112088 160303 112144
rect 156820 112086 160303 112088
rect 123437 112083 123503 112086
rect 160237 112083 160303 112086
rect 122977 111874 123043 111877
rect 119806 111872 123043 111874
rect 119806 111816 122982 111872
rect 123038 111816 123043 111872
rect 119806 111814 123043 111816
rect 122977 111811 123043 111814
rect 123161 111874 123227 111877
rect 160329 111874 160395 111877
rect 163966 111874 164026 112184
rect 123161 111872 127042 111874
rect 123161 111816 123166 111872
rect 123222 111816 127042 111872
rect 123161 111814 127042 111816
rect 123161 111811 123227 111814
rect 91470 111606 92052 111666
rect 88293 111602 88359 111605
rect 91470 111602 91530 111606
rect 88293 111600 91530 111602
rect 88293 111544 88298 111600
rect 88354 111544 91530 111600
rect 88293 111542 91530 111544
rect 88293 111539 88359 111542
rect 88109 111466 88175 111469
rect 84876 111464 88175 111466
rect 84876 111408 88114 111464
rect 88170 111408 88175 111464
rect 84876 111406 88175 111408
rect 88109 111403 88175 111406
rect 119806 111330 119866 111640
rect 126982 111504 127042 111814
rect 160329 111872 164026 111874
rect 160329 111816 160334 111872
rect 160390 111816 164026 111872
rect 160329 111814 164026 111816
rect 160329 111811 160395 111814
rect 160145 111466 160211 111469
rect 156820 111464 160211 111466
rect 156820 111408 160150 111464
rect 160206 111408 160211 111464
rect 156820 111406 160211 111408
rect 160145 111403 160211 111406
rect 121689 111330 121755 111333
rect 119806 111328 121755 111330
rect 119806 111272 121694 111328
rect 121750 111272 121755 111328
rect 119806 111270 121755 111272
rect 121689 111267 121755 111270
rect 51217 111194 51283 111197
rect 47862 111192 51283 111194
rect 47862 111136 51222 111192
rect 51278 111136 51283 111192
rect 47862 111134 51283 111136
rect 51217 111131 51283 111134
rect 160237 111194 160303 111197
rect 163966 111194 164026 111640
rect 160237 111192 164026 111194
rect 160237 111136 160242 111192
rect 160298 111136 164026 111192
rect 160237 111134 164026 111136
rect 160237 111131 160303 111134
rect 51217 111058 51283 111061
rect 47862 111056 51283 111058
rect 47862 111000 51222 111056
rect 51278 111000 51283 111056
rect 47862 110998 51283 111000
rect 47862 110960 47922 110998
rect 51217 110995 51283 110998
rect 88385 111058 88451 111061
rect 123161 111058 123227 111061
rect 88385 111056 91530 111058
rect 88385 111000 88390 111056
rect 88446 111000 91530 111056
rect 88385 110998 91530 111000
rect 88385 110995 88451 110998
rect 91470 110990 91530 110998
rect 119806 111056 123227 111058
rect 119806 111000 123166 111056
rect 123222 111000 123227 111056
rect 119806 110998 123227 111000
rect 91470 110930 92052 110990
rect 119806 110960 119866 110998
rect 123161 110995 123227 110998
rect 159869 111058 159935 111061
rect 159869 111056 164026 111058
rect 159869 111000 159874 111056
rect 159930 111000 164026 111056
rect 159869 110998 164026 111000
rect 159869 110995 159935 110998
rect 163966 110960 164026 110998
rect 51309 110922 51375 110925
rect 88017 110922 88083 110925
rect 51309 110920 55068 110922
rect 51309 110864 51314 110920
rect 51370 110864 55068 110920
rect 51309 110862 55068 110864
rect 84876 110920 88083 110922
rect 84876 110864 88022 110920
rect 88078 110864 88083 110920
rect 84876 110862 88083 110864
rect 51309 110859 51375 110862
rect 88017 110859 88083 110862
rect 123253 110922 123319 110925
rect 159961 110922 160027 110925
rect 123253 110920 127012 110922
rect 123253 110864 123258 110920
rect 123314 110864 127012 110920
rect 123253 110862 127012 110864
rect 156820 110920 160027 110922
rect 156820 110864 159966 110920
rect 160022 110864 160027 110920
rect 156820 110862 160027 110864
rect 123253 110859 123319 110862
rect 159961 110859 160027 110862
rect 51493 110786 51559 110789
rect 123345 110786 123411 110789
rect 51493 110784 55098 110786
rect 51493 110728 51498 110784
rect 51554 110728 55098 110784
rect 51493 110726 55098 110728
rect 51493 110723 51559 110726
rect 47862 110106 47922 110416
rect 55038 110280 55098 110726
rect 123345 110784 127042 110786
rect 123345 110728 123350 110784
rect 123406 110728 127042 110784
rect 123345 110726 127042 110728
rect 123345 110723 123411 110726
rect 91470 110382 92052 110442
rect 88569 110378 88635 110381
rect 91470 110378 91530 110382
rect 88569 110376 91530 110378
rect 88569 110320 88574 110376
rect 88630 110320 91530 110376
rect 88569 110318 91530 110320
rect 88569 110315 88635 110318
rect 88477 110242 88543 110245
rect 84876 110240 88543 110242
rect 84876 110184 88482 110240
rect 88538 110184 88543 110240
rect 84876 110182 88543 110184
rect 88477 110179 88543 110182
rect 51401 110106 51467 110109
rect 47862 110104 51467 110106
rect 47862 110048 51406 110104
rect 51462 110048 51467 110104
rect 47862 110046 51467 110048
rect 51401 110043 51467 110046
rect 51585 110106 51651 110109
rect 119806 110106 119866 110416
rect 126982 110280 127042 110726
rect 160053 110242 160119 110245
rect 156820 110240 160119 110242
rect 156820 110184 160058 110240
rect 160114 110184 160119 110240
rect 156820 110182 160119 110184
rect 160053 110179 160119 110182
rect 121689 110106 121755 110109
rect 51585 110104 55098 110106
rect 51585 110048 51590 110104
rect 51646 110048 55098 110104
rect 51585 110046 55098 110048
rect 119806 110104 121755 110106
rect 119806 110048 121694 110104
rect 121750 110048 121755 110104
rect 119806 110046 121755 110048
rect 51585 110043 51651 110046
rect 47862 109698 47922 109872
rect 55038 109736 55098 110046
rect 121689 110043 121755 110046
rect 123069 110106 123135 110109
rect 160145 110106 160211 110109
rect 163966 110106 164026 110416
rect 123069 110104 127042 110106
rect 123069 110048 123074 110104
rect 123130 110048 127042 110104
rect 123069 110046 127042 110048
rect 123069 110043 123135 110046
rect 91470 109838 92052 109898
rect 88201 109834 88267 109837
rect 91470 109834 91530 109838
rect 88201 109832 91530 109834
rect 88201 109776 88206 109832
rect 88262 109776 91530 109832
rect 88201 109774 91530 109776
rect 88201 109771 88267 109774
rect 51493 109698 51559 109701
rect 88661 109698 88727 109701
rect 47862 109696 51559 109698
rect 47862 109640 51498 109696
rect 51554 109640 51559 109696
rect 47862 109638 51559 109640
rect 84876 109696 88727 109698
rect 84876 109640 88666 109696
rect 88722 109640 88727 109696
rect 84876 109638 88727 109640
rect 119806 109698 119866 109872
rect 126982 109736 127042 110046
rect 160145 110104 164026 110106
rect 160145 110048 160150 110104
rect 160206 110048 164026 110104
rect 160145 110046 164026 110048
rect 160145 110043 160211 110046
rect 159961 109834 160027 109837
rect 163966 109834 164026 109872
rect 159961 109832 164026 109834
rect 159961 109776 159966 109832
rect 160022 109776 164026 109832
rect 159961 109774 164026 109776
rect 159961 109771 160027 109774
rect 122977 109698 123043 109701
rect 160329 109698 160395 109701
rect 119806 109696 123043 109698
rect 119806 109640 122982 109696
rect 123038 109640 123043 109696
rect 119806 109638 123043 109640
rect 156820 109696 160395 109698
rect 156820 109640 160334 109696
rect 160390 109640 160395 109696
rect 156820 109638 160395 109640
rect 51493 109635 51559 109638
rect 88661 109635 88727 109638
rect 122977 109635 123043 109638
rect 160329 109635 160395 109638
rect 51677 109562 51743 109565
rect 124265 109562 124331 109565
rect 51677 109560 55098 109562
rect 51677 109504 51682 109560
rect 51738 109504 55098 109560
rect 51677 109502 55098 109504
rect 51677 109499 51743 109502
rect 47862 108882 47922 109328
rect 55038 109192 55098 109502
rect 124265 109560 127042 109562
rect 124265 109504 124270 109560
rect 124326 109504 127042 109560
rect 124265 109502 127042 109504
rect 124265 109499 124331 109502
rect 91470 109294 92052 109354
rect 88109 109290 88175 109293
rect 91470 109290 91530 109294
rect 88109 109288 91530 109290
rect 88109 109232 88114 109288
rect 88170 109232 91530 109288
rect 88109 109230 91530 109232
rect 88109 109227 88175 109230
rect 88293 109154 88359 109157
rect 84876 109152 88359 109154
rect 84876 109096 88298 109152
rect 88354 109096 88359 109152
rect 84876 109094 88359 109096
rect 88293 109091 88359 109094
rect 51309 109018 51375 109021
rect 119806 109018 119866 109328
rect 126982 109192 127042 109502
rect 160237 109154 160303 109157
rect 156820 109152 160303 109154
rect 156820 109096 160242 109152
rect 160298 109096 160303 109152
rect 156820 109094 160303 109096
rect 160237 109091 160303 109094
rect 121689 109018 121755 109021
rect 51309 109016 55098 109018
rect 51309 108960 51314 109016
rect 51370 108960 55098 109016
rect 51309 108958 55098 108960
rect 119806 109016 121755 109018
rect 119806 108960 121694 109016
rect 121750 108960 121755 109016
rect 119806 108958 121755 108960
rect 51309 108955 51375 108958
rect 51217 108882 51283 108885
rect 47862 108880 51283 108882
rect 47862 108824 51222 108880
rect 51278 108824 51283 108880
rect 47862 108822 51283 108824
rect 51217 108819 51283 108822
rect 47862 108338 47922 108648
rect 55038 108512 55098 108958
rect 121689 108955 121755 108958
rect 123253 109018 123319 109021
rect 123253 109016 127042 109018
rect 123253 108960 123258 109016
rect 123314 108960 127042 109016
rect 123253 108958 127042 108960
rect 123253 108955 123319 108958
rect 91470 108614 92052 108674
rect 88293 108610 88359 108613
rect 91470 108610 91530 108614
rect 88293 108608 91530 108610
rect 88293 108552 88298 108608
rect 88354 108552 91530 108608
rect 88293 108550 91530 108552
rect 88293 108547 88359 108550
rect 88385 108474 88451 108477
rect 84876 108472 88451 108474
rect 84876 108416 88390 108472
rect 88446 108416 88451 108472
rect 84876 108414 88451 108416
rect 119806 108474 119866 108648
rect 126982 108512 127042 108958
rect 160053 108882 160119 108885
rect 163966 108882 164026 109328
rect 160053 108880 164026 108882
rect 160053 108824 160058 108880
rect 160114 108824 164026 108880
rect 160053 108822 164026 108824
rect 160053 108819 160119 108822
rect 123253 108474 123319 108477
rect 159869 108474 159935 108477
rect 119806 108472 123319 108474
rect 119806 108416 123258 108472
rect 123314 108416 123319 108472
rect 119806 108414 123319 108416
rect 156820 108472 159935 108474
rect 156820 108416 159874 108472
rect 159930 108416 159935 108472
rect 156820 108414 159935 108416
rect 88385 108411 88451 108414
rect 123253 108411 123319 108414
rect 159869 108411 159935 108414
rect 51217 108338 51283 108341
rect 47862 108336 51283 108338
rect 47862 108280 51222 108336
rect 51278 108280 51283 108336
rect 47862 108278 51283 108280
rect 51217 108275 51283 108278
rect 160237 108338 160303 108341
rect 163966 108338 164026 108648
rect 160237 108336 164026 108338
rect 160237 108280 160242 108336
rect 160298 108280 164026 108336
rect 160237 108278 164026 108280
rect 160237 108275 160303 108278
rect 51401 108202 51467 108205
rect 124357 108202 124423 108205
rect 51401 108200 55098 108202
rect 51401 108144 51406 108200
rect 51462 108144 55098 108200
rect 51401 108142 55098 108144
rect 51401 108139 51467 108142
rect 47862 107930 47922 108104
rect 55038 107968 55098 108142
rect 124357 108200 127042 108202
rect 124357 108144 124362 108200
rect 124418 108144 127042 108200
rect 124357 108142 127042 108144
rect 124357 108139 124423 108142
rect 91470 108070 92052 108130
rect 88569 108066 88635 108069
rect 91470 108066 91530 108070
rect 88569 108064 91530 108066
rect 88569 108008 88574 108064
rect 88630 108008 91530 108064
rect 88569 108006 91530 108008
rect 88569 108003 88635 108006
rect 51401 107930 51467 107933
rect 88477 107930 88543 107933
rect 47862 107928 51467 107930
rect 47862 107872 51406 107928
rect 51462 107872 51467 107928
rect 47862 107870 51467 107872
rect 84876 107928 88543 107930
rect 84876 107872 88482 107928
rect 88538 107872 88543 107928
rect 84876 107870 88543 107872
rect 51401 107867 51467 107870
rect 88477 107867 88543 107870
rect 51493 107794 51559 107797
rect 119806 107794 119866 108104
rect 126982 107968 127042 108142
rect 160145 107930 160211 107933
rect 156820 107928 160211 107930
rect 156820 107872 160150 107928
rect 160206 107872 160211 107928
rect 156820 107870 160211 107872
rect 160145 107867 160211 107870
rect 122977 107794 123043 107797
rect 51493 107792 55098 107794
rect 51493 107736 51498 107792
rect 51554 107736 55098 107792
rect 51493 107734 55098 107736
rect 119806 107792 123043 107794
rect 119806 107736 122982 107792
rect 123038 107736 123043 107792
rect 119806 107734 123043 107736
rect 51493 107731 51559 107734
rect 47862 107114 47922 107560
rect 55038 107288 55098 107734
rect 122977 107731 123043 107734
rect 123161 107794 123227 107797
rect 160329 107794 160395 107797
rect 163966 107794 164026 108104
rect 123161 107792 127042 107794
rect 123161 107736 123166 107792
rect 123222 107736 127042 107792
rect 123161 107734 127042 107736
rect 123161 107731 123227 107734
rect 91470 107526 92052 107586
rect 88017 107522 88083 107525
rect 91470 107522 91530 107526
rect 88017 107520 91530 107522
rect 88017 107464 88022 107520
rect 88078 107464 91530 107520
rect 88017 107462 91530 107464
rect 88017 107459 88083 107462
rect 88201 107250 88267 107253
rect 84876 107248 88267 107250
rect 84876 107192 88206 107248
rect 88262 107192 88267 107248
rect 84876 107190 88267 107192
rect 119806 107250 119866 107560
rect 126982 107288 127042 107734
rect 160329 107792 164026 107794
rect 160329 107736 160334 107792
rect 160390 107736 164026 107792
rect 160329 107734 164026 107736
rect 160329 107731 160395 107734
rect 121689 107250 121755 107253
rect 159961 107250 160027 107253
rect 119806 107248 121755 107250
rect 119806 107192 121694 107248
rect 121750 107192 121755 107248
rect 119806 107190 121755 107192
rect 156820 107248 160027 107250
rect 156820 107192 159966 107248
rect 160022 107192 160027 107248
rect 156820 107190 160027 107192
rect 88201 107187 88267 107190
rect 121689 107187 121755 107190
rect 159961 107187 160027 107190
rect 51217 107114 51283 107117
rect 47862 107112 51283 107114
rect 47862 107056 51222 107112
rect 51278 107056 51283 107112
rect 47862 107054 51283 107056
rect 51217 107051 51283 107054
rect 160145 107114 160211 107117
rect 163966 107114 164026 107560
rect 160145 107112 164026 107114
rect 160145 107056 160150 107112
rect 160206 107056 164026 107112
rect 160145 107054 164026 107056
rect 160145 107051 160211 107054
rect 47862 106842 47922 106880
rect 91470 106846 92052 106906
rect 51493 106842 51559 106845
rect 47862 106840 51559 106842
rect 47862 106784 51498 106840
rect 51554 106784 51559 106840
rect 47862 106782 51559 106784
rect 51493 106779 51559 106782
rect 85165 106844 85231 106845
rect 85165 106840 85212 106844
rect 85276 106842 85282 106844
rect 88477 106842 88543 106845
rect 91470 106842 91530 106846
rect 85165 106784 85170 106840
rect 85165 106780 85212 106784
rect 85276 106782 85322 106842
rect 88477 106840 91530 106842
rect 88477 106784 88482 106840
rect 88538 106784 91530 106840
rect 88477 106782 91530 106784
rect 119806 106842 119866 106880
rect 123069 106842 123135 106845
rect 119806 106840 123135 106842
rect 119806 106784 123074 106840
rect 123130 106784 123135 106840
rect 119806 106782 123135 106784
rect 85276 106780 85282 106782
rect 85165 106779 85231 106780
rect 88477 106779 88543 106782
rect 123069 106779 123135 106782
rect 159869 106842 159935 106845
rect 163966 106842 164026 106880
rect 159869 106840 164026 106842
rect 159869 106784 159874 106840
rect 159930 106784 164026 106840
rect 159869 106782 164026 106784
rect 159869 106779 159935 106782
rect 51585 106706 51651 106709
rect 88109 106706 88175 106709
rect 51585 106704 55068 106706
rect 51585 106648 51590 106704
rect 51646 106648 55068 106704
rect 51585 106646 55068 106648
rect 84876 106704 88175 106706
rect 84876 106648 88114 106704
rect 88170 106648 88175 106704
rect 84876 106646 88175 106648
rect 51585 106643 51651 106646
rect 88109 106643 88175 106646
rect 123437 106706 123503 106709
rect 160053 106706 160119 106709
rect 123437 106704 127012 106706
rect 123437 106648 123442 106704
rect 123498 106648 127012 106704
rect 123437 106646 127012 106648
rect 156820 106704 160119 106706
rect 156820 106648 160058 106704
rect 160114 106648 160119 106704
rect 156820 106646 160119 106648
rect 123437 106643 123503 106646
rect 160053 106643 160119 106646
rect 51309 106570 51375 106573
rect 123253 106570 123319 106573
rect 51309 106568 55098 106570
rect 51309 106512 51314 106568
rect 51370 106512 55098 106568
rect 51309 106510 55098 106512
rect 51309 106507 51375 106510
rect 19886 106100 19892 106164
rect 19956 106100 19962 106164
rect 19894 105520 19954 106100
rect 47862 106026 47922 106336
rect 55038 106200 55098 106510
rect 123253 106568 127042 106570
rect 123253 106512 123258 106568
rect 123314 106512 127042 106568
rect 123253 106510 127042 106512
rect 123253 106507 123319 106510
rect 91470 106302 92052 106362
rect 88385 106298 88451 106301
rect 91470 106298 91530 106302
rect 88385 106296 91530 106298
rect 88385 106240 88390 106296
rect 88446 106240 91530 106296
rect 88385 106238 91530 106240
rect 88385 106235 88451 106238
rect 88293 106162 88359 106165
rect 84876 106160 88359 106162
rect 84876 106104 88298 106160
rect 88354 106104 88359 106160
rect 84876 106102 88359 106104
rect 119806 106162 119866 106336
rect 126982 106200 127042 106510
rect 121689 106162 121755 106165
rect 160237 106162 160303 106165
rect 119806 106160 121755 106162
rect 119806 106104 121694 106160
rect 121750 106104 121755 106160
rect 119806 106102 121755 106104
rect 156820 106160 160303 106162
rect 156820 106104 160242 106160
rect 160298 106104 160303 106160
rect 156820 106102 160303 106104
rect 88293 106099 88359 106102
rect 121689 106099 121755 106102
rect 160237 106099 160303 106102
rect 51217 106026 51283 106029
rect 47862 106024 51283 106026
rect 47862 105968 51222 106024
rect 51278 105968 51283 106024
rect 47862 105966 51283 105968
rect 51217 105963 51283 105966
rect 51401 106026 51467 106029
rect 123161 106026 123227 106029
rect 160053 106026 160119 106029
rect 163966 106026 164026 106336
rect 193449 106162 193515 106165
rect 51401 106024 55098 106026
rect 51401 105968 51406 106024
rect 51462 105968 55098 106024
rect 51401 105966 55098 105968
rect 51401 105963 51467 105966
rect 47862 105482 47922 105792
rect 55038 105520 55098 105966
rect 123161 106024 127042 106026
rect 123161 105968 123166 106024
rect 123222 105968 127042 106024
rect 123161 105966 127042 105968
rect 123161 105963 123227 105966
rect 91470 105758 92052 105818
rect 88293 105754 88359 105757
rect 91470 105754 91530 105758
rect 88293 105752 91530 105754
rect 88293 105696 88298 105752
rect 88354 105696 91530 105752
rect 88293 105694 91530 105696
rect 119806 105754 119866 105792
rect 121689 105754 121755 105757
rect 119806 105752 121755 105754
rect 119806 105696 121694 105752
rect 121750 105696 121755 105752
rect 119806 105694 121755 105696
rect 88293 105691 88359 105694
rect 121689 105691 121755 105694
rect 126982 105520 127042 105966
rect 160053 106024 164026 106026
rect 160053 105968 160058 106024
rect 160114 105968 164026 106024
rect 160053 105966 164026 105968
rect 191750 106160 193515 106162
rect 191750 106104 193454 106160
rect 193510 106104 193515 106160
rect 191750 106102 193515 106104
rect 160053 105963 160119 105966
rect 159961 105618 160027 105621
rect 163966 105618 164026 105792
rect 159961 105616 164026 105618
rect 159961 105560 159966 105616
rect 160022 105560 164026 105616
rect 159961 105558 164026 105560
rect 159961 105555 160027 105558
rect 191750 105520 191810 106102
rect 193449 106099 193515 106102
rect 51401 105482 51467 105485
rect 88569 105482 88635 105485
rect 160237 105482 160303 105485
rect 47862 105480 51467 105482
rect 47862 105424 51406 105480
rect 51462 105424 51467 105480
rect 47862 105422 51467 105424
rect 84876 105480 88635 105482
rect 84876 105424 88574 105480
rect 88630 105424 88635 105480
rect 84876 105422 88635 105424
rect 156820 105480 160303 105482
rect 156820 105424 160242 105480
rect 160298 105424 160303 105480
rect 156820 105422 160303 105424
rect 51401 105419 51467 105422
rect 88569 105419 88635 105422
rect 160237 105419 160303 105422
rect 51309 105346 51375 105349
rect 124265 105346 124331 105349
rect 51309 105344 55098 105346
rect 51309 105288 51314 105344
rect 51370 105288 55098 105344
rect 51309 105286 55098 105288
rect 51309 105283 51375 105286
rect 47862 104802 47922 105248
rect 55038 104976 55098 105286
rect 124265 105344 127042 105346
rect 124265 105288 124270 105344
rect 124326 105288 127042 105344
rect 124265 105286 127042 105288
rect 124265 105283 124331 105286
rect 91470 105214 92052 105274
rect 88661 105210 88727 105213
rect 91470 105210 91530 105214
rect 88661 105208 91530 105210
rect 88661 105152 88666 105208
rect 88722 105152 91530 105208
rect 88661 105150 91530 105152
rect 88661 105147 88727 105150
rect 88017 104938 88083 104941
rect 84876 104936 88083 104938
rect 84876 104880 88022 104936
rect 88078 104880 88083 104936
rect 84876 104878 88083 104880
rect 88017 104875 88083 104878
rect 50665 104802 50731 104805
rect 47862 104800 50731 104802
rect 47862 104744 50670 104800
rect 50726 104744 50731 104800
rect 47862 104742 50731 104744
rect 50665 104739 50731 104742
rect 51493 104802 51559 104805
rect 119806 104802 119866 105248
rect 126982 104976 127042 105286
rect 160145 104938 160211 104941
rect 156820 104936 160211 104938
rect 156820 104880 160150 104936
rect 160206 104880 160211 104936
rect 156820 104878 160211 104880
rect 160145 104875 160211 104878
rect 121781 104802 121847 104805
rect 51493 104800 55098 104802
rect 51493 104744 51498 104800
rect 51554 104744 55098 104800
rect 51493 104742 55098 104744
rect 119806 104800 121847 104802
rect 119806 104744 121786 104800
rect 121842 104744 121847 104800
rect 119806 104742 121847 104744
rect 51493 104739 51559 104742
rect 47862 104258 47922 104568
rect 55038 104296 55098 104742
rect 121781 104739 121847 104742
rect 123069 104802 123135 104805
rect 161525 104802 161591 104805
rect 163966 104802 164026 105248
rect 123069 104800 127042 104802
rect 123069 104744 123074 104800
rect 123130 104744 127042 104800
rect 123069 104742 127042 104744
rect 123069 104739 123135 104742
rect 91470 104534 92052 104594
rect 88569 104530 88635 104533
rect 91470 104530 91530 104534
rect 88569 104528 91530 104530
rect 88569 104472 88574 104528
rect 88630 104472 91530 104528
rect 88569 104470 91530 104472
rect 88569 104467 88635 104470
rect 119806 104394 119866 104568
rect 121689 104394 121755 104397
rect 119806 104392 121755 104394
rect 119806 104336 121694 104392
rect 121750 104336 121755 104392
rect 119806 104334 121755 104336
rect 121689 104331 121755 104334
rect 126982 104296 127042 104742
rect 161525 104800 164026 104802
rect 161525 104744 161530 104800
rect 161586 104744 164026 104800
rect 161525 104742 164026 104744
rect 161525 104739 161591 104742
rect 50941 104258 51007 104261
rect 88477 104258 88543 104261
rect 159869 104258 159935 104261
rect 47862 104256 51007 104258
rect 47862 104200 50946 104256
rect 51002 104200 51007 104256
rect 47862 104198 51007 104200
rect 84876 104256 88543 104258
rect 84876 104200 88482 104256
rect 88538 104200 88543 104256
rect 84876 104198 88543 104200
rect 156820 104256 159935 104258
rect 156820 104200 159874 104256
rect 159930 104200 159935 104256
rect 156820 104198 159935 104200
rect 50941 104195 51007 104198
rect 88477 104195 88543 104198
rect 159869 104195 159935 104198
rect 160329 104258 160395 104261
rect 163966 104258 164026 104568
rect 160329 104256 164026 104258
rect 160329 104200 160334 104256
rect 160390 104200 164026 104256
rect 160329 104198 164026 104200
rect 160329 104195 160395 104198
rect 9896 104122 10376 104152
rect 13313 104122 13379 104125
rect 9896 104120 13379 104122
rect 9896 104064 13318 104120
rect 13374 104064 13379 104120
rect 9896 104062 13379 104064
rect 9896 104032 10376 104062
rect 13313 104059 13379 104062
rect 47862 103714 47922 104024
rect 91470 103990 92052 104050
rect 51309 103986 51375 103989
rect 88477 103986 88543 103989
rect 91470 103986 91530 103990
rect 51309 103984 55098 103986
rect 51309 103928 51314 103984
rect 51370 103928 55098 103984
rect 51309 103926 55098 103928
rect 51309 103923 51375 103926
rect 55038 103752 55098 103926
rect 88477 103984 91530 103986
rect 88477 103928 88482 103984
rect 88538 103928 91530 103984
rect 88477 103926 91530 103928
rect 88477 103923 88543 103926
rect 51217 103714 51283 103717
rect 88385 103714 88451 103717
rect 47862 103712 51283 103714
rect 47862 103656 51222 103712
rect 51278 103656 51283 103712
rect 47862 103654 51283 103656
rect 84876 103712 88451 103714
rect 84876 103656 88390 103712
rect 88446 103656 88451 103712
rect 84876 103654 88451 103656
rect 119806 103714 119866 104024
rect 124357 103986 124423 103989
rect 160053 103986 160119 103989
rect 124357 103984 127042 103986
rect 124357 103928 124362 103984
rect 124418 103928 127042 103984
rect 124357 103926 127042 103928
rect 124357 103923 124423 103926
rect 126982 103752 127042 103926
rect 156790 103984 160119 103986
rect 156790 103928 160058 103984
rect 160114 103928 160119 103984
rect 156790 103926 160119 103928
rect 121873 103714 121939 103717
rect 119806 103712 121939 103714
rect 119806 103656 121878 103712
rect 121934 103656 121939 103712
rect 156790 103684 156850 103926
rect 160053 103923 160119 103926
rect 160145 103714 160211 103717
rect 163966 103714 164026 104024
rect 160145 103712 164026 103714
rect 119806 103654 121939 103656
rect 51217 103651 51283 103654
rect 88385 103651 88451 103654
rect 121873 103651 121939 103654
rect 160145 103656 160150 103712
rect 160206 103656 164026 103712
rect 160145 103654 164026 103656
rect 160145 103651 160211 103654
rect 51401 103578 51467 103581
rect 124173 103578 124239 103581
rect 51401 103576 55098 103578
rect 51401 103520 51406 103576
rect 51462 103520 55098 103576
rect 51401 103518 55098 103520
rect 51401 103515 51467 103518
rect 47862 103170 47922 103480
rect 55038 103208 55098 103518
rect 124173 103576 127042 103578
rect 124173 103520 124178 103576
rect 124234 103520 127042 103576
rect 124173 103518 127042 103520
rect 124173 103515 124239 103518
rect 91470 103446 92052 103506
rect 88477 103442 88543 103445
rect 91470 103442 91530 103446
rect 88477 103440 91530 103442
rect 88477 103384 88482 103440
rect 88538 103384 91530 103440
rect 88477 103382 91530 103384
rect 88477 103379 88543 103382
rect 119806 103306 119866 103480
rect 121781 103306 121847 103309
rect 119806 103304 121847 103306
rect 119806 103248 121786 103304
rect 121842 103248 121847 103304
rect 119806 103246 121847 103248
rect 121781 103243 121847 103246
rect 126982 103208 127042 103518
rect 50757 103170 50823 103173
rect 88293 103170 88359 103173
rect 159961 103170 160027 103173
rect 47862 103168 50823 103170
rect 47862 103112 50762 103168
rect 50818 103112 50823 103168
rect 47862 103110 50823 103112
rect 84876 103168 88359 103170
rect 84876 103112 88298 103168
rect 88354 103112 88359 103168
rect 84876 103110 88359 103112
rect 156820 103168 160027 103170
rect 156820 103112 159966 103168
rect 160022 103112 160027 103168
rect 156820 103110 160027 103112
rect 50757 103107 50823 103110
rect 88293 103107 88359 103110
rect 159961 103107 160027 103110
rect 160237 103034 160303 103037
rect 163966 103034 164026 103480
rect 160237 103032 164026 103034
rect 160237 102976 160242 103032
rect 160298 102976 164026 103032
rect 160237 102974 164026 102976
rect 160237 102971 160303 102974
rect 121689 102898 121755 102901
rect 119806 102896 121755 102898
rect 119806 102840 121694 102896
rect 121750 102840 121755 102896
rect 119806 102838 121755 102840
rect 47862 102762 47922 102800
rect 91470 102766 92052 102826
rect 119806 102800 119866 102838
rect 121689 102835 121755 102838
rect 51401 102762 51467 102765
rect 47862 102760 51467 102762
rect 47862 102704 51406 102760
rect 51462 102704 51467 102760
rect 47862 102702 51467 102704
rect 51401 102699 51467 102702
rect 89673 102762 89739 102765
rect 91470 102762 91530 102766
rect 89673 102760 91530 102762
rect 89673 102704 89678 102760
rect 89734 102704 91530 102760
rect 89673 102702 91530 102704
rect 160513 102762 160579 102765
rect 163966 102762 164026 102800
rect 160513 102760 164026 102762
rect 160513 102704 160518 102760
rect 160574 102704 164026 102760
rect 160513 102702 164026 102704
rect 89673 102699 89739 102702
rect 160513 102699 160579 102702
rect 47862 101946 47922 102256
rect 91470 102222 92052 102282
rect 88661 102218 88727 102221
rect 91470 102218 91530 102222
rect 88661 102216 91530 102218
rect 88661 102160 88666 102216
rect 88722 102160 91530 102216
rect 88661 102158 91530 102160
rect 88661 102155 88727 102158
rect 51217 101946 51283 101949
rect 47862 101944 51283 101946
rect 47862 101888 51222 101944
rect 51278 101888 51283 101944
rect 47862 101886 51283 101888
rect 119806 101946 119866 102256
rect 123069 101946 123135 101949
rect 119806 101944 123135 101946
rect 119806 101888 123074 101944
rect 123130 101888 123135 101944
rect 119806 101886 123135 101888
rect 51217 101883 51283 101886
rect 123069 101883 123135 101886
rect 160329 101946 160395 101949
rect 163966 101946 164026 102256
rect 160329 101944 164026 101946
rect 160329 101888 160334 101944
rect 160390 101888 164026 101944
rect 160329 101886 164026 101888
rect 160329 101883 160395 101886
rect 47862 101402 47922 101712
rect 91470 101678 92052 101738
rect 88569 101674 88635 101677
rect 91470 101674 91530 101678
rect 88569 101672 91530 101674
rect 88569 101616 88574 101672
rect 88630 101616 91530 101672
rect 88569 101614 91530 101616
rect 88569 101611 88635 101614
rect 51309 101402 51375 101405
rect 47862 101400 51375 101402
rect 47862 101344 51314 101400
rect 51370 101344 51375 101400
rect 47862 101342 51375 101344
rect 119806 101402 119866 101712
rect 160421 101538 160487 101541
rect 163966 101538 164026 101712
rect 160421 101536 164026 101538
rect 160421 101480 160426 101536
rect 160482 101480 164026 101536
rect 160421 101478 164026 101480
rect 160421 101475 160487 101478
rect 123253 101402 123319 101405
rect 119806 101400 123319 101402
rect 119806 101344 123258 101400
rect 123314 101344 123319 101400
rect 119806 101342 123319 101344
rect 51309 101339 51375 101342
rect 123253 101339 123319 101342
rect 47862 101130 47922 101168
rect 50481 101130 50547 101133
rect 47862 101128 50547 101130
rect 47862 101072 50486 101128
rect 50542 101072 50547 101128
rect 47862 101070 50547 101072
rect 50481 101067 50547 101070
rect 55541 100994 55607 100997
rect 56737 100994 56803 100997
rect 48046 100992 56803 100994
rect 48046 100936 55546 100992
rect 55602 100936 56742 100992
rect 56798 100936 56803 100992
rect 48046 100934 56803 100936
rect 46382 100660 46388 100724
rect 46452 100722 46458 100724
rect 48046 100722 48106 100934
rect 55541 100931 55607 100934
rect 56737 100931 56803 100934
rect 46452 100662 48106 100722
rect 46452 100660 46458 100662
rect 88569 100586 88635 100589
rect 92022 100586 92082 101164
rect 116353 100722 116419 100725
rect 116854 100722 116860 100724
rect 116353 100720 116860 100722
rect 116353 100664 116358 100720
rect 116414 100664 116860 100720
rect 116353 100662 116860 100664
rect 116353 100659 116419 100662
rect 116854 100660 116860 100662
rect 116924 100660 116930 100724
rect 88569 100584 92082 100586
rect 88569 100528 88574 100584
rect 88630 100528 92082 100584
rect 88569 100526 92082 100528
rect 119806 100586 119866 101168
rect 122149 100586 122215 100589
rect 119806 100584 122215 100586
rect 119806 100528 122154 100584
rect 122210 100528 122215 100584
rect 119806 100526 122215 100528
rect 88569 100523 88635 100526
rect 122149 100523 122215 100526
rect 160329 100586 160395 100589
rect 163966 100586 164026 101168
rect 160329 100584 164026 100586
rect 160329 100528 160334 100584
rect 160390 100528 164026 100584
rect 160329 100526 164026 100528
rect 160329 100523 160395 100526
rect 20489 97866 20555 97869
rect 40310 97866 40316 97868
rect 20489 97864 40316 97866
rect 20489 97808 20494 97864
rect 20550 97808 40316 97864
rect 20489 97806 40316 97808
rect 20489 97803 20555 97806
rect 40310 97804 40316 97806
rect 40380 97804 40386 97868
rect 91697 93242 91763 93245
rect 164101 93242 164167 93245
rect 89844 93240 91763 93242
rect 89844 93184 91702 93240
rect 91758 93184 91763 93240
rect 89844 93182 91763 93184
rect 161788 93240 164167 93242
rect 161788 93184 164106 93240
rect 164162 93184 164167 93240
rect 161788 93182 164167 93184
rect 91697 93179 91763 93182
rect 164101 93179 164167 93182
rect 168517 92834 168583 92837
rect 168517 92832 170068 92834
rect 168517 92776 168522 92832
rect 168578 92776 170068 92832
rect 168517 92774 170068 92776
rect 168517 92771 168583 92774
rect 95285 92562 95351 92565
rect 95285 92560 97940 92562
rect 95285 92504 95290 92560
rect 95346 92504 97940 92560
rect 95285 92502 97940 92504
rect 95285 92499 95351 92502
rect 92249 92018 92315 92021
rect 163825 92018 163891 92021
rect 89844 92016 92315 92018
rect 89844 91960 92254 92016
rect 92310 91960 92315 92016
rect 89844 91958 92315 91960
rect 161788 92016 163891 92018
rect 161788 91960 163830 92016
rect 163886 91960 163891 92016
rect 161788 91958 163891 91960
rect 92249 91955 92315 91958
rect 163825 91955 163891 91958
rect 197589 91202 197655 91205
rect 201416 91202 201896 91232
rect 197589 91200 201896 91202
rect 197589 91144 197594 91200
rect 197650 91144 201896 91200
rect 197589 91142 201896 91144
rect 197589 91139 197655 91142
rect 201416 91112 201896 91142
rect 91513 90794 91579 90797
rect 163549 90794 163615 90797
rect 89844 90792 91579 90794
rect 89844 90736 91518 90792
rect 91574 90736 91579 90792
rect 89844 90734 91579 90736
rect 161788 90792 163615 90794
rect 161788 90736 163554 90792
rect 163610 90736 163615 90792
rect 161788 90734 163615 90736
rect 91513 90731 91579 90734
rect 163549 90731 163615 90734
rect 168374 90324 168380 90388
rect 168444 90386 168450 90388
rect 170038 90386 170098 90696
rect 188113 90522 188179 90525
rect 185892 90520 188179 90522
rect 185892 90464 188118 90520
rect 188174 90464 188179 90520
rect 185892 90462 188179 90464
rect 188113 90459 188179 90462
rect 168444 90326 170098 90386
rect 168444 90324 168450 90326
rect 95377 90250 95443 90253
rect 95377 90248 97940 90250
rect 95377 90192 95382 90248
rect 95438 90192 97940 90248
rect 95377 90190 97940 90192
rect 95377 90187 95443 90190
rect 22329 89842 22395 89845
rect 45053 89842 45119 89845
rect 22329 89840 25996 89842
rect 22329 89784 22334 89840
rect 22390 89784 25996 89840
rect 22329 89782 25996 89784
rect 41820 89840 45119 89842
rect 41820 89784 45058 89840
rect 45114 89784 45119 89840
rect 41820 89782 45119 89784
rect 22329 89779 22395 89782
rect 45053 89779 45119 89782
rect 92157 89570 92223 89573
rect 163825 89570 163891 89573
rect 89844 89568 92223 89570
rect 89844 89512 92162 89568
rect 92218 89512 92223 89568
rect 89844 89510 92223 89512
rect 161788 89568 163891 89570
rect 161788 89512 163830 89568
rect 163886 89512 163891 89568
rect 161788 89510 163891 89512
rect 92157 89507 92223 89510
rect 163825 89507 163891 89510
rect 92433 88346 92499 88349
rect 163457 88346 163523 88349
rect 89844 88344 92499 88346
rect 89844 88288 92438 88344
rect 92494 88288 92499 88344
rect 89844 88286 92499 88288
rect 161788 88344 163523 88346
rect 161788 88288 163462 88344
rect 163518 88288 163523 88344
rect 161788 88286 163523 88288
rect 92433 88283 92499 88286
rect 163457 88283 163523 88286
rect 167321 88074 167387 88077
rect 170038 88074 170098 88656
rect 167321 88072 170098 88074
rect 167321 88016 167326 88072
rect 167382 88016 170098 88072
rect 167321 88014 170098 88016
rect 167321 88011 167387 88014
rect 95377 87938 95443 87941
rect 95377 87936 97940 87938
rect 95377 87880 95382 87936
rect 95438 87880 97940 87936
rect 95377 87878 97940 87880
rect 95377 87875 95443 87878
rect 48406 87196 48412 87260
rect 48476 87258 48482 87260
rect 118929 87258 118995 87261
rect 48476 87198 49916 87258
rect 118929 87256 122044 87258
rect 118929 87200 118934 87256
rect 118990 87200 122044 87256
rect 118929 87198 122044 87200
rect 48476 87196 48482 87198
rect 118929 87195 118995 87198
rect 92801 87122 92867 87125
rect 163733 87122 163799 87125
rect 89844 87120 92867 87122
rect 89844 87064 92806 87120
rect 92862 87064 92867 87120
rect 89844 87062 92867 87064
rect 161788 87120 163799 87122
rect 161788 87064 163738 87120
rect 163794 87064 163799 87120
rect 161788 87062 163799 87064
rect 92801 87059 92867 87062
rect 163733 87059 163799 87062
rect 167873 86170 167939 86173
rect 170038 86170 170098 86752
rect 167873 86168 170098 86170
rect 167873 86112 167878 86168
rect 167934 86112 170098 86168
rect 167873 86110 170098 86112
rect 167873 86107 167939 86110
rect 91421 85898 91487 85901
rect 164561 85898 164627 85901
rect 89844 85896 91487 85898
rect 89844 85840 91426 85896
rect 91482 85840 91487 85896
rect 89844 85838 91487 85840
rect 161788 85896 164627 85898
rect 161788 85840 164566 85896
rect 164622 85840 164627 85896
rect 161788 85838 164627 85840
rect 91421 85835 91487 85838
rect 164561 85835 164627 85838
rect 94273 85490 94339 85493
rect 94273 85488 97940 85490
rect 94273 85432 94278 85488
rect 94334 85432 97940 85488
rect 94273 85430 97940 85432
rect 94273 85427 94339 85430
rect 167229 84810 167295 84813
rect 167229 84808 170068 84810
rect 167229 84752 167234 84808
rect 167290 84752 170068 84808
rect 167229 84750 170068 84752
rect 167229 84747 167295 84750
rect 91329 84674 91395 84677
rect 163089 84674 163155 84677
rect 89844 84672 91395 84674
rect 89844 84616 91334 84672
rect 91390 84616 91395 84672
rect 89844 84614 91395 84616
rect 161788 84672 163155 84674
rect 161788 84616 163094 84672
rect 163150 84616 163155 84672
rect 161788 84614 163155 84616
rect 91329 84611 91395 84614
rect 163089 84611 163155 84614
rect 116537 83858 116603 83861
rect 188113 83858 188179 83861
rect 113764 83856 116603 83858
rect 113764 83800 116542 83856
rect 116598 83800 116603 83856
rect 113764 83798 116603 83800
rect 185892 83856 188179 83858
rect 185892 83800 188118 83856
rect 188174 83800 188179 83856
rect 185892 83798 188179 83800
rect 116537 83795 116603 83798
rect 188113 83795 188179 83798
rect 91789 83450 91855 83453
rect 163917 83450 163983 83453
rect 89844 83448 91855 83450
rect 89844 83392 91794 83448
rect 91850 83392 91855 83448
rect 89844 83390 91855 83392
rect 161788 83448 163983 83450
rect 161788 83392 163922 83448
rect 163978 83392 163983 83448
rect 161788 83390 163983 83392
rect 91789 83387 91855 83390
rect 163917 83387 163983 83390
rect 95285 83178 95351 83181
rect 95285 83176 97940 83178
rect 95285 83120 95290 83176
rect 95346 83120 97940 83176
rect 95285 83118 97940 83120
rect 95285 83115 95351 83118
rect 9896 82906 10376 82936
rect 13221 82906 13287 82909
rect 9896 82904 13287 82906
rect 9896 82848 13226 82904
rect 13282 82848 13287 82904
rect 9896 82846 13287 82848
rect 9896 82816 10376 82846
rect 13221 82843 13287 82846
rect 92249 82226 92315 82229
rect 163917 82226 163983 82229
rect 89844 82224 92315 82226
rect 89844 82168 92254 82224
rect 92310 82168 92315 82224
rect 89844 82166 92315 82168
rect 161788 82224 163983 82226
rect 161788 82168 163922 82224
rect 163978 82168 163983 82224
rect 161788 82166 163983 82168
rect 92249 82163 92315 82166
rect 163917 82163 163983 82166
rect 167321 82090 167387 82093
rect 170038 82090 170098 82672
rect 167321 82088 170098 82090
rect 167321 82032 167326 82088
rect 167382 82032 170098 82088
rect 167321 82030 170098 82032
rect 167321 82027 167387 82030
rect 41598 81892 41604 81956
rect 41668 81892 41674 81956
rect 22329 81818 22395 81821
rect 22329 81816 25996 81818
rect 22329 81760 22334 81816
rect 22390 81760 25996 81816
rect 41606 81788 41666 81892
rect 22329 81758 25996 81760
rect 22329 81755 22395 81758
rect 92157 81138 92223 81141
rect 163549 81138 163615 81141
rect 89844 81136 92223 81138
rect 89844 81080 92162 81136
rect 92218 81080 92223 81136
rect 89844 81078 92223 81080
rect 161788 81136 163615 81138
rect 161788 81080 163554 81136
rect 163610 81080 163615 81136
rect 161788 81078 163615 81080
rect 92157 81075 92223 81078
rect 163549 81075 163615 81078
rect 95377 80866 95443 80869
rect 167229 80866 167295 80869
rect 95377 80864 97940 80866
rect 95377 80808 95382 80864
rect 95438 80808 97940 80864
rect 95377 80806 97940 80808
rect 167229 80864 170068 80866
rect 167229 80808 167234 80864
rect 167290 80808 170068 80864
rect 167229 80806 170068 80808
rect 95377 80803 95443 80806
rect 167229 80803 167295 80806
rect 91789 79914 91855 79917
rect 164101 79914 164167 79917
rect 89844 79912 91855 79914
rect 89844 79856 91794 79912
rect 91850 79856 91855 79912
rect 89844 79854 91855 79856
rect 161788 79912 164167 79914
rect 161788 79856 164106 79912
rect 164162 79856 164167 79912
rect 161788 79854 164167 79856
rect 91789 79851 91855 79854
rect 164101 79851 164167 79854
rect 91421 78690 91487 78693
rect 164377 78690 164443 78693
rect 89844 78688 91487 78690
rect 89844 78632 91426 78688
rect 91482 78632 91487 78688
rect 89844 78630 91487 78632
rect 161788 78688 164443 78690
rect 161788 78632 164382 78688
rect 164438 78632 164443 78688
rect 161788 78630 164443 78632
rect 91421 78627 91487 78630
rect 164377 78627 164443 78630
rect 94917 78418 94983 78421
rect 94917 78416 97940 78418
rect 94917 78360 94922 78416
rect 94978 78360 97940 78416
rect 94917 78358 97940 78360
rect 94917 78355 94983 78358
rect 167229 78146 167295 78149
rect 170038 78146 170098 78728
rect 167229 78144 170098 78146
rect 167229 78088 167234 78144
rect 167290 78088 170098 78144
rect 167229 78086 170098 78088
rect 167229 78083 167295 78086
rect 91697 77466 91763 77469
rect 164101 77466 164167 77469
rect 89844 77464 91763 77466
rect 89844 77408 91702 77464
rect 91758 77408 91763 77464
rect 89844 77406 91763 77408
rect 161788 77464 164167 77466
rect 161788 77408 164106 77464
rect 164162 77408 164167 77464
rect 161788 77406 164167 77408
rect 91697 77403 91763 77406
rect 164101 77403 164167 77406
rect 188573 77194 188639 77197
rect 185892 77192 188639 77194
rect 185892 77136 188578 77192
rect 188634 77136 188639 77192
rect 185892 77134 188639 77136
rect 188573 77131 188639 77134
rect 167229 76514 167295 76517
rect 170038 76514 170098 76688
rect 167229 76512 170098 76514
rect 167229 76456 167234 76512
rect 167290 76456 170098 76512
rect 167229 76454 170098 76456
rect 167229 76451 167295 76454
rect 91697 76242 91763 76245
rect 163733 76242 163799 76245
rect 89844 76240 91763 76242
rect 89844 76184 91702 76240
rect 91758 76184 91763 76240
rect 89844 76182 91763 76184
rect 161788 76240 163799 76242
rect 161788 76184 163738 76240
rect 163794 76184 163799 76240
rect 161788 76182 163799 76184
rect 91697 76179 91763 76182
rect 163733 76179 163799 76182
rect 98094 75154 98154 76076
rect 94046 75094 98154 75154
rect 94046 75018 94106 75094
rect 164101 75018 164167 75021
rect 89844 74958 94106 75018
rect 161788 75016 164167 75018
rect 161788 74960 164106 75016
rect 164162 74960 164167 75016
rect 161788 74958 164167 74960
rect 164101 74955 164167 74958
rect 167229 74882 167295 74885
rect 167229 74880 170068 74882
rect 167229 74824 167234 74880
rect 167290 74824 170068 74880
rect 167229 74822 170068 74824
rect 167229 74819 167295 74822
rect 47813 73930 47879 73933
rect 119573 73930 119639 73933
rect 47813 73928 49916 73930
rect 47813 73872 47818 73928
rect 47874 73872 49916 73928
rect 47813 73870 49916 73872
rect 119573 73928 122044 73930
rect 119573 73872 119578 73928
rect 119634 73872 122044 73928
rect 119573 73870 122044 73872
rect 47813 73867 47879 73870
rect 119573 73867 119639 73870
rect 22329 73794 22395 73797
rect 44358 73794 44364 73796
rect 22329 73792 25996 73794
rect 22329 73736 22334 73792
rect 22390 73736 25996 73792
rect 22329 73734 25996 73736
rect 41820 73734 44364 73794
rect 22329 73731 22395 73734
rect 44358 73732 44364 73734
rect 44428 73732 44434 73796
rect 164377 73794 164443 73797
rect 89844 73734 97940 73794
rect 161788 73792 164443 73794
rect 161788 73736 164382 73792
rect 164438 73736 164443 73792
rect 161788 73734 164443 73736
rect 164377 73731 164443 73734
rect 167137 72842 167203 72845
rect 167137 72840 170068 72842
rect 167137 72784 167142 72840
rect 167198 72784 170068 72840
rect 167137 72782 170068 72784
rect 167137 72779 167203 72782
rect 91697 72570 91763 72573
rect 164377 72570 164443 72573
rect 89844 72568 91763 72570
rect 89844 72512 91702 72568
rect 91758 72512 91763 72568
rect 89844 72510 91763 72512
rect 161788 72568 164443 72570
rect 161788 72512 164382 72568
rect 164438 72512 164443 72568
rect 161788 72510 164443 72512
rect 91697 72507 91763 72510
rect 164377 72507 164443 72510
rect 95377 71482 95443 71485
rect 95377 71480 97940 71482
rect 95377 71424 95382 71480
rect 95438 71424 97940 71480
rect 95377 71422 97940 71424
rect 95377 71419 95443 71422
rect 91697 71346 91763 71349
rect 164377 71346 164443 71349
rect 89844 71344 91763 71346
rect 89844 71288 91702 71344
rect 91758 71288 91763 71344
rect 89844 71286 91763 71288
rect 161788 71344 164443 71346
rect 161788 71288 164382 71344
rect 164438 71288 164443 71344
rect 161788 71286 164443 71288
rect 91697 71283 91763 71286
rect 164377 71283 164443 71286
rect 167229 70802 167295 70805
rect 167229 70800 170068 70802
rect 167229 70744 167234 70800
rect 167290 70744 170068 70800
rect 167229 70742 170068 70744
rect 167229 70739 167295 70742
rect 185862 70394 185922 70500
rect 186038 70394 186044 70396
rect 185862 70334 186044 70394
rect 186038 70332 186044 70334
rect 186108 70332 186114 70396
rect 91421 70122 91487 70125
rect 163549 70122 163615 70125
rect 89844 70120 91487 70122
rect 89844 70064 91426 70120
rect 91482 70064 91487 70120
rect 89844 70062 91487 70064
rect 161788 70120 163615 70122
rect 161788 70064 163554 70120
rect 163610 70064 163615 70120
rect 161788 70062 163615 70064
rect 91421 70059 91487 70062
rect 163549 70059 163615 70062
rect 95377 69034 95443 69037
rect 95377 69032 97940 69034
rect 95377 68976 95382 69032
rect 95438 68976 97940 69032
rect 95377 68974 97940 68976
rect 95377 68971 95443 68974
rect 91421 68898 91487 68901
rect 163733 68898 163799 68901
rect 89844 68896 91487 68898
rect 89844 68840 91426 68896
rect 91482 68840 91487 68896
rect 89844 68838 91487 68840
rect 161788 68896 163799 68898
rect 161788 68840 163738 68896
rect 163794 68840 163799 68896
rect 161788 68838 163799 68840
rect 91421 68835 91487 68838
rect 163733 68835 163799 68838
rect 167321 68762 167387 68765
rect 167321 68760 170068 68762
rect 167321 68704 167326 68760
rect 167382 68704 170068 68760
rect 167321 68702 170068 68704
rect 167321 68699 167387 68702
rect 91513 67810 91579 67813
rect 164377 67810 164443 67813
rect 89844 67808 91579 67810
rect 89844 67752 91518 67808
rect 91574 67752 91579 67808
rect 89844 67750 91579 67752
rect 161788 67808 164443 67810
rect 161788 67752 164382 67808
rect 164438 67752 164443 67808
rect 161788 67750 164443 67752
rect 91513 67747 91579 67750
rect 164377 67747 164443 67750
rect 197589 67674 197655 67677
rect 201416 67674 201896 67704
rect 197589 67672 201896 67674
rect 197589 67616 197594 67672
rect 197650 67616 201896 67672
rect 197589 67614 201896 67616
rect 197589 67611 197655 67614
rect 201416 67584 201896 67614
rect 167229 66858 167295 66861
rect 167229 66856 170068 66858
rect 167229 66800 167234 66856
rect 167290 66800 170068 66856
rect 167229 66798 170068 66800
rect 167229 66795 167295 66798
rect 95377 66722 95443 66725
rect 95377 66720 97940 66722
rect 95377 66664 95382 66720
rect 95438 66664 97940 66720
rect 95377 66662 97940 66664
rect 95377 66659 95443 66662
rect 92525 66586 92591 66589
rect 164377 66586 164443 66589
rect 89844 66584 92591 66586
rect 89844 66528 92530 66584
rect 92586 66528 92591 66584
rect 89844 66526 92591 66528
rect 161788 66584 164443 66586
rect 161788 66528 164382 66584
rect 164438 66528 164443 66584
rect 161788 66526 164443 66528
rect 92525 66523 92591 66526
rect 164377 66523 164443 66526
rect 22697 65770 22763 65773
rect 44409 65770 44475 65773
rect 22697 65768 25996 65770
rect 22697 65712 22702 65768
rect 22758 65712 25996 65768
rect 22697 65710 25996 65712
rect 41820 65768 44475 65770
rect 41820 65712 44414 65768
rect 44470 65712 44475 65768
rect 41820 65710 44475 65712
rect 22697 65707 22763 65710
rect 44409 65707 44475 65710
rect 93997 65498 94063 65501
rect 95377 65498 95443 65501
rect 93997 65496 95443 65498
rect 93997 65440 94002 65496
rect 94058 65440 95382 65496
rect 95438 65440 95443 65496
rect 93997 65438 95443 65440
rect 93997 65435 94063 65438
rect 95377 65435 95443 65438
rect 92341 65362 92407 65365
rect 164377 65362 164443 65365
rect 89844 65360 92407 65362
rect 89844 65304 92346 65360
rect 92402 65304 92407 65360
rect 89844 65302 92407 65304
rect 161788 65360 164443 65362
rect 161788 65304 164382 65360
rect 164438 65304 164443 65360
rect 161788 65302 164443 65304
rect 92341 65299 92407 65302
rect 164377 65299 164443 65302
rect 167321 64818 167387 64821
rect 167321 64816 170068 64818
rect 167321 64760 167326 64816
rect 167382 64760 170068 64816
rect 167321 64758 170068 64760
rect 167321 64755 167387 64758
rect 92617 64138 92683 64141
rect 89844 64136 92683 64138
rect 89844 64080 92622 64136
rect 92678 64080 92683 64136
rect 89844 64078 92683 64080
rect 92617 64075 92683 64078
rect 93905 64138 93971 64141
rect 97910 64138 97970 64380
rect 164377 64138 164443 64141
rect 93905 64136 97970 64138
rect 93905 64080 93910 64136
rect 93966 64080 97970 64136
rect 93905 64078 97970 64080
rect 161788 64136 164443 64138
rect 161788 64080 164382 64136
rect 164438 64080 164443 64136
rect 161788 64078 164443 64080
rect 93905 64075 93971 64078
rect 164377 64075 164443 64078
rect 187878 63866 187884 63868
rect 185892 63806 187884 63866
rect 187878 63804 187884 63806
rect 187948 63804 187954 63868
rect 113734 63186 113794 63768
rect 117457 63186 117523 63189
rect 113734 63184 117523 63186
rect 113734 63128 117462 63184
rect 117518 63128 117523 63184
rect 113734 63126 117523 63128
rect 117457 63123 117523 63126
rect 93353 62914 93419 62917
rect 163733 62914 163799 62917
rect 89844 62912 93419 62914
rect 89844 62856 93358 62912
rect 93414 62856 93419 62912
rect 89844 62854 93419 62856
rect 161788 62912 163799 62914
rect 161788 62856 163738 62912
rect 163794 62856 163799 62912
rect 161788 62854 163799 62856
rect 93353 62851 93419 62854
rect 163733 62851 163799 62854
rect 167873 62778 167939 62781
rect 167873 62776 170068 62778
rect 167873 62720 167878 62776
rect 167934 62720 170068 62776
rect 167873 62718 170068 62720
rect 167873 62715 167939 62718
rect 9896 61690 10376 61720
rect 13313 61690 13379 61693
rect 91421 61690 91487 61693
rect 9896 61688 13379 61690
rect 9896 61632 13318 61688
rect 13374 61632 13379 61688
rect 9896 61630 13379 61632
rect 89844 61688 91487 61690
rect 89844 61632 91426 61688
rect 91482 61632 91487 61688
rect 89844 61630 91487 61632
rect 9896 61600 10376 61630
rect 13313 61627 13379 61630
rect 91421 61627 91487 61630
rect 93629 61418 93695 61421
rect 97910 61418 97970 61932
rect 163825 61690 163891 61693
rect 161788 61688 163891 61690
rect 161788 61632 163830 61688
rect 163886 61632 163891 61688
rect 161788 61630 163891 61632
rect 163825 61627 163891 61630
rect 93629 61416 97970 61418
rect 93629 61360 93634 61416
rect 93690 61360 97970 61416
rect 93629 61358 97970 61360
rect 93629 61355 93695 61358
rect 167137 60874 167203 60877
rect 167137 60872 170068 60874
rect 167137 60816 167142 60872
rect 167198 60816 170068 60872
rect 167137 60814 170068 60816
rect 167137 60811 167203 60814
rect 47169 60602 47235 60605
rect 47537 60602 47603 60605
rect 119481 60602 119547 60605
rect 47169 60600 49916 60602
rect 47169 60544 47174 60600
rect 47230 60544 47542 60600
rect 47598 60544 49916 60600
rect 47169 60542 49916 60544
rect 119481 60600 122044 60602
rect 119481 60544 119486 60600
rect 119542 60572 122044 60600
rect 119542 60544 122074 60572
rect 119481 60542 122074 60544
rect 47169 60539 47235 60542
rect 47537 60539 47603 60542
rect 119481 60539 119547 60542
rect 94641 60466 94707 60469
rect 89844 60464 94707 60466
rect 89844 60408 94646 60464
rect 94702 60408 94707 60464
rect 89844 60406 94707 60408
rect 94641 60403 94707 60406
rect 122014 59924 122074 60542
rect 165113 60466 165179 60469
rect 161788 60464 165179 60466
rect 161788 60408 165118 60464
rect 165174 60408 165179 60464
rect 161788 60406 165179 60408
rect 165113 60403 165179 60406
rect 122006 59860 122012 59924
rect 122076 59860 122082 59924
rect 94089 59650 94155 59653
rect 94089 59648 97940 59650
rect 94089 59592 94094 59648
rect 94150 59592 97940 59648
rect 94089 59590 97940 59592
rect 94089 59587 94155 59590
rect 91513 59242 91579 59245
rect 164377 59242 164443 59245
rect 89844 59240 91579 59242
rect 89844 59184 91518 59240
rect 91574 59184 91579 59240
rect 89844 59182 91579 59184
rect 161788 59240 164443 59242
rect 161788 59184 164382 59240
rect 164438 59184 164443 59240
rect 161788 59182 164443 59184
rect 91513 59179 91579 59182
rect 164377 59179 164443 59182
rect 167045 58834 167111 58837
rect 167045 58832 170068 58834
rect 167045 58776 167050 58832
rect 167106 58776 170068 58832
rect 167045 58774 170068 58776
rect 167045 58771 167111 58774
rect 26142 58092 26148 58156
rect 26212 58092 26218 58156
rect 26150 57852 26210 58092
rect 92893 58018 92959 58021
rect 164377 58018 164443 58021
rect 89844 58016 92959 58018
rect 89844 57960 92898 58016
rect 92954 57960 92959 58016
rect 89844 57958 92959 57960
rect 161788 58016 164443 58018
rect 161788 57960 164382 58016
rect 164438 57960 164443 58016
rect 161788 57958 164443 57960
rect 92893 57955 92959 57958
rect 164377 57955 164443 57958
rect 44409 57882 44475 57885
rect 41820 57880 44475 57882
rect 41820 57824 44414 57880
rect 44470 57824 44475 57880
rect 41820 57822 44475 57824
rect 44409 57819 44475 57822
rect 161750 57412 161756 57476
rect 161820 57474 161826 57476
rect 170214 57474 170220 57476
rect 161820 57414 170220 57474
rect 161820 57412 161826 57414
rect 170214 57412 170220 57414
rect 170284 57412 170290 57476
rect 95193 57338 95259 57341
rect 95193 57336 97940 57338
rect 95193 57280 95198 57336
rect 95254 57280 97940 57336
rect 95193 57278 97940 57280
rect 95193 57275 95259 57278
rect 185854 57276 185860 57340
rect 185924 57338 185930 57340
rect 185924 57278 186106 57338
rect 185924 57276 185930 57278
rect 186046 57202 186106 57278
rect 187929 57202 187995 57205
rect 185892 57200 187995 57202
rect 185892 57144 187934 57200
rect 187990 57144 187995 57200
rect 185892 57142 187995 57144
rect 187929 57139 187995 57142
rect 91421 56794 91487 56797
rect 165021 56794 165087 56797
rect 89844 56792 91487 56794
rect 89844 56736 91426 56792
rect 91482 56736 91487 56792
rect 89844 56734 91487 56736
rect 161788 56792 165087 56794
rect 161788 56736 165026 56792
rect 165082 56736 165087 56792
rect 161788 56734 165087 56736
rect 91421 56731 91487 56734
rect 165021 56731 165087 56734
rect 166493 56794 166559 56797
rect 166493 56792 170068 56794
rect 166493 56736 166498 56792
rect 166554 56736 170068 56792
rect 166493 56734 170068 56736
rect 166493 56731 166559 56734
rect 92617 55570 92683 55573
rect 164561 55570 164627 55573
rect 89844 55568 92683 55570
rect 89844 55512 92622 55568
rect 92678 55512 92683 55568
rect 89844 55510 92683 55512
rect 161788 55568 164627 55570
rect 161788 55512 164566 55568
rect 164622 55512 164627 55568
rect 161788 55510 164627 55512
rect 92617 55507 92683 55510
rect 164561 55507 164627 55510
rect 93537 55026 93603 55029
rect 93537 55024 97940 55026
rect 93537 54968 93542 55024
rect 93598 54968 97940 55024
rect 93537 54966 97940 54968
rect 93537 54963 93603 54966
rect 91329 54482 91395 54485
rect 163089 54482 163155 54485
rect 89844 54480 91395 54482
rect 89844 54424 91334 54480
rect 91390 54424 91395 54480
rect 89844 54422 91395 54424
rect 161788 54480 163155 54482
rect 161788 54424 163094 54480
rect 163150 54424 163155 54480
rect 161788 54422 163155 54424
rect 91329 54419 91395 54422
rect 163089 54419 163155 54422
rect 168517 54482 168583 54485
rect 170038 54482 170098 54792
rect 168517 54480 170098 54482
rect 168517 54424 168522 54480
rect 168578 54424 170098 54480
rect 168517 54422 170098 54424
rect 168517 54419 168583 54422
rect 82129 51626 82195 51629
rect 83601 51628 83667 51629
rect 82262 51626 82268 51628
rect 82129 51624 82268 51626
rect 82129 51568 82134 51624
rect 82190 51568 82268 51624
rect 82129 51566 82268 51568
rect 82129 51563 82195 51566
rect 82262 51564 82268 51566
rect 82332 51564 82338 51628
rect 83550 51626 83556 51628
rect 83510 51566 83556 51626
rect 83620 51624 83667 51628
rect 83662 51568 83667 51624
rect 83550 51564 83556 51566
rect 83620 51564 83667 51568
rect 83601 51563 83667 51564
rect 53241 51490 53307 51493
rect 138750 51490 138756 51492
rect 53241 51488 138756 51490
rect 53241 51432 53246 51488
rect 53302 51432 138756 51488
rect 53241 51430 138756 51432
rect 53241 51427 53307 51430
rect 138750 51428 138756 51430
rect 138820 51428 138826 51492
rect 66581 50266 66647 50269
rect 66990 50266 66996 50268
rect 66581 50264 66996 50266
rect 66581 50208 66586 50264
rect 66642 50208 66996 50264
rect 66581 50206 66996 50208
rect 66581 50203 66647 50206
rect 66990 50204 66996 50206
rect 67060 50204 67066 50268
rect 47537 46866 47603 46869
rect 47494 46864 47603 46866
rect 47494 46808 47542 46864
rect 47598 46808 47603 46864
rect 47494 46803 47603 46808
rect 47494 46254 47554 46803
rect 129734 46668 129740 46732
rect 129804 46730 129810 46732
rect 142665 46730 142731 46733
rect 129804 46728 142731 46730
rect 129804 46672 142670 46728
rect 142726 46672 142731 46728
rect 129804 46670 142731 46672
rect 129804 46668 129810 46670
rect 142665 46667 142731 46670
rect 67726 46532 67732 46596
rect 67796 46594 67802 46596
rect 75045 46594 75111 46597
rect 67796 46592 75111 46594
rect 67796 46536 75050 46592
rect 75106 46536 75111 46592
rect 67796 46534 75111 46536
rect 67796 46532 67802 46534
rect 75045 46531 75111 46534
rect 138934 46532 138940 46596
rect 139004 46594 139010 46596
rect 145609 46594 145675 46597
rect 139004 46592 145675 46594
rect 139004 46536 145614 46592
rect 145670 46536 145675 46592
rect 139004 46534 145675 46536
rect 139004 46532 139010 46534
rect 145609 46531 145675 46534
rect 67174 46396 67180 46460
rect 67244 46458 67250 46460
rect 73573 46458 73639 46461
rect 67244 46456 73639 46458
rect 67244 46400 73578 46456
rect 73634 46400 73639 46456
rect 67244 46398 73639 46400
rect 67244 46396 67250 46398
rect 73573 46395 73639 46398
rect 67358 46260 67364 46324
rect 67428 46322 67434 46324
rect 72101 46322 72167 46325
rect 67428 46320 72167 46322
rect 67428 46264 72106 46320
rect 72162 46264 72167 46320
rect 67428 46262 72167 46264
rect 67428 46260 67434 46262
rect 72101 46259 72167 46262
rect 47494 46224 47892 46254
rect 47524 46194 47922 46224
rect 47862 46186 47922 46194
rect 50573 46186 50639 46189
rect 47862 46184 50639 46186
rect 47862 46128 50578 46184
rect 50634 46128 50639 46184
rect 47862 46126 50639 46128
rect 50573 46123 50639 46126
rect 67542 46124 67548 46188
rect 67612 46186 67618 46188
rect 70629 46186 70695 46189
rect 67612 46184 70695 46186
rect 67612 46128 70634 46184
rect 70690 46128 70695 46184
rect 67612 46126 70695 46128
rect 67612 46124 67618 46126
rect 70629 46123 70695 46126
rect 88385 46186 88451 46189
rect 92022 46186 92082 46496
rect 88385 46184 92082 46186
rect 88385 46128 88390 46184
rect 88446 46128 92082 46184
rect 88385 46126 92082 46128
rect 119806 46186 119866 46496
rect 138750 46396 138756 46460
rect 138820 46458 138826 46460
rect 147081 46458 147147 46461
rect 138820 46456 147147 46458
rect 138820 46400 147086 46456
rect 147142 46400 147147 46456
rect 138820 46398 147147 46400
rect 138820 46396 138826 46398
rect 147081 46395 147147 46398
rect 131206 46260 131212 46324
rect 131276 46322 131282 46324
rect 144137 46322 144203 46325
rect 131276 46320 144203 46322
rect 131276 46264 144142 46320
rect 144198 46264 144203 46320
rect 131276 46262 144203 46264
rect 131276 46260 131282 46262
rect 144137 46259 144203 46262
rect 122977 46186 123043 46189
rect 119806 46184 123043 46186
rect 119806 46128 122982 46184
rect 123038 46128 123043 46184
rect 119806 46126 123043 46128
rect 88385 46123 88451 46126
rect 122977 46123 123043 46126
rect 160237 46186 160303 46189
rect 163966 46186 164026 46496
rect 160237 46184 164026 46186
rect 160237 46128 160242 46184
rect 160298 46128 164026 46184
rect 160237 46126 164026 46128
rect 160237 46123 160303 46126
rect 47862 45234 47922 45680
rect 88569 45506 88635 45509
rect 92022 45506 92082 45952
rect 88569 45504 92082 45506
rect 88569 45448 88574 45504
rect 88630 45448 92082 45504
rect 88569 45446 92082 45448
rect 119806 45506 119866 45952
rect 122977 45506 123043 45509
rect 119806 45504 123043 45506
rect 119806 45448 122982 45504
rect 123038 45448 123043 45504
rect 119806 45446 123043 45448
rect 88569 45443 88635 45446
rect 122977 45443 123043 45446
rect 160329 45506 160395 45509
rect 163966 45506 164026 45952
rect 160329 45504 164026 45506
rect 160329 45448 160334 45504
rect 160390 45448 164026 45504
rect 160329 45446 164026 45448
rect 160329 45443 160395 45446
rect 49929 45234 49995 45237
rect 47862 45232 49995 45234
rect 47862 45176 49934 45232
rect 49990 45176 49995 45232
rect 47862 45174 49995 45176
rect 49929 45171 49995 45174
rect 47862 44962 47922 45000
rect 51309 44962 51375 44965
rect 47862 44960 51375 44962
rect 47862 44904 51314 44960
rect 51370 44904 51375 44960
rect 47862 44902 51375 44904
rect 51309 44899 51375 44902
rect 88109 44962 88175 44965
rect 92022 44962 92082 45272
rect 119806 45098 119866 45272
rect 121689 45098 121755 45101
rect 119806 45096 121755 45098
rect 119806 45040 121694 45096
rect 121750 45040 121755 45096
rect 119806 45038 121755 45040
rect 121689 45035 121755 45038
rect 88109 44960 92082 44962
rect 88109 44904 88114 44960
rect 88170 44904 92082 44960
rect 88109 44902 92082 44904
rect 160145 44962 160211 44965
rect 163966 44962 164026 45272
rect 160145 44960 164026 44962
rect 160145 44904 160150 44960
rect 160206 44904 164026 44960
rect 160145 44902 164026 44904
rect 88109 44899 88175 44902
rect 160145 44899 160211 44902
rect 49929 44826 49995 44829
rect 88477 44826 88543 44829
rect 121689 44826 121755 44829
rect 49929 44824 51418 44826
rect 49929 44768 49934 44824
rect 49990 44768 51418 44824
rect 49929 44766 51418 44768
rect 49929 44763 49995 44766
rect 51358 44690 51418 44766
rect 88477 44824 92082 44826
rect 88477 44768 88482 44824
rect 88538 44768 92082 44824
rect 88477 44766 92082 44768
rect 88477 44763 88543 44766
rect 92022 44732 92082 44766
rect 119806 44824 121755 44826
rect 119806 44768 121694 44824
rect 121750 44768 121755 44824
rect 119806 44766 121755 44768
rect 119806 44728 119866 44766
rect 121689 44763 121755 44766
rect 160053 44826 160119 44829
rect 160053 44824 164026 44826
rect 160053 44768 160058 44824
rect 160114 44768 164026 44824
rect 160053 44766 164026 44768
rect 160053 44763 160119 44766
rect 163966 44728 164026 44766
rect 51358 44630 55098 44690
rect 55038 44456 55098 44630
rect 67910 44628 67916 44692
rect 67980 44690 67986 44692
rect 68789 44690 68855 44693
rect 67980 44688 68855 44690
rect 67980 44632 68794 44688
rect 68850 44632 68855 44688
rect 67980 44630 68855 44632
rect 67980 44628 67986 44630
rect 68789 44627 68855 44630
rect 82865 44690 82931 44693
rect 139721 44692 139787 44693
rect 83550 44690 83556 44692
rect 82865 44688 83556 44690
rect 82865 44632 82870 44688
rect 82926 44632 83556 44688
rect 82865 44630 83556 44632
rect 82865 44627 82931 44630
rect 83550 44628 83556 44630
rect 83620 44628 83626 44692
rect 139670 44690 139676 44692
rect 139630 44630 139676 44690
rect 139740 44688 139787 44692
rect 139782 44632 139787 44688
rect 139670 44628 139676 44630
rect 139740 44628 139787 44632
rect 139721 44627 139787 44628
rect 140917 44692 140983 44693
rect 140917 44688 140964 44692
rect 141028 44690 141034 44692
rect 140917 44632 140922 44688
rect 140917 44628 140964 44632
rect 141028 44630 141074 44690
rect 141028 44628 141034 44630
rect 140917 44627 140983 44628
rect 47862 44146 47922 44456
rect 88385 44418 88451 44421
rect 84876 44416 88451 44418
rect 84876 44360 88390 44416
rect 88446 44360 88451 44416
rect 84876 44358 88451 44360
rect 88385 44355 88451 44358
rect 123161 44418 123227 44421
rect 160237 44418 160303 44421
rect 123161 44416 127012 44418
rect 123161 44360 123166 44416
rect 123222 44360 127012 44416
rect 123161 44358 127012 44360
rect 156820 44416 160303 44418
rect 156820 44360 160242 44416
rect 160298 44360 160303 44416
rect 156820 44358 160303 44360
rect 123161 44355 123227 44358
rect 160237 44355 160303 44358
rect 51309 44282 51375 44285
rect 123069 44282 123135 44285
rect 51309 44280 55098 44282
rect 51309 44224 51314 44280
rect 51370 44224 55098 44280
rect 51309 44222 55098 44224
rect 51309 44219 51375 44222
rect 51217 44146 51283 44149
rect 47862 44144 51283 44146
rect 47862 44088 51222 44144
rect 51278 44088 51283 44144
rect 47862 44086 51283 44088
rect 51217 44083 51283 44086
rect 55038 43912 55098 44222
rect 123069 44280 127042 44282
rect 123069 44224 123074 44280
rect 123130 44224 127042 44280
rect 123069 44222 127042 44224
rect 123069 44219 123135 44222
rect 47862 43466 47922 43912
rect 88477 43874 88543 43877
rect 84876 43872 88543 43874
rect 84876 43816 88482 43872
rect 88538 43816 88543 43872
rect 84876 43814 88543 43816
rect 88477 43811 88543 43814
rect 88569 43738 88635 43741
rect 92022 43738 92082 44048
rect 88569 43736 92082 43738
rect 88569 43680 88574 43736
rect 88630 43680 92082 43736
rect 88569 43678 92082 43680
rect 119806 43738 119866 44048
rect 126982 43912 127042 44222
rect 201269 44146 201335 44149
rect 201416 44146 201896 44176
rect 201269 44144 201896 44146
rect 201269 44088 201274 44144
rect 201330 44088 201896 44144
rect 201269 44086 201896 44088
rect 201269 44083 201335 44086
rect 201416 44056 201896 44086
rect 160237 43874 160303 43877
rect 156820 43872 160303 43874
rect 156820 43816 160242 43872
rect 160298 43816 160303 43872
rect 156820 43814 160303 43816
rect 160237 43811 160303 43814
rect 122977 43738 123043 43741
rect 119806 43736 123043 43738
rect 119806 43680 122982 43736
rect 123038 43680 123043 43736
rect 119806 43678 123043 43680
rect 88569 43675 88635 43678
rect 122977 43675 123043 43678
rect 160329 43738 160395 43741
rect 163966 43738 164026 44048
rect 201269 43874 201335 43877
rect 190646 43872 201335 43874
rect 190646 43816 201274 43872
rect 201330 43816 201335 43872
rect 190646 43814 201335 43816
rect 160329 43736 164026 43738
rect 160329 43680 160334 43736
rect 160390 43680 164026 43736
rect 160329 43678 164026 43680
rect 160329 43675 160395 43678
rect 187142 43676 187148 43740
rect 187212 43738 187218 43740
rect 190646 43738 190706 43814
rect 201269 43811 201335 43814
rect 187212 43678 190706 43738
rect 187212 43676 187218 43678
rect 88385 43466 88451 43469
rect 92022 43466 92082 43504
rect 47862 43406 51234 43466
rect 47862 42922 47922 43232
rect 51174 43194 51234 43406
rect 88385 43464 92082 43466
rect 88385 43408 88390 43464
rect 88446 43408 92082 43464
rect 88385 43406 92082 43408
rect 119806 43466 119866 43504
rect 121689 43466 121755 43469
rect 119806 43464 121755 43466
rect 119806 43408 121694 43464
rect 121750 43408 121755 43464
rect 119806 43406 121755 43408
rect 88385 43403 88451 43406
rect 121689 43403 121755 43406
rect 160145 43466 160211 43469
rect 163966 43466 164026 43504
rect 160145 43464 164026 43466
rect 160145 43408 160150 43464
rect 160206 43408 164026 43464
rect 160145 43406 164026 43408
rect 160145 43403 160211 43406
rect 51309 43330 51375 43333
rect 51309 43328 54546 43330
rect 51309 43272 51314 43328
rect 51370 43272 54546 43328
rect 51309 43270 54546 43272
rect 51309 43267 51375 43270
rect 54486 43262 54546 43270
rect 54486 43202 55068 43262
rect 88109 43194 88175 43197
rect 51174 43134 51372 43194
rect 84876 43192 88175 43194
rect 84876 43136 88114 43192
rect 88170 43136 88175 43192
rect 84876 43134 88175 43136
rect 51312 43058 51372 43134
rect 88109 43131 88175 43134
rect 123529 43194 123595 43197
rect 160053 43194 160119 43197
rect 123529 43192 127012 43194
rect 123529 43136 123534 43192
rect 123590 43136 127012 43192
rect 123529 43134 127012 43136
rect 156820 43192 160119 43194
rect 156820 43136 160058 43192
rect 160114 43136 160119 43192
rect 156820 43134 160119 43136
rect 123529 43131 123595 43134
rect 160053 43131 160119 43134
rect 123345 43058 123411 43061
rect 51312 42998 55098 43058
rect 47862 42862 48106 42922
rect 47862 42242 47922 42688
rect 48046 42514 48106 42862
rect 55038 42688 55098 42998
rect 123345 43056 127042 43058
rect 123345 43000 123350 43056
rect 123406 43000 127042 43056
rect 123345 42998 127042 43000
rect 123345 42995 123411 42998
rect 88293 42650 88359 42653
rect 84876 42648 88359 42650
rect 84876 42592 88298 42648
rect 88354 42592 88359 42648
rect 84876 42590 88359 42592
rect 88293 42587 88359 42590
rect 88661 42514 88727 42517
rect 92022 42514 92082 42824
rect 48046 42454 55098 42514
rect 47862 42182 51418 42242
rect 51217 42106 51283 42109
rect 47862 42104 51283 42106
rect 47862 42048 51222 42104
rect 51278 42048 51283 42104
rect 47862 42046 51283 42048
rect 47862 42008 47922 42046
rect 51217 42043 51283 42046
rect 51358 41970 51418 42182
rect 55038 42144 55098 42454
rect 88661 42512 92082 42514
rect 88661 42456 88666 42512
rect 88722 42456 92082 42512
rect 88661 42454 92082 42456
rect 119806 42514 119866 42824
rect 126982 42688 127042 42998
rect 159777 42650 159843 42653
rect 156820 42648 159843 42650
rect 156820 42592 159782 42648
rect 159838 42592 159843 42648
rect 156820 42590 159843 42592
rect 159777 42587 159843 42590
rect 122977 42514 123043 42517
rect 119806 42512 123043 42514
rect 119806 42456 122982 42512
rect 123038 42456 123043 42512
rect 119806 42454 123043 42456
rect 88661 42451 88727 42454
rect 122977 42451 123043 42454
rect 160329 42514 160395 42517
rect 163966 42514 164026 42824
rect 160329 42512 164026 42514
rect 160329 42456 160334 42512
rect 160390 42456 164026 42512
rect 160329 42454 164026 42456
rect 160329 42451 160395 42454
rect 123069 42378 123135 42381
rect 123069 42376 127042 42378
rect 123069 42320 123074 42376
rect 123130 42320 127042 42376
rect 123069 42318 127042 42320
rect 123069 42315 123135 42318
rect 88293 42242 88359 42245
rect 92022 42242 92082 42280
rect 88293 42240 92082 42242
rect 88293 42184 88298 42240
rect 88354 42184 92082 42240
rect 88293 42182 92082 42184
rect 119806 42242 119866 42280
rect 121689 42242 121755 42245
rect 119806 42240 121755 42242
rect 119806 42184 121694 42240
rect 121750 42184 121755 42240
rect 119806 42182 121755 42184
rect 88293 42179 88359 42182
rect 121689 42179 121755 42182
rect 126982 42144 127042 42318
rect 160053 42242 160119 42245
rect 163966 42242 164026 42280
rect 160053 42240 164026 42242
rect 160053 42184 160058 42240
rect 160114 42184 164026 42240
rect 160053 42182 164026 42184
rect 160053 42179 160119 42182
rect 88477 42106 88543 42109
rect 160237 42106 160303 42109
rect 84876 42104 88543 42106
rect 84876 42048 88482 42104
rect 88538 42048 88543 42104
rect 84876 42046 88543 42048
rect 156820 42104 160303 42106
rect 156820 42048 160242 42104
rect 160298 42048 160303 42104
rect 156820 42046 160303 42048
rect 88477 42043 88543 42046
rect 160237 42043 160303 42046
rect 124357 41970 124423 41973
rect 51358 41910 55098 41970
rect 55038 41464 55098 41910
rect 124357 41968 127042 41970
rect 124357 41912 124362 41968
rect 124418 41912 127042 41968
rect 124357 41910 127042 41912
rect 124357 41907 124423 41910
rect 47862 41154 47922 41464
rect 88385 41426 88451 41429
rect 84876 41424 88451 41426
rect 84876 41368 88390 41424
rect 88446 41368 88451 41424
rect 84876 41366 88451 41368
rect 88385 41363 88451 41366
rect 51309 41290 51375 41293
rect 88753 41290 88819 41293
rect 92022 41290 92082 41600
rect 51309 41288 55098 41290
rect 51309 41232 51314 41288
rect 51370 41232 55098 41288
rect 51309 41230 55098 41232
rect 51309 41227 51375 41230
rect 51217 41154 51283 41157
rect 47862 41152 51283 41154
rect 47862 41096 51222 41152
rect 51278 41096 51283 41152
rect 47862 41094 51283 41096
rect 51217 41091 51283 41094
rect 55038 40920 55098 41230
rect 88753 41288 92082 41290
rect 88753 41232 88758 41288
rect 88814 41232 92082 41288
rect 88753 41230 92082 41232
rect 119806 41290 119866 41600
rect 126982 41464 127042 41910
rect 160145 41426 160211 41429
rect 156820 41424 160211 41426
rect 156820 41368 160150 41424
rect 160206 41368 160211 41424
rect 156820 41366 160211 41368
rect 160145 41363 160211 41366
rect 122977 41290 123043 41293
rect 119806 41288 123043 41290
rect 119806 41232 122982 41288
rect 123038 41232 123043 41288
rect 119806 41230 123043 41232
rect 88753 41227 88819 41230
rect 122977 41227 123043 41230
rect 123161 41290 123227 41293
rect 160421 41290 160487 41293
rect 163966 41290 164026 41600
rect 123161 41288 127042 41290
rect 123161 41232 123166 41288
rect 123222 41232 127042 41288
rect 123161 41230 127042 41232
rect 123161 41227 123227 41230
rect 47862 40610 47922 40920
rect 88477 40882 88543 40885
rect 84876 40880 88543 40882
rect 84876 40824 88482 40880
rect 88538 40824 88543 40880
rect 84876 40822 88543 40824
rect 88477 40819 88543 40822
rect 88385 40610 88451 40613
rect 92022 40610 92082 41056
rect 119806 40882 119866 41056
rect 126982 40920 127042 41230
rect 160421 41288 164026 41290
rect 160421 41232 160426 41288
rect 160482 41232 164026 41288
rect 160421 41230 164026 41232
rect 160421 41227 160487 41230
rect 121689 40882 121755 40885
rect 160237 40882 160303 40885
rect 119806 40880 121755 40882
rect 119806 40824 121694 40880
rect 121750 40824 121755 40880
rect 119806 40822 121755 40824
rect 156820 40880 160303 40882
rect 156820 40824 160242 40880
rect 160298 40824 160303 40880
rect 156820 40822 160303 40824
rect 121689 40819 121755 40822
rect 160237 40819 160303 40822
rect 47862 40550 51234 40610
rect 9896 40474 10376 40504
rect 13313 40474 13379 40477
rect 9896 40472 13379 40474
rect 9896 40416 13318 40472
rect 13374 40416 13379 40472
rect 9896 40414 13379 40416
rect 9896 40384 10376 40414
rect 13313 40411 13379 40414
rect 51174 40338 51234 40550
rect 88385 40608 92082 40610
rect 88385 40552 88390 40608
rect 88446 40552 92082 40608
rect 88385 40550 92082 40552
rect 160237 40610 160303 40613
rect 163966 40610 164026 41056
rect 160237 40608 164026 40610
rect 160237 40552 160242 40608
rect 160298 40552 164026 40608
rect 160237 40550 164026 40552
rect 88385 40547 88451 40550
rect 160237 40547 160303 40550
rect 51309 40474 51375 40477
rect 124265 40474 124331 40477
rect 51309 40472 55098 40474
rect 51309 40416 51314 40472
rect 51370 40416 55098 40472
rect 51309 40414 55098 40416
rect 51309 40411 51375 40414
rect 51174 40278 51418 40338
rect 18005 40202 18071 40205
rect 18005 40200 19954 40202
rect 18005 40144 18010 40200
rect 18066 40144 19954 40200
rect 18005 40142 19954 40144
rect 18005 40139 18071 40142
rect 19894 39560 19954 40142
rect 47862 39930 47922 40240
rect 51358 40066 51418 40278
rect 55038 40240 55098 40414
rect 124265 40472 127042 40474
rect 124265 40416 124270 40472
rect 124326 40416 127042 40472
rect 124265 40414 127042 40416
rect 124265 40411 124331 40414
rect 88293 40202 88359 40205
rect 84876 40200 88359 40202
rect 84876 40144 88298 40200
rect 88354 40144 88359 40200
rect 84876 40142 88359 40144
rect 88293 40139 88359 40142
rect 88569 40066 88635 40069
rect 92022 40066 92082 40376
rect 51358 40006 55098 40066
rect 51217 39930 51283 39933
rect 47862 39928 51283 39930
rect 47862 39872 51222 39928
rect 51278 39872 51283 39928
rect 47862 39870 51283 39872
rect 51217 39867 51283 39870
rect 55038 39696 55098 40006
rect 88569 40064 92082 40066
rect 88569 40008 88574 40064
rect 88630 40008 92082 40064
rect 88569 40006 92082 40008
rect 119806 40066 119866 40376
rect 126982 40240 127042 40414
rect 160053 40202 160119 40205
rect 156820 40200 160119 40202
rect 156820 40144 160058 40200
rect 160114 40144 160119 40200
rect 156820 40142 160119 40144
rect 160053 40139 160119 40142
rect 123161 40066 123227 40069
rect 119806 40064 123227 40066
rect 119806 40008 123166 40064
rect 123222 40008 123227 40064
rect 119806 40006 123227 40008
rect 88569 40003 88635 40006
rect 123161 40003 123227 40006
rect 160329 40066 160395 40069
rect 163966 40066 164026 40376
rect 160329 40064 164026 40066
rect 160329 40008 160334 40064
rect 160390 40008 164026 40064
rect 160329 40006 164026 40008
rect 160329 40003 160395 40006
rect 123069 39930 123135 39933
rect 123069 39928 127042 39930
rect 123069 39872 123074 39928
rect 123130 39872 127042 39928
rect 123069 39870 127042 39872
rect 123069 39867 123135 39870
rect 47862 39386 47922 39696
rect 88477 39658 88543 39661
rect 84876 39656 88543 39658
rect 84876 39600 88482 39656
rect 88538 39600 88543 39656
rect 84876 39598 88543 39600
rect 88477 39595 88543 39598
rect 88661 39386 88727 39389
rect 92022 39386 92082 39832
rect 47862 39326 51234 39386
rect 47862 38706 47922 39152
rect 51174 38978 51234 39326
rect 88661 39384 92082 39386
rect 88661 39328 88666 39384
rect 88722 39328 92082 39384
rect 88661 39326 92082 39328
rect 119806 39386 119866 39832
rect 126982 39696 127042 39870
rect 160421 39658 160487 39661
rect 156820 39656 160487 39658
rect 156820 39600 160426 39656
rect 160482 39600 160487 39656
rect 156820 39598 160487 39600
rect 160421 39595 160487 39598
rect 122977 39386 123043 39389
rect 119806 39384 123043 39386
rect 119806 39328 122982 39384
rect 123038 39328 123043 39384
rect 119806 39326 123043 39328
rect 88661 39323 88727 39326
rect 122977 39323 123043 39326
rect 160513 39386 160579 39389
rect 163966 39386 164026 39832
rect 160513 39384 164026 39386
rect 160513 39328 160518 39384
rect 160574 39328 164026 39384
rect 160513 39326 164026 39328
rect 160513 39323 160579 39326
rect 51309 39114 51375 39117
rect 88385 39114 88451 39117
rect 51309 39112 55068 39114
rect 51309 39056 51314 39112
rect 51370 39056 55068 39112
rect 51309 39054 55068 39056
rect 84876 39112 88451 39114
rect 84876 39056 88390 39112
rect 88446 39056 88451 39112
rect 84876 39054 88451 39056
rect 51309 39051 51375 39054
rect 88385 39051 88451 39054
rect 51174 38918 55098 38978
rect 47862 38646 48106 38706
rect 47862 38162 47922 38472
rect 48046 38298 48106 38646
rect 55038 38472 55098 38918
rect 88753 38842 88819 38845
rect 92022 38842 92082 39152
rect 88753 38840 92082 38842
rect 88753 38784 88758 38840
rect 88814 38784 92082 38840
rect 88753 38782 92082 38784
rect 119806 38842 119866 39152
rect 124357 39114 124423 39117
rect 160237 39114 160303 39117
rect 124357 39112 127012 39114
rect 124357 39056 124362 39112
rect 124418 39056 127012 39112
rect 124357 39054 127012 39056
rect 156820 39112 160303 39114
rect 156820 39056 160242 39112
rect 160298 39056 160303 39112
rect 156820 39054 160303 39056
rect 124357 39051 124423 39054
rect 160237 39051 160303 39054
rect 123161 38978 123227 38981
rect 123161 38976 127042 38978
rect 123161 38920 123166 38976
rect 123222 38920 127042 38976
rect 123161 38918 127042 38920
rect 123161 38915 123227 38918
rect 121781 38842 121847 38845
rect 119806 38840 121847 38842
rect 119806 38784 121786 38840
rect 121842 38784 121847 38840
rect 119806 38782 121847 38784
rect 88753 38779 88819 38782
rect 121781 38779 121847 38782
rect 88477 38434 88543 38437
rect 84876 38432 88543 38434
rect 84876 38376 88482 38432
rect 88538 38376 88543 38432
rect 84876 38374 88543 38376
rect 88477 38371 88543 38374
rect 88477 38298 88543 38301
rect 48046 38238 55098 38298
rect 47862 38102 51418 38162
rect 51217 38026 51283 38029
rect 47862 38024 51283 38026
rect 47862 37968 51222 38024
rect 51278 37968 51283 38024
rect 47862 37966 51283 37968
rect 47862 37928 47922 37966
rect 51217 37963 51283 37966
rect 51358 37754 51418 38102
rect 55038 37928 55098 38238
rect 84846 38296 88543 38298
rect 84846 38240 88482 38296
rect 88538 38240 88543 38296
rect 84846 38238 88543 38240
rect 84846 37860 84906 38238
rect 88477 38235 88543 38238
rect 88569 38162 88635 38165
rect 92022 38162 92082 38608
rect 119806 38434 119866 38608
rect 126982 38472 127042 38918
rect 160421 38842 160487 38845
rect 163966 38842 164026 39152
rect 160421 38840 164026 38842
rect 160421 38784 160426 38840
rect 160482 38784 164026 38840
rect 160421 38782 164026 38784
rect 160421 38779 160487 38782
rect 121689 38434 121755 38437
rect 160237 38434 160303 38437
rect 119806 38432 121755 38434
rect 119806 38376 121694 38432
rect 121750 38376 121755 38432
rect 119806 38374 121755 38376
rect 156820 38432 160303 38434
rect 156820 38376 160242 38432
rect 160298 38376 160303 38432
rect 156820 38374 160303 38376
rect 121689 38371 121755 38374
rect 160237 38371 160303 38374
rect 123069 38298 123135 38301
rect 160329 38298 160395 38301
rect 163966 38298 164026 38608
rect 123069 38296 127042 38298
rect 123069 38240 123074 38296
rect 123130 38240 127042 38296
rect 123069 38238 127042 38240
rect 123069 38235 123135 38238
rect 88569 38160 92082 38162
rect 88569 38104 88574 38160
rect 88630 38104 92082 38160
rect 88569 38102 92082 38104
rect 88569 38099 88635 38102
rect 126982 37928 127042 38238
rect 160329 38296 164026 38298
rect 160329 38240 160334 38296
rect 160390 38240 164026 38296
rect 160329 38238 164026 38240
rect 160329 38235 160395 38238
rect 160145 38026 160211 38029
rect 160145 38024 160714 38026
rect 160145 37968 160150 38024
rect 160206 37968 160714 38024
rect 160145 37966 160714 37968
rect 160145 37963 160211 37966
rect 88477 37890 88543 37893
rect 92022 37890 92082 37928
rect 88477 37888 92082 37890
rect 88477 37832 88482 37888
rect 88538 37832 92082 37888
rect 88477 37830 92082 37832
rect 119806 37890 119866 37928
rect 121689 37890 121755 37893
rect 159041 37890 159107 37893
rect 160421 37890 160487 37893
rect 119806 37888 121755 37890
rect 119806 37832 121694 37888
rect 121750 37832 121755 37888
rect 119806 37830 121755 37832
rect 156820 37888 159107 37890
rect 156820 37832 159046 37888
rect 159102 37832 159107 37888
rect 156820 37830 159107 37832
rect 88477 37827 88543 37830
rect 121689 37827 121755 37830
rect 159041 37827 159107 37830
rect 160240 37888 160487 37890
rect 160240 37832 160426 37888
rect 160482 37832 160487 37888
rect 160240 37830 160487 37832
rect 160654 37890 160714 37966
rect 163966 37890 164026 37928
rect 160654 37830 164026 37890
rect 123897 37754 123963 37757
rect 160240 37754 160300 37830
rect 160421 37827 160487 37830
rect 51358 37694 55098 37754
rect 55038 37248 55098 37694
rect 123897 37752 127042 37754
rect 123897 37696 123902 37752
rect 123958 37696 127042 37752
rect 123897 37694 127042 37696
rect 123897 37691 123963 37694
rect 47862 36938 47922 37248
rect 88201 37210 88267 37213
rect 84876 37208 88267 37210
rect 84876 37152 88206 37208
rect 88262 37152 88267 37208
rect 84876 37150 88267 37152
rect 88201 37147 88267 37150
rect 51309 37074 51375 37077
rect 51309 37072 55098 37074
rect 51309 37016 51314 37072
rect 51370 37016 55098 37072
rect 51309 37014 55098 37016
rect 51309 37011 51375 37014
rect 51217 36938 51283 36941
rect 47862 36936 51283 36938
rect 47862 36880 51222 36936
rect 51278 36880 51283 36936
rect 47862 36878 51283 36880
rect 51217 36875 51283 36878
rect 55038 36704 55098 37014
rect 88661 36938 88727 36941
rect 92022 36938 92082 37384
rect 88661 36936 92082 36938
rect 88661 36880 88666 36936
rect 88722 36880 92082 36936
rect 88661 36878 92082 36880
rect 119806 36938 119866 37384
rect 126982 37248 127042 37694
rect 156790 37694 160300 37754
rect 156790 37180 156850 37694
rect 123437 37074 123503 37077
rect 123437 37072 127042 37074
rect 123437 37016 123442 37072
rect 123498 37016 127042 37072
rect 123437 37014 127042 37016
rect 123437 37011 123503 37014
rect 122977 36938 123043 36941
rect 119806 36936 123043 36938
rect 119806 36880 122982 36936
rect 123038 36880 123043 36936
rect 119806 36878 123043 36880
rect 88661 36875 88727 36878
rect 122977 36875 123043 36878
rect 126982 36704 127042 37014
rect 160329 36938 160395 36941
rect 163966 36938 164026 37384
rect 160329 36936 164026 36938
rect 160329 36880 160334 36936
rect 160390 36880 164026 36936
rect 160329 36878 164026 36880
rect 160329 36875 160395 36878
rect 47862 36666 47922 36704
rect 51217 36666 51283 36669
rect 88569 36666 88635 36669
rect 47862 36664 51283 36666
rect 47862 36608 51222 36664
rect 51278 36608 51283 36664
rect 47862 36606 51283 36608
rect 84876 36664 88635 36666
rect 84876 36608 88574 36664
rect 88630 36608 88635 36664
rect 84876 36606 88635 36608
rect 51217 36603 51283 36606
rect 88569 36603 88635 36606
rect 88385 36530 88451 36533
rect 92022 36530 92082 36704
rect 88385 36528 92082 36530
rect 88385 36472 88390 36528
rect 88446 36472 92082 36528
rect 88385 36470 92082 36472
rect 119806 36530 119866 36704
rect 160237 36666 160303 36669
rect 156820 36664 160303 36666
rect 156820 36608 160242 36664
rect 160298 36608 160303 36664
rect 156820 36606 160303 36608
rect 160237 36603 160303 36606
rect 123253 36530 123319 36533
rect 119806 36528 123319 36530
rect 119806 36472 123258 36528
rect 123314 36472 123319 36528
rect 119806 36470 123319 36472
rect 88385 36467 88451 36470
rect 123253 36467 123319 36470
rect 160237 36530 160303 36533
rect 163966 36530 164026 36704
rect 160237 36528 164026 36530
rect 160237 36472 160242 36528
rect 160298 36472 164026 36528
rect 160237 36470 164026 36472
rect 160237 36467 160303 36470
rect 51401 36394 51467 36397
rect 124357 36394 124423 36397
rect 51401 36392 55098 36394
rect 51401 36336 51406 36392
rect 51462 36336 55098 36392
rect 51401 36334 55098 36336
rect 51401 36331 51467 36334
rect 55038 36160 55098 36334
rect 124357 36392 127042 36394
rect 124357 36336 124362 36392
rect 124418 36336 127042 36392
rect 124357 36334 127042 36336
rect 124357 36331 124423 36334
rect 126982 36160 127042 36334
rect 47862 35714 47922 36160
rect 88477 36122 88543 36125
rect 84876 36120 88543 36122
rect 84876 36064 88482 36120
rect 88538 36064 88543 36120
rect 84876 36062 88543 36064
rect 88477 36059 88543 36062
rect 51309 35986 51375 35989
rect 51309 35984 55098 35986
rect 51309 35928 51314 35984
rect 51370 35928 55098 35984
rect 51309 35926 55098 35928
rect 51309 35923 51375 35926
rect 47862 35654 51234 35714
rect 47862 35170 47922 35480
rect 51174 35306 51234 35654
rect 55038 35480 55098 35926
rect 88661 35714 88727 35717
rect 92022 35714 92082 36160
rect 88661 35712 92082 35714
rect 88661 35656 88666 35712
rect 88722 35656 92082 35712
rect 88661 35654 92082 35656
rect 119806 35714 119866 36160
rect 160145 36122 160211 36125
rect 156820 36120 160211 36122
rect 156820 36064 160150 36120
rect 160206 36064 160211 36120
rect 156820 36062 160211 36064
rect 160145 36059 160211 36062
rect 123069 35986 123135 35989
rect 123069 35984 127042 35986
rect 123069 35928 123074 35984
rect 123130 35928 127042 35984
rect 123069 35926 127042 35928
rect 123069 35923 123135 35926
rect 122977 35714 123043 35717
rect 119806 35712 123043 35714
rect 119806 35656 122982 35712
rect 123038 35656 123043 35712
rect 119806 35654 123043 35656
rect 88661 35651 88727 35654
rect 122977 35651 123043 35654
rect 126982 35480 127042 35926
rect 160421 35714 160487 35717
rect 163966 35714 164026 36160
rect 160421 35712 164026 35714
rect 160421 35656 160426 35712
rect 160482 35656 164026 35712
rect 160421 35654 164026 35656
rect 160421 35651 160487 35654
rect 88477 35442 88543 35445
rect 84876 35440 88543 35442
rect 84876 35384 88482 35440
rect 88538 35384 88543 35440
rect 84876 35382 88543 35384
rect 88477 35379 88543 35382
rect 88293 35306 88359 35309
rect 92022 35306 92082 35480
rect 51174 35246 51418 35306
rect 47862 35110 51234 35170
rect 47862 34490 47922 34936
rect 51174 34898 51234 35110
rect 51358 35034 51418 35246
rect 88293 35304 92082 35306
rect 88293 35248 88298 35304
rect 88354 35248 92082 35304
rect 88293 35246 92082 35248
rect 119806 35306 119866 35480
rect 160329 35442 160395 35445
rect 156820 35440 160395 35442
rect 156820 35384 160334 35440
rect 160390 35384 160395 35440
rect 156820 35382 160395 35384
rect 160329 35379 160395 35382
rect 121689 35306 121755 35309
rect 119806 35304 121755 35306
rect 119806 35248 121694 35304
rect 121750 35248 121755 35304
rect 119806 35246 121755 35248
rect 88293 35243 88359 35246
rect 121689 35243 121755 35246
rect 160053 35170 160119 35173
rect 163966 35170 164026 35480
rect 160053 35168 164026 35170
rect 160053 35112 160058 35168
rect 160114 35112 164026 35168
rect 160053 35110 164026 35112
rect 160053 35107 160119 35110
rect 51358 34974 54546 35034
rect 54486 34966 54546 34974
rect 54486 34906 55068 34966
rect 88385 34898 88451 34901
rect 51174 34838 51418 34898
rect 84876 34896 88451 34898
rect 84876 34840 88390 34896
rect 88446 34840 88451 34896
rect 84876 34838 88451 34840
rect 51358 34762 51418 34838
rect 88385 34835 88451 34838
rect 51358 34702 55098 34762
rect 51217 34490 51283 34493
rect 47862 34488 51283 34490
rect 47862 34432 51222 34488
rect 51278 34432 51283 34488
rect 47862 34430 51283 34432
rect 51217 34427 51283 34430
rect 55038 34256 55098 34702
rect 88569 34490 88635 34493
rect 92022 34490 92082 34936
rect 88569 34488 92082 34490
rect 88569 34432 88574 34488
rect 88630 34432 92082 34488
rect 88569 34430 92082 34432
rect 119806 34490 119866 34936
rect 123253 34898 123319 34901
rect 160237 34898 160303 34901
rect 123253 34896 127012 34898
rect 123253 34840 123258 34896
rect 123314 34840 127012 34896
rect 123253 34838 127012 34840
rect 156820 34896 160303 34898
rect 156820 34840 160242 34896
rect 160298 34840 160303 34896
rect 156820 34838 160303 34840
rect 123253 34835 123319 34838
rect 160237 34835 160303 34838
rect 123161 34626 123227 34629
rect 123161 34624 127042 34626
rect 123161 34568 123166 34624
rect 123222 34568 127042 34624
rect 123161 34566 127042 34568
rect 123161 34563 123227 34566
rect 121689 34490 121755 34493
rect 119806 34488 121755 34490
rect 119806 34432 121694 34488
rect 121750 34432 121755 34488
rect 119806 34430 121755 34432
rect 88569 34427 88635 34430
rect 121689 34427 121755 34430
rect 126982 34256 127042 34566
rect 160329 34490 160395 34493
rect 163966 34490 164026 34936
rect 160329 34488 164026 34490
rect 160329 34432 160334 34488
rect 160390 34432 164026 34488
rect 160329 34430 164026 34432
rect 160329 34427 160395 34430
rect 47862 34218 47922 34256
rect 50481 34218 50547 34221
rect 88661 34218 88727 34221
rect 47862 34216 50547 34218
rect 47862 34160 50486 34216
rect 50542 34160 50547 34216
rect 47862 34158 50547 34160
rect 84876 34216 88727 34218
rect 84876 34160 88666 34216
rect 88722 34160 88727 34216
rect 84876 34158 88727 34160
rect 50481 34155 50547 34158
rect 88661 34155 88727 34158
rect 51217 34082 51283 34085
rect 47678 34080 51283 34082
rect 47678 34024 51222 34080
rect 51278 34024 51283 34080
rect 47678 34022 51283 34024
rect 47678 33712 47738 34022
rect 51217 34019 51283 34022
rect 88569 33946 88635 33949
rect 92022 33946 92082 34256
rect 88569 33944 92082 33946
rect 88569 33888 88574 33944
rect 88630 33888 92082 33944
rect 88569 33886 92082 33888
rect 119806 33946 119866 34256
rect 160421 34218 160487 34221
rect 156820 34216 160487 34218
rect 156820 34160 160426 34216
rect 160482 34160 160487 34216
rect 156820 34158 160487 34160
rect 160421 34155 160487 34158
rect 122977 33946 123043 33949
rect 119806 33944 123043 33946
rect 119806 33888 122982 33944
rect 123038 33888 123043 33944
rect 119806 33886 123043 33888
rect 88569 33883 88635 33886
rect 122977 33883 123043 33886
rect 160421 33946 160487 33949
rect 163966 33946 164026 34256
rect 160421 33944 164026 33946
rect 160421 33888 160426 33944
rect 160482 33888 164026 33944
rect 160421 33886 164026 33888
rect 160421 33883 160487 33886
rect 50481 33810 50547 33813
rect 88385 33810 88451 33813
rect 121689 33810 121755 33813
rect 50481 33808 51372 33810
rect 50481 33752 50486 33808
rect 50542 33752 51372 33808
rect 50481 33750 51372 33752
rect 50481 33747 50547 33750
rect 51312 33538 51372 33750
rect 88385 33808 92082 33810
rect 88385 33752 88390 33808
rect 88446 33752 92082 33808
rect 88385 33750 92082 33752
rect 88385 33747 88451 33750
rect 92022 33716 92082 33750
rect 119806 33808 121755 33810
rect 119806 33752 121694 33808
rect 121750 33752 121755 33808
rect 119806 33750 121755 33752
rect 119806 33712 119866 33750
rect 121689 33747 121755 33750
rect 160145 33810 160211 33813
rect 160145 33808 164026 33810
rect 160145 33752 160150 33808
rect 160206 33752 164026 33808
rect 160145 33750 164026 33752
rect 160145 33747 160211 33750
rect 163966 33712 164026 33750
rect 51493 33674 51559 33677
rect 88293 33674 88359 33677
rect 51493 33672 55068 33674
rect 51493 33616 51498 33672
rect 51554 33616 55068 33672
rect 51493 33614 55068 33616
rect 84876 33672 88359 33674
rect 84876 33616 88298 33672
rect 88354 33616 88359 33672
rect 84876 33614 88359 33616
rect 51493 33611 51559 33614
rect 88293 33611 88359 33614
rect 123621 33674 123687 33677
rect 160053 33674 160119 33677
rect 123621 33672 127012 33674
rect 123621 33616 123626 33672
rect 123682 33616 127012 33672
rect 123621 33614 127012 33616
rect 156820 33672 160119 33674
rect 156820 33616 160058 33672
rect 160114 33616 160119 33672
rect 156820 33614 160119 33616
rect 123621 33611 123687 33614
rect 160053 33611 160119 33614
rect 124357 33538 124423 33541
rect 51312 33478 55098 33538
rect 55038 33168 55098 33478
rect 124357 33536 127042 33538
rect 124357 33480 124362 33536
rect 124418 33480 127042 33536
rect 124357 33478 127042 33480
rect 124357 33475 124423 33478
rect 126982 33168 127042 33478
rect 47862 32722 47922 33168
rect 88477 33130 88543 33133
rect 84876 33128 88543 33130
rect 84876 33072 88482 33128
rect 88538 33072 88543 33128
rect 84876 33070 88543 33072
rect 88477 33067 88543 33070
rect 51309 32994 51375 32997
rect 51309 32992 55098 32994
rect 51309 32936 51314 32992
rect 51370 32936 55098 32992
rect 51309 32934 55098 32936
rect 51309 32931 51375 32934
rect 50481 32722 50547 32725
rect 47862 32720 50547 32722
rect 47862 32664 50486 32720
rect 50542 32664 50547 32720
rect 47862 32662 50547 32664
rect 50481 32659 50547 32662
rect 55038 32488 55098 32934
rect 88661 32722 88727 32725
rect 92022 32722 92082 33168
rect 119806 32858 119866 33168
rect 160237 33130 160303 33133
rect 156820 33128 160303 33130
rect 156820 33072 160242 33128
rect 160298 33072 160303 33128
rect 156820 33070 160303 33072
rect 160237 33067 160303 33070
rect 123069 32994 123135 32997
rect 123069 32992 127042 32994
rect 123069 32936 123074 32992
rect 123130 32936 127042 32992
rect 123069 32934 127042 32936
rect 123069 32931 123135 32934
rect 122977 32858 123043 32861
rect 119806 32856 123043 32858
rect 119806 32800 122982 32856
rect 123038 32800 123043 32856
rect 119806 32798 123043 32800
rect 122977 32795 123043 32798
rect 88661 32720 92082 32722
rect 88661 32664 88666 32720
rect 88722 32664 92082 32720
rect 88661 32662 92082 32664
rect 88661 32659 88727 32662
rect 126982 32488 127042 32934
rect 160513 32722 160579 32725
rect 163966 32722 164026 33168
rect 160513 32720 164026 32722
rect 160513 32664 160518 32720
rect 160574 32664 164026 32720
rect 160513 32662 164026 32664
rect 160513 32659 160579 32662
rect 47862 32450 47922 32488
rect 51217 32450 51283 32453
rect 88477 32450 88543 32453
rect 47862 32448 51283 32450
rect 47862 32392 51222 32448
rect 51278 32392 51283 32448
rect 47862 32390 51283 32392
rect 84876 32448 88543 32450
rect 84876 32392 88482 32448
rect 88538 32392 88543 32448
rect 84876 32390 88543 32392
rect 51217 32387 51283 32390
rect 88477 32387 88543 32390
rect 50481 32314 50547 32317
rect 88477 32314 88543 32317
rect 92022 32314 92082 32488
rect 119806 32450 119866 32488
rect 121689 32450 121755 32453
rect 160237 32450 160303 32453
rect 119806 32448 121755 32450
rect 119806 32392 121694 32448
rect 121750 32392 121755 32448
rect 119806 32390 121755 32392
rect 156820 32448 160303 32450
rect 156820 32392 160242 32448
rect 160298 32392 160303 32448
rect 156820 32390 160303 32392
rect 121689 32387 121755 32390
rect 160237 32387 160303 32390
rect 50481 32312 51372 32314
rect 50481 32256 50486 32312
rect 50542 32256 51372 32312
rect 50481 32254 51372 32256
rect 50481 32251 50547 32254
rect 51312 32178 51372 32254
rect 88477 32312 92082 32314
rect 88477 32256 88482 32312
rect 88538 32256 92082 32312
rect 88477 32254 92082 32256
rect 160053 32314 160119 32317
rect 163966 32314 164026 32488
rect 160053 32312 164026 32314
rect 160053 32256 160058 32312
rect 160114 32256 164026 32312
rect 160053 32254 164026 32256
rect 88477 32251 88543 32254
rect 160053 32251 160119 32254
rect 124265 32178 124331 32181
rect 51312 32118 55098 32178
rect 55038 31944 55098 32118
rect 124265 32176 127042 32178
rect 124265 32120 124270 32176
rect 124326 32120 127042 32176
rect 124265 32118 127042 32120
rect 124265 32115 124331 32118
rect 126982 31944 127042 32118
rect 47862 31634 47922 31944
rect 88385 31906 88451 31909
rect 84876 31904 88451 31906
rect 84876 31848 88390 31904
rect 88446 31848 88451 31904
rect 84876 31846 88451 31848
rect 88385 31843 88451 31846
rect 51309 31770 51375 31773
rect 51309 31768 55098 31770
rect 51309 31712 51314 31768
rect 51370 31712 55098 31768
rect 51309 31710 55098 31712
rect 51309 31707 51375 31710
rect 51217 31634 51283 31637
rect 47862 31632 51283 31634
rect 47862 31576 51222 31632
rect 51278 31576 51283 31632
rect 47862 31574 51283 31576
rect 51217 31571 51283 31574
rect 47862 30954 47922 31400
rect 55038 31264 55098 31710
rect 88569 31498 88635 31501
rect 92022 31498 92082 31944
rect 88569 31496 92082 31498
rect 88569 31440 88574 31496
rect 88630 31440 92082 31496
rect 88569 31438 92082 31440
rect 119806 31498 119866 31944
rect 160145 31906 160211 31909
rect 156820 31904 160211 31906
rect 156820 31848 160150 31904
rect 160206 31848 160211 31904
rect 156820 31846 160211 31848
rect 160145 31843 160211 31846
rect 123069 31770 123135 31773
rect 123069 31768 127042 31770
rect 123069 31712 123074 31768
rect 123130 31712 127042 31768
rect 123069 31710 127042 31712
rect 123069 31707 123135 31710
rect 122977 31498 123043 31501
rect 119806 31496 123043 31498
rect 119806 31440 122982 31496
rect 123038 31440 123043 31496
rect 119806 31438 123043 31440
rect 88569 31435 88635 31438
rect 122977 31435 123043 31438
rect 126982 31264 127042 31710
rect 160329 31498 160395 31501
rect 163966 31498 164026 31944
rect 160329 31496 164026 31498
rect 160329 31440 160334 31496
rect 160390 31440 164026 31496
rect 160329 31438 164026 31440
rect 160329 31435 160395 31438
rect 88661 31226 88727 31229
rect 84876 31224 88727 31226
rect 84876 31168 88666 31224
rect 88722 31168 88727 31224
rect 84876 31166 88727 31168
rect 88661 31163 88727 31166
rect 88385 30954 88451 30957
rect 92022 30954 92082 31264
rect 119806 31226 119866 31264
rect 121689 31226 121755 31229
rect 160237 31226 160303 31229
rect 119806 31224 121755 31226
rect 119806 31168 121694 31224
rect 121750 31168 121755 31224
rect 119806 31166 121755 31168
rect 156820 31224 160303 31226
rect 156820 31168 160242 31224
rect 160298 31168 160303 31224
rect 156820 31166 160303 31168
rect 121689 31163 121755 31166
rect 160237 31163 160303 31166
rect 47862 30894 51234 30954
rect 47862 30410 47922 30720
rect 51174 30682 51234 30894
rect 88385 30952 92082 30954
rect 88385 30896 88390 30952
rect 88446 30896 92082 30952
rect 88385 30894 92082 30896
rect 160145 30954 160211 30957
rect 163966 30954 164026 31264
rect 160145 30952 164026 30954
rect 160145 30896 160150 30952
rect 160206 30896 164026 30952
rect 160145 30894 164026 30896
rect 88385 30891 88451 30894
rect 160145 30891 160211 30894
rect 51309 30818 51375 30821
rect 51309 30816 54546 30818
rect 51309 30760 51314 30816
rect 51370 30760 54546 30816
rect 51309 30758 54546 30760
rect 51309 30755 51375 30758
rect 54486 30750 54546 30758
rect 54486 30690 55068 30750
rect 88477 30682 88543 30685
rect 51174 30622 51372 30682
rect 84876 30680 88543 30682
rect 84876 30624 88482 30680
rect 88538 30624 88543 30680
rect 84876 30622 88543 30624
rect 51312 30546 51372 30622
rect 88477 30619 88543 30622
rect 51312 30486 55098 30546
rect 51217 30410 51283 30413
rect 47862 30408 51283 30410
rect 47862 30352 51222 30408
rect 51278 30352 51283 30408
rect 47862 30350 51283 30352
rect 51217 30347 51283 30350
rect 55038 30176 55098 30486
rect 88661 30274 88727 30277
rect 92022 30274 92082 30720
rect 88661 30272 92082 30274
rect 88661 30216 88666 30272
rect 88722 30216 92082 30272
rect 88661 30214 92082 30216
rect 119806 30274 119866 30720
rect 123989 30682 124055 30685
rect 160053 30682 160119 30685
rect 123989 30680 127012 30682
rect 123989 30624 123994 30680
rect 124050 30624 127012 30680
rect 123989 30622 127012 30624
rect 156820 30680 160119 30682
rect 156820 30624 160058 30680
rect 160114 30624 160119 30680
rect 156820 30622 160119 30624
rect 123989 30619 124055 30622
rect 160053 30619 160119 30622
rect 123069 30546 123135 30549
rect 123069 30544 127042 30546
rect 123069 30488 123074 30544
rect 123130 30488 127042 30544
rect 123069 30486 127042 30488
rect 123069 30483 123135 30486
rect 123161 30274 123227 30277
rect 119806 30272 123227 30274
rect 119806 30216 123166 30272
rect 123222 30216 123227 30272
rect 119806 30214 123227 30216
rect 88661 30211 88727 30214
rect 123161 30211 123227 30214
rect 126982 30176 127042 30486
rect 160421 30274 160487 30277
rect 163966 30274 164026 30720
rect 160421 30272 164026 30274
rect 160421 30216 160426 30272
rect 160482 30216 164026 30272
rect 160421 30214 164026 30216
rect 160421 30211 160487 30214
rect 47862 29730 47922 30176
rect 88477 30138 88543 30141
rect 160237 30138 160303 30141
rect 84876 30136 88543 30138
rect 84876 30080 88482 30136
rect 88538 30080 88543 30136
rect 84876 30078 88543 30080
rect 156820 30136 160303 30138
rect 156820 30080 160242 30136
rect 160298 30080 160303 30136
rect 156820 30078 160303 30080
rect 88477 30075 88543 30078
rect 160237 30075 160303 30078
rect 88569 29730 88635 29733
rect 92022 29730 92082 30040
rect 47862 29670 51234 29730
rect 47862 29186 47922 29496
rect 51174 29322 51234 29670
rect 88569 29728 92082 29730
rect 88569 29672 88574 29728
rect 88630 29672 92082 29728
rect 88569 29670 92082 29672
rect 119806 29730 119866 30040
rect 122977 29730 123043 29733
rect 119806 29728 123043 29730
rect 119806 29672 122982 29728
rect 123038 29672 123043 29728
rect 119806 29670 123043 29672
rect 88569 29667 88635 29670
rect 122977 29667 123043 29670
rect 160329 29730 160395 29733
rect 163966 29730 164026 30040
rect 160329 29728 164026 29730
rect 160329 29672 160334 29728
rect 160390 29672 164026 29728
rect 160329 29670 164026 29672
rect 160329 29667 160395 29670
rect 51309 29458 51375 29461
rect 88385 29458 88451 29461
rect 51309 29456 55068 29458
rect 51309 29400 51314 29456
rect 51370 29400 55068 29456
rect 51309 29398 55068 29400
rect 84876 29456 88451 29458
rect 84876 29400 88390 29456
rect 88446 29400 88451 29456
rect 84876 29398 88451 29400
rect 51309 29395 51375 29398
rect 88385 29395 88451 29398
rect 51174 29262 55098 29322
rect 47862 29126 48106 29186
rect 47862 28642 47922 28952
rect 48046 28778 48106 29126
rect 55038 28952 55098 29262
rect 88753 29050 88819 29053
rect 92022 29050 92082 29496
rect 119806 29186 119866 29496
rect 124357 29458 124423 29461
rect 160145 29458 160211 29461
rect 124357 29456 127012 29458
rect 124357 29400 124362 29456
rect 124418 29400 127012 29456
rect 124357 29398 127012 29400
rect 156820 29456 160211 29458
rect 156820 29400 160150 29456
rect 160206 29400 160211 29456
rect 156820 29398 160211 29400
rect 124357 29395 124423 29398
rect 160145 29395 160211 29398
rect 123161 29322 123227 29325
rect 123161 29320 127042 29322
rect 123161 29264 123166 29320
rect 123222 29264 127042 29320
rect 123161 29262 127042 29264
rect 123161 29259 123227 29262
rect 121689 29186 121755 29189
rect 119806 29184 121755 29186
rect 119806 29128 121694 29184
rect 121750 29128 121755 29184
rect 119806 29126 121755 29128
rect 121689 29123 121755 29126
rect 88753 29048 92082 29050
rect 88753 28992 88758 29048
rect 88814 28992 92082 29048
rect 88753 28990 92082 28992
rect 88753 28987 88819 28990
rect 126982 28952 127042 29262
rect 160513 29050 160579 29053
rect 163966 29050 164026 29496
rect 160513 29048 164026 29050
rect 160513 28992 160518 29048
rect 160574 28992 164026 29048
rect 160513 28990 164026 28992
rect 160513 28987 160579 28990
rect 88477 28914 88543 28917
rect 160237 28914 160303 28917
rect 84876 28912 88543 28914
rect 84876 28856 88482 28912
rect 88538 28856 88543 28912
rect 84876 28854 88543 28856
rect 156820 28912 160303 28914
rect 156820 28856 160242 28912
rect 160298 28856 160303 28912
rect 156820 28854 160303 28856
rect 88477 28851 88543 28854
rect 160237 28851 160303 28854
rect 88385 28778 88451 28781
rect 48046 28718 55098 28778
rect 51217 28642 51283 28645
rect 47862 28640 51283 28642
rect 47862 28584 51222 28640
rect 51278 28584 51283 28640
rect 47862 28582 51283 28584
rect 51217 28579 51283 28582
rect 47862 28370 47922 28408
rect 51217 28370 51283 28373
rect 47862 28368 51283 28370
rect 47862 28312 51222 28368
rect 51278 28312 51283 28368
rect 47862 28310 51283 28312
rect 51217 28307 51283 28310
rect 55038 28272 55098 28718
rect 84846 28776 88451 28778
rect 84846 28720 88390 28776
rect 88446 28720 88451 28776
rect 84846 28718 88451 28720
rect 84846 28204 84906 28718
rect 88385 28715 88451 28718
rect 88569 28506 88635 28509
rect 92022 28506 92082 28816
rect 119806 28642 119866 28816
rect 123069 28778 123135 28781
rect 123069 28776 127042 28778
rect 123069 28720 123074 28776
rect 123130 28720 127042 28776
rect 123069 28718 127042 28720
rect 123069 28715 123135 28718
rect 121689 28642 121755 28645
rect 119806 28640 121755 28642
rect 119806 28584 121694 28640
rect 121750 28584 121755 28640
rect 119806 28582 121755 28584
rect 121689 28579 121755 28582
rect 88569 28504 92082 28506
rect 88569 28448 88574 28504
rect 88630 28448 92082 28504
rect 88569 28446 92082 28448
rect 88569 28443 88635 28446
rect 126982 28272 127042 28718
rect 160329 28506 160395 28509
rect 163966 28506 164026 28816
rect 160329 28504 164026 28506
rect 160329 28448 160334 28504
rect 160390 28448 164026 28504
rect 160329 28446 164026 28448
rect 160329 28443 160395 28446
rect 88385 28234 88451 28237
rect 92022 28234 92082 28272
rect 88385 28232 92082 28234
rect 88385 28176 88390 28232
rect 88446 28176 92082 28232
rect 88385 28174 92082 28176
rect 119806 28234 119866 28272
rect 121689 28234 121755 28237
rect 160145 28234 160211 28237
rect 160513 28234 160579 28237
rect 119806 28232 121755 28234
rect 119806 28176 121694 28232
rect 121750 28176 121755 28232
rect 119806 28174 121755 28176
rect 156820 28232 160211 28234
rect 156820 28176 160150 28232
rect 160206 28176 160211 28232
rect 156820 28174 160211 28176
rect 88385 28171 88451 28174
rect 121689 28171 121755 28174
rect 160145 28171 160211 28174
rect 160286 28232 160579 28234
rect 160286 28176 160518 28232
rect 160574 28176 160579 28232
rect 160286 28174 160579 28176
rect 51401 28098 51467 28101
rect 123529 28098 123595 28101
rect 160286 28098 160346 28174
rect 160513 28171 160579 28174
rect 160697 28234 160763 28237
rect 163966 28234 164026 28272
rect 160697 28232 164026 28234
rect 160697 28176 160702 28232
rect 160758 28176 164026 28232
rect 160697 28174 164026 28176
rect 160697 28171 160763 28174
rect 51401 28096 55098 28098
rect 51401 28040 51406 28096
rect 51462 28040 55098 28096
rect 51401 28038 55098 28040
rect 51401 28035 51467 28038
rect 55038 27728 55098 28038
rect 123529 28096 127042 28098
rect 123529 28040 123534 28096
rect 123590 28040 127042 28096
rect 123529 28038 127042 28040
rect 123529 28035 123595 28038
rect 126982 27728 127042 28038
rect 156790 28038 160346 28098
rect 47862 27418 47922 27728
rect 88293 27690 88359 27693
rect 84876 27688 88359 27690
rect 84876 27632 88298 27688
rect 88354 27632 88359 27688
rect 156790 27660 156850 28038
rect 84876 27630 88359 27632
rect 88293 27627 88359 27630
rect 51309 27554 51375 27557
rect 51309 27552 55098 27554
rect 51309 27496 51314 27552
rect 51370 27496 55098 27552
rect 51309 27494 55098 27496
rect 51309 27491 51375 27494
rect 51217 27418 51283 27421
rect 47862 27416 51283 27418
rect 47862 27360 51222 27416
rect 51278 27360 51283 27416
rect 47862 27358 51283 27360
rect 51217 27355 51283 27358
rect 55038 27184 55098 27494
rect 88569 27282 88635 27285
rect 92022 27282 92082 27592
rect 88569 27280 92082 27282
rect 88569 27224 88574 27280
rect 88630 27224 92082 27280
rect 88569 27222 92082 27224
rect 119806 27282 119866 27592
rect 124357 27554 124423 27557
rect 124357 27552 127042 27554
rect 124357 27496 124362 27552
rect 124418 27496 127042 27552
rect 124357 27494 127042 27496
rect 124357 27491 124423 27494
rect 122977 27282 123043 27285
rect 119806 27280 123043 27282
rect 119806 27224 122982 27280
rect 123038 27224 123043 27280
rect 119806 27222 123043 27224
rect 88569 27219 88635 27222
rect 122977 27219 123043 27222
rect 126982 27184 127042 27494
rect 160329 27282 160395 27285
rect 163966 27282 164026 27592
rect 160329 27280 164026 27282
rect 160329 27224 160334 27280
rect 160390 27224 164026 27280
rect 160329 27222 164026 27224
rect 160329 27219 160395 27222
rect 47862 26874 47922 27184
rect 88477 27146 88543 27149
rect 160237 27146 160303 27149
rect 84876 27144 88543 27146
rect 84876 27088 88482 27144
rect 88538 27088 88543 27144
rect 84876 27086 88543 27088
rect 156820 27144 160303 27146
rect 156820 27088 160242 27144
rect 160298 27088 160303 27144
rect 156820 27086 160303 27088
rect 88477 27083 88543 27086
rect 160237 27083 160303 27086
rect 88293 26874 88359 26877
rect 92022 26874 92082 27048
rect 47862 26814 51234 26874
rect 51174 26602 51234 26814
rect 88293 26872 92082 26874
rect 88293 26816 88298 26872
rect 88354 26816 92082 26872
rect 88293 26814 92082 26816
rect 119806 26874 119866 27048
rect 123253 26874 123319 26877
rect 119806 26872 123319 26874
rect 119806 26816 123258 26872
rect 123314 26816 123319 26872
rect 119806 26814 123319 26816
rect 88293 26811 88359 26814
rect 123253 26811 123319 26814
rect 160145 26874 160211 26877
rect 163966 26874 164026 27048
rect 160145 26872 164026 26874
rect 160145 26816 160150 26872
rect 160206 26816 164026 26872
rect 160145 26814 164026 26816
rect 160145 26811 160211 26814
rect 51309 26738 51375 26741
rect 124081 26738 124147 26741
rect 51309 26736 55098 26738
rect 51309 26680 51314 26736
rect 51370 26680 55098 26736
rect 51309 26678 55098 26680
rect 51309 26675 51375 26678
rect 51174 26542 51418 26602
rect 47862 26194 47922 26504
rect 51358 26330 51418 26542
rect 55038 26504 55098 26678
rect 124081 26736 127042 26738
rect 124081 26680 124086 26736
rect 124142 26680 127042 26736
rect 124081 26678 127042 26680
rect 124081 26675 124147 26678
rect 126982 26504 127042 26678
rect 88385 26466 88451 26469
rect 159041 26466 159107 26469
rect 84876 26464 88451 26466
rect 84876 26408 88390 26464
rect 88446 26408 88451 26464
rect 84876 26406 88451 26408
rect 156820 26464 159107 26466
rect 156820 26408 159046 26464
rect 159102 26408 159107 26464
rect 156820 26406 159107 26408
rect 88385 26403 88451 26406
rect 159041 26403 159107 26406
rect 51358 26270 55098 26330
rect 51401 26194 51467 26197
rect 47862 26192 51467 26194
rect 47862 26136 51406 26192
rect 51462 26136 51467 26192
rect 47862 26134 51467 26136
rect 51401 26131 51467 26134
rect 55038 25960 55098 26270
rect 88661 26058 88727 26061
rect 92022 26058 92082 26368
rect 88661 26056 92082 26058
rect 88661 26000 88666 26056
rect 88722 26000 92082 26056
rect 88661 25998 92082 26000
rect 119806 26058 119866 26368
rect 123069 26330 123135 26333
rect 123069 26328 127042 26330
rect 123069 26272 123074 26328
rect 123130 26272 127042 26328
rect 123069 26270 127042 26272
rect 123069 26267 123135 26270
rect 123161 26058 123227 26061
rect 119806 26056 123227 26058
rect 119806 26000 123166 26056
rect 123222 26000 123227 26056
rect 119806 25998 123227 26000
rect 88661 25995 88727 25998
rect 123161 25995 123227 25998
rect 126982 25960 127042 26270
rect 160421 26058 160487 26061
rect 163966 26058 164026 26368
rect 160421 26056 164026 26058
rect 160421 26000 160426 26056
rect 160482 26000 164026 26056
rect 160421 25998 164026 26000
rect 160421 25995 160487 25998
rect 47862 25650 47922 25960
rect 88477 25922 88543 25925
rect 160237 25922 160303 25925
rect 84876 25920 88543 25922
rect 84876 25864 88482 25920
rect 88538 25864 88543 25920
rect 84876 25862 88543 25864
rect 156820 25920 160303 25922
rect 156820 25864 160242 25920
rect 160298 25864 160303 25920
rect 156820 25862 160303 25864
rect 88477 25859 88543 25862
rect 160237 25859 160303 25862
rect 51309 25650 51375 25653
rect 47862 25648 51375 25650
rect 47862 25592 51314 25648
rect 51370 25592 51375 25648
rect 47862 25590 51375 25592
rect 51309 25587 51375 25590
rect 88569 25650 88635 25653
rect 92022 25650 92082 25824
rect 88569 25648 92082 25650
rect 88569 25592 88574 25648
rect 88630 25592 92082 25648
rect 88569 25590 92082 25592
rect 88569 25587 88635 25590
rect 18097 25514 18163 25517
rect 19894 25514 19954 25552
rect 51217 25514 51283 25517
rect 51401 25514 51467 25517
rect 18097 25512 19954 25514
rect 18097 25456 18102 25512
rect 18158 25456 19954 25512
rect 18097 25454 19954 25456
rect 47862 25512 51283 25514
rect 47862 25456 51222 25512
rect 51278 25456 51283 25512
rect 47862 25454 51283 25456
rect 18097 25451 18163 25454
rect 47862 25416 47922 25454
rect 51217 25451 51283 25454
rect 51358 25512 51467 25514
rect 51358 25456 51406 25512
rect 51462 25456 51467 25512
rect 51358 25451 51467 25456
rect 119806 25514 119866 25824
rect 122977 25514 123043 25517
rect 119806 25512 123043 25514
rect 119806 25456 122982 25512
rect 123038 25456 123043 25512
rect 119806 25454 123043 25456
rect 122977 25451 123043 25454
rect 160329 25514 160395 25517
rect 163966 25514 164026 25824
rect 160329 25512 164026 25514
rect 160329 25456 160334 25512
rect 160390 25456 164026 25512
rect 160329 25454 164026 25456
rect 160329 25451 160395 25454
rect 51358 25378 51418 25451
rect 51358 25318 54546 25378
rect 54486 25310 54546 25318
rect 54486 25250 55068 25310
rect 88293 25242 88359 25245
rect 84876 25240 88359 25242
rect 84876 25184 88298 25240
rect 88354 25184 88359 25240
rect 84876 25182 88359 25184
rect 88293 25179 88359 25182
rect 123253 25242 123319 25245
rect 160145 25242 160211 25245
rect 123253 25240 127012 25242
rect 123253 25184 123258 25240
rect 123314 25184 127012 25240
rect 123253 25182 127012 25184
rect 156820 25240 160211 25242
rect 156820 25184 160150 25240
rect 160206 25184 160211 25240
rect 156820 25182 160211 25184
rect 123253 25179 123319 25182
rect 160145 25179 160211 25182
rect 51309 25106 51375 25109
rect 88477 25106 88543 25109
rect 51309 25104 55098 25106
rect 51309 25048 51314 25104
rect 51370 25048 55098 25104
rect 51309 25046 55098 25048
rect 51309 25043 51375 25046
rect 55038 24736 55098 25046
rect 84846 25104 88543 25106
rect 84846 25048 88482 25104
rect 88538 25048 88543 25104
rect 84846 25046 88543 25048
rect 47862 24426 47922 24736
rect 84846 24668 84906 25046
rect 88477 25043 88543 25046
rect 88569 24834 88635 24837
rect 92022 24834 92082 25144
rect 88569 24832 92082 24834
rect 88569 24776 88574 24832
rect 88630 24776 92082 24832
rect 88569 24774 92082 24776
rect 119806 24834 119866 25144
rect 123161 25106 123227 25109
rect 160237 25106 160303 25109
rect 123161 25104 127042 25106
rect 123161 25048 123166 25104
rect 123222 25048 127042 25104
rect 123161 25046 127042 25048
rect 123161 25043 123227 25046
rect 121689 24834 121755 24837
rect 119806 24832 121755 24834
rect 119806 24776 121694 24832
rect 121750 24776 121755 24832
rect 119806 24774 121755 24776
rect 88569 24771 88635 24774
rect 121689 24771 121755 24774
rect 126982 24736 127042 25046
rect 156790 25104 160303 25106
rect 156790 25048 160242 25104
rect 160298 25048 160303 25104
rect 156790 25046 160303 25048
rect 156790 24668 156850 25046
rect 160237 25043 160303 25046
rect 160329 24834 160395 24837
rect 163966 24834 164026 25144
rect 160329 24832 164026 24834
rect 160329 24776 160334 24832
rect 160390 24776 164026 24832
rect 160329 24774 164026 24776
rect 160329 24771 160395 24774
rect 51309 24562 51375 24565
rect 51309 24560 55098 24562
rect 51309 24504 51314 24560
rect 51370 24504 55098 24560
rect 51309 24502 55098 24504
rect 51309 24499 51375 24502
rect 47862 24366 51280 24426
rect 47862 24154 47922 24192
rect 51033 24154 51099 24157
rect 47862 24152 51099 24154
rect 47862 24096 51038 24152
rect 51094 24096 51099 24152
rect 47862 24094 51099 24096
rect 51033 24091 51099 24094
rect 51220 24018 51280 24366
rect 55038 24192 55098 24502
rect 88385 24154 88451 24157
rect 92022 24154 92082 24600
rect 84876 24152 88451 24154
rect 84876 24096 88390 24152
rect 88446 24096 88451 24152
rect 84876 24094 88451 24096
rect 88385 24091 88451 24094
rect 88526 24094 92082 24154
rect 119806 24154 119866 24600
rect 123069 24562 123135 24565
rect 123069 24560 127042 24562
rect 123069 24504 123074 24560
rect 123130 24504 127042 24560
rect 123069 24502 127042 24504
rect 123069 24499 123135 24502
rect 126982 24192 127042 24502
rect 160421 24290 160487 24293
rect 163966 24290 164026 24600
rect 160421 24288 164026 24290
rect 160421 24232 160426 24288
rect 160482 24232 164026 24288
rect 160421 24230 164026 24232
rect 160421 24227 160487 24230
rect 122977 24154 123043 24157
rect 158949 24154 159015 24157
rect 119806 24152 123043 24154
rect 119806 24096 122982 24152
rect 123038 24096 123043 24152
rect 119806 24094 123043 24096
rect 156820 24152 159015 24154
rect 156820 24096 158954 24152
rect 159010 24096 159015 24152
rect 156820 24094 159015 24096
rect 87925 24018 87991 24021
rect 88526 24018 88586 24094
rect 122977 24091 123043 24094
rect 158949 24091 159015 24094
rect 51220 23958 55098 24018
rect 47862 23202 47922 23648
rect 55038 23512 55098 23958
rect 87925 24016 88586 24018
rect 87925 23960 87930 24016
rect 87986 23960 88586 24016
rect 87925 23958 88586 23960
rect 87925 23955 87991 23958
rect 88661 23610 88727 23613
rect 92022 23610 92082 23920
rect 88661 23608 92082 23610
rect 88661 23552 88666 23608
rect 88722 23552 92082 23608
rect 88661 23550 92082 23552
rect 119806 23610 119866 23920
rect 123437 23882 123503 23885
rect 123437 23880 127042 23882
rect 123437 23824 123442 23880
rect 123498 23824 127042 23880
rect 123437 23822 127042 23824
rect 123437 23819 123503 23822
rect 123253 23610 123319 23613
rect 119806 23608 123319 23610
rect 119806 23552 123258 23608
rect 123314 23552 123319 23608
rect 119806 23550 123319 23552
rect 88661 23547 88727 23550
rect 123253 23547 123319 23550
rect 126982 23512 127042 23822
rect 160513 23610 160579 23613
rect 163966 23610 164026 23920
rect 160513 23608 164026 23610
rect 160513 23552 160518 23608
rect 160574 23552 164026 23608
rect 160513 23550 164026 23552
rect 160513 23547 160579 23550
rect 88477 23474 88543 23477
rect 160237 23474 160303 23477
rect 84876 23472 88543 23474
rect 84876 23416 88482 23472
rect 88538 23416 88543 23472
rect 84876 23414 88543 23416
rect 156820 23472 160303 23474
rect 156820 23416 160242 23472
rect 160298 23416 160303 23472
rect 156820 23414 160303 23416
rect 88477 23411 88543 23414
rect 160237 23411 160303 23414
rect 51309 23338 51375 23341
rect 51309 23336 55098 23338
rect 51309 23280 51314 23336
rect 51370 23280 55098 23336
rect 51309 23278 55098 23280
rect 51309 23275 51375 23278
rect 51217 23202 51283 23205
rect 47862 23200 51283 23202
rect 47862 23144 51222 23200
rect 51278 23144 51283 23200
rect 47862 23142 51283 23144
rect 51217 23139 51283 23142
rect 55038 22968 55098 23278
rect 47862 22658 47922 22968
rect 87925 22930 87991 22933
rect 84876 22928 87991 22930
rect 84876 22872 87930 22928
rect 87986 22872 87991 22928
rect 84876 22870 87991 22872
rect 87925 22867 87991 22870
rect 88569 22930 88635 22933
rect 92022 22930 92082 23376
rect 119806 23066 119866 23376
rect 123069 23338 123135 23341
rect 123069 23336 127042 23338
rect 123069 23280 123074 23336
rect 123130 23280 127042 23336
rect 123069 23278 127042 23280
rect 123069 23275 123135 23278
rect 122977 23066 123043 23069
rect 119806 23064 123043 23066
rect 119806 23008 122982 23064
rect 123038 23008 123043 23064
rect 119806 23006 123043 23008
rect 122977 23003 123043 23006
rect 126982 22968 127042 23278
rect 160237 22930 160303 22933
rect 88569 22928 92082 22930
rect 88569 22872 88574 22928
rect 88630 22872 92082 22928
rect 88569 22870 92082 22872
rect 156820 22928 160303 22930
rect 156820 22872 160242 22928
rect 160298 22872 160303 22928
rect 156820 22870 160303 22872
rect 88569 22867 88635 22870
rect 160237 22867 160303 22870
rect 160605 22930 160671 22933
rect 163966 22930 164026 23376
rect 160605 22928 164026 22930
rect 160605 22872 160610 22928
rect 160666 22872 164026 22928
rect 160605 22870 164026 22872
rect 160605 22867 160671 22870
rect 88477 22658 88543 22661
rect 92022 22658 92082 22696
rect 47862 22598 51372 22658
rect 47862 21978 47922 22424
rect 51312 22114 51372 22598
rect 88477 22656 92082 22658
rect 88477 22600 88482 22656
rect 88538 22600 92082 22656
rect 88477 22598 92082 22600
rect 119806 22658 119866 22696
rect 123161 22658 123227 22661
rect 160513 22658 160579 22661
rect 119806 22656 123227 22658
rect 119806 22600 123166 22656
rect 123222 22600 123227 22656
rect 119806 22598 123227 22600
rect 88477 22595 88543 22598
rect 123161 22595 123227 22598
rect 160286 22656 160579 22658
rect 160286 22600 160518 22656
rect 160574 22600 160579 22656
rect 160286 22598 160579 22600
rect 51493 22522 51559 22525
rect 88753 22522 88819 22525
rect 122885 22522 122951 22525
rect 51493 22520 55098 22522
rect 51493 22464 51498 22520
rect 51554 22464 55098 22520
rect 51493 22462 55098 22464
rect 51493 22459 51559 22462
rect 55038 22288 55098 22462
rect 88753 22520 92082 22522
rect 88753 22464 88758 22520
rect 88814 22464 92082 22520
rect 88753 22462 92082 22464
rect 88753 22459 88819 22462
rect 88661 22250 88727 22253
rect 84876 22248 88727 22250
rect 84876 22192 88666 22248
rect 88722 22192 88727 22248
rect 84876 22190 88727 22192
rect 88661 22187 88727 22190
rect 92022 22156 92082 22462
rect 119806 22520 122951 22522
rect 119806 22464 122890 22520
rect 122946 22464 122951 22520
rect 119806 22462 122951 22464
rect 119806 22152 119866 22462
rect 122885 22459 122951 22462
rect 123253 22522 123319 22525
rect 160286 22522 160346 22598
rect 160513 22595 160579 22598
rect 160697 22658 160763 22661
rect 163966 22658 164026 22696
rect 160697 22656 164026 22658
rect 160697 22600 160702 22656
rect 160758 22600 164026 22656
rect 160697 22598 164026 22600
rect 160697 22595 160763 22598
rect 123253 22520 127042 22522
rect 123253 22464 123258 22520
rect 123314 22464 127042 22520
rect 123253 22462 127042 22464
rect 123253 22459 123319 22462
rect 126982 22288 127042 22462
rect 156790 22462 160346 22522
rect 160421 22522 160487 22525
rect 160421 22520 164026 22522
rect 160421 22464 160426 22520
rect 160482 22464 164026 22520
rect 160421 22462 164026 22464
rect 156790 22220 156850 22462
rect 160421 22459 160487 22462
rect 163966 22152 164026 22462
rect 123069 22114 123135 22117
rect 51312 22054 55098 22114
rect 51217 21978 51283 21981
rect 47862 21976 51283 21978
rect 47862 21920 51222 21976
rect 51278 21920 51283 21976
rect 47862 21918 51283 21920
rect 51217 21915 51283 21918
rect 50941 21842 51007 21845
rect 47862 21840 51007 21842
rect 47862 21784 50946 21840
rect 51002 21784 51007 21840
rect 47862 21782 51007 21784
rect 47862 21744 47922 21782
rect 50941 21779 51007 21782
rect 55038 21744 55098 22054
rect 123069 22112 127042 22114
rect 123069 22056 123074 22112
rect 123130 22056 127042 22112
rect 123069 22054 127042 22056
rect 123069 22051 123135 22054
rect 88518 21916 88524 21980
rect 88588 21978 88594 21980
rect 122701 21978 122767 21981
rect 88588 21918 92082 21978
rect 88588 21916 88594 21918
rect 88569 21706 88635 21709
rect 84876 21704 88635 21706
rect 84876 21648 88574 21704
rect 88630 21648 88635 21704
rect 84876 21646 88635 21648
rect 88569 21643 88635 21646
rect 92022 21476 92082 21918
rect 119806 21976 122767 21978
rect 119806 21920 122706 21976
rect 122762 21920 122767 21976
rect 119806 21918 122767 21920
rect 119806 21472 119866 21918
rect 122701 21915 122767 21918
rect 126982 21744 127042 22054
rect 160513 21978 160579 21981
rect 160513 21976 164026 21978
rect 160513 21920 160518 21976
rect 160574 21920 164026 21976
rect 160513 21918 164026 21920
rect 160513 21915 160579 21918
rect 160237 21706 160303 21709
rect 156820 21704 160303 21706
rect 156820 21648 160242 21704
rect 160298 21648 160303 21704
rect 156820 21646 160303 21648
rect 160237 21643 160303 21646
rect 163966 21472 164026 21918
rect 47862 21162 47922 21200
rect 50757 21162 50823 21165
rect 47862 21160 50823 21162
rect 47862 21104 50762 21160
rect 50818 21104 50823 21160
rect 47862 21102 50823 21104
rect 50757 21099 50823 21102
rect 51309 21162 51375 21165
rect 88477 21162 88543 21165
rect 122609 21162 122675 21165
rect 51309 21160 55068 21162
rect 51309 21104 51314 21160
rect 51370 21104 55068 21160
rect 51309 21102 55068 21104
rect 84876 21160 88543 21162
rect 84876 21104 88482 21160
rect 88538 21104 88543 21160
rect 84876 21102 88543 21104
rect 51309 21099 51375 21102
rect 88477 21099 88543 21102
rect 119806 21160 122675 21162
rect 119806 21104 122614 21160
rect 122670 21104 122675 21160
rect 119806 21102 122675 21104
rect 51125 21026 51191 21029
rect 47862 21024 51191 21026
rect 47862 20968 51130 21024
rect 51186 20968 51191 21024
rect 47862 20966 51191 20968
rect 47862 20656 47922 20966
rect 51125 20963 51191 20966
rect 58761 21026 58827 21029
rect 67358 21026 67364 21028
rect 58761 21024 67364 21026
rect 58761 20968 58766 21024
rect 58822 20968 67364 21024
rect 58761 20966 67364 20968
rect 58761 20963 58827 20966
rect 67358 20964 67364 20966
rect 67428 20964 67434 21028
rect 88017 21026 88083 21029
rect 88017 21024 92082 21026
rect 88017 20968 88022 21024
rect 88078 20968 92082 21024
rect 88017 20966 92082 20968
rect 88017 20963 88083 20966
rect 92022 20932 92082 20966
rect 119806 20928 119866 21102
rect 122609 21099 122675 21102
rect 123161 21162 123227 21165
rect 159041 21162 159107 21165
rect 123161 21160 127012 21162
rect 123161 21104 123166 21160
rect 123222 21104 127012 21160
rect 123161 21102 127012 21104
rect 156820 21160 159107 21162
rect 156820 21104 159046 21160
rect 159102 21104 159107 21160
rect 156820 21102 159107 21104
rect 123161 21099 123227 21102
rect 159041 21099 159107 21102
rect 160329 21162 160395 21165
rect 160329 21160 164026 21162
rect 160329 21104 160334 21160
rect 160390 21104 164026 21160
rect 160329 21102 164026 21104
rect 160329 21099 160395 21102
rect 129693 21028 129759 21029
rect 129693 21026 129740 21028
rect 129648 21024 129740 21026
rect 129648 20968 129698 21024
rect 129648 20966 129740 20968
rect 129693 20964 129740 20966
rect 129804 20964 129810 21028
rect 130705 21026 130771 21029
rect 131206 21026 131212 21028
rect 130705 21024 131212 21026
rect 130705 20968 130710 21024
rect 130766 20968 131212 21024
rect 130705 20966 131212 20968
rect 129693 20963 129759 20964
rect 130705 20963 130771 20966
rect 131206 20964 131212 20966
rect 131276 20964 131282 21028
rect 163966 20928 164026 21102
rect 60785 20890 60851 20893
rect 67726 20890 67732 20892
rect 60785 20888 67732 20890
rect 60785 20832 60790 20888
rect 60846 20832 67732 20888
rect 60785 20830 67732 20832
rect 60785 20827 60851 20830
rect 67726 20828 67732 20830
rect 67796 20828 67802 20892
rect 135857 20890 135923 20893
rect 136726 20890 136732 20892
rect 135857 20888 136732 20890
rect 135857 20832 135862 20888
rect 135918 20832 136732 20888
rect 135857 20830 136732 20832
rect 135857 20827 135923 20830
rect 136726 20828 136732 20830
rect 136796 20828 136802 20892
rect 59497 20754 59563 20757
rect 67174 20754 67180 20756
rect 59497 20752 67180 20754
rect 59497 20696 59502 20752
rect 59558 20696 67180 20752
rect 59497 20694 67180 20696
rect 59497 20691 59563 20694
rect 67174 20692 67180 20694
rect 67244 20692 67250 20756
rect 88569 20754 88635 20757
rect 122425 20754 122491 20757
rect 88569 20752 92082 20754
rect 88569 20696 88574 20752
rect 88630 20696 92082 20752
rect 88569 20694 92082 20696
rect 88569 20691 88635 20694
rect 50849 20482 50915 20485
rect 47862 20480 50915 20482
rect 47862 20424 50854 20480
rect 50910 20424 50915 20480
rect 47862 20422 50915 20424
rect 47862 19976 47922 20422
rect 50849 20419 50915 20422
rect 92022 20252 92082 20694
rect 119806 20752 122491 20754
rect 119806 20696 122430 20752
rect 122486 20696 122491 20752
rect 119806 20694 122491 20696
rect 119806 20248 119866 20694
rect 122425 20691 122491 20694
rect 159685 20754 159751 20757
rect 159685 20752 164026 20754
rect 159685 20696 159690 20752
rect 159746 20696 164026 20752
rect 159685 20694 164026 20696
rect 159685 20691 159751 20694
rect 163966 20248 164026 20694
rect 196853 20618 196919 20621
rect 201416 20618 201896 20648
rect 196853 20616 201896 20618
rect 196853 20560 196858 20616
rect 196914 20560 201896 20616
rect 196853 20558 201896 20560
rect 196853 20555 196919 20558
rect 201416 20528 201896 20558
rect 50573 19802 50639 19805
rect 47862 19800 50639 19802
rect 47862 19744 50578 19800
rect 50634 19744 50639 19800
rect 47862 19742 50639 19744
rect 47862 19432 47922 19742
rect 50573 19739 50639 19742
rect 88569 19802 88635 19805
rect 122517 19802 122583 19805
rect 88569 19800 92082 19802
rect 88569 19744 88574 19800
rect 88630 19744 92082 19800
rect 88569 19742 92082 19744
rect 88569 19739 88635 19742
rect 92022 19708 92082 19742
rect 119806 19800 122583 19802
rect 119806 19744 122522 19800
rect 122578 19744 122583 19800
rect 119806 19742 122583 19744
rect 119806 19704 119866 19742
rect 122517 19739 122583 19742
rect 159593 19802 159659 19805
rect 159593 19800 164026 19802
rect 159593 19744 159598 19800
rect 159654 19744 164026 19800
rect 159593 19742 164026 19744
rect 159593 19739 159659 19742
rect 163966 19704 164026 19742
rect 87833 19530 87899 19533
rect 122333 19530 122399 19533
rect 87833 19528 92082 19530
rect 87833 19472 87838 19528
rect 87894 19472 92082 19528
rect 87833 19470 92082 19472
rect 87833 19467 87899 19470
rect 9896 19394 10376 19424
rect 13129 19394 13195 19397
rect 9896 19392 13195 19394
rect 9896 19336 13134 19392
rect 13190 19336 13195 19392
rect 9896 19334 13195 19336
rect 9896 19304 10376 19334
rect 13129 19331 13195 19334
rect 50665 19258 50731 19261
rect 47862 19256 50731 19258
rect 47862 19200 50670 19256
rect 50726 19200 50731 19256
rect 47862 19198 50731 19200
rect 47862 18888 47922 19198
rect 50665 19195 50731 19198
rect 66489 19258 66555 19261
rect 66990 19258 66996 19260
rect 66489 19256 66996 19258
rect 66489 19200 66494 19256
rect 66550 19200 66996 19256
rect 66489 19198 66996 19200
rect 66489 19195 66555 19198
rect 66990 19196 66996 19198
rect 67060 19196 67066 19260
rect 92022 19164 92082 19470
rect 119806 19528 122399 19530
rect 119806 19472 122338 19528
rect 122394 19472 122399 19528
rect 119806 19470 122399 19472
rect 119806 19160 119866 19470
rect 122333 19467 122399 19470
rect 160329 19530 160395 19533
rect 160329 19528 164026 19530
rect 160329 19472 160334 19528
rect 160390 19472 164026 19528
rect 160329 19470 164026 19472
rect 160329 19467 160395 19470
rect 163966 19160 164026 19470
rect 127393 18306 127459 18309
rect 139670 18306 139676 18308
rect 127393 18304 139676 18306
rect 127393 18248 127398 18304
rect 127454 18248 139676 18304
rect 127393 18246 139676 18248
rect 127393 18243 127459 18246
rect 139670 18244 139676 18246
rect 139740 18244 139746 18308
rect 132545 18170 132611 18173
rect 138750 18170 138756 18172
rect 132545 18168 138756 18170
rect 132545 18112 132550 18168
rect 132606 18112 138756 18168
rect 132545 18110 138756 18112
rect 132545 18107 132611 18110
rect 138750 18108 138756 18110
rect 138820 18108 138826 18172
rect 56369 18034 56435 18037
rect 67910 18034 67916 18036
rect 56369 18032 67916 18034
rect 56369 17976 56374 18032
rect 56430 17976 67916 18032
rect 56369 17974 67916 17976
rect 56369 17971 56435 17974
rect 67910 17972 67916 17974
rect 67980 17972 67986 18036
rect 128405 18034 128471 18037
rect 140958 18034 140964 18036
rect 128405 18032 140964 18034
rect 128405 17976 128410 18032
rect 128466 17976 140964 18032
rect 128405 17974 140964 17976
rect 128405 17971 128471 17974
rect 140958 17972 140964 17974
rect 141028 17972 141034 18036
rect 57381 17898 57447 17901
rect 67542 17898 67548 17900
rect 57381 17896 67548 17898
rect 57381 17840 57386 17896
rect 57442 17840 67548 17896
rect 57381 17838 67548 17840
rect 57381 17835 57447 17838
rect 67542 17836 67548 17838
rect 67612 17836 67618 17900
rect 131441 17898 131507 17901
rect 138934 17898 138940 17900
rect 131441 17896 138940 17898
rect 131441 17840 131446 17896
rect 131502 17840 138940 17896
rect 131441 17838 138940 17840
rect 131441 17835 131507 17838
rect 138934 17836 138940 17838
rect 139004 17836 139010 17900
rect 177809 17082 177875 17085
rect 187878 17082 187884 17084
rect 177809 17080 187884 17082
rect 177809 17024 177814 17080
rect 177870 17024 187884 17080
rect 177809 17022 187884 17024
rect 177809 17019 177875 17022
rect 187878 17020 187884 17022
rect 187948 17020 187954 17084
<< via3 >>
rect 23572 213132 23636 213196
rect 187148 213132 187212 213196
rect 190644 210684 190708 210748
rect 81716 210276 81780 210340
rect 153476 210276 153540 210340
rect 191564 197356 191628 197420
rect 81716 184980 81780 185044
rect 153476 184980 153540 185044
rect 40316 180492 40380 180556
rect 89076 177228 89140 177292
rect 138756 177228 138820 177292
rect 168380 172060 168444 172124
rect 23572 171788 23636 171852
rect 41604 164172 41668 164236
rect 191196 159140 191260 159204
rect 44364 155740 44428 155804
rect 186044 152476 186108 152540
rect 190644 145812 190708 145876
rect 46388 142548 46452 142612
rect 116860 142608 116924 142612
rect 116860 142552 116874 142608
rect 116874 142552 116924 142608
rect 116860 142548 116924 142552
rect 89628 141732 89692 141796
rect 26148 140372 26212 140436
rect 82268 133028 82332 133092
rect 83556 133088 83620 133092
rect 83556 133032 83606 133088
rect 83606 133032 83620 133088
rect 83556 133028 83620 133032
rect 191564 114940 191628 115004
rect 191748 114532 191812 114596
rect 85212 106840 85276 106844
rect 85212 106784 85226 106840
rect 85226 106784 85276 106840
rect 85212 106780 85276 106784
rect 19892 106100 19956 106164
rect 46388 100660 46452 100724
rect 116860 100660 116924 100724
rect 40316 97804 40380 97868
rect 168380 90324 168444 90388
rect 48412 87196 48476 87260
rect 41604 81892 41668 81956
rect 44364 73732 44428 73796
rect 186044 70332 186108 70396
rect 187884 63804 187948 63868
rect 122012 59860 122076 59924
rect 26148 58092 26212 58156
rect 161756 57412 161820 57476
rect 170220 57412 170284 57476
rect 185860 57276 185924 57340
rect 82268 51564 82332 51628
rect 83556 51624 83620 51628
rect 83556 51568 83606 51624
rect 83606 51568 83620 51624
rect 83556 51564 83620 51568
rect 138756 51428 138820 51492
rect 66996 50204 67060 50268
rect 129740 46668 129804 46732
rect 67732 46532 67796 46596
rect 138940 46532 139004 46596
rect 67180 46396 67244 46460
rect 67364 46260 67428 46324
rect 67548 46124 67612 46188
rect 138756 46396 138820 46460
rect 131212 46260 131276 46324
rect 67916 44628 67980 44692
rect 83556 44628 83620 44692
rect 139676 44688 139740 44692
rect 139676 44632 139726 44688
rect 139726 44632 139740 44688
rect 139676 44628 139740 44632
rect 140964 44688 141028 44692
rect 140964 44632 140978 44688
rect 140978 44632 141028 44688
rect 140964 44628 141028 44632
rect 187148 43676 187212 43740
rect 88524 21916 88588 21980
rect 67364 20964 67428 21028
rect 129740 21024 129804 21028
rect 129740 20968 129754 21024
rect 129754 20968 129804 21024
rect 129740 20964 129804 20968
rect 131212 20964 131276 21028
rect 67732 20828 67796 20892
rect 136732 20828 136796 20892
rect 67180 20692 67244 20756
rect 66996 19196 67060 19260
rect 139676 18244 139740 18308
rect 138756 18108 138820 18172
rect 67916 17972 67980 18036
rect 140964 17972 141028 18036
rect 67548 17836 67612 17900
rect 138940 17836 139004 17900
rect 187884 17020 187948 17084
<< metal4 >>
rect 0 229142 4000 229264
rect 0 228906 122 229142
rect 358 228906 442 229142
rect 678 228906 762 229142
rect 998 228906 1082 229142
rect 1318 228906 1402 229142
rect 1638 228906 1722 229142
rect 1958 228906 2042 229142
rect 2278 228906 2362 229142
rect 2598 228906 2682 229142
rect 2918 228906 3002 229142
rect 3238 228906 3322 229142
rect 3558 228906 3642 229142
rect 3878 228906 4000 229142
rect 0 228822 4000 228906
rect 0 228586 122 228822
rect 358 228586 442 228822
rect 678 228586 762 228822
rect 998 228586 1082 228822
rect 1318 228586 1402 228822
rect 1638 228586 1722 228822
rect 1958 228586 2042 228822
rect 2278 228586 2362 228822
rect 2598 228586 2682 228822
rect 2918 228586 3002 228822
rect 3238 228586 3322 228822
rect 3558 228586 3642 228822
rect 3878 228586 4000 228822
rect 0 228502 4000 228586
rect 0 228266 122 228502
rect 358 228266 442 228502
rect 678 228266 762 228502
rect 998 228266 1082 228502
rect 1318 228266 1402 228502
rect 1638 228266 1722 228502
rect 1958 228266 2042 228502
rect 2278 228266 2362 228502
rect 2598 228266 2682 228502
rect 2918 228266 3002 228502
rect 3238 228266 3322 228502
rect 3558 228266 3642 228502
rect 3878 228266 4000 228502
rect 0 228182 4000 228266
rect 0 227946 122 228182
rect 358 227946 442 228182
rect 678 227946 762 228182
rect 998 227946 1082 228182
rect 1318 227946 1402 228182
rect 1638 227946 1722 228182
rect 1958 227946 2042 228182
rect 2278 227946 2362 228182
rect 2598 227946 2682 228182
rect 2918 227946 3002 228182
rect 3238 227946 3322 228182
rect 3558 227946 3642 228182
rect 3878 227946 4000 228182
rect 0 227862 4000 227946
rect 0 227626 122 227862
rect 358 227626 442 227862
rect 678 227626 762 227862
rect 998 227626 1082 227862
rect 1318 227626 1402 227862
rect 1638 227626 1722 227862
rect 1958 227626 2042 227862
rect 2278 227626 2362 227862
rect 2598 227626 2682 227862
rect 2918 227626 3002 227862
rect 3238 227626 3322 227862
rect 3558 227626 3642 227862
rect 3878 227626 4000 227862
rect 0 227542 4000 227626
rect 0 227306 122 227542
rect 358 227306 442 227542
rect 678 227306 762 227542
rect 998 227306 1082 227542
rect 1318 227306 1402 227542
rect 1638 227306 1722 227542
rect 1958 227306 2042 227542
rect 2278 227306 2362 227542
rect 2598 227306 2682 227542
rect 2918 227306 3002 227542
rect 3238 227306 3322 227542
rect 3558 227306 3642 227542
rect 3878 227306 4000 227542
rect 0 227222 4000 227306
rect 0 226986 122 227222
rect 358 226986 442 227222
rect 678 226986 762 227222
rect 998 226986 1082 227222
rect 1318 226986 1402 227222
rect 1638 226986 1722 227222
rect 1958 226986 2042 227222
rect 2278 226986 2362 227222
rect 2598 226986 2682 227222
rect 2918 226986 3002 227222
rect 3238 226986 3322 227222
rect 3558 226986 3642 227222
rect 3878 226986 4000 227222
rect 0 226902 4000 226986
rect 0 226666 122 226902
rect 358 226666 442 226902
rect 678 226666 762 226902
rect 998 226666 1082 226902
rect 1318 226666 1402 226902
rect 1638 226666 1722 226902
rect 1958 226666 2042 226902
rect 2278 226666 2362 226902
rect 2598 226666 2682 226902
rect 2918 226666 3002 226902
rect 3238 226666 3322 226902
rect 3558 226666 3642 226902
rect 3878 226666 4000 226902
rect 0 226582 4000 226666
rect 0 226346 122 226582
rect 358 226346 442 226582
rect 678 226346 762 226582
rect 998 226346 1082 226582
rect 1318 226346 1402 226582
rect 1638 226346 1722 226582
rect 1958 226346 2042 226582
rect 2278 226346 2362 226582
rect 2598 226346 2682 226582
rect 2918 226346 3002 226582
rect 3238 226346 3322 226582
rect 3558 226346 3642 226582
rect 3878 226346 4000 226582
rect 0 226262 4000 226346
rect 0 226026 122 226262
rect 358 226026 442 226262
rect 678 226026 762 226262
rect 998 226026 1082 226262
rect 1318 226026 1402 226262
rect 1638 226026 1722 226262
rect 1958 226026 2042 226262
rect 2278 226026 2362 226262
rect 2598 226026 2682 226262
rect 2918 226026 3002 226262
rect 3238 226026 3322 226262
rect 3558 226026 3642 226262
rect 3878 226026 4000 226262
rect 0 225942 4000 226026
rect 0 225706 122 225942
rect 358 225706 442 225942
rect 678 225706 762 225942
rect 998 225706 1082 225942
rect 1318 225706 1402 225942
rect 1638 225706 1722 225942
rect 1958 225706 2042 225942
rect 2278 225706 2362 225942
rect 2598 225706 2682 225942
rect 2918 225706 3002 225942
rect 3238 225706 3322 225942
rect 3558 225706 3642 225942
rect 3878 225706 4000 225942
rect 0 225622 4000 225706
rect 0 225386 122 225622
rect 358 225386 442 225622
rect 678 225386 762 225622
rect 998 225386 1082 225622
rect 1318 225386 1402 225622
rect 1638 225386 1722 225622
rect 1958 225386 2042 225622
rect 2278 225386 2362 225622
rect 2598 225386 2682 225622
rect 2918 225386 3002 225622
rect 3238 225386 3322 225622
rect 3558 225386 3642 225622
rect 3878 225386 4000 225622
rect 0 206518 4000 225386
rect 207704 229142 211704 229264
rect 207704 228906 207826 229142
rect 208062 228906 208146 229142
rect 208382 228906 208466 229142
rect 208702 228906 208786 229142
rect 209022 228906 209106 229142
rect 209342 228906 209426 229142
rect 209662 228906 209746 229142
rect 209982 228906 210066 229142
rect 210302 228906 210386 229142
rect 210622 228906 210706 229142
rect 210942 228906 211026 229142
rect 211262 228906 211346 229142
rect 211582 228906 211704 229142
rect 207704 228822 211704 228906
rect 207704 228586 207826 228822
rect 208062 228586 208146 228822
rect 208382 228586 208466 228822
rect 208702 228586 208786 228822
rect 209022 228586 209106 228822
rect 209342 228586 209426 228822
rect 209662 228586 209746 228822
rect 209982 228586 210066 228822
rect 210302 228586 210386 228822
rect 210622 228586 210706 228822
rect 210942 228586 211026 228822
rect 211262 228586 211346 228822
rect 211582 228586 211704 228822
rect 207704 228502 211704 228586
rect 207704 228266 207826 228502
rect 208062 228266 208146 228502
rect 208382 228266 208466 228502
rect 208702 228266 208786 228502
rect 209022 228266 209106 228502
rect 209342 228266 209426 228502
rect 209662 228266 209746 228502
rect 209982 228266 210066 228502
rect 210302 228266 210386 228502
rect 210622 228266 210706 228502
rect 210942 228266 211026 228502
rect 211262 228266 211346 228502
rect 211582 228266 211704 228502
rect 207704 228182 211704 228266
rect 207704 227946 207826 228182
rect 208062 227946 208146 228182
rect 208382 227946 208466 228182
rect 208702 227946 208786 228182
rect 209022 227946 209106 228182
rect 209342 227946 209426 228182
rect 209662 227946 209746 228182
rect 209982 227946 210066 228182
rect 210302 227946 210386 228182
rect 210622 227946 210706 228182
rect 210942 227946 211026 228182
rect 211262 227946 211346 228182
rect 211582 227946 211704 228182
rect 207704 227862 211704 227946
rect 207704 227626 207826 227862
rect 208062 227626 208146 227862
rect 208382 227626 208466 227862
rect 208702 227626 208786 227862
rect 209022 227626 209106 227862
rect 209342 227626 209426 227862
rect 209662 227626 209746 227862
rect 209982 227626 210066 227862
rect 210302 227626 210386 227862
rect 210622 227626 210706 227862
rect 210942 227626 211026 227862
rect 211262 227626 211346 227862
rect 211582 227626 211704 227862
rect 207704 227542 211704 227626
rect 207704 227306 207826 227542
rect 208062 227306 208146 227542
rect 208382 227306 208466 227542
rect 208702 227306 208786 227542
rect 209022 227306 209106 227542
rect 209342 227306 209426 227542
rect 209662 227306 209746 227542
rect 209982 227306 210066 227542
rect 210302 227306 210386 227542
rect 210622 227306 210706 227542
rect 210942 227306 211026 227542
rect 211262 227306 211346 227542
rect 211582 227306 211704 227542
rect 207704 227222 211704 227306
rect 207704 226986 207826 227222
rect 208062 226986 208146 227222
rect 208382 226986 208466 227222
rect 208702 226986 208786 227222
rect 209022 226986 209106 227222
rect 209342 226986 209426 227222
rect 209662 226986 209746 227222
rect 209982 226986 210066 227222
rect 210302 226986 210386 227222
rect 210622 226986 210706 227222
rect 210942 226986 211026 227222
rect 211262 226986 211346 227222
rect 211582 226986 211704 227222
rect 207704 226902 211704 226986
rect 207704 226666 207826 226902
rect 208062 226666 208146 226902
rect 208382 226666 208466 226902
rect 208702 226666 208786 226902
rect 209022 226666 209106 226902
rect 209342 226666 209426 226902
rect 209662 226666 209746 226902
rect 209982 226666 210066 226902
rect 210302 226666 210386 226902
rect 210622 226666 210706 226902
rect 210942 226666 211026 226902
rect 211262 226666 211346 226902
rect 211582 226666 211704 226902
rect 207704 226582 211704 226666
rect 207704 226346 207826 226582
rect 208062 226346 208146 226582
rect 208382 226346 208466 226582
rect 208702 226346 208786 226582
rect 209022 226346 209106 226582
rect 209342 226346 209426 226582
rect 209662 226346 209746 226582
rect 209982 226346 210066 226582
rect 210302 226346 210386 226582
rect 210622 226346 210706 226582
rect 210942 226346 211026 226582
rect 211262 226346 211346 226582
rect 211582 226346 211704 226582
rect 207704 226262 211704 226346
rect 207704 226026 207826 226262
rect 208062 226026 208146 226262
rect 208382 226026 208466 226262
rect 208702 226026 208786 226262
rect 209022 226026 209106 226262
rect 209342 226026 209426 226262
rect 209662 226026 209746 226262
rect 209982 226026 210066 226262
rect 210302 226026 210386 226262
rect 210622 226026 210706 226262
rect 210942 226026 211026 226262
rect 211262 226026 211346 226262
rect 211582 226026 211704 226262
rect 207704 225942 211704 226026
rect 207704 225706 207826 225942
rect 208062 225706 208146 225942
rect 208382 225706 208466 225942
rect 208702 225706 208786 225942
rect 209022 225706 209106 225942
rect 209342 225706 209426 225942
rect 209662 225706 209746 225942
rect 209982 225706 210066 225942
rect 210302 225706 210386 225942
rect 210622 225706 210706 225942
rect 210942 225706 211026 225942
rect 211262 225706 211346 225942
rect 211582 225706 211704 225942
rect 207704 225622 211704 225706
rect 207704 225386 207826 225622
rect 208062 225386 208146 225622
rect 208382 225386 208466 225622
rect 208702 225386 208786 225622
rect 209022 225386 209106 225622
rect 209342 225386 209426 225622
rect 209662 225386 209746 225622
rect 209982 225386 210066 225622
rect 210302 225386 210386 225622
rect 210622 225386 210706 225622
rect 210942 225386 211026 225622
rect 211262 225386 211346 225622
rect 211582 225386 211704 225622
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 4000 206518
rect 0 184118 4000 206282
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 4000 184118
rect 0 161718 4000 183882
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 4000 161718
rect 0 139318 4000 161482
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 4000 139318
rect 0 116918 4000 139082
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 4000 116918
rect 0 94518 4000 116682
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 4000 94518
rect 0 72118 4000 94282
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 4000 72118
rect 0 49718 4000 71882
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 4000 49718
rect 0 27318 4000 49482
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 4000 27318
rect 0 3878 4000 27082
rect 5000 224142 9000 224264
rect 5000 223906 5122 224142
rect 5358 223906 5442 224142
rect 5678 223906 5762 224142
rect 5998 223906 6082 224142
rect 6318 223906 6402 224142
rect 6638 223906 6722 224142
rect 6958 223906 7042 224142
rect 7278 223906 7362 224142
rect 7598 223906 7682 224142
rect 7918 223906 8002 224142
rect 8238 223906 8322 224142
rect 8558 223906 8642 224142
rect 8878 223906 9000 224142
rect 5000 223822 9000 223906
rect 5000 223586 5122 223822
rect 5358 223586 5442 223822
rect 5678 223586 5762 223822
rect 5998 223586 6082 223822
rect 6318 223586 6402 223822
rect 6638 223586 6722 223822
rect 6958 223586 7042 223822
rect 7278 223586 7362 223822
rect 7598 223586 7682 223822
rect 7918 223586 8002 223822
rect 8238 223586 8322 223822
rect 8558 223586 8642 223822
rect 8878 223586 9000 223822
rect 5000 223502 9000 223586
rect 5000 223266 5122 223502
rect 5358 223266 5442 223502
rect 5678 223266 5762 223502
rect 5998 223266 6082 223502
rect 6318 223266 6402 223502
rect 6638 223266 6722 223502
rect 6958 223266 7042 223502
rect 7278 223266 7362 223502
rect 7598 223266 7682 223502
rect 7918 223266 8002 223502
rect 8238 223266 8322 223502
rect 8558 223266 8642 223502
rect 8878 223266 9000 223502
rect 5000 223182 9000 223266
rect 5000 222946 5122 223182
rect 5358 222946 5442 223182
rect 5678 222946 5762 223182
rect 5998 222946 6082 223182
rect 6318 222946 6402 223182
rect 6638 222946 6722 223182
rect 6958 222946 7042 223182
rect 7278 222946 7362 223182
rect 7598 222946 7682 223182
rect 7918 222946 8002 223182
rect 8238 222946 8322 223182
rect 8558 222946 8642 223182
rect 8878 222946 9000 223182
rect 5000 222862 9000 222946
rect 5000 222626 5122 222862
rect 5358 222626 5442 222862
rect 5678 222626 5762 222862
rect 5998 222626 6082 222862
rect 6318 222626 6402 222862
rect 6638 222626 6722 222862
rect 6958 222626 7042 222862
rect 7278 222626 7362 222862
rect 7598 222626 7682 222862
rect 7918 222626 8002 222862
rect 8238 222626 8322 222862
rect 8558 222626 8642 222862
rect 8878 222626 9000 222862
rect 5000 222542 9000 222626
rect 5000 222306 5122 222542
rect 5358 222306 5442 222542
rect 5678 222306 5762 222542
rect 5998 222306 6082 222542
rect 6318 222306 6402 222542
rect 6638 222306 6722 222542
rect 6958 222306 7042 222542
rect 7278 222306 7362 222542
rect 7598 222306 7682 222542
rect 7918 222306 8002 222542
rect 8238 222306 8322 222542
rect 8558 222306 8642 222542
rect 8878 222306 9000 222542
rect 5000 222222 9000 222306
rect 5000 221986 5122 222222
rect 5358 221986 5442 222222
rect 5678 221986 5762 222222
rect 5998 221986 6082 222222
rect 6318 221986 6402 222222
rect 6638 221986 6722 222222
rect 6958 221986 7042 222222
rect 7278 221986 7362 222222
rect 7598 221986 7682 222222
rect 7918 221986 8002 222222
rect 8238 221986 8322 222222
rect 8558 221986 8642 222222
rect 8878 221986 9000 222222
rect 5000 221902 9000 221986
rect 5000 221666 5122 221902
rect 5358 221666 5442 221902
rect 5678 221666 5762 221902
rect 5998 221666 6082 221902
rect 6318 221666 6402 221902
rect 6638 221666 6722 221902
rect 6958 221666 7042 221902
rect 7278 221666 7362 221902
rect 7598 221666 7682 221902
rect 7918 221666 8002 221902
rect 8238 221666 8322 221902
rect 8558 221666 8642 221902
rect 8878 221666 9000 221902
rect 5000 221582 9000 221666
rect 5000 221346 5122 221582
rect 5358 221346 5442 221582
rect 5678 221346 5762 221582
rect 5998 221346 6082 221582
rect 6318 221346 6402 221582
rect 6638 221346 6722 221582
rect 6958 221346 7042 221582
rect 7278 221346 7362 221582
rect 7598 221346 7682 221582
rect 7918 221346 8002 221582
rect 8238 221346 8322 221582
rect 8558 221346 8642 221582
rect 8878 221346 9000 221582
rect 5000 221262 9000 221346
rect 5000 221026 5122 221262
rect 5358 221026 5442 221262
rect 5678 221026 5762 221262
rect 5998 221026 6082 221262
rect 6318 221026 6402 221262
rect 6638 221026 6722 221262
rect 6958 221026 7042 221262
rect 7278 221026 7362 221262
rect 7598 221026 7682 221262
rect 7918 221026 8002 221262
rect 8238 221026 8322 221262
rect 8558 221026 8642 221262
rect 8878 221026 9000 221262
rect 5000 220942 9000 221026
rect 5000 220706 5122 220942
rect 5358 220706 5442 220942
rect 5678 220706 5762 220942
rect 5998 220706 6082 220942
rect 6318 220706 6402 220942
rect 6638 220706 6722 220942
rect 6958 220706 7042 220942
rect 7278 220706 7362 220942
rect 7598 220706 7682 220942
rect 7918 220706 8002 220942
rect 8238 220706 8322 220942
rect 8558 220706 8642 220942
rect 8878 220706 9000 220942
rect 5000 220622 9000 220706
rect 5000 220386 5122 220622
rect 5358 220386 5442 220622
rect 5678 220386 5762 220622
rect 5998 220386 6082 220622
rect 6318 220386 6402 220622
rect 6638 220386 6722 220622
rect 6958 220386 7042 220622
rect 7278 220386 7362 220622
rect 7598 220386 7682 220622
rect 7918 220386 8002 220622
rect 8238 220386 8322 220622
rect 8558 220386 8642 220622
rect 8878 220386 9000 220622
rect 5000 217718 9000 220386
rect 5000 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 9000 217718
rect 5000 195318 9000 217482
rect 202704 224142 206704 224264
rect 202704 223906 202826 224142
rect 203062 223906 203146 224142
rect 203382 223906 203466 224142
rect 203702 223906 203786 224142
rect 204022 223906 204106 224142
rect 204342 223906 204426 224142
rect 204662 223906 204746 224142
rect 204982 223906 205066 224142
rect 205302 223906 205386 224142
rect 205622 223906 205706 224142
rect 205942 223906 206026 224142
rect 206262 223906 206346 224142
rect 206582 223906 206704 224142
rect 202704 223822 206704 223906
rect 202704 223586 202826 223822
rect 203062 223586 203146 223822
rect 203382 223586 203466 223822
rect 203702 223586 203786 223822
rect 204022 223586 204106 223822
rect 204342 223586 204426 223822
rect 204662 223586 204746 223822
rect 204982 223586 205066 223822
rect 205302 223586 205386 223822
rect 205622 223586 205706 223822
rect 205942 223586 206026 223822
rect 206262 223586 206346 223822
rect 206582 223586 206704 223822
rect 202704 223502 206704 223586
rect 202704 223266 202826 223502
rect 203062 223266 203146 223502
rect 203382 223266 203466 223502
rect 203702 223266 203786 223502
rect 204022 223266 204106 223502
rect 204342 223266 204426 223502
rect 204662 223266 204746 223502
rect 204982 223266 205066 223502
rect 205302 223266 205386 223502
rect 205622 223266 205706 223502
rect 205942 223266 206026 223502
rect 206262 223266 206346 223502
rect 206582 223266 206704 223502
rect 202704 223182 206704 223266
rect 202704 222946 202826 223182
rect 203062 222946 203146 223182
rect 203382 222946 203466 223182
rect 203702 222946 203786 223182
rect 204022 222946 204106 223182
rect 204342 222946 204426 223182
rect 204662 222946 204746 223182
rect 204982 222946 205066 223182
rect 205302 222946 205386 223182
rect 205622 222946 205706 223182
rect 205942 222946 206026 223182
rect 206262 222946 206346 223182
rect 206582 222946 206704 223182
rect 202704 222862 206704 222946
rect 202704 222626 202826 222862
rect 203062 222626 203146 222862
rect 203382 222626 203466 222862
rect 203702 222626 203786 222862
rect 204022 222626 204106 222862
rect 204342 222626 204426 222862
rect 204662 222626 204746 222862
rect 204982 222626 205066 222862
rect 205302 222626 205386 222862
rect 205622 222626 205706 222862
rect 205942 222626 206026 222862
rect 206262 222626 206346 222862
rect 206582 222626 206704 222862
rect 202704 222542 206704 222626
rect 202704 222306 202826 222542
rect 203062 222306 203146 222542
rect 203382 222306 203466 222542
rect 203702 222306 203786 222542
rect 204022 222306 204106 222542
rect 204342 222306 204426 222542
rect 204662 222306 204746 222542
rect 204982 222306 205066 222542
rect 205302 222306 205386 222542
rect 205622 222306 205706 222542
rect 205942 222306 206026 222542
rect 206262 222306 206346 222542
rect 206582 222306 206704 222542
rect 202704 222222 206704 222306
rect 202704 221986 202826 222222
rect 203062 221986 203146 222222
rect 203382 221986 203466 222222
rect 203702 221986 203786 222222
rect 204022 221986 204106 222222
rect 204342 221986 204426 222222
rect 204662 221986 204746 222222
rect 204982 221986 205066 222222
rect 205302 221986 205386 222222
rect 205622 221986 205706 222222
rect 205942 221986 206026 222222
rect 206262 221986 206346 222222
rect 206582 221986 206704 222222
rect 202704 221902 206704 221986
rect 202704 221666 202826 221902
rect 203062 221666 203146 221902
rect 203382 221666 203466 221902
rect 203702 221666 203786 221902
rect 204022 221666 204106 221902
rect 204342 221666 204426 221902
rect 204662 221666 204746 221902
rect 204982 221666 205066 221902
rect 205302 221666 205386 221902
rect 205622 221666 205706 221902
rect 205942 221666 206026 221902
rect 206262 221666 206346 221902
rect 206582 221666 206704 221902
rect 202704 221582 206704 221666
rect 202704 221346 202826 221582
rect 203062 221346 203146 221582
rect 203382 221346 203466 221582
rect 203702 221346 203786 221582
rect 204022 221346 204106 221582
rect 204342 221346 204426 221582
rect 204662 221346 204746 221582
rect 204982 221346 205066 221582
rect 205302 221346 205386 221582
rect 205622 221346 205706 221582
rect 205942 221346 206026 221582
rect 206262 221346 206346 221582
rect 206582 221346 206704 221582
rect 202704 221262 206704 221346
rect 202704 221026 202826 221262
rect 203062 221026 203146 221262
rect 203382 221026 203466 221262
rect 203702 221026 203786 221262
rect 204022 221026 204106 221262
rect 204342 221026 204426 221262
rect 204662 221026 204746 221262
rect 204982 221026 205066 221262
rect 205302 221026 205386 221262
rect 205622 221026 205706 221262
rect 205942 221026 206026 221262
rect 206262 221026 206346 221262
rect 206582 221026 206704 221262
rect 202704 220942 206704 221026
rect 202704 220706 202826 220942
rect 203062 220706 203146 220942
rect 203382 220706 203466 220942
rect 203702 220706 203786 220942
rect 204022 220706 204106 220942
rect 204342 220706 204426 220942
rect 204662 220706 204746 220942
rect 204982 220706 205066 220942
rect 205302 220706 205386 220942
rect 205622 220706 205706 220942
rect 205942 220706 206026 220942
rect 206262 220706 206346 220942
rect 206582 220706 206704 220942
rect 202704 220622 206704 220706
rect 202704 220386 202826 220622
rect 203062 220386 203146 220622
rect 203382 220386 203466 220622
rect 203702 220386 203786 220622
rect 204022 220386 204106 220622
rect 204342 220386 204426 220622
rect 204662 220386 204746 220622
rect 204982 220386 205066 220622
rect 205302 220386 205386 220622
rect 205622 220386 205706 220622
rect 205942 220386 206026 220622
rect 206262 220386 206346 220622
rect 206582 220386 206704 220622
rect 202704 217718 206704 220386
rect 202704 217482 202826 217718
rect 203062 217482 203146 217718
rect 203382 217482 203466 217718
rect 203702 217482 203786 217718
rect 204022 217482 204106 217718
rect 204342 217482 204426 217718
rect 204662 217482 204746 217718
rect 204982 217482 205066 217718
rect 205302 217482 205386 217718
rect 205622 217482 205706 217718
rect 205942 217482 206026 217718
rect 206262 217482 206346 217718
rect 206582 217482 206704 217718
rect 23571 213196 23637 213197
rect 23571 213132 23572 213196
rect 23636 213132 23637 213196
rect 23571 213131 23637 213132
rect 187147 213196 187213 213197
rect 187147 213132 187148 213196
rect 187212 213132 187213 213196
rect 187147 213131 187213 213132
rect 5000 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 9000 195318
rect 5000 172918 9000 195082
rect 5000 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 9000 172918
rect 5000 150518 9000 172682
rect 23574 171853 23634 213131
rect 81715 210340 81781 210341
rect 81715 210276 81716 210340
rect 81780 210276 81781 210340
rect 81715 210275 81781 210276
rect 153475 210340 153541 210341
rect 153475 210276 153476 210340
rect 153540 210276 153541 210340
rect 153475 210275 153541 210276
rect 29148 206518 29469 206560
rect 29148 206282 29190 206518
rect 29426 206282 29469 206518
rect 29148 206240 29469 206282
rect 65104 206518 65424 206560
rect 65104 206282 65146 206518
rect 65382 206282 65424 206518
rect 65104 206240 65424 206282
rect 24850 195318 25171 195360
rect 24850 195082 24892 195318
rect 25128 195082 25171 195318
rect 24850 195040 25171 195082
rect 60472 195318 60792 195360
rect 60472 195082 60514 195318
rect 60750 195082 60792 195318
rect 60472 195040 60792 195082
rect 81718 185045 81778 210275
rect 101437 206518 101757 206560
rect 101437 206282 101479 206518
rect 101715 206282 101757 206518
rect 101437 206240 101757 206282
rect 137104 206518 137424 206560
rect 137104 206282 137146 206518
rect 137382 206282 137424 206518
rect 137104 206240 137424 206282
rect 97139 195318 97459 195360
rect 97139 195082 97181 195318
rect 97417 195082 97459 195318
rect 97139 195040 97459 195082
rect 132472 195318 132792 195360
rect 132472 195082 132514 195318
rect 132750 195082 132792 195318
rect 132472 195040 132792 195082
rect 153478 185045 153538 210275
rect 173437 206518 173757 206560
rect 173437 206282 173479 206518
rect 173715 206282 173757 206518
rect 173437 206240 173757 206282
rect 169139 195318 169459 195360
rect 169139 195082 169181 195318
rect 169417 195082 169459 195318
rect 169139 195040 169459 195082
rect 81715 185044 81781 185045
rect 81715 184980 81716 185044
rect 81780 184980 81781 185044
rect 81715 184979 81781 184980
rect 153475 185044 153541 185045
rect 153475 184980 153476 185044
rect 153540 184980 153541 185044
rect 153475 184979 153541 184980
rect 40315 180556 40381 180557
rect 40315 180492 40316 180556
rect 40380 180492 40381 180556
rect 40315 180491 40381 180492
rect 29139 172918 29459 172960
rect 29139 172682 29181 172918
rect 29417 172682 29459 172918
rect 29139 172640 29459 172682
rect 23571 171852 23637 171853
rect 23571 171788 23572 171852
rect 23636 171788 23637 171852
rect 23571 171787 23637 171788
rect 40318 164234 40378 180491
rect 89075 177292 89141 177293
rect 89075 177228 89076 177292
rect 89140 177228 89141 177292
rect 89075 177227 89141 177228
rect 138755 177292 138821 177293
rect 138755 177228 138756 177292
rect 138820 177228 138821 177292
rect 138755 177227 138821 177228
rect 54104 172918 54424 172960
rect 54104 172682 54146 172918
rect 54382 172682 54424 172918
rect 54104 172640 54424 172682
rect 41603 164236 41669 164237
rect 41603 164234 41604 164236
rect 40318 164174 41604 164234
rect 41603 164172 41604 164174
rect 41668 164172 41669 164236
rect 41603 164171 41669 164172
rect 31437 161718 31757 161760
rect 31437 161482 31479 161718
rect 31715 161482 31757 161718
rect 31437 161440 31757 161482
rect 69464 161718 69784 161760
rect 69464 161482 69506 161718
rect 69742 161482 69784 161718
rect 69464 161440 69784 161482
rect 44363 155804 44429 155805
rect 44363 155740 44364 155804
rect 44428 155740 44429 155804
rect 44363 155739 44429 155740
rect 5000 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 9000 150518
rect 5000 128118 9000 150282
rect 29139 150518 29459 150560
rect 29139 150282 29181 150518
rect 29417 150282 29459 150518
rect 29139 150240 29459 150282
rect 44366 140522 44426 155739
rect 54104 150518 54424 150560
rect 54104 150282 54146 150518
rect 54382 150282 54424 150518
rect 54104 150240 54424 150282
rect 46387 142612 46453 142613
rect 46387 142548 46388 142612
rect 46452 142548 46453 142612
rect 46387 142547 46453 142548
rect 31437 139318 31757 139360
rect 31437 139082 31479 139318
rect 31715 139082 31757 139318
rect 31437 139040 31757 139082
rect 5000 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 9000 128118
rect 5000 105718 9000 127882
rect 29437 116918 29757 116960
rect 29437 116682 29479 116918
rect 29715 116682 29757 116918
rect 29437 116640 29757 116682
rect 46390 106522 46450 142547
rect 89078 141794 89138 177227
rect 101139 172918 101459 172960
rect 101139 172682 101181 172918
rect 101417 172682 101459 172918
rect 101139 172640 101459 172682
rect 126104 172918 126424 172960
rect 126104 172682 126146 172918
rect 126382 172682 126424 172918
rect 126104 172640 126424 172682
rect 103437 161718 103757 161760
rect 103437 161482 103479 161718
rect 103715 161482 103757 161718
rect 103437 161440 103757 161482
rect 101139 150518 101459 150560
rect 101139 150282 101181 150518
rect 101417 150282 101459 150518
rect 101139 150240 101459 150282
rect 126104 150518 126424 150560
rect 126104 150282 126146 150518
rect 126382 150282 126424 150518
rect 126104 150240 126424 150282
rect 116859 142612 116925 142613
rect 116859 142548 116860 142612
rect 116924 142548 116925 142612
rect 116859 142547 116925 142548
rect 89627 141796 89693 141797
rect 89627 141794 89628 141796
rect 89078 141734 89628 141794
rect 89627 141732 89628 141734
rect 89692 141732 89693 141796
rect 89627 141731 89693 141732
rect 69464 139318 69784 139360
rect 69464 139082 69506 139318
rect 69742 139082 69784 139318
rect 69464 139040 69784 139082
rect 103437 139318 103757 139360
rect 103437 139082 103479 139318
rect 103715 139082 103757 139318
rect 103437 139040 103757 139082
rect 82267 133092 82333 133093
rect 82267 133028 82268 133092
rect 82332 133028 82333 133092
rect 82267 133027 82333 133028
rect 83555 133092 83621 133093
rect 83555 133028 83556 133092
rect 83620 133028 83621 133092
rect 83555 133027 83621 133028
rect 65104 116918 65424 116960
rect 65104 116682 65146 116918
rect 65382 116682 65424 116918
rect 65104 116640 65424 116682
rect 19894 106165 19954 106286
rect 19891 106164 19957 106165
rect 19891 106100 19892 106164
rect 19956 106100 19957 106164
rect 19891 106099 19957 106100
rect 5000 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 9000 105718
rect 5000 83318 9000 105482
rect 25139 105718 25459 105760
rect 25139 105482 25181 105718
rect 25417 105482 25459 105718
rect 25139 105440 25459 105482
rect 46390 100725 46450 106286
rect 60472 105718 60792 105760
rect 60472 105482 60514 105718
rect 60750 105482 60792 105718
rect 60472 105440 60792 105482
rect 46387 100724 46453 100725
rect 46387 100660 46388 100724
rect 46452 100660 46453 100724
rect 46387 100659 46453 100660
rect 40315 97868 40381 97869
rect 40315 97804 40316 97868
rect 40380 97804 40381 97868
rect 40315 97803 40381 97804
rect 5000 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 9000 83318
rect 5000 60918 9000 83082
rect 29139 83318 29459 83360
rect 29139 83082 29181 83318
rect 29417 83082 29459 83318
rect 29139 83040 29459 83082
rect 40318 81954 40378 97803
rect 48414 87261 48474 92006
rect 48411 87260 48477 87261
rect 48411 87196 48412 87260
rect 48476 87196 48477 87260
rect 48411 87195 48477 87196
rect 54104 83318 54424 83360
rect 54104 83082 54146 83318
rect 54382 83082 54424 83318
rect 54104 83040 54424 83082
rect 41603 81956 41669 81957
rect 41603 81954 41604 81956
rect 40318 81894 41604 81954
rect 41603 81892 41604 81894
rect 41668 81892 41669 81956
rect 41603 81891 41669 81892
rect 44363 73796 44429 73797
rect 44363 73732 44364 73796
rect 44428 73732 44429 73796
rect 44363 73731 44429 73732
rect 31437 72118 31757 72160
rect 31437 71882 31479 72118
rect 31715 71882 31757 72118
rect 31437 71840 31757 71882
rect 5000 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 9000 60918
rect 5000 38518 9000 60682
rect 29139 60918 29459 60960
rect 29139 60682 29181 60918
rect 29417 60682 29459 60918
rect 29139 60640 29459 60682
rect 44366 58242 44426 73731
rect 69464 72118 69784 72160
rect 69464 71882 69506 72118
rect 69742 71882 69784 72118
rect 69464 71840 69784 71882
rect 54104 60918 54424 60960
rect 54104 60682 54146 60918
rect 54382 60682 54424 60918
rect 54104 60640 54424 60682
rect 82270 51629 82330 133027
rect 83558 51629 83618 133027
rect 101437 116918 101757 116960
rect 101437 116682 101479 116918
rect 101715 116682 101757 116918
rect 101437 116640 101757 116682
rect 85211 106844 85277 106845
rect 85211 106780 85212 106844
rect 85276 106780 85277 106844
rect 85211 106779 85277 106780
rect 85214 92242 85274 106779
rect 97139 105718 97459 105760
rect 97139 105482 97181 105718
rect 97417 105482 97459 105718
rect 97139 105440 97459 105482
rect 116862 100725 116922 142547
rect 137104 116918 137424 116960
rect 137104 116682 137146 116918
rect 137382 116682 137424 116918
rect 137104 116640 137424 116682
rect 132472 105718 132792 105760
rect 132472 105482 132514 105718
rect 132750 105482 132792 105718
rect 132472 105440 132792 105482
rect 116859 100724 116925 100725
rect 116859 100660 116860 100724
rect 116924 100660 116925 100724
rect 116859 100659 116925 100660
rect 101139 83318 101459 83360
rect 101139 83082 101181 83318
rect 101417 83082 101459 83318
rect 101139 83040 101459 83082
rect 126104 83318 126424 83360
rect 126104 83082 126146 83318
rect 126382 83082 126424 83318
rect 126104 83040 126424 83082
rect 103437 72118 103757 72160
rect 103437 71882 103479 72118
rect 103715 71882 103757 72118
rect 103437 71840 103757 71882
rect 101139 60918 101459 60960
rect 101139 60682 101181 60918
rect 101417 60682 101459 60918
rect 101139 60640 101459 60682
rect 126104 60918 126424 60960
rect 126104 60682 126146 60918
rect 126382 60682 126424 60918
rect 126104 60640 126424 60682
rect 122011 59924 122077 59925
rect 122011 59860 122012 59924
rect 122076 59860 122077 59924
rect 122011 59859 122077 59860
rect 122014 59602 122074 59859
rect 136734 56202 136794 58686
rect 82267 51628 82333 51629
rect 82267 51564 82268 51628
rect 82332 51564 82333 51628
rect 82267 51563 82333 51564
rect 83555 51628 83621 51629
rect 83555 51564 83556 51628
rect 83620 51564 83621 51628
rect 83555 51563 83621 51564
rect 66995 50268 67061 50269
rect 66995 50204 66996 50268
rect 67060 50204 67061 50268
rect 66995 50203 67061 50204
rect 5000 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 9000 38518
rect 5000 16118 9000 38282
rect 25139 38518 25459 38560
rect 25139 38282 25181 38518
rect 25417 38282 25459 38518
rect 25139 38240 25459 38282
rect 60472 38518 60792 38560
rect 60472 38282 60514 38518
rect 60750 38282 60792 38518
rect 60472 38240 60792 38282
rect 29437 27318 29757 27360
rect 29437 27082 29479 27318
rect 29715 27082 29757 27318
rect 29437 27040 29757 27082
rect 65104 27318 65424 27360
rect 65104 27082 65146 27318
rect 65382 27082 65424 27318
rect 65104 27040 65424 27082
rect 66998 19261 67058 50203
rect 129739 46732 129805 46733
rect 129739 46668 129740 46732
rect 129804 46668 129805 46732
rect 129739 46667 129805 46668
rect 67731 46596 67797 46597
rect 67731 46532 67732 46596
rect 67796 46532 67797 46596
rect 67731 46531 67797 46532
rect 67179 46460 67245 46461
rect 67179 46396 67180 46460
rect 67244 46396 67245 46460
rect 67179 46395 67245 46396
rect 67182 20757 67242 46395
rect 67363 46324 67429 46325
rect 67363 46260 67364 46324
rect 67428 46260 67429 46324
rect 67363 46259 67429 46260
rect 67366 21029 67426 46259
rect 67547 46188 67613 46189
rect 67547 46124 67548 46188
rect 67612 46124 67613 46188
rect 67547 46123 67613 46124
rect 67363 21028 67429 21029
rect 67363 20964 67364 21028
rect 67428 20964 67429 21028
rect 67363 20963 67429 20964
rect 67179 20756 67245 20757
rect 67179 20692 67180 20756
rect 67244 20692 67245 20756
rect 67179 20691 67245 20692
rect 66995 19260 67061 19261
rect 66995 19196 66996 19260
rect 67060 19196 67061 19260
rect 66995 19195 67061 19196
rect 67550 17901 67610 46123
rect 67734 20893 67794 46531
rect 67915 44692 67981 44693
rect 67915 44628 67916 44692
rect 67980 44628 67981 44692
rect 67915 44627 67981 44628
rect 83555 44692 83621 44693
rect 83555 44628 83556 44692
rect 83620 44628 83621 44692
rect 83555 44627 83621 44628
rect 67731 20892 67797 20893
rect 67731 20828 67732 20892
rect 67796 20828 67797 20892
rect 67731 20827 67797 20828
rect 67918 18037 67978 44627
rect 83558 22202 83618 44627
rect 97139 38518 97459 38560
rect 97139 38282 97181 38518
rect 97417 38282 97459 38518
rect 97139 38240 97459 38282
rect 101437 27318 101757 27360
rect 101437 27082 101479 27318
rect 101715 27082 101757 27318
rect 101437 27040 101757 27082
rect 88523 21916 88524 21966
rect 88588 21916 88589 21966
rect 88523 21915 88589 21916
rect 129742 21029 129802 46667
rect 131211 46324 131277 46325
rect 131211 46260 131212 46324
rect 131276 46260 131277 46324
rect 131211 46259 131277 46260
rect 131214 21029 131274 46259
rect 132472 38518 132792 38560
rect 132472 38282 132514 38518
rect 132750 38282 132792 38518
rect 132472 38240 132792 38282
rect 129739 21028 129805 21029
rect 129739 20964 129740 21028
rect 129804 20964 129805 21028
rect 129739 20963 129805 20964
rect 131211 21028 131277 21029
rect 131211 20964 131212 21028
rect 131276 20964 131277 21028
rect 131211 20963 131277 20964
rect 136734 20893 136794 55966
rect 138758 51493 138818 177227
rect 173139 172918 173459 172960
rect 173139 172682 173181 172918
rect 173417 172682 173459 172918
rect 173139 172640 173459 172682
rect 168379 172124 168445 172125
rect 168379 172060 168380 172124
rect 168444 172060 168445 172124
rect 168379 172059 168445 172060
rect 141464 161718 141784 161760
rect 141464 161482 141506 161718
rect 141742 161482 141784 161718
rect 141464 161440 141784 161482
rect 168382 153442 168442 172059
rect 175437 161718 175757 161760
rect 175437 161482 175479 161718
rect 175715 161482 175757 161718
rect 175437 161440 175757 161482
rect 186046 152541 186106 153206
rect 186043 152540 186109 152541
rect 186043 152476 186044 152540
rect 186108 152476 186109 152540
rect 186043 152475 186109 152476
rect 173139 150518 173459 150560
rect 173139 150282 173181 150518
rect 173417 150282 173459 150518
rect 173139 150240 173459 150282
rect 141464 139318 141784 139360
rect 141464 139082 141506 139318
rect 141742 139082 141784 139318
rect 141464 139040 141784 139082
rect 175437 139318 175757 139360
rect 175437 139082 175479 139318
rect 175715 139082 175757 139318
rect 175437 139040 175757 139082
rect 173437 116918 173757 116960
rect 173437 116682 173479 116918
rect 173715 116682 173757 116918
rect 173437 116640 173757 116682
rect 169139 105718 169459 105760
rect 169139 105482 169181 105718
rect 169417 105482 169459 105718
rect 169139 105440 169459 105482
rect 168379 90388 168445 90389
rect 168379 90324 168380 90388
rect 168444 90324 168445 90388
rect 168379 90323 168445 90324
rect 141464 72118 141784 72160
rect 141464 71882 141506 72118
rect 141742 71882 141784 72118
rect 141464 71840 141784 71882
rect 168382 70482 168442 90323
rect 173139 83318 173459 83360
rect 173139 83082 173181 83318
rect 173417 83082 173459 83318
rect 173139 83040 173459 83082
rect 175437 72118 175757 72160
rect 175437 71882 175479 72118
rect 175715 71882 175757 72118
rect 175437 71840 175757 71882
rect 173139 60918 173459 60960
rect 173139 60682 173181 60918
rect 173417 60682 173459 60918
rect 173139 60640 173459 60682
rect 161755 57476 161821 57477
rect 161755 57412 161756 57476
rect 161820 57412 161821 57476
rect 161755 57411 161821 57412
rect 170219 57476 170285 57477
rect 170219 57412 170220 57476
rect 170284 57474 170285 57476
rect 170284 57414 171054 57474
rect 170284 57412 170285 57414
rect 170219 57411 170285 57412
rect 161758 56882 161818 57411
rect 185859 57276 185860 57326
rect 185924 57276 185925 57326
rect 185859 57275 185925 57276
rect 138755 51492 138821 51493
rect 138755 51428 138756 51492
rect 138820 51428 138821 51492
rect 138755 51427 138821 51428
rect 138939 46596 139005 46597
rect 138939 46532 138940 46596
rect 139004 46532 139005 46596
rect 138939 46531 139005 46532
rect 138755 46460 138821 46461
rect 138755 46396 138756 46460
rect 138820 46396 138821 46460
rect 138755 46395 138821 46396
rect 137104 27318 137424 27360
rect 137104 27082 137146 27318
rect 137382 27082 137424 27318
rect 137104 27040 137424 27082
rect 136731 20892 136797 20893
rect 136731 20828 136732 20892
rect 136796 20828 136797 20892
rect 136731 20827 136797 20828
rect 138758 18173 138818 46395
rect 138755 18172 138821 18173
rect 138755 18108 138756 18172
rect 138820 18108 138821 18172
rect 138755 18107 138821 18108
rect 67915 18036 67981 18037
rect 67915 17972 67916 18036
rect 67980 17972 67981 18036
rect 67915 17971 67981 17972
rect 138942 17901 139002 46531
rect 139675 44692 139741 44693
rect 139675 44628 139676 44692
rect 139740 44628 139741 44692
rect 139675 44627 139741 44628
rect 140963 44692 141029 44693
rect 140963 44628 140964 44692
rect 141028 44628 141029 44692
rect 140963 44627 141029 44628
rect 139678 18309 139738 44627
rect 139675 18308 139741 18309
rect 139675 18244 139676 18308
rect 139740 18244 139741 18308
rect 139675 18243 139741 18244
rect 140966 18037 141026 44627
rect 187150 43741 187210 213131
rect 190643 210748 190709 210749
rect 190643 210684 190644 210748
rect 190708 210684 190709 210748
rect 190643 210683 190709 210684
rect 190646 199594 190706 210683
rect 190646 199534 191626 199594
rect 191566 197421 191626 199534
rect 191563 197420 191629 197421
rect 191563 197356 191564 197420
rect 191628 197356 191629 197420
rect 191563 197355 191629 197356
rect 202704 195318 206704 217482
rect 202704 195082 202826 195318
rect 203062 195082 203146 195318
rect 203382 195082 203466 195318
rect 203702 195082 203786 195318
rect 204022 195082 204106 195318
rect 204342 195082 204426 195318
rect 204662 195082 204746 195318
rect 204982 195082 205066 195318
rect 205302 195082 205386 195318
rect 205622 195082 205706 195318
rect 205942 195082 206026 195318
rect 206262 195082 206346 195318
rect 206582 195082 206704 195318
rect 202704 172918 206704 195082
rect 202704 172682 202826 172918
rect 203062 172682 203146 172918
rect 203382 172682 203466 172918
rect 203702 172682 203786 172918
rect 204022 172682 204106 172918
rect 204342 172682 204426 172918
rect 204662 172682 204746 172918
rect 204982 172682 205066 172918
rect 205302 172682 205386 172918
rect 205622 172682 205706 172918
rect 205942 172682 206026 172918
rect 206262 172682 206346 172918
rect 206582 172682 206704 172918
rect 191195 159204 191261 159205
rect 191195 159140 191196 159204
rect 191260 159140 191261 159204
rect 191195 159139 191261 159140
rect 190643 145876 190709 145877
rect 190643 145812 190644 145876
rect 190708 145812 190709 145876
rect 190643 145811 190709 145812
rect 190646 118674 190706 145811
rect 191198 119354 191258 159139
rect 202704 150518 206704 172682
rect 202704 150282 202826 150518
rect 203062 150282 203146 150518
rect 203382 150282 203466 150518
rect 203702 150282 203786 150518
rect 204022 150282 204106 150518
rect 204342 150282 204426 150518
rect 204662 150282 204746 150518
rect 204982 150282 205066 150518
rect 205302 150282 205386 150518
rect 205622 150282 205706 150518
rect 205942 150282 206026 150518
rect 206262 150282 206346 150518
rect 206582 150282 206704 150518
rect 202704 128118 206704 150282
rect 202704 127882 202826 128118
rect 203062 127882 203146 128118
rect 203382 127882 203466 128118
rect 203702 127882 203786 128118
rect 204022 127882 204106 128118
rect 204342 127882 204426 128118
rect 204662 127882 204746 128118
rect 204982 127882 205066 128118
rect 205302 127882 205386 128118
rect 205622 127882 205706 128118
rect 205942 127882 206026 128118
rect 206262 127882 206346 128118
rect 206582 127882 206704 128118
rect 191198 119294 191810 119354
rect 190646 118614 191626 118674
rect 191566 115005 191626 118614
rect 191563 115004 191629 115005
rect 191563 114940 191564 115004
rect 191628 114940 191629 115004
rect 191563 114939 191629 114940
rect 191750 114597 191810 119294
rect 191747 114596 191813 114597
rect 191747 114532 191748 114596
rect 191812 114532 191813 114596
rect 191747 114531 191813 114532
rect 202704 105718 206704 127882
rect 202704 105482 202826 105718
rect 203062 105482 203146 105718
rect 203382 105482 203466 105718
rect 203702 105482 203786 105718
rect 204022 105482 204106 105718
rect 204342 105482 204426 105718
rect 204662 105482 204746 105718
rect 204982 105482 205066 105718
rect 205302 105482 205386 105718
rect 205622 105482 205706 105718
rect 205942 105482 206026 105718
rect 206262 105482 206346 105718
rect 206582 105482 206704 105718
rect 202704 83318 206704 105482
rect 202704 83082 202826 83318
rect 203062 83082 203146 83318
rect 203382 83082 203466 83318
rect 203702 83082 203786 83318
rect 204022 83082 204106 83318
rect 204342 83082 204426 83318
rect 204662 83082 204746 83318
rect 204982 83082 205066 83318
rect 205302 83082 205386 83318
rect 205622 83082 205706 83318
rect 205942 83082 206026 83318
rect 206262 83082 206346 83318
rect 206582 83082 206704 83318
rect 187883 63868 187949 63869
rect 187883 63804 187884 63868
rect 187948 63804 187949 63868
rect 187883 63803 187949 63804
rect 187147 43740 187213 43741
rect 187147 43676 187148 43740
rect 187212 43676 187213 43740
rect 187147 43675 187213 43676
rect 169139 38518 169459 38560
rect 169139 38282 169181 38518
rect 169417 38282 169459 38518
rect 169139 38240 169459 38282
rect 173437 27318 173757 27360
rect 173437 27082 173479 27318
rect 173715 27082 173757 27318
rect 173437 27040 173757 27082
rect 140963 18036 141029 18037
rect 140963 17972 140964 18036
rect 141028 17972 141029 18036
rect 140963 17971 141029 17972
rect 67547 17900 67613 17901
rect 67547 17836 67548 17900
rect 67612 17836 67613 17900
rect 67547 17835 67613 17836
rect 138939 17900 139005 17901
rect 138939 17836 138940 17900
rect 139004 17836 139005 17900
rect 138939 17835 139005 17836
rect 187886 17085 187946 63803
rect 202704 60918 206704 83082
rect 202704 60682 202826 60918
rect 203062 60682 203146 60918
rect 203382 60682 203466 60918
rect 203702 60682 203786 60918
rect 204022 60682 204106 60918
rect 204342 60682 204426 60918
rect 204662 60682 204746 60918
rect 204982 60682 205066 60918
rect 205302 60682 205386 60918
rect 205622 60682 205706 60918
rect 205942 60682 206026 60918
rect 206262 60682 206346 60918
rect 206582 60682 206704 60918
rect 202704 38518 206704 60682
rect 202704 38282 202826 38518
rect 203062 38282 203146 38518
rect 203382 38282 203466 38518
rect 203702 38282 203786 38518
rect 204022 38282 204106 38518
rect 204342 38282 204426 38518
rect 204662 38282 204746 38518
rect 204982 38282 205066 38518
rect 205302 38282 205386 38518
rect 205622 38282 205706 38518
rect 205942 38282 206026 38518
rect 206262 38282 206346 38518
rect 206582 38282 206704 38518
rect 187883 17084 187949 17085
rect 187883 17020 187884 17084
rect 187948 17020 187949 17084
rect 187883 17019 187949 17020
rect 5000 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 9000 16118
rect 5000 8878 9000 15882
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 202704 16118 206704 38282
rect 202704 15882 202826 16118
rect 203062 15882 203146 16118
rect 203382 15882 203466 16118
rect 203702 15882 203786 16118
rect 204022 15882 204106 16118
rect 204342 15882 204426 16118
rect 204662 15882 204746 16118
rect 204982 15882 205066 16118
rect 205302 15882 205386 16118
rect 205622 15882 205706 16118
rect 205942 15882 206026 16118
rect 206262 15882 206346 16118
rect 206582 15882 206704 16118
rect 202704 8878 206704 15882
rect 202704 8642 202826 8878
rect 203062 8642 203146 8878
rect 203382 8642 203466 8878
rect 203702 8642 203786 8878
rect 204022 8642 204106 8878
rect 204342 8642 204426 8878
rect 204662 8642 204746 8878
rect 204982 8642 205066 8878
rect 205302 8642 205386 8878
rect 205622 8642 205706 8878
rect 205942 8642 206026 8878
rect 206262 8642 206346 8878
rect 206582 8642 206704 8878
rect 202704 8558 206704 8642
rect 202704 8322 202826 8558
rect 203062 8322 203146 8558
rect 203382 8322 203466 8558
rect 203702 8322 203786 8558
rect 204022 8322 204106 8558
rect 204342 8322 204426 8558
rect 204662 8322 204746 8558
rect 204982 8322 205066 8558
rect 205302 8322 205386 8558
rect 205622 8322 205706 8558
rect 205942 8322 206026 8558
rect 206262 8322 206346 8558
rect 206582 8322 206704 8558
rect 202704 8238 206704 8322
rect 202704 8002 202826 8238
rect 203062 8002 203146 8238
rect 203382 8002 203466 8238
rect 203702 8002 203786 8238
rect 204022 8002 204106 8238
rect 204342 8002 204426 8238
rect 204662 8002 204746 8238
rect 204982 8002 205066 8238
rect 205302 8002 205386 8238
rect 205622 8002 205706 8238
rect 205942 8002 206026 8238
rect 206262 8002 206346 8238
rect 206582 8002 206704 8238
rect 202704 7918 206704 8002
rect 202704 7682 202826 7918
rect 203062 7682 203146 7918
rect 203382 7682 203466 7918
rect 203702 7682 203786 7918
rect 204022 7682 204106 7918
rect 204342 7682 204426 7918
rect 204662 7682 204746 7918
rect 204982 7682 205066 7918
rect 205302 7682 205386 7918
rect 205622 7682 205706 7918
rect 205942 7682 206026 7918
rect 206262 7682 206346 7918
rect 206582 7682 206704 7918
rect 202704 7598 206704 7682
rect 202704 7362 202826 7598
rect 203062 7362 203146 7598
rect 203382 7362 203466 7598
rect 203702 7362 203786 7598
rect 204022 7362 204106 7598
rect 204342 7362 204426 7598
rect 204662 7362 204746 7598
rect 204982 7362 205066 7598
rect 205302 7362 205386 7598
rect 205622 7362 205706 7598
rect 205942 7362 206026 7598
rect 206262 7362 206346 7598
rect 206582 7362 206704 7598
rect 202704 7278 206704 7362
rect 202704 7042 202826 7278
rect 203062 7042 203146 7278
rect 203382 7042 203466 7278
rect 203702 7042 203786 7278
rect 204022 7042 204106 7278
rect 204342 7042 204426 7278
rect 204662 7042 204746 7278
rect 204982 7042 205066 7278
rect 205302 7042 205386 7278
rect 205622 7042 205706 7278
rect 205942 7042 206026 7278
rect 206262 7042 206346 7278
rect 206582 7042 206704 7278
rect 202704 6958 206704 7042
rect 202704 6722 202826 6958
rect 203062 6722 203146 6958
rect 203382 6722 203466 6958
rect 203702 6722 203786 6958
rect 204022 6722 204106 6958
rect 204342 6722 204426 6958
rect 204662 6722 204746 6958
rect 204982 6722 205066 6958
rect 205302 6722 205386 6958
rect 205622 6722 205706 6958
rect 205942 6722 206026 6958
rect 206262 6722 206346 6958
rect 206582 6722 206704 6958
rect 202704 6638 206704 6722
rect 202704 6402 202826 6638
rect 203062 6402 203146 6638
rect 203382 6402 203466 6638
rect 203702 6402 203786 6638
rect 204022 6402 204106 6638
rect 204342 6402 204426 6638
rect 204662 6402 204746 6638
rect 204982 6402 205066 6638
rect 205302 6402 205386 6638
rect 205622 6402 205706 6638
rect 205942 6402 206026 6638
rect 206262 6402 206346 6638
rect 206582 6402 206704 6638
rect 202704 6318 206704 6402
rect 202704 6082 202826 6318
rect 203062 6082 203146 6318
rect 203382 6082 203466 6318
rect 203702 6082 203786 6318
rect 204022 6082 204106 6318
rect 204342 6082 204426 6318
rect 204662 6082 204746 6318
rect 204982 6082 205066 6318
rect 205302 6082 205386 6318
rect 205622 6082 205706 6318
rect 205942 6082 206026 6318
rect 206262 6082 206346 6318
rect 206582 6082 206704 6318
rect 202704 5998 206704 6082
rect 202704 5762 202826 5998
rect 203062 5762 203146 5998
rect 203382 5762 203466 5998
rect 203702 5762 203786 5998
rect 204022 5762 204106 5998
rect 204342 5762 204426 5998
rect 204662 5762 204746 5998
rect 204982 5762 205066 5998
rect 205302 5762 205386 5998
rect 205622 5762 205706 5998
rect 205942 5762 206026 5998
rect 206262 5762 206346 5998
rect 206582 5762 206704 5998
rect 202704 5678 206704 5762
rect 202704 5442 202826 5678
rect 203062 5442 203146 5678
rect 203382 5442 203466 5678
rect 203702 5442 203786 5678
rect 204022 5442 204106 5678
rect 204342 5442 204426 5678
rect 204662 5442 204746 5678
rect 204982 5442 205066 5678
rect 205302 5442 205386 5678
rect 205622 5442 205706 5678
rect 205942 5442 206026 5678
rect 206262 5442 206346 5678
rect 206582 5442 206704 5678
rect 202704 5358 206704 5442
rect 202704 5122 202826 5358
rect 203062 5122 203146 5358
rect 203382 5122 203466 5358
rect 203702 5122 203786 5358
rect 204022 5122 204106 5358
rect 204342 5122 204426 5358
rect 204662 5122 204746 5358
rect 204982 5122 205066 5358
rect 205302 5122 205386 5358
rect 205622 5122 205706 5358
rect 205942 5122 206026 5358
rect 206262 5122 206346 5358
rect 206582 5122 206704 5358
rect 202704 5000 206704 5122
rect 207704 206518 211704 225386
rect 207704 206282 207826 206518
rect 208062 206282 208146 206518
rect 208382 206282 208466 206518
rect 208702 206282 208786 206518
rect 209022 206282 209106 206518
rect 209342 206282 209426 206518
rect 209662 206282 209746 206518
rect 209982 206282 210066 206518
rect 210302 206282 210386 206518
rect 210622 206282 210706 206518
rect 210942 206282 211026 206518
rect 211262 206282 211346 206518
rect 211582 206282 211704 206518
rect 207704 184118 211704 206282
rect 207704 183882 207826 184118
rect 208062 183882 208146 184118
rect 208382 183882 208466 184118
rect 208702 183882 208786 184118
rect 209022 183882 209106 184118
rect 209342 183882 209426 184118
rect 209662 183882 209746 184118
rect 209982 183882 210066 184118
rect 210302 183882 210386 184118
rect 210622 183882 210706 184118
rect 210942 183882 211026 184118
rect 211262 183882 211346 184118
rect 211582 183882 211704 184118
rect 207704 161718 211704 183882
rect 207704 161482 207826 161718
rect 208062 161482 208146 161718
rect 208382 161482 208466 161718
rect 208702 161482 208786 161718
rect 209022 161482 209106 161718
rect 209342 161482 209426 161718
rect 209662 161482 209746 161718
rect 209982 161482 210066 161718
rect 210302 161482 210386 161718
rect 210622 161482 210706 161718
rect 210942 161482 211026 161718
rect 211262 161482 211346 161718
rect 211582 161482 211704 161718
rect 207704 139318 211704 161482
rect 207704 139082 207826 139318
rect 208062 139082 208146 139318
rect 208382 139082 208466 139318
rect 208702 139082 208786 139318
rect 209022 139082 209106 139318
rect 209342 139082 209426 139318
rect 209662 139082 209746 139318
rect 209982 139082 210066 139318
rect 210302 139082 210386 139318
rect 210622 139082 210706 139318
rect 210942 139082 211026 139318
rect 211262 139082 211346 139318
rect 211582 139082 211704 139318
rect 207704 116918 211704 139082
rect 207704 116682 207826 116918
rect 208062 116682 208146 116918
rect 208382 116682 208466 116918
rect 208702 116682 208786 116918
rect 209022 116682 209106 116918
rect 209342 116682 209426 116918
rect 209662 116682 209746 116918
rect 209982 116682 210066 116918
rect 210302 116682 210386 116918
rect 210622 116682 210706 116918
rect 210942 116682 211026 116918
rect 211262 116682 211346 116918
rect 211582 116682 211704 116918
rect 207704 94518 211704 116682
rect 207704 94282 207826 94518
rect 208062 94282 208146 94518
rect 208382 94282 208466 94518
rect 208702 94282 208786 94518
rect 209022 94282 209106 94518
rect 209342 94282 209426 94518
rect 209662 94282 209746 94518
rect 209982 94282 210066 94518
rect 210302 94282 210386 94518
rect 210622 94282 210706 94518
rect 210942 94282 211026 94518
rect 211262 94282 211346 94518
rect 211582 94282 211704 94518
rect 207704 72118 211704 94282
rect 207704 71882 207826 72118
rect 208062 71882 208146 72118
rect 208382 71882 208466 72118
rect 208702 71882 208786 72118
rect 209022 71882 209106 72118
rect 209342 71882 209426 72118
rect 209662 71882 209746 72118
rect 209982 71882 210066 72118
rect 210302 71882 210386 72118
rect 210622 71882 210706 72118
rect 210942 71882 211026 72118
rect 211262 71882 211346 72118
rect 211582 71882 211704 72118
rect 207704 49718 211704 71882
rect 207704 49482 207826 49718
rect 208062 49482 208146 49718
rect 208382 49482 208466 49718
rect 208702 49482 208786 49718
rect 209022 49482 209106 49718
rect 209342 49482 209426 49718
rect 209662 49482 209746 49718
rect 209982 49482 210066 49718
rect 210302 49482 210386 49718
rect 210622 49482 210706 49718
rect 210942 49482 211026 49718
rect 211262 49482 211346 49718
rect 211582 49482 211704 49718
rect 207704 27318 211704 49482
rect 207704 27082 207826 27318
rect 208062 27082 208146 27318
rect 208382 27082 208466 27318
rect 208702 27082 208786 27318
rect 209022 27082 209106 27318
rect 209342 27082 209426 27318
rect 209662 27082 209746 27318
rect 209982 27082 210066 27318
rect 210302 27082 210386 27318
rect 210622 27082 210706 27318
rect 210942 27082 211026 27318
rect 211262 27082 211346 27318
rect 211582 27082 211704 27318
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 207704 3878 211704 27082
rect 207704 3642 207826 3878
rect 208062 3642 208146 3878
rect 208382 3642 208466 3878
rect 208702 3642 208786 3878
rect 209022 3642 209106 3878
rect 209342 3642 209426 3878
rect 209662 3642 209746 3878
rect 209982 3642 210066 3878
rect 210302 3642 210386 3878
rect 210622 3642 210706 3878
rect 210942 3642 211026 3878
rect 211262 3642 211346 3878
rect 211582 3642 211704 3878
rect 207704 3558 211704 3642
rect 207704 3322 207826 3558
rect 208062 3322 208146 3558
rect 208382 3322 208466 3558
rect 208702 3322 208786 3558
rect 209022 3322 209106 3558
rect 209342 3322 209426 3558
rect 209662 3322 209746 3558
rect 209982 3322 210066 3558
rect 210302 3322 210386 3558
rect 210622 3322 210706 3558
rect 210942 3322 211026 3558
rect 211262 3322 211346 3558
rect 211582 3322 211704 3558
rect 207704 3238 211704 3322
rect 207704 3002 207826 3238
rect 208062 3002 208146 3238
rect 208382 3002 208466 3238
rect 208702 3002 208786 3238
rect 209022 3002 209106 3238
rect 209342 3002 209426 3238
rect 209662 3002 209746 3238
rect 209982 3002 210066 3238
rect 210302 3002 210386 3238
rect 210622 3002 210706 3238
rect 210942 3002 211026 3238
rect 211262 3002 211346 3238
rect 211582 3002 211704 3238
rect 207704 2918 211704 3002
rect 207704 2682 207826 2918
rect 208062 2682 208146 2918
rect 208382 2682 208466 2918
rect 208702 2682 208786 2918
rect 209022 2682 209106 2918
rect 209342 2682 209426 2918
rect 209662 2682 209746 2918
rect 209982 2682 210066 2918
rect 210302 2682 210386 2918
rect 210622 2682 210706 2918
rect 210942 2682 211026 2918
rect 211262 2682 211346 2918
rect 211582 2682 211704 2918
rect 207704 2598 211704 2682
rect 207704 2362 207826 2598
rect 208062 2362 208146 2598
rect 208382 2362 208466 2598
rect 208702 2362 208786 2598
rect 209022 2362 209106 2598
rect 209342 2362 209426 2598
rect 209662 2362 209746 2598
rect 209982 2362 210066 2598
rect 210302 2362 210386 2598
rect 210622 2362 210706 2598
rect 210942 2362 211026 2598
rect 211262 2362 211346 2598
rect 211582 2362 211704 2598
rect 207704 2278 211704 2362
rect 207704 2042 207826 2278
rect 208062 2042 208146 2278
rect 208382 2042 208466 2278
rect 208702 2042 208786 2278
rect 209022 2042 209106 2278
rect 209342 2042 209426 2278
rect 209662 2042 209746 2278
rect 209982 2042 210066 2278
rect 210302 2042 210386 2278
rect 210622 2042 210706 2278
rect 210942 2042 211026 2278
rect 211262 2042 211346 2278
rect 211582 2042 211704 2278
rect 207704 1958 211704 2042
rect 207704 1722 207826 1958
rect 208062 1722 208146 1958
rect 208382 1722 208466 1958
rect 208702 1722 208786 1958
rect 209022 1722 209106 1958
rect 209342 1722 209426 1958
rect 209662 1722 209746 1958
rect 209982 1722 210066 1958
rect 210302 1722 210386 1958
rect 210622 1722 210706 1958
rect 210942 1722 211026 1958
rect 211262 1722 211346 1958
rect 211582 1722 211704 1958
rect 207704 1638 211704 1722
rect 207704 1402 207826 1638
rect 208062 1402 208146 1638
rect 208382 1402 208466 1638
rect 208702 1402 208786 1638
rect 209022 1402 209106 1638
rect 209342 1402 209426 1638
rect 209662 1402 209746 1638
rect 209982 1402 210066 1638
rect 210302 1402 210386 1638
rect 210622 1402 210706 1638
rect 210942 1402 211026 1638
rect 211262 1402 211346 1638
rect 211582 1402 211704 1638
rect 207704 1318 211704 1402
rect 207704 1082 207826 1318
rect 208062 1082 208146 1318
rect 208382 1082 208466 1318
rect 208702 1082 208786 1318
rect 209022 1082 209106 1318
rect 209342 1082 209426 1318
rect 209662 1082 209746 1318
rect 209982 1082 210066 1318
rect 210302 1082 210386 1318
rect 210622 1082 210706 1318
rect 210942 1082 211026 1318
rect 211262 1082 211346 1318
rect 211582 1082 211704 1318
rect 207704 998 211704 1082
rect 207704 762 207826 998
rect 208062 762 208146 998
rect 208382 762 208466 998
rect 208702 762 208786 998
rect 209022 762 209106 998
rect 209342 762 209426 998
rect 209662 762 209746 998
rect 209982 762 210066 998
rect 210302 762 210386 998
rect 210622 762 210706 998
rect 210942 762 211026 998
rect 211262 762 211346 998
rect 211582 762 211704 998
rect 207704 678 211704 762
rect 207704 442 207826 678
rect 208062 442 208146 678
rect 208382 442 208466 678
rect 208702 442 208786 678
rect 209022 442 209106 678
rect 209342 442 209426 678
rect 209662 442 209746 678
rect 209982 442 210066 678
rect 210302 442 210386 678
rect 210622 442 210706 678
rect 210942 442 211026 678
rect 211262 442 211346 678
rect 211582 442 211704 678
rect 207704 358 211704 442
rect 207704 122 207826 358
rect 208062 122 208146 358
rect 208382 122 208466 358
rect 208702 122 208786 358
rect 209022 122 209106 358
rect 209342 122 209426 358
rect 209662 122 209746 358
rect 209982 122 210066 358
rect 210302 122 210386 358
rect 210622 122 210706 358
rect 210942 122 211026 358
rect 211262 122 211346 358
rect 211582 122 211704 358
rect 207704 0 211704 122
<< via4 >>
rect 122 228906 358 229142
rect 442 228906 678 229142
rect 762 228906 998 229142
rect 1082 228906 1318 229142
rect 1402 228906 1638 229142
rect 1722 228906 1958 229142
rect 2042 228906 2278 229142
rect 2362 228906 2598 229142
rect 2682 228906 2918 229142
rect 3002 228906 3238 229142
rect 3322 228906 3558 229142
rect 3642 228906 3878 229142
rect 122 228586 358 228822
rect 442 228586 678 228822
rect 762 228586 998 228822
rect 1082 228586 1318 228822
rect 1402 228586 1638 228822
rect 1722 228586 1958 228822
rect 2042 228586 2278 228822
rect 2362 228586 2598 228822
rect 2682 228586 2918 228822
rect 3002 228586 3238 228822
rect 3322 228586 3558 228822
rect 3642 228586 3878 228822
rect 122 228266 358 228502
rect 442 228266 678 228502
rect 762 228266 998 228502
rect 1082 228266 1318 228502
rect 1402 228266 1638 228502
rect 1722 228266 1958 228502
rect 2042 228266 2278 228502
rect 2362 228266 2598 228502
rect 2682 228266 2918 228502
rect 3002 228266 3238 228502
rect 3322 228266 3558 228502
rect 3642 228266 3878 228502
rect 122 227946 358 228182
rect 442 227946 678 228182
rect 762 227946 998 228182
rect 1082 227946 1318 228182
rect 1402 227946 1638 228182
rect 1722 227946 1958 228182
rect 2042 227946 2278 228182
rect 2362 227946 2598 228182
rect 2682 227946 2918 228182
rect 3002 227946 3238 228182
rect 3322 227946 3558 228182
rect 3642 227946 3878 228182
rect 122 227626 358 227862
rect 442 227626 678 227862
rect 762 227626 998 227862
rect 1082 227626 1318 227862
rect 1402 227626 1638 227862
rect 1722 227626 1958 227862
rect 2042 227626 2278 227862
rect 2362 227626 2598 227862
rect 2682 227626 2918 227862
rect 3002 227626 3238 227862
rect 3322 227626 3558 227862
rect 3642 227626 3878 227862
rect 122 227306 358 227542
rect 442 227306 678 227542
rect 762 227306 998 227542
rect 1082 227306 1318 227542
rect 1402 227306 1638 227542
rect 1722 227306 1958 227542
rect 2042 227306 2278 227542
rect 2362 227306 2598 227542
rect 2682 227306 2918 227542
rect 3002 227306 3238 227542
rect 3322 227306 3558 227542
rect 3642 227306 3878 227542
rect 122 226986 358 227222
rect 442 226986 678 227222
rect 762 226986 998 227222
rect 1082 226986 1318 227222
rect 1402 226986 1638 227222
rect 1722 226986 1958 227222
rect 2042 226986 2278 227222
rect 2362 226986 2598 227222
rect 2682 226986 2918 227222
rect 3002 226986 3238 227222
rect 3322 226986 3558 227222
rect 3642 226986 3878 227222
rect 122 226666 358 226902
rect 442 226666 678 226902
rect 762 226666 998 226902
rect 1082 226666 1318 226902
rect 1402 226666 1638 226902
rect 1722 226666 1958 226902
rect 2042 226666 2278 226902
rect 2362 226666 2598 226902
rect 2682 226666 2918 226902
rect 3002 226666 3238 226902
rect 3322 226666 3558 226902
rect 3642 226666 3878 226902
rect 122 226346 358 226582
rect 442 226346 678 226582
rect 762 226346 998 226582
rect 1082 226346 1318 226582
rect 1402 226346 1638 226582
rect 1722 226346 1958 226582
rect 2042 226346 2278 226582
rect 2362 226346 2598 226582
rect 2682 226346 2918 226582
rect 3002 226346 3238 226582
rect 3322 226346 3558 226582
rect 3642 226346 3878 226582
rect 122 226026 358 226262
rect 442 226026 678 226262
rect 762 226026 998 226262
rect 1082 226026 1318 226262
rect 1402 226026 1638 226262
rect 1722 226026 1958 226262
rect 2042 226026 2278 226262
rect 2362 226026 2598 226262
rect 2682 226026 2918 226262
rect 3002 226026 3238 226262
rect 3322 226026 3558 226262
rect 3642 226026 3878 226262
rect 122 225706 358 225942
rect 442 225706 678 225942
rect 762 225706 998 225942
rect 1082 225706 1318 225942
rect 1402 225706 1638 225942
rect 1722 225706 1958 225942
rect 2042 225706 2278 225942
rect 2362 225706 2598 225942
rect 2682 225706 2918 225942
rect 3002 225706 3238 225942
rect 3322 225706 3558 225942
rect 3642 225706 3878 225942
rect 122 225386 358 225622
rect 442 225386 678 225622
rect 762 225386 998 225622
rect 1082 225386 1318 225622
rect 1402 225386 1638 225622
rect 1722 225386 1958 225622
rect 2042 225386 2278 225622
rect 2362 225386 2598 225622
rect 2682 225386 2918 225622
rect 3002 225386 3238 225622
rect 3322 225386 3558 225622
rect 3642 225386 3878 225622
rect 207826 228906 208062 229142
rect 208146 228906 208382 229142
rect 208466 228906 208702 229142
rect 208786 228906 209022 229142
rect 209106 228906 209342 229142
rect 209426 228906 209662 229142
rect 209746 228906 209982 229142
rect 210066 228906 210302 229142
rect 210386 228906 210622 229142
rect 210706 228906 210942 229142
rect 211026 228906 211262 229142
rect 211346 228906 211582 229142
rect 207826 228586 208062 228822
rect 208146 228586 208382 228822
rect 208466 228586 208702 228822
rect 208786 228586 209022 228822
rect 209106 228586 209342 228822
rect 209426 228586 209662 228822
rect 209746 228586 209982 228822
rect 210066 228586 210302 228822
rect 210386 228586 210622 228822
rect 210706 228586 210942 228822
rect 211026 228586 211262 228822
rect 211346 228586 211582 228822
rect 207826 228266 208062 228502
rect 208146 228266 208382 228502
rect 208466 228266 208702 228502
rect 208786 228266 209022 228502
rect 209106 228266 209342 228502
rect 209426 228266 209662 228502
rect 209746 228266 209982 228502
rect 210066 228266 210302 228502
rect 210386 228266 210622 228502
rect 210706 228266 210942 228502
rect 211026 228266 211262 228502
rect 211346 228266 211582 228502
rect 207826 227946 208062 228182
rect 208146 227946 208382 228182
rect 208466 227946 208702 228182
rect 208786 227946 209022 228182
rect 209106 227946 209342 228182
rect 209426 227946 209662 228182
rect 209746 227946 209982 228182
rect 210066 227946 210302 228182
rect 210386 227946 210622 228182
rect 210706 227946 210942 228182
rect 211026 227946 211262 228182
rect 211346 227946 211582 228182
rect 207826 227626 208062 227862
rect 208146 227626 208382 227862
rect 208466 227626 208702 227862
rect 208786 227626 209022 227862
rect 209106 227626 209342 227862
rect 209426 227626 209662 227862
rect 209746 227626 209982 227862
rect 210066 227626 210302 227862
rect 210386 227626 210622 227862
rect 210706 227626 210942 227862
rect 211026 227626 211262 227862
rect 211346 227626 211582 227862
rect 207826 227306 208062 227542
rect 208146 227306 208382 227542
rect 208466 227306 208702 227542
rect 208786 227306 209022 227542
rect 209106 227306 209342 227542
rect 209426 227306 209662 227542
rect 209746 227306 209982 227542
rect 210066 227306 210302 227542
rect 210386 227306 210622 227542
rect 210706 227306 210942 227542
rect 211026 227306 211262 227542
rect 211346 227306 211582 227542
rect 207826 226986 208062 227222
rect 208146 226986 208382 227222
rect 208466 226986 208702 227222
rect 208786 226986 209022 227222
rect 209106 226986 209342 227222
rect 209426 226986 209662 227222
rect 209746 226986 209982 227222
rect 210066 226986 210302 227222
rect 210386 226986 210622 227222
rect 210706 226986 210942 227222
rect 211026 226986 211262 227222
rect 211346 226986 211582 227222
rect 207826 226666 208062 226902
rect 208146 226666 208382 226902
rect 208466 226666 208702 226902
rect 208786 226666 209022 226902
rect 209106 226666 209342 226902
rect 209426 226666 209662 226902
rect 209746 226666 209982 226902
rect 210066 226666 210302 226902
rect 210386 226666 210622 226902
rect 210706 226666 210942 226902
rect 211026 226666 211262 226902
rect 211346 226666 211582 226902
rect 207826 226346 208062 226582
rect 208146 226346 208382 226582
rect 208466 226346 208702 226582
rect 208786 226346 209022 226582
rect 209106 226346 209342 226582
rect 209426 226346 209662 226582
rect 209746 226346 209982 226582
rect 210066 226346 210302 226582
rect 210386 226346 210622 226582
rect 210706 226346 210942 226582
rect 211026 226346 211262 226582
rect 211346 226346 211582 226582
rect 207826 226026 208062 226262
rect 208146 226026 208382 226262
rect 208466 226026 208702 226262
rect 208786 226026 209022 226262
rect 209106 226026 209342 226262
rect 209426 226026 209662 226262
rect 209746 226026 209982 226262
rect 210066 226026 210302 226262
rect 210386 226026 210622 226262
rect 210706 226026 210942 226262
rect 211026 226026 211262 226262
rect 211346 226026 211582 226262
rect 207826 225706 208062 225942
rect 208146 225706 208382 225942
rect 208466 225706 208702 225942
rect 208786 225706 209022 225942
rect 209106 225706 209342 225942
rect 209426 225706 209662 225942
rect 209746 225706 209982 225942
rect 210066 225706 210302 225942
rect 210386 225706 210622 225942
rect 210706 225706 210942 225942
rect 211026 225706 211262 225942
rect 211346 225706 211582 225942
rect 207826 225386 208062 225622
rect 208146 225386 208382 225622
rect 208466 225386 208702 225622
rect 208786 225386 209022 225622
rect 209106 225386 209342 225622
rect 209426 225386 209662 225622
rect 209746 225386 209982 225622
rect 210066 225386 210302 225622
rect 210386 225386 210622 225622
rect 210706 225386 210942 225622
rect 211026 225386 211262 225622
rect 211346 225386 211582 225622
rect 122 206282 358 206518
rect 442 206282 678 206518
rect 762 206282 998 206518
rect 1082 206282 1318 206518
rect 1402 206282 1638 206518
rect 1722 206282 1958 206518
rect 2042 206282 2278 206518
rect 2362 206282 2598 206518
rect 2682 206282 2918 206518
rect 3002 206282 3238 206518
rect 3322 206282 3558 206518
rect 3642 206282 3878 206518
rect 122 183882 358 184118
rect 442 183882 678 184118
rect 762 183882 998 184118
rect 1082 183882 1318 184118
rect 1402 183882 1638 184118
rect 1722 183882 1958 184118
rect 2042 183882 2278 184118
rect 2362 183882 2598 184118
rect 2682 183882 2918 184118
rect 3002 183882 3238 184118
rect 3322 183882 3558 184118
rect 3642 183882 3878 184118
rect 122 161482 358 161718
rect 442 161482 678 161718
rect 762 161482 998 161718
rect 1082 161482 1318 161718
rect 1402 161482 1638 161718
rect 1722 161482 1958 161718
rect 2042 161482 2278 161718
rect 2362 161482 2598 161718
rect 2682 161482 2918 161718
rect 3002 161482 3238 161718
rect 3322 161482 3558 161718
rect 3642 161482 3878 161718
rect 122 139082 358 139318
rect 442 139082 678 139318
rect 762 139082 998 139318
rect 1082 139082 1318 139318
rect 1402 139082 1638 139318
rect 1722 139082 1958 139318
rect 2042 139082 2278 139318
rect 2362 139082 2598 139318
rect 2682 139082 2918 139318
rect 3002 139082 3238 139318
rect 3322 139082 3558 139318
rect 3642 139082 3878 139318
rect 122 116682 358 116918
rect 442 116682 678 116918
rect 762 116682 998 116918
rect 1082 116682 1318 116918
rect 1402 116682 1638 116918
rect 1722 116682 1958 116918
rect 2042 116682 2278 116918
rect 2362 116682 2598 116918
rect 2682 116682 2918 116918
rect 3002 116682 3238 116918
rect 3322 116682 3558 116918
rect 3642 116682 3878 116918
rect 122 94282 358 94518
rect 442 94282 678 94518
rect 762 94282 998 94518
rect 1082 94282 1318 94518
rect 1402 94282 1638 94518
rect 1722 94282 1958 94518
rect 2042 94282 2278 94518
rect 2362 94282 2598 94518
rect 2682 94282 2918 94518
rect 3002 94282 3238 94518
rect 3322 94282 3558 94518
rect 3642 94282 3878 94518
rect 122 71882 358 72118
rect 442 71882 678 72118
rect 762 71882 998 72118
rect 1082 71882 1318 72118
rect 1402 71882 1638 72118
rect 1722 71882 1958 72118
rect 2042 71882 2278 72118
rect 2362 71882 2598 72118
rect 2682 71882 2918 72118
rect 3002 71882 3238 72118
rect 3322 71882 3558 72118
rect 3642 71882 3878 72118
rect 122 49482 358 49718
rect 442 49482 678 49718
rect 762 49482 998 49718
rect 1082 49482 1318 49718
rect 1402 49482 1638 49718
rect 1722 49482 1958 49718
rect 2042 49482 2278 49718
rect 2362 49482 2598 49718
rect 2682 49482 2918 49718
rect 3002 49482 3238 49718
rect 3322 49482 3558 49718
rect 3642 49482 3878 49718
rect 122 27082 358 27318
rect 442 27082 678 27318
rect 762 27082 998 27318
rect 1082 27082 1318 27318
rect 1402 27082 1638 27318
rect 1722 27082 1958 27318
rect 2042 27082 2278 27318
rect 2362 27082 2598 27318
rect 2682 27082 2918 27318
rect 3002 27082 3238 27318
rect 3322 27082 3558 27318
rect 3642 27082 3878 27318
rect 5122 223906 5358 224142
rect 5442 223906 5678 224142
rect 5762 223906 5998 224142
rect 6082 223906 6318 224142
rect 6402 223906 6638 224142
rect 6722 223906 6958 224142
rect 7042 223906 7278 224142
rect 7362 223906 7598 224142
rect 7682 223906 7918 224142
rect 8002 223906 8238 224142
rect 8322 223906 8558 224142
rect 8642 223906 8878 224142
rect 5122 223586 5358 223822
rect 5442 223586 5678 223822
rect 5762 223586 5998 223822
rect 6082 223586 6318 223822
rect 6402 223586 6638 223822
rect 6722 223586 6958 223822
rect 7042 223586 7278 223822
rect 7362 223586 7598 223822
rect 7682 223586 7918 223822
rect 8002 223586 8238 223822
rect 8322 223586 8558 223822
rect 8642 223586 8878 223822
rect 5122 223266 5358 223502
rect 5442 223266 5678 223502
rect 5762 223266 5998 223502
rect 6082 223266 6318 223502
rect 6402 223266 6638 223502
rect 6722 223266 6958 223502
rect 7042 223266 7278 223502
rect 7362 223266 7598 223502
rect 7682 223266 7918 223502
rect 8002 223266 8238 223502
rect 8322 223266 8558 223502
rect 8642 223266 8878 223502
rect 5122 222946 5358 223182
rect 5442 222946 5678 223182
rect 5762 222946 5998 223182
rect 6082 222946 6318 223182
rect 6402 222946 6638 223182
rect 6722 222946 6958 223182
rect 7042 222946 7278 223182
rect 7362 222946 7598 223182
rect 7682 222946 7918 223182
rect 8002 222946 8238 223182
rect 8322 222946 8558 223182
rect 8642 222946 8878 223182
rect 5122 222626 5358 222862
rect 5442 222626 5678 222862
rect 5762 222626 5998 222862
rect 6082 222626 6318 222862
rect 6402 222626 6638 222862
rect 6722 222626 6958 222862
rect 7042 222626 7278 222862
rect 7362 222626 7598 222862
rect 7682 222626 7918 222862
rect 8002 222626 8238 222862
rect 8322 222626 8558 222862
rect 8642 222626 8878 222862
rect 5122 222306 5358 222542
rect 5442 222306 5678 222542
rect 5762 222306 5998 222542
rect 6082 222306 6318 222542
rect 6402 222306 6638 222542
rect 6722 222306 6958 222542
rect 7042 222306 7278 222542
rect 7362 222306 7598 222542
rect 7682 222306 7918 222542
rect 8002 222306 8238 222542
rect 8322 222306 8558 222542
rect 8642 222306 8878 222542
rect 5122 221986 5358 222222
rect 5442 221986 5678 222222
rect 5762 221986 5998 222222
rect 6082 221986 6318 222222
rect 6402 221986 6638 222222
rect 6722 221986 6958 222222
rect 7042 221986 7278 222222
rect 7362 221986 7598 222222
rect 7682 221986 7918 222222
rect 8002 221986 8238 222222
rect 8322 221986 8558 222222
rect 8642 221986 8878 222222
rect 5122 221666 5358 221902
rect 5442 221666 5678 221902
rect 5762 221666 5998 221902
rect 6082 221666 6318 221902
rect 6402 221666 6638 221902
rect 6722 221666 6958 221902
rect 7042 221666 7278 221902
rect 7362 221666 7598 221902
rect 7682 221666 7918 221902
rect 8002 221666 8238 221902
rect 8322 221666 8558 221902
rect 8642 221666 8878 221902
rect 5122 221346 5358 221582
rect 5442 221346 5678 221582
rect 5762 221346 5998 221582
rect 6082 221346 6318 221582
rect 6402 221346 6638 221582
rect 6722 221346 6958 221582
rect 7042 221346 7278 221582
rect 7362 221346 7598 221582
rect 7682 221346 7918 221582
rect 8002 221346 8238 221582
rect 8322 221346 8558 221582
rect 8642 221346 8878 221582
rect 5122 221026 5358 221262
rect 5442 221026 5678 221262
rect 5762 221026 5998 221262
rect 6082 221026 6318 221262
rect 6402 221026 6638 221262
rect 6722 221026 6958 221262
rect 7042 221026 7278 221262
rect 7362 221026 7598 221262
rect 7682 221026 7918 221262
rect 8002 221026 8238 221262
rect 8322 221026 8558 221262
rect 8642 221026 8878 221262
rect 5122 220706 5358 220942
rect 5442 220706 5678 220942
rect 5762 220706 5998 220942
rect 6082 220706 6318 220942
rect 6402 220706 6638 220942
rect 6722 220706 6958 220942
rect 7042 220706 7278 220942
rect 7362 220706 7598 220942
rect 7682 220706 7918 220942
rect 8002 220706 8238 220942
rect 8322 220706 8558 220942
rect 8642 220706 8878 220942
rect 5122 220386 5358 220622
rect 5442 220386 5678 220622
rect 5762 220386 5998 220622
rect 6082 220386 6318 220622
rect 6402 220386 6638 220622
rect 6722 220386 6958 220622
rect 7042 220386 7278 220622
rect 7362 220386 7598 220622
rect 7682 220386 7918 220622
rect 8002 220386 8238 220622
rect 8322 220386 8558 220622
rect 8642 220386 8878 220622
rect 5122 217482 5358 217718
rect 5442 217482 5678 217718
rect 5762 217482 5998 217718
rect 6082 217482 6318 217718
rect 6402 217482 6638 217718
rect 6722 217482 6958 217718
rect 7042 217482 7278 217718
rect 7362 217482 7598 217718
rect 7682 217482 7918 217718
rect 8002 217482 8238 217718
rect 8322 217482 8558 217718
rect 8642 217482 8878 217718
rect 202826 223906 203062 224142
rect 203146 223906 203382 224142
rect 203466 223906 203702 224142
rect 203786 223906 204022 224142
rect 204106 223906 204342 224142
rect 204426 223906 204662 224142
rect 204746 223906 204982 224142
rect 205066 223906 205302 224142
rect 205386 223906 205622 224142
rect 205706 223906 205942 224142
rect 206026 223906 206262 224142
rect 206346 223906 206582 224142
rect 202826 223586 203062 223822
rect 203146 223586 203382 223822
rect 203466 223586 203702 223822
rect 203786 223586 204022 223822
rect 204106 223586 204342 223822
rect 204426 223586 204662 223822
rect 204746 223586 204982 223822
rect 205066 223586 205302 223822
rect 205386 223586 205622 223822
rect 205706 223586 205942 223822
rect 206026 223586 206262 223822
rect 206346 223586 206582 223822
rect 202826 223266 203062 223502
rect 203146 223266 203382 223502
rect 203466 223266 203702 223502
rect 203786 223266 204022 223502
rect 204106 223266 204342 223502
rect 204426 223266 204662 223502
rect 204746 223266 204982 223502
rect 205066 223266 205302 223502
rect 205386 223266 205622 223502
rect 205706 223266 205942 223502
rect 206026 223266 206262 223502
rect 206346 223266 206582 223502
rect 202826 222946 203062 223182
rect 203146 222946 203382 223182
rect 203466 222946 203702 223182
rect 203786 222946 204022 223182
rect 204106 222946 204342 223182
rect 204426 222946 204662 223182
rect 204746 222946 204982 223182
rect 205066 222946 205302 223182
rect 205386 222946 205622 223182
rect 205706 222946 205942 223182
rect 206026 222946 206262 223182
rect 206346 222946 206582 223182
rect 202826 222626 203062 222862
rect 203146 222626 203382 222862
rect 203466 222626 203702 222862
rect 203786 222626 204022 222862
rect 204106 222626 204342 222862
rect 204426 222626 204662 222862
rect 204746 222626 204982 222862
rect 205066 222626 205302 222862
rect 205386 222626 205622 222862
rect 205706 222626 205942 222862
rect 206026 222626 206262 222862
rect 206346 222626 206582 222862
rect 202826 222306 203062 222542
rect 203146 222306 203382 222542
rect 203466 222306 203702 222542
rect 203786 222306 204022 222542
rect 204106 222306 204342 222542
rect 204426 222306 204662 222542
rect 204746 222306 204982 222542
rect 205066 222306 205302 222542
rect 205386 222306 205622 222542
rect 205706 222306 205942 222542
rect 206026 222306 206262 222542
rect 206346 222306 206582 222542
rect 202826 221986 203062 222222
rect 203146 221986 203382 222222
rect 203466 221986 203702 222222
rect 203786 221986 204022 222222
rect 204106 221986 204342 222222
rect 204426 221986 204662 222222
rect 204746 221986 204982 222222
rect 205066 221986 205302 222222
rect 205386 221986 205622 222222
rect 205706 221986 205942 222222
rect 206026 221986 206262 222222
rect 206346 221986 206582 222222
rect 202826 221666 203062 221902
rect 203146 221666 203382 221902
rect 203466 221666 203702 221902
rect 203786 221666 204022 221902
rect 204106 221666 204342 221902
rect 204426 221666 204662 221902
rect 204746 221666 204982 221902
rect 205066 221666 205302 221902
rect 205386 221666 205622 221902
rect 205706 221666 205942 221902
rect 206026 221666 206262 221902
rect 206346 221666 206582 221902
rect 202826 221346 203062 221582
rect 203146 221346 203382 221582
rect 203466 221346 203702 221582
rect 203786 221346 204022 221582
rect 204106 221346 204342 221582
rect 204426 221346 204662 221582
rect 204746 221346 204982 221582
rect 205066 221346 205302 221582
rect 205386 221346 205622 221582
rect 205706 221346 205942 221582
rect 206026 221346 206262 221582
rect 206346 221346 206582 221582
rect 202826 221026 203062 221262
rect 203146 221026 203382 221262
rect 203466 221026 203702 221262
rect 203786 221026 204022 221262
rect 204106 221026 204342 221262
rect 204426 221026 204662 221262
rect 204746 221026 204982 221262
rect 205066 221026 205302 221262
rect 205386 221026 205622 221262
rect 205706 221026 205942 221262
rect 206026 221026 206262 221262
rect 206346 221026 206582 221262
rect 202826 220706 203062 220942
rect 203146 220706 203382 220942
rect 203466 220706 203702 220942
rect 203786 220706 204022 220942
rect 204106 220706 204342 220942
rect 204426 220706 204662 220942
rect 204746 220706 204982 220942
rect 205066 220706 205302 220942
rect 205386 220706 205622 220942
rect 205706 220706 205942 220942
rect 206026 220706 206262 220942
rect 206346 220706 206582 220942
rect 202826 220386 203062 220622
rect 203146 220386 203382 220622
rect 203466 220386 203702 220622
rect 203786 220386 204022 220622
rect 204106 220386 204342 220622
rect 204426 220386 204662 220622
rect 204746 220386 204982 220622
rect 205066 220386 205302 220622
rect 205386 220386 205622 220622
rect 205706 220386 205942 220622
rect 206026 220386 206262 220622
rect 206346 220386 206582 220622
rect 202826 217482 203062 217718
rect 203146 217482 203382 217718
rect 203466 217482 203702 217718
rect 203786 217482 204022 217718
rect 204106 217482 204342 217718
rect 204426 217482 204662 217718
rect 204746 217482 204982 217718
rect 205066 217482 205302 217718
rect 205386 217482 205622 217718
rect 205706 217482 205942 217718
rect 206026 217482 206262 217718
rect 206346 217482 206582 217718
rect 5122 195082 5358 195318
rect 5442 195082 5678 195318
rect 5762 195082 5998 195318
rect 6082 195082 6318 195318
rect 6402 195082 6638 195318
rect 6722 195082 6958 195318
rect 7042 195082 7278 195318
rect 7362 195082 7598 195318
rect 7682 195082 7918 195318
rect 8002 195082 8238 195318
rect 8322 195082 8558 195318
rect 8642 195082 8878 195318
rect 5122 172682 5358 172918
rect 5442 172682 5678 172918
rect 5762 172682 5998 172918
rect 6082 172682 6318 172918
rect 6402 172682 6638 172918
rect 6722 172682 6958 172918
rect 7042 172682 7278 172918
rect 7362 172682 7598 172918
rect 7682 172682 7918 172918
rect 8002 172682 8238 172918
rect 8322 172682 8558 172918
rect 8642 172682 8878 172918
rect 29190 206282 29426 206518
rect 65146 206282 65382 206518
rect 24892 195082 25128 195318
rect 60514 195082 60750 195318
rect 101479 206282 101715 206518
rect 137146 206282 137382 206518
rect 97181 195082 97417 195318
rect 132514 195082 132750 195318
rect 173479 206282 173715 206518
rect 169181 195082 169417 195318
rect 29181 172682 29417 172918
rect 54146 172682 54382 172918
rect 31479 161482 31715 161718
rect 69506 161482 69742 161718
rect 5122 150282 5358 150518
rect 5442 150282 5678 150518
rect 5762 150282 5998 150518
rect 6082 150282 6318 150518
rect 6402 150282 6638 150518
rect 6722 150282 6958 150518
rect 7042 150282 7278 150518
rect 7362 150282 7598 150518
rect 7682 150282 7918 150518
rect 8002 150282 8238 150518
rect 8322 150282 8558 150518
rect 8642 150282 8878 150518
rect 29181 150282 29417 150518
rect 54146 150282 54382 150518
rect 26062 140436 26298 140522
rect 26062 140372 26148 140436
rect 26148 140372 26212 140436
rect 26212 140372 26298 140436
rect 26062 140286 26298 140372
rect 44278 140286 44514 140522
rect 31479 139082 31715 139318
rect 5122 127882 5358 128118
rect 5442 127882 5678 128118
rect 5762 127882 5998 128118
rect 6082 127882 6318 128118
rect 6402 127882 6638 128118
rect 6722 127882 6958 128118
rect 7042 127882 7278 128118
rect 7362 127882 7598 128118
rect 7682 127882 7918 128118
rect 8002 127882 8238 128118
rect 8322 127882 8558 128118
rect 8642 127882 8878 128118
rect 29479 116682 29715 116918
rect 101181 172682 101417 172918
rect 126146 172682 126382 172918
rect 103479 161482 103715 161718
rect 101181 150282 101417 150518
rect 126146 150282 126382 150518
rect 69506 139082 69742 139318
rect 103479 139082 103715 139318
rect 65146 116682 65382 116918
rect 19806 106286 20042 106522
rect 46302 106286 46538 106522
rect 5122 105482 5358 105718
rect 5442 105482 5678 105718
rect 5762 105482 5998 105718
rect 6082 105482 6318 105718
rect 6402 105482 6638 105718
rect 6722 105482 6958 105718
rect 7042 105482 7278 105718
rect 7362 105482 7598 105718
rect 7682 105482 7918 105718
rect 8002 105482 8238 105718
rect 8322 105482 8558 105718
rect 8642 105482 8878 105718
rect 25181 105482 25417 105718
rect 60514 105482 60750 105718
rect 5122 83082 5358 83318
rect 5442 83082 5678 83318
rect 5762 83082 5998 83318
rect 6082 83082 6318 83318
rect 6402 83082 6638 83318
rect 6722 83082 6958 83318
rect 7042 83082 7278 83318
rect 7362 83082 7598 83318
rect 7682 83082 7918 83318
rect 8002 83082 8238 83318
rect 8322 83082 8558 83318
rect 8642 83082 8878 83318
rect 29181 83082 29417 83318
rect 48326 92006 48562 92242
rect 54146 83082 54382 83318
rect 31479 71882 31715 72118
rect 5122 60682 5358 60918
rect 5442 60682 5678 60918
rect 5762 60682 5998 60918
rect 6082 60682 6318 60918
rect 6402 60682 6638 60918
rect 6722 60682 6958 60918
rect 7042 60682 7278 60918
rect 7362 60682 7598 60918
rect 7682 60682 7918 60918
rect 8002 60682 8238 60918
rect 8322 60682 8558 60918
rect 8642 60682 8878 60918
rect 29181 60682 29417 60918
rect 69506 71882 69742 72118
rect 54146 60682 54382 60918
rect 26062 58156 26298 58242
rect 26062 58092 26148 58156
rect 26148 58092 26212 58156
rect 26212 58092 26298 58156
rect 26062 58006 26298 58092
rect 44278 58006 44514 58242
rect 101479 116682 101715 116918
rect 97181 105482 97417 105718
rect 137146 116682 137382 116918
rect 132514 105482 132750 105718
rect 85126 92006 85362 92242
rect 101181 83082 101417 83318
rect 126146 83082 126382 83318
rect 103479 71882 103715 72118
rect 101181 60682 101417 60918
rect 126146 60682 126382 60918
rect 121926 59366 122162 59602
rect 136646 58686 136882 58922
rect 136646 55966 136882 56202
rect 5122 38282 5358 38518
rect 5442 38282 5678 38518
rect 5762 38282 5998 38518
rect 6082 38282 6318 38518
rect 6402 38282 6638 38518
rect 6722 38282 6958 38518
rect 7042 38282 7278 38518
rect 7362 38282 7598 38518
rect 7682 38282 7918 38518
rect 8002 38282 8238 38518
rect 8322 38282 8558 38518
rect 8642 38282 8878 38518
rect 25181 38282 25417 38518
rect 60514 38282 60750 38518
rect 29479 27082 29715 27318
rect 65146 27082 65382 27318
rect 97181 38282 97417 38518
rect 101479 27082 101715 27318
rect 83470 21966 83706 22202
rect 88438 21980 88674 22202
rect 88438 21966 88524 21980
rect 88524 21966 88588 21980
rect 88588 21966 88674 21980
rect 132514 38282 132750 38518
rect 173181 172682 173417 172918
rect 141506 161482 141742 161718
rect 175479 161482 175715 161718
rect 168294 153206 168530 153442
rect 185958 153206 186194 153442
rect 173181 150282 173417 150518
rect 141506 139082 141742 139318
rect 175479 139082 175715 139318
rect 173479 116682 173715 116918
rect 169181 105482 169417 105718
rect 141506 71882 141742 72118
rect 173181 83082 173417 83318
rect 175479 71882 175715 72118
rect 168294 70246 168530 70482
rect 185958 70396 186194 70482
rect 185958 70332 186044 70396
rect 186044 70332 186108 70396
rect 186108 70332 186194 70396
rect 185958 70246 186194 70332
rect 173181 60682 173417 60918
rect 171054 57326 171290 57562
rect 185774 57340 186010 57562
rect 185774 57326 185860 57340
rect 185860 57326 185924 57340
rect 185924 57326 186010 57340
rect 161670 56646 161906 56882
rect 137146 27082 137382 27318
rect 202826 195082 203062 195318
rect 203146 195082 203382 195318
rect 203466 195082 203702 195318
rect 203786 195082 204022 195318
rect 204106 195082 204342 195318
rect 204426 195082 204662 195318
rect 204746 195082 204982 195318
rect 205066 195082 205302 195318
rect 205386 195082 205622 195318
rect 205706 195082 205942 195318
rect 206026 195082 206262 195318
rect 206346 195082 206582 195318
rect 202826 172682 203062 172918
rect 203146 172682 203382 172918
rect 203466 172682 203702 172918
rect 203786 172682 204022 172918
rect 204106 172682 204342 172918
rect 204426 172682 204662 172918
rect 204746 172682 204982 172918
rect 205066 172682 205302 172918
rect 205386 172682 205622 172918
rect 205706 172682 205942 172918
rect 206026 172682 206262 172918
rect 206346 172682 206582 172918
rect 202826 150282 203062 150518
rect 203146 150282 203382 150518
rect 203466 150282 203702 150518
rect 203786 150282 204022 150518
rect 204106 150282 204342 150518
rect 204426 150282 204662 150518
rect 204746 150282 204982 150518
rect 205066 150282 205302 150518
rect 205386 150282 205622 150518
rect 205706 150282 205942 150518
rect 206026 150282 206262 150518
rect 206346 150282 206582 150518
rect 202826 127882 203062 128118
rect 203146 127882 203382 128118
rect 203466 127882 203702 128118
rect 203786 127882 204022 128118
rect 204106 127882 204342 128118
rect 204426 127882 204662 128118
rect 204746 127882 204982 128118
rect 205066 127882 205302 128118
rect 205386 127882 205622 128118
rect 205706 127882 205942 128118
rect 206026 127882 206262 128118
rect 206346 127882 206582 128118
rect 202826 105482 203062 105718
rect 203146 105482 203382 105718
rect 203466 105482 203702 105718
rect 203786 105482 204022 105718
rect 204106 105482 204342 105718
rect 204426 105482 204662 105718
rect 204746 105482 204982 105718
rect 205066 105482 205302 105718
rect 205386 105482 205622 105718
rect 205706 105482 205942 105718
rect 206026 105482 206262 105718
rect 206346 105482 206582 105718
rect 202826 83082 203062 83318
rect 203146 83082 203382 83318
rect 203466 83082 203702 83318
rect 203786 83082 204022 83318
rect 204106 83082 204342 83318
rect 204426 83082 204662 83318
rect 204746 83082 204982 83318
rect 205066 83082 205302 83318
rect 205386 83082 205622 83318
rect 205706 83082 205942 83318
rect 206026 83082 206262 83318
rect 206346 83082 206582 83318
rect 169181 38282 169417 38518
rect 173479 27082 173715 27318
rect 202826 60682 203062 60918
rect 203146 60682 203382 60918
rect 203466 60682 203702 60918
rect 203786 60682 204022 60918
rect 204106 60682 204342 60918
rect 204426 60682 204662 60918
rect 204746 60682 204982 60918
rect 205066 60682 205302 60918
rect 205386 60682 205622 60918
rect 205706 60682 205942 60918
rect 206026 60682 206262 60918
rect 206346 60682 206582 60918
rect 202826 38282 203062 38518
rect 203146 38282 203382 38518
rect 203466 38282 203702 38518
rect 203786 38282 204022 38518
rect 204106 38282 204342 38518
rect 204426 38282 204662 38518
rect 204746 38282 204982 38518
rect 205066 38282 205302 38518
rect 205386 38282 205622 38518
rect 205706 38282 205942 38518
rect 206026 38282 206262 38518
rect 206346 38282 206582 38518
rect 5122 15882 5358 16118
rect 5442 15882 5678 16118
rect 5762 15882 5998 16118
rect 6082 15882 6318 16118
rect 6402 15882 6638 16118
rect 6722 15882 6958 16118
rect 7042 15882 7278 16118
rect 7362 15882 7598 16118
rect 7682 15882 7918 16118
rect 8002 15882 8238 16118
rect 8322 15882 8558 16118
rect 8642 15882 8878 16118
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 202826 15882 203062 16118
rect 203146 15882 203382 16118
rect 203466 15882 203702 16118
rect 203786 15882 204022 16118
rect 204106 15882 204342 16118
rect 204426 15882 204662 16118
rect 204746 15882 204982 16118
rect 205066 15882 205302 16118
rect 205386 15882 205622 16118
rect 205706 15882 205942 16118
rect 206026 15882 206262 16118
rect 206346 15882 206582 16118
rect 202826 8642 203062 8878
rect 203146 8642 203382 8878
rect 203466 8642 203702 8878
rect 203786 8642 204022 8878
rect 204106 8642 204342 8878
rect 204426 8642 204662 8878
rect 204746 8642 204982 8878
rect 205066 8642 205302 8878
rect 205386 8642 205622 8878
rect 205706 8642 205942 8878
rect 206026 8642 206262 8878
rect 206346 8642 206582 8878
rect 202826 8322 203062 8558
rect 203146 8322 203382 8558
rect 203466 8322 203702 8558
rect 203786 8322 204022 8558
rect 204106 8322 204342 8558
rect 204426 8322 204662 8558
rect 204746 8322 204982 8558
rect 205066 8322 205302 8558
rect 205386 8322 205622 8558
rect 205706 8322 205942 8558
rect 206026 8322 206262 8558
rect 206346 8322 206582 8558
rect 202826 8002 203062 8238
rect 203146 8002 203382 8238
rect 203466 8002 203702 8238
rect 203786 8002 204022 8238
rect 204106 8002 204342 8238
rect 204426 8002 204662 8238
rect 204746 8002 204982 8238
rect 205066 8002 205302 8238
rect 205386 8002 205622 8238
rect 205706 8002 205942 8238
rect 206026 8002 206262 8238
rect 206346 8002 206582 8238
rect 202826 7682 203062 7918
rect 203146 7682 203382 7918
rect 203466 7682 203702 7918
rect 203786 7682 204022 7918
rect 204106 7682 204342 7918
rect 204426 7682 204662 7918
rect 204746 7682 204982 7918
rect 205066 7682 205302 7918
rect 205386 7682 205622 7918
rect 205706 7682 205942 7918
rect 206026 7682 206262 7918
rect 206346 7682 206582 7918
rect 202826 7362 203062 7598
rect 203146 7362 203382 7598
rect 203466 7362 203702 7598
rect 203786 7362 204022 7598
rect 204106 7362 204342 7598
rect 204426 7362 204662 7598
rect 204746 7362 204982 7598
rect 205066 7362 205302 7598
rect 205386 7362 205622 7598
rect 205706 7362 205942 7598
rect 206026 7362 206262 7598
rect 206346 7362 206582 7598
rect 202826 7042 203062 7278
rect 203146 7042 203382 7278
rect 203466 7042 203702 7278
rect 203786 7042 204022 7278
rect 204106 7042 204342 7278
rect 204426 7042 204662 7278
rect 204746 7042 204982 7278
rect 205066 7042 205302 7278
rect 205386 7042 205622 7278
rect 205706 7042 205942 7278
rect 206026 7042 206262 7278
rect 206346 7042 206582 7278
rect 202826 6722 203062 6958
rect 203146 6722 203382 6958
rect 203466 6722 203702 6958
rect 203786 6722 204022 6958
rect 204106 6722 204342 6958
rect 204426 6722 204662 6958
rect 204746 6722 204982 6958
rect 205066 6722 205302 6958
rect 205386 6722 205622 6958
rect 205706 6722 205942 6958
rect 206026 6722 206262 6958
rect 206346 6722 206582 6958
rect 202826 6402 203062 6638
rect 203146 6402 203382 6638
rect 203466 6402 203702 6638
rect 203786 6402 204022 6638
rect 204106 6402 204342 6638
rect 204426 6402 204662 6638
rect 204746 6402 204982 6638
rect 205066 6402 205302 6638
rect 205386 6402 205622 6638
rect 205706 6402 205942 6638
rect 206026 6402 206262 6638
rect 206346 6402 206582 6638
rect 202826 6082 203062 6318
rect 203146 6082 203382 6318
rect 203466 6082 203702 6318
rect 203786 6082 204022 6318
rect 204106 6082 204342 6318
rect 204426 6082 204662 6318
rect 204746 6082 204982 6318
rect 205066 6082 205302 6318
rect 205386 6082 205622 6318
rect 205706 6082 205942 6318
rect 206026 6082 206262 6318
rect 206346 6082 206582 6318
rect 202826 5762 203062 5998
rect 203146 5762 203382 5998
rect 203466 5762 203702 5998
rect 203786 5762 204022 5998
rect 204106 5762 204342 5998
rect 204426 5762 204662 5998
rect 204746 5762 204982 5998
rect 205066 5762 205302 5998
rect 205386 5762 205622 5998
rect 205706 5762 205942 5998
rect 206026 5762 206262 5998
rect 206346 5762 206582 5998
rect 202826 5442 203062 5678
rect 203146 5442 203382 5678
rect 203466 5442 203702 5678
rect 203786 5442 204022 5678
rect 204106 5442 204342 5678
rect 204426 5442 204662 5678
rect 204746 5442 204982 5678
rect 205066 5442 205302 5678
rect 205386 5442 205622 5678
rect 205706 5442 205942 5678
rect 206026 5442 206262 5678
rect 206346 5442 206582 5678
rect 202826 5122 203062 5358
rect 203146 5122 203382 5358
rect 203466 5122 203702 5358
rect 203786 5122 204022 5358
rect 204106 5122 204342 5358
rect 204426 5122 204662 5358
rect 204746 5122 204982 5358
rect 205066 5122 205302 5358
rect 205386 5122 205622 5358
rect 205706 5122 205942 5358
rect 206026 5122 206262 5358
rect 206346 5122 206582 5358
rect 207826 206282 208062 206518
rect 208146 206282 208382 206518
rect 208466 206282 208702 206518
rect 208786 206282 209022 206518
rect 209106 206282 209342 206518
rect 209426 206282 209662 206518
rect 209746 206282 209982 206518
rect 210066 206282 210302 206518
rect 210386 206282 210622 206518
rect 210706 206282 210942 206518
rect 211026 206282 211262 206518
rect 211346 206282 211582 206518
rect 207826 183882 208062 184118
rect 208146 183882 208382 184118
rect 208466 183882 208702 184118
rect 208786 183882 209022 184118
rect 209106 183882 209342 184118
rect 209426 183882 209662 184118
rect 209746 183882 209982 184118
rect 210066 183882 210302 184118
rect 210386 183882 210622 184118
rect 210706 183882 210942 184118
rect 211026 183882 211262 184118
rect 211346 183882 211582 184118
rect 207826 161482 208062 161718
rect 208146 161482 208382 161718
rect 208466 161482 208702 161718
rect 208786 161482 209022 161718
rect 209106 161482 209342 161718
rect 209426 161482 209662 161718
rect 209746 161482 209982 161718
rect 210066 161482 210302 161718
rect 210386 161482 210622 161718
rect 210706 161482 210942 161718
rect 211026 161482 211262 161718
rect 211346 161482 211582 161718
rect 207826 139082 208062 139318
rect 208146 139082 208382 139318
rect 208466 139082 208702 139318
rect 208786 139082 209022 139318
rect 209106 139082 209342 139318
rect 209426 139082 209662 139318
rect 209746 139082 209982 139318
rect 210066 139082 210302 139318
rect 210386 139082 210622 139318
rect 210706 139082 210942 139318
rect 211026 139082 211262 139318
rect 211346 139082 211582 139318
rect 207826 116682 208062 116918
rect 208146 116682 208382 116918
rect 208466 116682 208702 116918
rect 208786 116682 209022 116918
rect 209106 116682 209342 116918
rect 209426 116682 209662 116918
rect 209746 116682 209982 116918
rect 210066 116682 210302 116918
rect 210386 116682 210622 116918
rect 210706 116682 210942 116918
rect 211026 116682 211262 116918
rect 211346 116682 211582 116918
rect 207826 94282 208062 94518
rect 208146 94282 208382 94518
rect 208466 94282 208702 94518
rect 208786 94282 209022 94518
rect 209106 94282 209342 94518
rect 209426 94282 209662 94518
rect 209746 94282 209982 94518
rect 210066 94282 210302 94518
rect 210386 94282 210622 94518
rect 210706 94282 210942 94518
rect 211026 94282 211262 94518
rect 211346 94282 211582 94518
rect 207826 71882 208062 72118
rect 208146 71882 208382 72118
rect 208466 71882 208702 72118
rect 208786 71882 209022 72118
rect 209106 71882 209342 72118
rect 209426 71882 209662 72118
rect 209746 71882 209982 72118
rect 210066 71882 210302 72118
rect 210386 71882 210622 72118
rect 210706 71882 210942 72118
rect 211026 71882 211262 72118
rect 211346 71882 211582 72118
rect 207826 49482 208062 49718
rect 208146 49482 208382 49718
rect 208466 49482 208702 49718
rect 208786 49482 209022 49718
rect 209106 49482 209342 49718
rect 209426 49482 209662 49718
rect 209746 49482 209982 49718
rect 210066 49482 210302 49718
rect 210386 49482 210622 49718
rect 210706 49482 210942 49718
rect 211026 49482 211262 49718
rect 211346 49482 211582 49718
rect 207826 27082 208062 27318
rect 208146 27082 208382 27318
rect 208466 27082 208702 27318
rect 208786 27082 209022 27318
rect 209106 27082 209342 27318
rect 209426 27082 209662 27318
rect 209746 27082 209982 27318
rect 210066 27082 210302 27318
rect 210386 27082 210622 27318
rect 210706 27082 210942 27318
rect 211026 27082 211262 27318
rect 211346 27082 211582 27318
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 207826 3642 208062 3878
rect 208146 3642 208382 3878
rect 208466 3642 208702 3878
rect 208786 3642 209022 3878
rect 209106 3642 209342 3878
rect 209426 3642 209662 3878
rect 209746 3642 209982 3878
rect 210066 3642 210302 3878
rect 210386 3642 210622 3878
rect 210706 3642 210942 3878
rect 211026 3642 211262 3878
rect 211346 3642 211582 3878
rect 207826 3322 208062 3558
rect 208146 3322 208382 3558
rect 208466 3322 208702 3558
rect 208786 3322 209022 3558
rect 209106 3322 209342 3558
rect 209426 3322 209662 3558
rect 209746 3322 209982 3558
rect 210066 3322 210302 3558
rect 210386 3322 210622 3558
rect 210706 3322 210942 3558
rect 211026 3322 211262 3558
rect 211346 3322 211582 3558
rect 207826 3002 208062 3238
rect 208146 3002 208382 3238
rect 208466 3002 208702 3238
rect 208786 3002 209022 3238
rect 209106 3002 209342 3238
rect 209426 3002 209662 3238
rect 209746 3002 209982 3238
rect 210066 3002 210302 3238
rect 210386 3002 210622 3238
rect 210706 3002 210942 3238
rect 211026 3002 211262 3238
rect 211346 3002 211582 3238
rect 207826 2682 208062 2918
rect 208146 2682 208382 2918
rect 208466 2682 208702 2918
rect 208786 2682 209022 2918
rect 209106 2682 209342 2918
rect 209426 2682 209662 2918
rect 209746 2682 209982 2918
rect 210066 2682 210302 2918
rect 210386 2682 210622 2918
rect 210706 2682 210942 2918
rect 211026 2682 211262 2918
rect 211346 2682 211582 2918
rect 207826 2362 208062 2598
rect 208146 2362 208382 2598
rect 208466 2362 208702 2598
rect 208786 2362 209022 2598
rect 209106 2362 209342 2598
rect 209426 2362 209662 2598
rect 209746 2362 209982 2598
rect 210066 2362 210302 2598
rect 210386 2362 210622 2598
rect 210706 2362 210942 2598
rect 211026 2362 211262 2598
rect 211346 2362 211582 2598
rect 207826 2042 208062 2278
rect 208146 2042 208382 2278
rect 208466 2042 208702 2278
rect 208786 2042 209022 2278
rect 209106 2042 209342 2278
rect 209426 2042 209662 2278
rect 209746 2042 209982 2278
rect 210066 2042 210302 2278
rect 210386 2042 210622 2278
rect 210706 2042 210942 2278
rect 211026 2042 211262 2278
rect 211346 2042 211582 2278
rect 207826 1722 208062 1958
rect 208146 1722 208382 1958
rect 208466 1722 208702 1958
rect 208786 1722 209022 1958
rect 209106 1722 209342 1958
rect 209426 1722 209662 1958
rect 209746 1722 209982 1958
rect 210066 1722 210302 1958
rect 210386 1722 210622 1958
rect 210706 1722 210942 1958
rect 211026 1722 211262 1958
rect 211346 1722 211582 1958
rect 207826 1402 208062 1638
rect 208146 1402 208382 1638
rect 208466 1402 208702 1638
rect 208786 1402 209022 1638
rect 209106 1402 209342 1638
rect 209426 1402 209662 1638
rect 209746 1402 209982 1638
rect 210066 1402 210302 1638
rect 210386 1402 210622 1638
rect 210706 1402 210942 1638
rect 211026 1402 211262 1638
rect 211346 1402 211582 1638
rect 207826 1082 208062 1318
rect 208146 1082 208382 1318
rect 208466 1082 208702 1318
rect 208786 1082 209022 1318
rect 209106 1082 209342 1318
rect 209426 1082 209662 1318
rect 209746 1082 209982 1318
rect 210066 1082 210302 1318
rect 210386 1082 210622 1318
rect 210706 1082 210942 1318
rect 211026 1082 211262 1318
rect 211346 1082 211582 1318
rect 207826 762 208062 998
rect 208146 762 208382 998
rect 208466 762 208702 998
rect 208786 762 209022 998
rect 209106 762 209342 998
rect 209426 762 209662 998
rect 209746 762 209982 998
rect 210066 762 210302 998
rect 210386 762 210622 998
rect 210706 762 210942 998
rect 211026 762 211262 998
rect 211346 762 211582 998
rect 207826 442 208062 678
rect 208146 442 208382 678
rect 208466 442 208702 678
rect 208786 442 209022 678
rect 209106 442 209342 678
rect 209426 442 209662 678
rect 209746 442 209982 678
rect 210066 442 210302 678
rect 210386 442 210622 678
rect 210706 442 210942 678
rect 211026 442 211262 678
rect 211346 442 211582 678
rect 207826 122 208062 358
rect 208146 122 208382 358
rect 208466 122 208702 358
rect 208786 122 209022 358
rect 209106 122 209342 358
rect 209426 122 209662 358
rect 209746 122 209982 358
rect 210066 122 210302 358
rect 210386 122 210622 358
rect 210706 122 210942 358
rect 211026 122 211262 358
rect 211346 122 211582 358
<< metal5 >>
rect 0 229142 211704 229264
rect 0 228906 122 229142
rect 358 228906 442 229142
rect 678 228906 762 229142
rect 998 228906 1082 229142
rect 1318 228906 1402 229142
rect 1638 228906 1722 229142
rect 1958 228906 2042 229142
rect 2278 228906 2362 229142
rect 2598 228906 2682 229142
rect 2918 228906 3002 229142
rect 3238 228906 3322 229142
rect 3558 228906 3642 229142
rect 3878 228906 207826 229142
rect 208062 228906 208146 229142
rect 208382 228906 208466 229142
rect 208702 228906 208786 229142
rect 209022 228906 209106 229142
rect 209342 228906 209426 229142
rect 209662 228906 209746 229142
rect 209982 228906 210066 229142
rect 210302 228906 210386 229142
rect 210622 228906 210706 229142
rect 210942 228906 211026 229142
rect 211262 228906 211346 229142
rect 211582 228906 211704 229142
rect 0 228822 211704 228906
rect 0 228586 122 228822
rect 358 228586 442 228822
rect 678 228586 762 228822
rect 998 228586 1082 228822
rect 1318 228586 1402 228822
rect 1638 228586 1722 228822
rect 1958 228586 2042 228822
rect 2278 228586 2362 228822
rect 2598 228586 2682 228822
rect 2918 228586 3002 228822
rect 3238 228586 3322 228822
rect 3558 228586 3642 228822
rect 3878 228586 207826 228822
rect 208062 228586 208146 228822
rect 208382 228586 208466 228822
rect 208702 228586 208786 228822
rect 209022 228586 209106 228822
rect 209342 228586 209426 228822
rect 209662 228586 209746 228822
rect 209982 228586 210066 228822
rect 210302 228586 210386 228822
rect 210622 228586 210706 228822
rect 210942 228586 211026 228822
rect 211262 228586 211346 228822
rect 211582 228586 211704 228822
rect 0 228502 211704 228586
rect 0 228266 122 228502
rect 358 228266 442 228502
rect 678 228266 762 228502
rect 998 228266 1082 228502
rect 1318 228266 1402 228502
rect 1638 228266 1722 228502
rect 1958 228266 2042 228502
rect 2278 228266 2362 228502
rect 2598 228266 2682 228502
rect 2918 228266 3002 228502
rect 3238 228266 3322 228502
rect 3558 228266 3642 228502
rect 3878 228266 207826 228502
rect 208062 228266 208146 228502
rect 208382 228266 208466 228502
rect 208702 228266 208786 228502
rect 209022 228266 209106 228502
rect 209342 228266 209426 228502
rect 209662 228266 209746 228502
rect 209982 228266 210066 228502
rect 210302 228266 210386 228502
rect 210622 228266 210706 228502
rect 210942 228266 211026 228502
rect 211262 228266 211346 228502
rect 211582 228266 211704 228502
rect 0 228182 211704 228266
rect 0 227946 122 228182
rect 358 227946 442 228182
rect 678 227946 762 228182
rect 998 227946 1082 228182
rect 1318 227946 1402 228182
rect 1638 227946 1722 228182
rect 1958 227946 2042 228182
rect 2278 227946 2362 228182
rect 2598 227946 2682 228182
rect 2918 227946 3002 228182
rect 3238 227946 3322 228182
rect 3558 227946 3642 228182
rect 3878 227946 207826 228182
rect 208062 227946 208146 228182
rect 208382 227946 208466 228182
rect 208702 227946 208786 228182
rect 209022 227946 209106 228182
rect 209342 227946 209426 228182
rect 209662 227946 209746 228182
rect 209982 227946 210066 228182
rect 210302 227946 210386 228182
rect 210622 227946 210706 228182
rect 210942 227946 211026 228182
rect 211262 227946 211346 228182
rect 211582 227946 211704 228182
rect 0 227862 211704 227946
rect 0 227626 122 227862
rect 358 227626 442 227862
rect 678 227626 762 227862
rect 998 227626 1082 227862
rect 1318 227626 1402 227862
rect 1638 227626 1722 227862
rect 1958 227626 2042 227862
rect 2278 227626 2362 227862
rect 2598 227626 2682 227862
rect 2918 227626 3002 227862
rect 3238 227626 3322 227862
rect 3558 227626 3642 227862
rect 3878 227626 207826 227862
rect 208062 227626 208146 227862
rect 208382 227626 208466 227862
rect 208702 227626 208786 227862
rect 209022 227626 209106 227862
rect 209342 227626 209426 227862
rect 209662 227626 209746 227862
rect 209982 227626 210066 227862
rect 210302 227626 210386 227862
rect 210622 227626 210706 227862
rect 210942 227626 211026 227862
rect 211262 227626 211346 227862
rect 211582 227626 211704 227862
rect 0 227542 211704 227626
rect 0 227306 122 227542
rect 358 227306 442 227542
rect 678 227306 762 227542
rect 998 227306 1082 227542
rect 1318 227306 1402 227542
rect 1638 227306 1722 227542
rect 1958 227306 2042 227542
rect 2278 227306 2362 227542
rect 2598 227306 2682 227542
rect 2918 227306 3002 227542
rect 3238 227306 3322 227542
rect 3558 227306 3642 227542
rect 3878 227306 207826 227542
rect 208062 227306 208146 227542
rect 208382 227306 208466 227542
rect 208702 227306 208786 227542
rect 209022 227306 209106 227542
rect 209342 227306 209426 227542
rect 209662 227306 209746 227542
rect 209982 227306 210066 227542
rect 210302 227306 210386 227542
rect 210622 227306 210706 227542
rect 210942 227306 211026 227542
rect 211262 227306 211346 227542
rect 211582 227306 211704 227542
rect 0 227222 211704 227306
rect 0 226986 122 227222
rect 358 226986 442 227222
rect 678 226986 762 227222
rect 998 226986 1082 227222
rect 1318 226986 1402 227222
rect 1638 226986 1722 227222
rect 1958 226986 2042 227222
rect 2278 226986 2362 227222
rect 2598 226986 2682 227222
rect 2918 226986 3002 227222
rect 3238 226986 3322 227222
rect 3558 226986 3642 227222
rect 3878 226986 207826 227222
rect 208062 226986 208146 227222
rect 208382 226986 208466 227222
rect 208702 226986 208786 227222
rect 209022 226986 209106 227222
rect 209342 226986 209426 227222
rect 209662 226986 209746 227222
rect 209982 226986 210066 227222
rect 210302 226986 210386 227222
rect 210622 226986 210706 227222
rect 210942 226986 211026 227222
rect 211262 226986 211346 227222
rect 211582 226986 211704 227222
rect 0 226902 211704 226986
rect 0 226666 122 226902
rect 358 226666 442 226902
rect 678 226666 762 226902
rect 998 226666 1082 226902
rect 1318 226666 1402 226902
rect 1638 226666 1722 226902
rect 1958 226666 2042 226902
rect 2278 226666 2362 226902
rect 2598 226666 2682 226902
rect 2918 226666 3002 226902
rect 3238 226666 3322 226902
rect 3558 226666 3642 226902
rect 3878 226666 207826 226902
rect 208062 226666 208146 226902
rect 208382 226666 208466 226902
rect 208702 226666 208786 226902
rect 209022 226666 209106 226902
rect 209342 226666 209426 226902
rect 209662 226666 209746 226902
rect 209982 226666 210066 226902
rect 210302 226666 210386 226902
rect 210622 226666 210706 226902
rect 210942 226666 211026 226902
rect 211262 226666 211346 226902
rect 211582 226666 211704 226902
rect 0 226582 211704 226666
rect 0 226346 122 226582
rect 358 226346 442 226582
rect 678 226346 762 226582
rect 998 226346 1082 226582
rect 1318 226346 1402 226582
rect 1638 226346 1722 226582
rect 1958 226346 2042 226582
rect 2278 226346 2362 226582
rect 2598 226346 2682 226582
rect 2918 226346 3002 226582
rect 3238 226346 3322 226582
rect 3558 226346 3642 226582
rect 3878 226346 207826 226582
rect 208062 226346 208146 226582
rect 208382 226346 208466 226582
rect 208702 226346 208786 226582
rect 209022 226346 209106 226582
rect 209342 226346 209426 226582
rect 209662 226346 209746 226582
rect 209982 226346 210066 226582
rect 210302 226346 210386 226582
rect 210622 226346 210706 226582
rect 210942 226346 211026 226582
rect 211262 226346 211346 226582
rect 211582 226346 211704 226582
rect 0 226262 211704 226346
rect 0 226026 122 226262
rect 358 226026 442 226262
rect 678 226026 762 226262
rect 998 226026 1082 226262
rect 1318 226026 1402 226262
rect 1638 226026 1722 226262
rect 1958 226026 2042 226262
rect 2278 226026 2362 226262
rect 2598 226026 2682 226262
rect 2918 226026 3002 226262
rect 3238 226026 3322 226262
rect 3558 226026 3642 226262
rect 3878 226026 207826 226262
rect 208062 226026 208146 226262
rect 208382 226026 208466 226262
rect 208702 226026 208786 226262
rect 209022 226026 209106 226262
rect 209342 226026 209426 226262
rect 209662 226026 209746 226262
rect 209982 226026 210066 226262
rect 210302 226026 210386 226262
rect 210622 226026 210706 226262
rect 210942 226026 211026 226262
rect 211262 226026 211346 226262
rect 211582 226026 211704 226262
rect 0 225942 211704 226026
rect 0 225706 122 225942
rect 358 225706 442 225942
rect 678 225706 762 225942
rect 998 225706 1082 225942
rect 1318 225706 1402 225942
rect 1638 225706 1722 225942
rect 1958 225706 2042 225942
rect 2278 225706 2362 225942
rect 2598 225706 2682 225942
rect 2918 225706 3002 225942
rect 3238 225706 3322 225942
rect 3558 225706 3642 225942
rect 3878 225706 207826 225942
rect 208062 225706 208146 225942
rect 208382 225706 208466 225942
rect 208702 225706 208786 225942
rect 209022 225706 209106 225942
rect 209342 225706 209426 225942
rect 209662 225706 209746 225942
rect 209982 225706 210066 225942
rect 210302 225706 210386 225942
rect 210622 225706 210706 225942
rect 210942 225706 211026 225942
rect 211262 225706 211346 225942
rect 211582 225706 211704 225942
rect 0 225622 211704 225706
rect 0 225386 122 225622
rect 358 225386 442 225622
rect 678 225386 762 225622
rect 998 225386 1082 225622
rect 1318 225386 1402 225622
rect 1638 225386 1722 225622
rect 1958 225386 2042 225622
rect 2278 225386 2362 225622
rect 2598 225386 2682 225622
rect 2918 225386 3002 225622
rect 3238 225386 3322 225622
rect 3558 225386 3642 225622
rect 3878 225386 207826 225622
rect 208062 225386 208146 225622
rect 208382 225386 208466 225622
rect 208702 225386 208786 225622
rect 209022 225386 209106 225622
rect 209342 225386 209426 225622
rect 209662 225386 209746 225622
rect 209982 225386 210066 225622
rect 210302 225386 210386 225622
rect 210622 225386 210706 225622
rect 210942 225386 211026 225622
rect 211262 225386 211346 225622
rect 211582 225386 211704 225622
rect 0 225264 211704 225386
rect 5000 224142 206704 224264
rect 5000 223906 5122 224142
rect 5358 223906 5442 224142
rect 5678 223906 5762 224142
rect 5998 223906 6082 224142
rect 6318 223906 6402 224142
rect 6638 223906 6722 224142
rect 6958 223906 7042 224142
rect 7278 223906 7362 224142
rect 7598 223906 7682 224142
rect 7918 223906 8002 224142
rect 8238 223906 8322 224142
rect 8558 223906 8642 224142
rect 8878 223906 202826 224142
rect 203062 223906 203146 224142
rect 203382 223906 203466 224142
rect 203702 223906 203786 224142
rect 204022 223906 204106 224142
rect 204342 223906 204426 224142
rect 204662 223906 204746 224142
rect 204982 223906 205066 224142
rect 205302 223906 205386 224142
rect 205622 223906 205706 224142
rect 205942 223906 206026 224142
rect 206262 223906 206346 224142
rect 206582 223906 206704 224142
rect 5000 223822 206704 223906
rect 5000 223586 5122 223822
rect 5358 223586 5442 223822
rect 5678 223586 5762 223822
rect 5998 223586 6082 223822
rect 6318 223586 6402 223822
rect 6638 223586 6722 223822
rect 6958 223586 7042 223822
rect 7278 223586 7362 223822
rect 7598 223586 7682 223822
rect 7918 223586 8002 223822
rect 8238 223586 8322 223822
rect 8558 223586 8642 223822
rect 8878 223586 202826 223822
rect 203062 223586 203146 223822
rect 203382 223586 203466 223822
rect 203702 223586 203786 223822
rect 204022 223586 204106 223822
rect 204342 223586 204426 223822
rect 204662 223586 204746 223822
rect 204982 223586 205066 223822
rect 205302 223586 205386 223822
rect 205622 223586 205706 223822
rect 205942 223586 206026 223822
rect 206262 223586 206346 223822
rect 206582 223586 206704 223822
rect 5000 223502 206704 223586
rect 5000 223266 5122 223502
rect 5358 223266 5442 223502
rect 5678 223266 5762 223502
rect 5998 223266 6082 223502
rect 6318 223266 6402 223502
rect 6638 223266 6722 223502
rect 6958 223266 7042 223502
rect 7278 223266 7362 223502
rect 7598 223266 7682 223502
rect 7918 223266 8002 223502
rect 8238 223266 8322 223502
rect 8558 223266 8642 223502
rect 8878 223266 202826 223502
rect 203062 223266 203146 223502
rect 203382 223266 203466 223502
rect 203702 223266 203786 223502
rect 204022 223266 204106 223502
rect 204342 223266 204426 223502
rect 204662 223266 204746 223502
rect 204982 223266 205066 223502
rect 205302 223266 205386 223502
rect 205622 223266 205706 223502
rect 205942 223266 206026 223502
rect 206262 223266 206346 223502
rect 206582 223266 206704 223502
rect 5000 223182 206704 223266
rect 5000 222946 5122 223182
rect 5358 222946 5442 223182
rect 5678 222946 5762 223182
rect 5998 222946 6082 223182
rect 6318 222946 6402 223182
rect 6638 222946 6722 223182
rect 6958 222946 7042 223182
rect 7278 222946 7362 223182
rect 7598 222946 7682 223182
rect 7918 222946 8002 223182
rect 8238 222946 8322 223182
rect 8558 222946 8642 223182
rect 8878 222946 202826 223182
rect 203062 222946 203146 223182
rect 203382 222946 203466 223182
rect 203702 222946 203786 223182
rect 204022 222946 204106 223182
rect 204342 222946 204426 223182
rect 204662 222946 204746 223182
rect 204982 222946 205066 223182
rect 205302 222946 205386 223182
rect 205622 222946 205706 223182
rect 205942 222946 206026 223182
rect 206262 222946 206346 223182
rect 206582 222946 206704 223182
rect 5000 222862 206704 222946
rect 5000 222626 5122 222862
rect 5358 222626 5442 222862
rect 5678 222626 5762 222862
rect 5998 222626 6082 222862
rect 6318 222626 6402 222862
rect 6638 222626 6722 222862
rect 6958 222626 7042 222862
rect 7278 222626 7362 222862
rect 7598 222626 7682 222862
rect 7918 222626 8002 222862
rect 8238 222626 8322 222862
rect 8558 222626 8642 222862
rect 8878 222626 202826 222862
rect 203062 222626 203146 222862
rect 203382 222626 203466 222862
rect 203702 222626 203786 222862
rect 204022 222626 204106 222862
rect 204342 222626 204426 222862
rect 204662 222626 204746 222862
rect 204982 222626 205066 222862
rect 205302 222626 205386 222862
rect 205622 222626 205706 222862
rect 205942 222626 206026 222862
rect 206262 222626 206346 222862
rect 206582 222626 206704 222862
rect 5000 222542 206704 222626
rect 5000 222306 5122 222542
rect 5358 222306 5442 222542
rect 5678 222306 5762 222542
rect 5998 222306 6082 222542
rect 6318 222306 6402 222542
rect 6638 222306 6722 222542
rect 6958 222306 7042 222542
rect 7278 222306 7362 222542
rect 7598 222306 7682 222542
rect 7918 222306 8002 222542
rect 8238 222306 8322 222542
rect 8558 222306 8642 222542
rect 8878 222306 202826 222542
rect 203062 222306 203146 222542
rect 203382 222306 203466 222542
rect 203702 222306 203786 222542
rect 204022 222306 204106 222542
rect 204342 222306 204426 222542
rect 204662 222306 204746 222542
rect 204982 222306 205066 222542
rect 205302 222306 205386 222542
rect 205622 222306 205706 222542
rect 205942 222306 206026 222542
rect 206262 222306 206346 222542
rect 206582 222306 206704 222542
rect 5000 222222 206704 222306
rect 5000 221986 5122 222222
rect 5358 221986 5442 222222
rect 5678 221986 5762 222222
rect 5998 221986 6082 222222
rect 6318 221986 6402 222222
rect 6638 221986 6722 222222
rect 6958 221986 7042 222222
rect 7278 221986 7362 222222
rect 7598 221986 7682 222222
rect 7918 221986 8002 222222
rect 8238 221986 8322 222222
rect 8558 221986 8642 222222
rect 8878 221986 202826 222222
rect 203062 221986 203146 222222
rect 203382 221986 203466 222222
rect 203702 221986 203786 222222
rect 204022 221986 204106 222222
rect 204342 221986 204426 222222
rect 204662 221986 204746 222222
rect 204982 221986 205066 222222
rect 205302 221986 205386 222222
rect 205622 221986 205706 222222
rect 205942 221986 206026 222222
rect 206262 221986 206346 222222
rect 206582 221986 206704 222222
rect 5000 221902 206704 221986
rect 5000 221666 5122 221902
rect 5358 221666 5442 221902
rect 5678 221666 5762 221902
rect 5998 221666 6082 221902
rect 6318 221666 6402 221902
rect 6638 221666 6722 221902
rect 6958 221666 7042 221902
rect 7278 221666 7362 221902
rect 7598 221666 7682 221902
rect 7918 221666 8002 221902
rect 8238 221666 8322 221902
rect 8558 221666 8642 221902
rect 8878 221666 202826 221902
rect 203062 221666 203146 221902
rect 203382 221666 203466 221902
rect 203702 221666 203786 221902
rect 204022 221666 204106 221902
rect 204342 221666 204426 221902
rect 204662 221666 204746 221902
rect 204982 221666 205066 221902
rect 205302 221666 205386 221902
rect 205622 221666 205706 221902
rect 205942 221666 206026 221902
rect 206262 221666 206346 221902
rect 206582 221666 206704 221902
rect 5000 221582 206704 221666
rect 5000 221346 5122 221582
rect 5358 221346 5442 221582
rect 5678 221346 5762 221582
rect 5998 221346 6082 221582
rect 6318 221346 6402 221582
rect 6638 221346 6722 221582
rect 6958 221346 7042 221582
rect 7278 221346 7362 221582
rect 7598 221346 7682 221582
rect 7918 221346 8002 221582
rect 8238 221346 8322 221582
rect 8558 221346 8642 221582
rect 8878 221346 202826 221582
rect 203062 221346 203146 221582
rect 203382 221346 203466 221582
rect 203702 221346 203786 221582
rect 204022 221346 204106 221582
rect 204342 221346 204426 221582
rect 204662 221346 204746 221582
rect 204982 221346 205066 221582
rect 205302 221346 205386 221582
rect 205622 221346 205706 221582
rect 205942 221346 206026 221582
rect 206262 221346 206346 221582
rect 206582 221346 206704 221582
rect 5000 221262 206704 221346
rect 5000 221026 5122 221262
rect 5358 221026 5442 221262
rect 5678 221026 5762 221262
rect 5998 221026 6082 221262
rect 6318 221026 6402 221262
rect 6638 221026 6722 221262
rect 6958 221026 7042 221262
rect 7278 221026 7362 221262
rect 7598 221026 7682 221262
rect 7918 221026 8002 221262
rect 8238 221026 8322 221262
rect 8558 221026 8642 221262
rect 8878 221026 202826 221262
rect 203062 221026 203146 221262
rect 203382 221026 203466 221262
rect 203702 221026 203786 221262
rect 204022 221026 204106 221262
rect 204342 221026 204426 221262
rect 204662 221026 204746 221262
rect 204982 221026 205066 221262
rect 205302 221026 205386 221262
rect 205622 221026 205706 221262
rect 205942 221026 206026 221262
rect 206262 221026 206346 221262
rect 206582 221026 206704 221262
rect 5000 220942 206704 221026
rect 5000 220706 5122 220942
rect 5358 220706 5442 220942
rect 5678 220706 5762 220942
rect 5998 220706 6082 220942
rect 6318 220706 6402 220942
rect 6638 220706 6722 220942
rect 6958 220706 7042 220942
rect 7278 220706 7362 220942
rect 7598 220706 7682 220942
rect 7918 220706 8002 220942
rect 8238 220706 8322 220942
rect 8558 220706 8642 220942
rect 8878 220706 202826 220942
rect 203062 220706 203146 220942
rect 203382 220706 203466 220942
rect 203702 220706 203786 220942
rect 204022 220706 204106 220942
rect 204342 220706 204426 220942
rect 204662 220706 204746 220942
rect 204982 220706 205066 220942
rect 205302 220706 205386 220942
rect 205622 220706 205706 220942
rect 205942 220706 206026 220942
rect 206262 220706 206346 220942
rect 206582 220706 206704 220942
rect 5000 220622 206704 220706
rect 5000 220386 5122 220622
rect 5358 220386 5442 220622
rect 5678 220386 5762 220622
rect 5998 220386 6082 220622
rect 6318 220386 6402 220622
rect 6638 220386 6722 220622
rect 6958 220386 7042 220622
rect 7278 220386 7362 220622
rect 7598 220386 7682 220622
rect 7918 220386 8002 220622
rect 8238 220386 8322 220622
rect 8558 220386 8642 220622
rect 8878 220386 202826 220622
rect 203062 220386 203146 220622
rect 203382 220386 203466 220622
rect 203702 220386 203786 220622
rect 204022 220386 204106 220622
rect 204342 220386 204426 220622
rect 204662 220386 204746 220622
rect 204982 220386 205066 220622
rect 205302 220386 205386 220622
rect 205622 220386 205706 220622
rect 205942 220386 206026 220622
rect 206262 220386 206346 220622
rect 206582 220386 206704 220622
rect 5000 220264 206704 220386
rect 0 217718 211704 217760
rect 0 217482 5122 217718
rect 5358 217482 5442 217718
rect 5678 217482 5762 217718
rect 5998 217482 6082 217718
rect 6318 217482 6402 217718
rect 6638 217482 6722 217718
rect 6958 217482 7042 217718
rect 7278 217482 7362 217718
rect 7598 217482 7682 217718
rect 7918 217482 8002 217718
rect 8238 217482 8322 217718
rect 8558 217482 8642 217718
rect 8878 217482 202826 217718
rect 203062 217482 203146 217718
rect 203382 217482 203466 217718
rect 203702 217482 203786 217718
rect 204022 217482 204106 217718
rect 204342 217482 204426 217718
rect 204662 217482 204746 217718
rect 204982 217482 205066 217718
rect 205302 217482 205386 217718
rect 205622 217482 205706 217718
rect 205942 217482 206026 217718
rect 206262 217482 206346 217718
rect 206582 217482 211704 217718
rect 0 217440 211704 217482
rect 0 206518 211704 206560
rect 0 206282 122 206518
rect 358 206282 442 206518
rect 678 206282 762 206518
rect 998 206282 1082 206518
rect 1318 206282 1402 206518
rect 1638 206282 1722 206518
rect 1958 206282 2042 206518
rect 2278 206282 2362 206518
rect 2598 206282 2682 206518
rect 2918 206282 3002 206518
rect 3238 206282 3322 206518
rect 3558 206282 3642 206518
rect 3878 206282 29190 206518
rect 29426 206282 65146 206518
rect 65382 206282 101479 206518
rect 101715 206282 137146 206518
rect 137382 206282 173479 206518
rect 173715 206282 207826 206518
rect 208062 206282 208146 206518
rect 208382 206282 208466 206518
rect 208702 206282 208786 206518
rect 209022 206282 209106 206518
rect 209342 206282 209426 206518
rect 209662 206282 209746 206518
rect 209982 206282 210066 206518
rect 210302 206282 210386 206518
rect 210622 206282 210706 206518
rect 210942 206282 211026 206518
rect 211262 206282 211346 206518
rect 211582 206282 211704 206518
rect 0 206240 211704 206282
rect 0 195318 211704 195360
rect 0 195082 5122 195318
rect 5358 195082 5442 195318
rect 5678 195082 5762 195318
rect 5998 195082 6082 195318
rect 6318 195082 6402 195318
rect 6638 195082 6722 195318
rect 6958 195082 7042 195318
rect 7278 195082 7362 195318
rect 7598 195082 7682 195318
rect 7918 195082 8002 195318
rect 8238 195082 8322 195318
rect 8558 195082 8642 195318
rect 8878 195082 24892 195318
rect 25128 195082 60514 195318
rect 60750 195082 97181 195318
rect 97417 195082 132514 195318
rect 132750 195082 169181 195318
rect 169417 195082 202826 195318
rect 203062 195082 203146 195318
rect 203382 195082 203466 195318
rect 203702 195082 203786 195318
rect 204022 195082 204106 195318
rect 204342 195082 204426 195318
rect 204662 195082 204746 195318
rect 204982 195082 205066 195318
rect 205302 195082 205386 195318
rect 205622 195082 205706 195318
rect 205942 195082 206026 195318
rect 206262 195082 206346 195318
rect 206582 195082 211704 195318
rect 0 195040 211704 195082
rect 0 184118 211704 184160
rect 0 183882 122 184118
rect 358 183882 442 184118
rect 678 183882 762 184118
rect 998 183882 1082 184118
rect 1318 183882 1402 184118
rect 1638 183882 1722 184118
rect 1958 183882 2042 184118
rect 2278 183882 2362 184118
rect 2598 183882 2682 184118
rect 2918 183882 3002 184118
rect 3238 183882 3322 184118
rect 3558 183882 3642 184118
rect 3878 183882 207826 184118
rect 208062 183882 208146 184118
rect 208382 183882 208466 184118
rect 208702 183882 208786 184118
rect 209022 183882 209106 184118
rect 209342 183882 209426 184118
rect 209662 183882 209746 184118
rect 209982 183882 210066 184118
rect 210302 183882 210386 184118
rect 210622 183882 210706 184118
rect 210942 183882 211026 184118
rect 211262 183882 211346 184118
rect 211582 183882 211704 184118
rect 0 183840 211704 183882
rect 0 172918 211704 172960
rect 0 172682 5122 172918
rect 5358 172682 5442 172918
rect 5678 172682 5762 172918
rect 5998 172682 6082 172918
rect 6318 172682 6402 172918
rect 6638 172682 6722 172918
rect 6958 172682 7042 172918
rect 7278 172682 7362 172918
rect 7598 172682 7682 172918
rect 7918 172682 8002 172918
rect 8238 172682 8322 172918
rect 8558 172682 8642 172918
rect 8878 172682 29181 172918
rect 29417 172682 54146 172918
rect 54382 172682 101181 172918
rect 101417 172682 126146 172918
rect 126382 172682 173181 172918
rect 173417 172682 202826 172918
rect 203062 172682 203146 172918
rect 203382 172682 203466 172918
rect 203702 172682 203786 172918
rect 204022 172682 204106 172918
rect 204342 172682 204426 172918
rect 204662 172682 204746 172918
rect 204982 172682 205066 172918
rect 205302 172682 205386 172918
rect 205622 172682 205706 172918
rect 205942 172682 206026 172918
rect 206262 172682 206346 172918
rect 206582 172682 211704 172918
rect 0 172640 211704 172682
rect 0 161718 211704 161760
rect 0 161482 122 161718
rect 358 161482 442 161718
rect 678 161482 762 161718
rect 998 161482 1082 161718
rect 1318 161482 1402 161718
rect 1638 161482 1722 161718
rect 1958 161482 2042 161718
rect 2278 161482 2362 161718
rect 2598 161482 2682 161718
rect 2918 161482 3002 161718
rect 3238 161482 3322 161718
rect 3558 161482 3642 161718
rect 3878 161482 31479 161718
rect 31715 161482 69506 161718
rect 69742 161482 103479 161718
rect 103715 161482 141506 161718
rect 141742 161482 175479 161718
rect 175715 161482 207826 161718
rect 208062 161482 208146 161718
rect 208382 161482 208466 161718
rect 208702 161482 208786 161718
rect 209022 161482 209106 161718
rect 209342 161482 209426 161718
rect 209662 161482 209746 161718
rect 209982 161482 210066 161718
rect 210302 161482 210386 161718
rect 210622 161482 210706 161718
rect 210942 161482 211026 161718
rect 211262 161482 211346 161718
rect 211582 161482 211704 161718
rect 0 161440 211704 161482
rect 168252 153442 186236 153484
rect 168252 153206 168294 153442
rect 168530 153206 185958 153442
rect 186194 153206 186236 153442
rect 168252 153164 186236 153206
rect 0 150518 211704 150560
rect 0 150282 5122 150518
rect 5358 150282 5442 150518
rect 5678 150282 5762 150518
rect 5998 150282 6082 150518
rect 6318 150282 6402 150518
rect 6638 150282 6722 150518
rect 6958 150282 7042 150518
rect 7278 150282 7362 150518
rect 7598 150282 7682 150518
rect 7918 150282 8002 150518
rect 8238 150282 8322 150518
rect 8558 150282 8642 150518
rect 8878 150282 29181 150518
rect 29417 150282 54146 150518
rect 54382 150282 101181 150518
rect 101417 150282 126146 150518
rect 126382 150282 173181 150518
rect 173417 150282 202826 150518
rect 203062 150282 203146 150518
rect 203382 150282 203466 150518
rect 203702 150282 203786 150518
rect 204022 150282 204106 150518
rect 204342 150282 204426 150518
rect 204662 150282 204746 150518
rect 204982 150282 205066 150518
rect 205302 150282 205386 150518
rect 205622 150282 205706 150518
rect 205942 150282 206026 150518
rect 206262 150282 206346 150518
rect 206582 150282 211704 150518
rect 0 150240 211704 150282
rect 26020 140522 44556 140564
rect 26020 140286 26062 140522
rect 26298 140286 44278 140522
rect 44514 140286 44556 140522
rect 26020 140244 44556 140286
rect 0 139318 211704 139360
rect 0 139082 122 139318
rect 358 139082 442 139318
rect 678 139082 762 139318
rect 998 139082 1082 139318
rect 1318 139082 1402 139318
rect 1638 139082 1722 139318
rect 1958 139082 2042 139318
rect 2278 139082 2362 139318
rect 2598 139082 2682 139318
rect 2918 139082 3002 139318
rect 3238 139082 3322 139318
rect 3558 139082 3642 139318
rect 3878 139082 31479 139318
rect 31715 139082 69506 139318
rect 69742 139082 103479 139318
rect 103715 139082 141506 139318
rect 141742 139082 175479 139318
rect 175715 139082 207826 139318
rect 208062 139082 208146 139318
rect 208382 139082 208466 139318
rect 208702 139082 208786 139318
rect 209022 139082 209106 139318
rect 209342 139082 209426 139318
rect 209662 139082 209746 139318
rect 209982 139082 210066 139318
rect 210302 139082 210386 139318
rect 210622 139082 210706 139318
rect 210942 139082 211026 139318
rect 211262 139082 211346 139318
rect 211582 139082 211704 139318
rect 0 139040 211704 139082
rect 0 128118 211704 128160
rect 0 127882 5122 128118
rect 5358 127882 5442 128118
rect 5678 127882 5762 128118
rect 5998 127882 6082 128118
rect 6318 127882 6402 128118
rect 6638 127882 6722 128118
rect 6958 127882 7042 128118
rect 7278 127882 7362 128118
rect 7598 127882 7682 128118
rect 7918 127882 8002 128118
rect 8238 127882 8322 128118
rect 8558 127882 8642 128118
rect 8878 127882 202826 128118
rect 203062 127882 203146 128118
rect 203382 127882 203466 128118
rect 203702 127882 203786 128118
rect 204022 127882 204106 128118
rect 204342 127882 204426 128118
rect 204662 127882 204746 128118
rect 204982 127882 205066 128118
rect 205302 127882 205386 128118
rect 205622 127882 205706 128118
rect 205942 127882 206026 128118
rect 206262 127882 206346 128118
rect 206582 127882 211704 128118
rect 0 127840 211704 127882
rect 0 116918 211704 116960
rect 0 116682 122 116918
rect 358 116682 442 116918
rect 678 116682 762 116918
rect 998 116682 1082 116918
rect 1318 116682 1402 116918
rect 1638 116682 1722 116918
rect 1958 116682 2042 116918
rect 2278 116682 2362 116918
rect 2598 116682 2682 116918
rect 2918 116682 3002 116918
rect 3238 116682 3322 116918
rect 3558 116682 3642 116918
rect 3878 116682 29479 116918
rect 29715 116682 65146 116918
rect 65382 116682 101479 116918
rect 101715 116682 137146 116918
rect 137382 116682 173479 116918
rect 173715 116682 207826 116918
rect 208062 116682 208146 116918
rect 208382 116682 208466 116918
rect 208702 116682 208786 116918
rect 209022 116682 209106 116918
rect 209342 116682 209426 116918
rect 209662 116682 209746 116918
rect 209982 116682 210066 116918
rect 210302 116682 210386 116918
rect 210622 116682 210706 116918
rect 210942 116682 211026 116918
rect 211262 116682 211346 116918
rect 211582 116682 211704 116918
rect 0 116640 211704 116682
rect 19764 106522 46580 106564
rect 19764 106286 19806 106522
rect 20042 106286 46302 106522
rect 46538 106286 46580 106522
rect 19764 106244 46580 106286
rect 0 105718 211704 105760
rect 0 105482 5122 105718
rect 5358 105482 5442 105718
rect 5678 105482 5762 105718
rect 5998 105482 6082 105718
rect 6318 105482 6402 105718
rect 6638 105482 6722 105718
rect 6958 105482 7042 105718
rect 7278 105482 7362 105718
rect 7598 105482 7682 105718
rect 7918 105482 8002 105718
rect 8238 105482 8322 105718
rect 8558 105482 8642 105718
rect 8878 105482 25181 105718
rect 25417 105482 60514 105718
rect 60750 105482 97181 105718
rect 97417 105482 132514 105718
rect 132750 105482 169181 105718
rect 169417 105482 202826 105718
rect 203062 105482 203146 105718
rect 203382 105482 203466 105718
rect 203702 105482 203786 105718
rect 204022 105482 204106 105718
rect 204342 105482 204426 105718
rect 204662 105482 204746 105718
rect 204982 105482 205066 105718
rect 205302 105482 205386 105718
rect 205622 105482 205706 105718
rect 205942 105482 206026 105718
rect 206262 105482 206346 105718
rect 206582 105482 211704 105718
rect 0 105440 211704 105482
rect 0 94518 211704 94560
rect 0 94282 122 94518
rect 358 94282 442 94518
rect 678 94282 762 94518
rect 998 94282 1082 94518
rect 1318 94282 1402 94518
rect 1638 94282 1722 94518
rect 1958 94282 2042 94518
rect 2278 94282 2362 94518
rect 2598 94282 2682 94518
rect 2918 94282 3002 94518
rect 3238 94282 3322 94518
rect 3558 94282 3642 94518
rect 3878 94282 207826 94518
rect 208062 94282 208146 94518
rect 208382 94282 208466 94518
rect 208702 94282 208786 94518
rect 209022 94282 209106 94518
rect 209342 94282 209426 94518
rect 209662 94282 209746 94518
rect 209982 94282 210066 94518
rect 210302 94282 210386 94518
rect 210622 94282 210706 94518
rect 210942 94282 211026 94518
rect 211262 94282 211346 94518
rect 211582 94282 211704 94518
rect 0 94240 211704 94282
rect 48284 92242 85404 92284
rect 48284 92006 48326 92242
rect 48562 92006 85126 92242
rect 85362 92006 85404 92242
rect 48284 91964 85404 92006
rect 0 83318 211704 83360
rect 0 83082 5122 83318
rect 5358 83082 5442 83318
rect 5678 83082 5762 83318
rect 5998 83082 6082 83318
rect 6318 83082 6402 83318
rect 6638 83082 6722 83318
rect 6958 83082 7042 83318
rect 7278 83082 7362 83318
rect 7598 83082 7682 83318
rect 7918 83082 8002 83318
rect 8238 83082 8322 83318
rect 8558 83082 8642 83318
rect 8878 83082 29181 83318
rect 29417 83082 54146 83318
rect 54382 83082 101181 83318
rect 101417 83082 126146 83318
rect 126382 83082 173181 83318
rect 173417 83082 202826 83318
rect 203062 83082 203146 83318
rect 203382 83082 203466 83318
rect 203702 83082 203786 83318
rect 204022 83082 204106 83318
rect 204342 83082 204426 83318
rect 204662 83082 204746 83318
rect 204982 83082 205066 83318
rect 205302 83082 205386 83318
rect 205622 83082 205706 83318
rect 205942 83082 206026 83318
rect 206262 83082 206346 83318
rect 206582 83082 211704 83318
rect 0 83040 211704 83082
rect 0 72118 211704 72160
rect 0 71882 122 72118
rect 358 71882 442 72118
rect 678 71882 762 72118
rect 998 71882 1082 72118
rect 1318 71882 1402 72118
rect 1638 71882 1722 72118
rect 1958 71882 2042 72118
rect 2278 71882 2362 72118
rect 2598 71882 2682 72118
rect 2918 71882 3002 72118
rect 3238 71882 3322 72118
rect 3558 71882 3642 72118
rect 3878 71882 31479 72118
rect 31715 71882 69506 72118
rect 69742 71882 103479 72118
rect 103715 71882 141506 72118
rect 141742 71882 175479 72118
rect 175715 71882 207826 72118
rect 208062 71882 208146 72118
rect 208382 71882 208466 72118
rect 208702 71882 208786 72118
rect 209022 71882 209106 72118
rect 209342 71882 209426 72118
rect 209662 71882 209746 72118
rect 209982 71882 210066 72118
rect 210302 71882 210386 72118
rect 210622 71882 210706 72118
rect 210942 71882 211026 72118
rect 211262 71882 211346 72118
rect 211582 71882 211704 72118
rect 0 71840 211704 71882
rect 168252 70482 186236 70524
rect 168252 70246 168294 70482
rect 168530 70246 185958 70482
rect 186194 70246 186236 70482
rect 168252 70204 186236 70246
rect 0 60918 211704 60960
rect 0 60682 5122 60918
rect 5358 60682 5442 60918
rect 5678 60682 5762 60918
rect 5998 60682 6082 60918
rect 6318 60682 6402 60918
rect 6638 60682 6722 60918
rect 6958 60682 7042 60918
rect 7278 60682 7362 60918
rect 7598 60682 7682 60918
rect 7918 60682 8002 60918
rect 8238 60682 8322 60918
rect 8558 60682 8642 60918
rect 8878 60682 29181 60918
rect 29417 60682 54146 60918
rect 54382 60682 101181 60918
rect 101417 60682 126146 60918
rect 126382 60682 173181 60918
rect 173417 60682 202826 60918
rect 203062 60682 203146 60918
rect 203382 60682 203466 60918
rect 203702 60682 203786 60918
rect 204022 60682 204106 60918
rect 204342 60682 204426 60918
rect 204662 60682 204746 60918
rect 204982 60682 205066 60918
rect 205302 60682 205386 60918
rect 205622 60682 205706 60918
rect 205942 60682 206026 60918
rect 206262 60682 206346 60918
rect 206582 60682 211704 60918
rect 0 60640 211704 60682
rect 121884 59602 128460 59644
rect 121884 59366 121926 59602
rect 122162 59366 128460 59602
rect 121884 59324 128460 59366
rect 128140 58284 128460 59324
rect 172668 59324 182372 59644
rect 129060 58922 136924 58964
rect 129060 58686 136646 58922
rect 136882 58686 136924 58922
rect 129060 58644 136924 58686
rect 129060 58284 129380 58644
rect 172668 58284 172988 59324
rect 26020 58242 44556 58284
rect 26020 58006 26062 58242
rect 26298 58006 44278 58242
rect 44514 58006 44556 58242
rect 26020 57964 44556 58006
rect 128140 57964 129380 58284
rect 172484 57964 172988 58284
rect 172484 57604 172804 57964
rect 182052 57604 182372 59324
rect 153348 57284 157716 57604
rect 171012 57562 172804 57604
rect 171012 57326 171054 57562
rect 171290 57326 172804 57562
rect 171012 57284 172804 57326
rect 181868 57284 182372 57604
rect 185732 57562 186052 57604
rect 185732 57326 185774 57562
rect 186010 57326 186052 57562
rect 153348 56924 153668 57284
rect 143596 56604 153668 56924
rect 157396 56924 157716 57284
rect 181868 56924 182188 57284
rect 185732 56924 186052 57326
rect 157396 56882 161948 56924
rect 157396 56646 161670 56882
rect 161906 56646 161948 56882
rect 157396 56604 161948 56646
rect 181868 56604 186052 56924
rect 143596 56244 143916 56604
rect 136604 56202 143916 56244
rect 136604 55966 136646 56202
rect 136882 55966 143916 56202
rect 136604 55924 143916 55966
rect 0 49718 211704 49760
rect 0 49482 122 49718
rect 358 49482 442 49718
rect 678 49482 762 49718
rect 998 49482 1082 49718
rect 1318 49482 1402 49718
rect 1638 49482 1722 49718
rect 1958 49482 2042 49718
rect 2278 49482 2362 49718
rect 2598 49482 2682 49718
rect 2918 49482 3002 49718
rect 3238 49482 3322 49718
rect 3558 49482 3642 49718
rect 3878 49482 207826 49718
rect 208062 49482 208146 49718
rect 208382 49482 208466 49718
rect 208702 49482 208786 49718
rect 209022 49482 209106 49718
rect 209342 49482 209426 49718
rect 209662 49482 209746 49718
rect 209982 49482 210066 49718
rect 210302 49482 210386 49718
rect 210622 49482 210706 49718
rect 210942 49482 211026 49718
rect 211262 49482 211346 49718
rect 211582 49482 211704 49718
rect 0 49440 211704 49482
rect 0 38518 211704 38560
rect 0 38282 5122 38518
rect 5358 38282 5442 38518
rect 5678 38282 5762 38518
rect 5998 38282 6082 38518
rect 6318 38282 6402 38518
rect 6638 38282 6722 38518
rect 6958 38282 7042 38518
rect 7278 38282 7362 38518
rect 7598 38282 7682 38518
rect 7918 38282 8002 38518
rect 8238 38282 8322 38518
rect 8558 38282 8642 38518
rect 8878 38282 25181 38518
rect 25417 38282 60514 38518
rect 60750 38282 97181 38518
rect 97417 38282 132514 38518
rect 132750 38282 169181 38518
rect 169417 38282 202826 38518
rect 203062 38282 203146 38518
rect 203382 38282 203466 38518
rect 203702 38282 203786 38518
rect 204022 38282 204106 38518
rect 204342 38282 204426 38518
rect 204662 38282 204746 38518
rect 204982 38282 205066 38518
rect 205302 38282 205386 38518
rect 205622 38282 205706 38518
rect 205942 38282 206026 38518
rect 206262 38282 206346 38518
rect 206582 38282 211704 38518
rect 0 38240 211704 38282
rect 0 27318 211704 27360
rect 0 27082 122 27318
rect 358 27082 442 27318
rect 678 27082 762 27318
rect 998 27082 1082 27318
rect 1318 27082 1402 27318
rect 1638 27082 1722 27318
rect 1958 27082 2042 27318
rect 2278 27082 2362 27318
rect 2598 27082 2682 27318
rect 2918 27082 3002 27318
rect 3238 27082 3322 27318
rect 3558 27082 3642 27318
rect 3878 27082 29479 27318
rect 29715 27082 65146 27318
rect 65382 27082 101479 27318
rect 101715 27082 137146 27318
rect 137382 27082 173479 27318
rect 173715 27082 207826 27318
rect 208062 27082 208146 27318
rect 208382 27082 208466 27318
rect 208702 27082 208786 27318
rect 209022 27082 209106 27318
rect 209342 27082 209426 27318
rect 209662 27082 209746 27318
rect 209982 27082 210066 27318
rect 210302 27082 210386 27318
rect 210622 27082 210706 27318
rect 210942 27082 211026 27318
rect 211262 27082 211346 27318
rect 211582 27082 211704 27318
rect 0 27040 211704 27082
rect 83428 22202 88716 22244
rect 83428 21966 83470 22202
rect 83706 21966 88438 22202
rect 88674 21966 88716 22202
rect 83428 21924 88716 21966
rect 0 16118 211704 16160
rect 0 15882 5122 16118
rect 5358 15882 5442 16118
rect 5678 15882 5762 16118
rect 5998 15882 6082 16118
rect 6318 15882 6402 16118
rect 6638 15882 6722 16118
rect 6958 15882 7042 16118
rect 7278 15882 7362 16118
rect 7598 15882 7682 16118
rect 7918 15882 8002 16118
rect 8238 15882 8322 16118
rect 8558 15882 8642 16118
rect 8878 15882 202826 16118
rect 203062 15882 203146 16118
rect 203382 15882 203466 16118
rect 203702 15882 203786 16118
rect 204022 15882 204106 16118
rect 204342 15882 204426 16118
rect 204662 15882 204746 16118
rect 204982 15882 205066 16118
rect 205302 15882 205386 16118
rect 205622 15882 205706 16118
rect 205942 15882 206026 16118
rect 206262 15882 206346 16118
rect 206582 15882 211704 16118
rect 0 15840 211704 15882
rect 5000 8878 206704 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 202826 8878
rect 203062 8642 203146 8878
rect 203382 8642 203466 8878
rect 203702 8642 203786 8878
rect 204022 8642 204106 8878
rect 204342 8642 204426 8878
rect 204662 8642 204746 8878
rect 204982 8642 205066 8878
rect 205302 8642 205386 8878
rect 205622 8642 205706 8878
rect 205942 8642 206026 8878
rect 206262 8642 206346 8878
rect 206582 8642 206704 8878
rect 5000 8558 206704 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 202826 8558
rect 203062 8322 203146 8558
rect 203382 8322 203466 8558
rect 203702 8322 203786 8558
rect 204022 8322 204106 8558
rect 204342 8322 204426 8558
rect 204662 8322 204746 8558
rect 204982 8322 205066 8558
rect 205302 8322 205386 8558
rect 205622 8322 205706 8558
rect 205942 8322 206026 8558
rect 206262 8322 206346 8558
rect 206582 8322 206704 8558
rect 5000 8238 206704 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 202826 8238
rect 203062 8002 203146 8238
rect 203382 8002 203466 8238
rect 203702 8002 203786 8238
rect 204022 8002 204106 8238
rect 204342 8002 204426 8238
rect 204662 8002 204746 8238
rect 204982 8002 205066 8238
rect 205302 8002 205386 8238
rect 205622 8002 205706 8238
rect 205942 8002 206026 8238
rect 206262 8002 206346 8238
rect 206582 8002 206704 8238
rect 5000 7918 206704 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 202826 7918
rect 203062 7682 203146 7918
rect 203382 7682 203466 7918
rect 203702 7682 203786 7918
rect 204022 7682 204106 7918
rect 204342 7682 204426 7918
rect 204662 7682 204746 7918
rect 204982 7682 205066 7918
rect 205302 7682 205386 7918
rect 205622 7682 205706 7918
rect 205942 7682 206026 7918
rect 206262 7682 206346 7918
rect 206582 7682 206704 7918
rect 5000 7598 206704 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 202826 7598
rect 203062 7362 203146 7598
rect 203382 7362 203466 7598
rect 203702 7362 203786 7598
rect 204022 7362 204106 7598
rect 204342 7362 204426 7598
rect 204662 7362 204746 7598
rect 204982 7362 205066 7598
rect 205302 7362 205386 7598
rect 205622 7362 205706 7598
rect 205942 7362 206026 7598
rect 206262 7362 206346 7598
rect 206582 7362 206704 7598
rect 5000 7278 206704 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 202826 7278
rect 203062 7042 203146 7278
rect 203382 7042 203466 7278
rect 203702 7042 203786 7278
rect 204022 7042 204106 7278
rect 204342 7042 204426 7278
rect 204662 7042 204746 7278
rect 204982 7042 205066 7278
rect 205302 7042 205386 7278
rect 205622 7042 205706 7278
rect 205942 7042 206026 7278
rect 206262 7042 206346 7278
rect 206582 7042 206704 7278
rect 5000 6958 206704 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 202826 6958
rect 203062 6722 203146 6958
rect 203382 6722 203466 6958
rect 203702 6722 203786 6958
rect 204022 6722 204106 6958
rect 204342 6722 204426 6958
rect 204662 6722 204746 6958
rect 204982 6722 205066 6958
rect 205302 6722 205386 6958
rect 205622 6722 205706 6958
rect 205942 6722 206026 6958
rect 206262 6722 206346 6958
rect 206582 6722 206704 6958
rect 5000 6638 206704 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 202826 6638
rect 203062 6402 203146 6638
rect 203382 6402 203466 6638
rect 203702 6402 203786 6638
rect 204022 6402 204106 6638
rect 204342 6402 204426 6638
rect 204662 6402 204746 6638
rect 204982 6402 205066 6638
rect 205302 6402 205386 6638
rect 205622 6402 205706 6638
rect 205942 6402 206026 6638
rect 206262 6402 206346 6638
rect 206582 6402 206704 6638
rect 5000 6318 206704 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 202826 6318
rect 203062 6082 203146 6318
rect 203382 6082 203466 6318
rect 203702 6082 203786 6318
rect 204022 6082 204106 6318
rect 204342 6082 204426 6318
rect 204662 6082 204746 6318
rect 204982 6082 205066 6318
rect 205302 6082 205386 6318
rect 205622 6082 205706 6318
rect 205942 6082 206026 6318
rect 206262 6082 206346 6318
rect 206582 6082 206704 6318
rect 5000 5998 206704 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 202826 5998
rect 203062 5762 203146 5998
rect 203382 5762 203466 5998
rect 203702 5762 203786 5998
rect 204022 5762 204106 5998
rect 204342 5762 204426 5998
rect 204662 5762 204746 5998
rect 204982 5762 205066 5998
rect 205302 5762 205386 5998
rect 205622 5762 205706 5998
rect 205942 5762 206026 5998
rect 206262 5762 206346 5998
rect 206582 5762 206704 5998
rect 5000 5678 206704 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 202826 5678
rect 203062 5442 203146 5678
rect 203382 5442 203466 5678
rect 203702 5442 203786 5678
rect 204022 5442 204106 5678
rect 204342 5442 204426 5678
rect 204662 5442 204746 5678
rect 204982 5442 205066 5678
rect 205302 5442 205386 5678
rect 205622 5442 205706 5678
rect 205942 5442 206026 5678
rect 206262 5442 206346 5678
rect 206582 5442 206704 5678
rect 5000 5358 206704 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 202826 5358
rect 203062 5122 203146 5358
rect 203382 5122 203466 5358
rect 203702 5122 203786 5358
rect 204022 5122 204106 5358
rect 204342 5122 204426 5358
rect 204662 5122 204746 5358
rect 204982 5122 205066 5358
rect 205302 5122 205386 5358
rect 205622 5122 205706 5358
rect 205942 5122 206026 5358
rect 206262 5122 206346 5358
rect 206582 5122 206704 5358
rect 5000 5000 206704 5122
rect 0 3878 211704 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 207826 3878
rect 208062 3642 208146 3878
rect 208382 3642 208466 3878
rect 208702 3642 208786 3878
rect 209022 3642 209106 3878
rect 209342 3642 209426 3878
rect 209662 3642 209746 3878
rect 209982 3642 210066 3878
rect 210302 3642 210386 3878
rect 210622 3642 210706 3878
rect 210942 3642 211026 3878
rect 211262 3642 211346 3878
rect 211582 3642 211704 3878
rect 0 3558 211704 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 207826 3558
rect 208062 3322 208146 3558
rect 208382 3322 208466 3558
rect 208702 3322 208786 3558
rect 209022 3322 209106 3558
rect 209342 3322 209426 3558
rect 209662 3322 209746 3558
rect 209982 3322 210066 3558
rect 210302 3322 210386 3558
rect 210622 3322 210706 3558
rect 210942 3322 211026 3558
rect 211262 3322 211346 3558
rect 211582 3322 211704 3558
rect 0 3238 211704 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 207826 3238
rect 208062 3002 208146 3238
rect 208382 3002 208466 3238
rect 208702 3002 208786 3238
rect 209022 3002 209106 3238
rect 209342 3002 209426 3238
rect 209662 3002 209746 3238
rect 209982 3002 210066 3238
rect 210302 3002 210386 3238
rect 210622 3002 210706 3238
rect 210942 3002 211026 3238
rect 211262 3002 211346 3238
rect 211582 3002 211704 3238
rect 0 2918 211704 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 207826 2918
rect 208062 2682 208146 2918
rect 208382 2682 208466 2918
rect 208702 2682 208786 2918
rect 209022 2682 209106 2918
rect 209342 2682 209426 2918
rect 209662 2682 209746 2918
rect 209982 2682 210066 2918
rect 210302 2682 210386 2918
rect 210622 2682 210706 2918
rect 210942 2682 211026 2918
rect 211262 2682 211346 2918
rect 211582 2682 211704 2918
rect 0 2598 211704 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 207826 2598
rect 208062 2362 208146 2598
rect 208382 2362 208466 2598
rect 208702 2362 208786 2598
rect 209022 2362 209106 2598
rect 209342 2362 209426 2598
rect 209662 2362 209746 2598
rect 209982 2362 210066 2598
rect 210302 2362 210386 2598
rect 210622 2362 210706 2598
rect 210942 2362 211026 2598
rect 211262 2362 211346 2598
rect 211582 2362 211704 2598
rect 0 2278 211704 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 207826 2278
rect 208062 2042 208146 2278
rect 208382 2042 208466 2278
rect 208702 2042 208786 2278
rect 209022 2042 209106 2278
rect 209342 2042 209426 2278
rect 209662 2042 209746 2278
rect 209982 2042 210066 2278
rect 210302 2042 210386 2278
rect 210622 2042 210706 2278
rect 210942 2042 211026 2278
rect 211262 2042 211346 2278
rect 211582 2042 211704 2278
rect 0 1958 211704 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 207826 1958
rect 208062 1722 208146 1958
rect 208382 1722 208466 1958
rect 208702 1722 208786 1958
rect 209022 1722 209106 1958
rect 209342 1722 209426 1958
rect 209662 1722 209746 1958
rect 209982 1722 210066 1958
rect 210302 1722 210386 1958
rect 210622 1722 210706 1958
rect 210942 1722 211026 1958
rect 211262 1722 211346 1958
rect 211582 1722 211704 1958
rect 0 1638 211704 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 207826 1638
rect 208062 1402 208146 1638
rect 208382 1402 208466 1638
rect 208702 1402 208786 1638
rect 209022 1402 209106 1638
rect 209342 1402 209426 1638
rect 209662 1402 209746 1638
rect 209982 1402 210066 1638
rect 210302 1402 210386 1638
rect 210622 1402 210706 1638
rect 210942 1402 211026 1638
rect 211262 1402 211346 1638
rect 211582 1402 211704 1638
rect 0 1318 211704 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 207826 1318
rect 208062 1082 208146 1318
rect 208382 1082 208466 1318
rect 208702 1082 208786 1318
rect 209022 1082 209106 1318
rect 209342 1082 209426 1318
rect 209662 1082 209746 1318
rect 209982 1082 210066 1318
rect 210302 1082 210386 1318
rect 210622 1082 210706 1318
rect 210942 1082 211026 1318
rect 211262 1082 211346 1318
rect 211582 1082 211704 1318
rect 0 998 211704 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 207826 998
rect 208062 762 208146 998
rect 208382 762 208466 998
rect 208702 762 208786 998
rect 209022 762 209106 998
rect 209342 762 209426 998
rect 209662 762 209746 998
rect 209982 762 210066 998
rect 210302 762 210386 998
rect 210622 762 210706 998
rect 210942 762 211026 998
rect 211262 762 211346 998
rect 211582 762 211704 998
rect 0 678 211704 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 207826 678
rect 208062 442 208146 678
rect 208382 442 208466 678
rect 208702 442 208786 678
rect 209022 442 209106 678
rect 209342 442 209426 678
rect 209662 442 209746 678
rect 209982 442 210066 678
rect 210302 442 210386 678
rect 210622 442 210706 678
rect 210942 442 211026 678
rect 211262 442 211346 678
rect 211582 442 211704 678
rect 0 358 211704 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 207826 358
rect 208062 122 208146 358
rect 208382 122 208466 358
rect 208702 122 208786 358
rect 209022 122 209106 358
rect 209342 122 209426 358
rect 209662 122 209746 358
rect 209982 122 210066 358
rect 210302 122 210386 358
rect 210622 122 210706 358
rect 210942 122 211026 358
rect 211262 122 211346 358
rect 211582 122 211704 358
rect 0 0 211704 122
use grid_clb  grid_clb_1__1_
timestamp 1606150568
transform 1 0 49896 0 1 53824
box 0 0 40000 40000
use sb_0__0_  sb_0__0_
timestamp 1606150568
transform 1 0 19896 0 1 18824
box 0 0 28000 27720
use cby_0__1_  cby_0__1_
timestamp 1606150568
transform 1 0 25896 0 1 53824
box 0 0 16000 40000
use cbx_1__0_  cbx_1__0_
timestamp 1606150568
transform 1 0 54896 0 1 20824
box 0 0 30000 24000
use sb_1__0_  sb_1__0_
timestamp 1606150568
transform 1 0 91896 0 1 18824
box 0 0 28000 28000
use cby_1__1_  cby_1__1_
timestamp 1606150568
transform 1 0 97896 0 1 53824
box 0 0 16000 40000
use grid_clb  grid_clb_2__1_
timestamp 1606150568
transform 1 0 121896 0 1 53824
box 0 0 40000 40000
use cbx_1__0_  cbx_2__0_
timestamp 1606150568
transform 1 0 126896 0 1 20824
box 0 0 30000 24000
use sb_2__0_  sb_2__0_
timestamp 1606150568
transform 1 0 163896 0 1 18824
box 0 0 27678 28000
use cby_2__1_  cby_2__1_
timestamp 1606150568
transform 1 0 169896 0 1 53824
box 0 0 16000 40000
use grid_clb  grid_clb_1__2_
timestamp 1606150568
transform 1 0 49896 0 1 135824
box 0 0 40000 40000
use sb_0__1_  sb_0__1_
timestamp 1606150568
transform 1 0 19896 0 1 100824
box 0 0 28000 28000
use cby_0__1_  cby_0__2_
timestamp 1606150568
transform 1 0 25896 0 1 135824
box 0 0 16000 40000
use cbx_1__1_  cbx_1__1_
timestamp 1606150568
transform 1 0 54896 0 1 102824
box 0 0 30000 24000
use sky130_fd_sc_hd__conb_1  _5_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606150568
transform 1 0 84968 0 -1 107288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _6_
timestamp 1606150568
transform 1 0 77884 0 1 134488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _8_
timestamp 1606150568
transform 1 0 90856 0 -1 105112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _9_
timestamp 1606150568
transform 1 0 91224 0 1 133400
box -38 -48 314 592
use sb_1__1_  sb_1__1_
timestamp 1606150568
transform 1 0 91896 0 1 100824
box 0 0 28000 28000
use cby_1__1_  cby_1__2_
timestamp 1606150568
transform 1 0 97896 0 1 135824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1606150568
transform 1 0 121896 0 1 135824
box 0 0 40000 40000
use cbx_1__1_  cbx_2__1_
timestamp 1606150568
transform 1 0 126896 0 1 102824
box 0 0 30000 24000
use sb_2__1_  sb_2__1_
timestamp 1606150568
transform 1 0 163896 0 1 100824
box 0 0 28000 28000
use cby_2__1_  cby_2__2_
timestamp 1606150568
transform 1 0 169896 0 1 135824
box 0 0 16000 40000
use sky130_fd_sc_hd__conb_1  _7_
timestamp 1606150568
transform 1 0 91500 0 1 141016
box -38 -48 314 592
use sb_0__2_  sb_0__2_
timestamp 1606150568
transform 1 0 19895 0 1 182824
box 1 0 27712 28000
use cbx_1__2_  cbx_1__2_
timestamp 1606150568
transform 1 0 54896 0 1 184824
box 0 0 30000 24000
use sb_1__2_  sb_1__2_
timestamp 1606150568
transform 1 0 91896 0 1 182824
box 0 0 28000 28000
use cbx_1__2_  cbx_2__2_
timestamp 1606150568
transform 1 0 126896 0 1 184824
box 0 0 30000 24000
use sb_2__2_  sb_2__2_
timestamp 1606150568
transform 1 0 163896 0 1 182824
box 0 0 28000 27736
<< labels >>
rlabel metal3 s 9896 19304 10376 19424 6 Test_en
port 0 nsew default input
rlabel metal3 s 201416 20528 201896 20648 6 ccff_head
port 1 nsew default input
rlabel metal3 s 9896 188896 10376 189016 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 9896 40384 10376 40504 6 clk
port 3 nsew default input
rlabel metal2 s 25830 220344 25886 220824 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
port 4 nsew default tristate
rlabel metal2 s 108446 8824 108502 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
port 5 nsew default tristate
rlabel metal2 s 113782 8824 113838 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
port 6 nsew default tristate
rlabel metal2 s 119118 8824 119174 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
port 7 nsew default tristate
rlabel metal2 s 124454 8824 124510 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
port 8 nsew default tristate
rlabel metal2 s 129790 8824 129846 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
port 9 nsew default tristate
rlabel metal2 s 135126 8824 135182 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
port 10 nsew default tristate
rlabel metal3 s 9896 61600 10376 61720 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
port 11 nsew default tristate
rlabel metal3 s 9896 125248 10376 125368 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
port 12 nsew default tristate
rlabel metal2 s 57754 220344 57810 220824 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
port 13 nsew default tristate
rlabel metal3 s 201416 91112 201896 91232 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
port 14 nsew default tristate
rlabel metal3 s 201416 114640 201896 114760 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
port 15 nsew default tristate
rlabel metal2 s 12490 8824 12546 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
port 16 nsew default tristate
rlabel metal2 s 17734 8824 17790 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
port 17 nsew default tristate
rlabel metal2 s 23070 8824 23126 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
port 18 nsew default tristate
rlabel metal2 s 28406 8824 28462 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
port 19 nsew default tristate
rlabel metal2 s 33742 8824 33798 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
port 20 nsew default tristate
rlabel metal2 s 39078 8824 39134 9304 6 gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
port 21 nsew default tristate
rlabel metal2 s 89770 220344 89826 220824 6 gfpga_pad_EMBEDDED_IO_SOC_IN[0]
port 22 nsew default input
rlabel metal2 s 140462 8824 140518 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[10]
port 23 nsew default input
rlabel metal2 s 145798 8824 145854 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[11]
port 24 nsew default input
rlabel metal2 s 151134 8824 151190 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[12]
port 25 nsew default input
rlabel metal2 s 156470 8824 156526 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[13]
port 26 nsew default input
rlabel metal2 s 161806 8824 161862 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[14]
port 27 nsew default input
rlabel metal2 s 167142 8824 167198 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[15]
port 28 nsew default input
rlabel metal3 s 9896 82816 10376 82936 6 gfpga_pad_EMBEDDED_IO_SOC_IN[16]
port 29 nsew default input
rlabel metal3 s 9896 146464 10376 146584 6 gfpga_pad_EMBEDDED_IO_SOC_IN[17]
port 30 nsew default input
rlabel metal2 s 121786 220344 121842 220824 6 gfpga_pad_EMBEDDED_IO_SOC_IN[1]
port 31 nsew default input
rlabel metal3 s 201416 138304 201896 138424 6 gfpga_pad_EMBEDDED_IO_SOC_IN[2]
port 32 nsew default input
rlabel metal3 s 201416 161832 201896 161952 6 gfpga_pad_EMBEDDED_IO_SOC_IN[3]
port 33 nsew default input
rlabel metal2 s 44414 8824 44470 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[4]
port 34 nsew default input
rlabel metal2 s 49750 8824 49806 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[5]
port 35 nsew default input
rlabel metal2 s 55086 8824 55142 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[6]
port 36 nsew default input
rlabel metal2 s 60422 8824 60478 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[7]
port 37 nsew default input
rlabel metal2 s 65758 8824 65814 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[8]
port 38 nsew default input
rlabel metal2 s 71094 8824 71150 9304 6 gfpga_pad_EMBEDDED_IO_SOC_IN[9]
port 39 nsew default input
rlabel metal2 s 153802 220344 153858 220824 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
port 40 nsew default tristate
rlabel metal2 s 172478 8824 172534 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
port 41 nsew default tristate
rlabel metal2 s 177814 8824 177870 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
port 42 nsew default tristate
rlabel metal2 s 183150 8824 183206 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
port 43 nsew default tristate
rlabel metal2 s 188486 8824 188542 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
port 44 nsew default tristate
rlabel metal2 s 193822 8824 193878 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
port 45 nsew default tristate
rlabel metal2 s 199158 8824 199214 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
port 46 nsew default tristate
rlabel metal3 s 9896 104032 10376 104152 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
port 47 nsew default tristate
rlabel metal3 s 9896 167680 10376 167800 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
port 48 nsew default tristate
rlabel metal2 s 185818 220344 185874 220824 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
port 49 nsew default tristate
rlabel metal3 s 201416 185360 201896 185480 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
port 50 nsew default tristate
rlabel metal3 s 201416 208888 201896 209008 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
port 51 nsew default tristate
rlabel metal2 s 76430 8824 76486 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
port 52 nsew default tristate
rlabel metal2 s 81766 8824 81822 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
port 53 nsew default tristate
rlabel metal2 s 87102 8824 87158 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
port 54 nsew default tristate
rlabel metal2 s 92438 8824 92494 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
port 55 nsew default tristate
rlabel metal2 s 97774 8824 97830 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
port 56 nsew default tristate
rlabel metal2 s 103110 8824 103166 9304 6 gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
port 57 nsew default tristate
rlabel metal3 s 201416 67584 201896 67704 6 prog_clk
port 58 nsew default input
rlabel metal3 s 201416 44056 201896 44176 6 sc_head
port 59 nsew default input
rlabel metal3 s 9896 210112 10376 210232 6 sc_tail
port 60 nsew default tristate
rlabel metal5 s 5000 5000 206704 9000 8 VPWR
port 61 nsew default input
rlabel metal5 s 0 0 211704 4000 8 VGND
port 62 nsew default input
<< properties >>
string FIXED_BBOX 0 0 211704 229264
<< end >>
