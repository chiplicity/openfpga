magic
tech EFS8A
magscale 1 2
timestamp 1604338020
<< viali >>
rect 16727 11849 16761 11883
rect 14933 11645 14967 11679
rect 16656 11645 16690 11679
rect 15117 11509 15151 11543
rect 15577 11509 15611 11543
rect 17141 11509 17175 11543
rect 16589 9469 16623 9503
rect 17141 9469 17175 9503
rect 16773 9333 16807 9367
rect 16282 5797 16316 5831
rect 16037 5661 16071 5695
rect 17417 5593 17451 5627
rect 16405 5321 16439 5355
rect 16129 5253 16163 5287
rect 20085 2601 20119 2635
rect 19901 2465 19935 2499
rect 20545 2465 20579 2499
rect 21557 2465 21591 2499
rect 22201 2329 22235 2363
rect 21741 2261 21775 2295
<< metal1 >>
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 16758 11889 16764 11892
rect 16715 11883 16764 11889
rect 16715 11849 16727 11883
rect 16761 11849 16764 11883
rect 16715 11843 16764 11849
rect 16758 11840 16764 11843
rect 16816 11840 16822 11892
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 16644 11679 16702 11685
rect 14967 11648 15608 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 15102 11540 15108 11552
rect 15063 11512 15108 11540
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15580 11549 15608 11648
rect 16644 11645 16656 11679
rect 16690 11676 16702 11679
rect 16690 11645 16712 11676
rect 16644 11639 16712 11645
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 16684 11540 16712 11639
rect 17129 11543 17187 11549
rect 17129 11540 17141 11543
rect 15611 11512 17141 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 17129 11509 17141 11512
rect 17175 11540 17187 11543
rect 17402 11540 17408 11552
rect 17175 11512 17408 11540
rect 17175 11509 17187 11512
rect 17129 11503 17187 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 16632 9472 17141 9500
rect 16632 9460 16638 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 16758 9364 16764 9376
rect 16719 9336 16764 9364
rect 16758 9324 16764 9336
rect 16816 9324 16822 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 16206 5788 16212 5840
rect 16264 5837 16270 5840
rect 16264 5831 16328 5837
rect 16264 5797 16282 5831
rect 16316 5797 16328 5831
rect 16264 5791 16328 5797
rect 16264 5788 16270 5791
rect 16022 5692 16028 5704
rect 15983 5664 16028 5692
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 17402 5624 17408 5636
rect 17363 5596 17408 5624
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 16080 5324 16405 5352
rect 16080 5312 16086 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 16393 5315 16451 5321
rect 16117 5287 16175 5293
rect 16117 5253 16129 5287
rect 16163 5284 16175 5287
rect 16206 5284 16212 5296
rect 16163 5256 16212 5284
rect 16163 5253 16175 5256
rect 16117 5247 16175 5253
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 20070 2632 20076 2644
rect 20031 2604 20076 2632
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 19935 2468 20545 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20533 2465 20545 2468
rect 20579 2496 20591 2499
rect 21545 2499 21603 2505
rect 21545 2496 21557 2499
rect 20579 2468 21557 2496
rect 20579 2465 20591 2468
rect 20533 2459 20591 2465
rect 21545 2465 21557 2468
rect 21591 2496 21603 2499
rect 21591 2468 22232 2496
rect 21591 2465 21603 2468
rect 21545 2459 21603 2465
rect 22204 2372 22232 2468
rect 22186 2360 22192 2372
rect 22147 2332 22192 2360
rect 22186 2320 22192 2332
rect 22244 2320 22250 2372
rect 21726 2292 21732 2304
rect 21687 2264 21732 2292
rect 21726 2252 21732 2264
rect 21784 2252 21790 2304
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 16764 11840 16816 11892
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 17408 11500 17460 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 16580 9503 16632 9512
rect 16580 9469 16589 9503
rect 16589 9469 16623 9503
rect 16623 9469 16632 9503
rect 16580 9460 16632 9469
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 16212 5788 16264 5840
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 16028 5312 16080 5364
rect 16212 5244 16264 5296
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 20076 2635 20128 2644
rect 20076 2601 20085 2635
rect 20085 2601 20119 2635
rect 20119 2601 20128 2635
rect 20076 2592 20128 2601
rect 22192 2363 22244 2372
rect 22192 2329 22201 2363
rect 22201 2329 22235 2363
rect 22235 2329 22244 2363
rect 22192 2320 22244 2329
rect 21732 2295 21784 2304
rect 21732 2261 21741 2295
rect 21741 2261 21775 2295
rect 21775 2261 21784 2295
rect 21732 2252 21784 2261
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
<< metal2 >>
rect 6642 15520 6698 16000
rect 19982 15520 20038 16000
rect 33322 15520 33378 16000
rect 6656 11665 6684 15520
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 19996 11937 20024 15520
rect 33336 15450 33364 15520
rect 33152 15422 33364 15450
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 16762 11928 16818 11937
rect 16762 11863 16764 11872
rect 16816 11863 16818 11872
rect 19982 11928 20038 11937
rect 20956 11920 21252 11940
rect 19982 11863 20038 11872
rect 16764 11834 16816 11840
rect 6642 11656 6698 11665
rect 6642 11591 6698 11600
rect 15106 11656 15162 11665
rect 15106 11591 15162 11600
rect 15120 11558 15148 11591
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16762 9480 16818 9489
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 16592 9081 16620 9454
rect 16762 9415 16818 9424
rect 16776 9382 16804 9415
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 4986 9072 5042 9081
rect 4986 9007 5042 9016
rect 16578 9072 16634 9081
rect 16578 9007 16634 9016
rect 2962 8120 3018 8129
rect 2962 8055 3018 8064
rect 2976 5817 3004 8055
rect 2962 5808 3018 5817
rect 2962 5743 3018 5752
rect 5000 480 5028 9007
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 16212 5840 16264 5846
rect 16210 5808 16212 5817
rect 16264 5808 16266 5817
rect 16210 5743 16266 5752
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 16040 5370 16068 5646
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16040 5137 16068 5306
rect 16224 5302 16252 5743
rect 17420 5681 17448 11494
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 33152 6882 33180 15422
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 34702 12064 34758 12073
rect 34289 11996 34585 12016
rect 34702 11999 34758 12008
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34716 9489 34744 11999
rect 34702 9480 34758 9489
rect 34702 9415 34758 9424
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 33152 6854 33364 6882
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 17406 5672 17462 5681
rect 17406 5607 17408 5616
rect 17460 5607 17462 5616
rect 17408 5578 17460 5584
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16026 5128 16082 5137
rect 16026 5063 16082 5072
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 14922 2952 14978 2961
rect 14922 2887 14978 2896
rect 20074 2952 20130 2961
rect 20074 2887 20130 2896
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 14936 480 14964 2887
rect 20088 2650 20116 2887
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 33336 2417 33364 6854
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34610 5672 34666 5681
rect 34610 5607 34666 5616
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 34624 4049 34652 5607
rect 34978 5128 35034 5137
rect 34978 5063 35034 5072
rect 34610 4040 34666 4049
rect 34610 3975 34666 3984
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 22190 2408 22246 2417
rect 22190 2343 22192 2352
rect 22244 2343 22246 2352
rect 33322 2408 33378 2417
rect 33322 2343 33378 2352
rect 22192 2314 22244 2320
rect 21732 2304 21784 2310
rect 21732 2246 21784 2252
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 21744 1465 21772 2246
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 21730 1456 21786 1465
rect 21730 1391 21786 1400
rect 24950 1456 25006 1465
rect 24950 1391 25006 1400
rect 24964 480 24992 1391
rect 34992 480 35020 5063
rect 4986 0 5042 480
rect 14922 0 14978 480
rect 24950 0 25006 480
rect 34978 0 35034 480
<< via2 >>
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 16762 11892 16818 11928
rect 16762 11872 16764 11892
rect 16764 11872 16816 11892
rect 16816 11872 16818 11892
rect 19982 11872 20038 11928
rect 6642 11600 6698 11656
rect 15106 11600 15162 11656
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 16762 9424 16818 9480
rect 4986 9016 5042 9072
rect 16578 9016 16634 9072
rect 2962 8064 3018 8120
rect 2962 5752 3018 5808
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 16210 5788 16212 5808
rect 16212 5788 16264 5808
rect 16264 5788 16266 5808
rect 16210 5752 16266 5788
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34702 12008 34758 12064
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34702 9424 34758 9480
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 17406 5636 17462 5672
rect 17406 5616 17408 5636
rect 17408 5616 17460 5636
rect 17460 5616 17462 5636
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 16026 5072 16082 5128
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 14922 2896 14978 2952
rect 20074 2896 20130 2952
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 34610 5616 34666 5672
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 34978 5072 35034 5128
rect 34610 3984 34666 4040
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 22190 2372 22246 2408
rect 22190 2352 22192 2372
rect 22192 2352 22244 2372
rect 22244 2352 22246 2372
rect 33322 2352 33378 2408
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 21730 1400 21786 1456
rect 24950 1400 25006 1456
<< metal3 >>
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 34697 12066 34763 12069
rect 39520 12066 40000 12096
rect 34697 12064 40000 12066
rect 34697 12008 34702 12064
rect 34758 12008 40000 12064
rect 34697 12006 40000 12008
rect 34697 12003 34763 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12006
rect 34277 11935 34597 11936
rect 16757 11930 16823 11933
rect 19977 11930 20043 11933
rect 16757 11928 20043 11930
rect 16757 11872 16762 11928
rect 16818 11872 19982 11928
rect 20038 11872 20043 11928
rect 16757 11870 20043 11872
rect 16757 11867 16823 11870
rect 19977 11867 20043 11870
rect 6637 11658 6703 11661
rect 15101 11658 15167 11661
rect 6637 11656 15167 11658
rect 6637 11600 6642 11656
rect 6698 11600 15106 11656
rect 15162 11600 15167 11656
rect 6637 11598 15167 11600
rect 6637 11595 6703 11598
rect 15101 11595 15167 11598
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 16757 9482 16823 9485
rect 34697 9482 34763 9485
rect 16757 9480 34763 9482
rect 16757 9424 16762 9480
rect 16818 9424 34702 9480
rect 34758 9424 34763 9480
rect 16757 9422 34763 9424
rect 16757 9419 16823 9422
rect 34697 9419 34763 9422
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 9215 27930 9216
rect 4981 9074 5047 9077
rect 16573 9074 16639 9077
rect 4981 9072 16639 9074
rect 4981 9016 4986 9072
rect 5042 9016 16578 9072
rect 16634 9016 16639 9072
rect 4981 9014 16639 9016
rect 4981 9011 5047 9014
rect 16573 9011 16639 9014
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 14277 8192 14597 8193
rect 0 8122 480 8152
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 2957 8122 3023 8125
rect 0 8120 3023 8122
rect 0 8064 2962 8120
rect 3018 8064 3023 8120
rect 0 8062 3023 8064
rect 0 8032 480 8062
rect 2957 8059 3023 8062
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 2957 5810 3023 5813
rect 16205 5810 16271 5813
rect 2957 5808 16271 5810
rect 2957 5752 2962 5808
rect 3018 5752 16210 5808
rect 16266 5752 16271 5808
rect 2957 5750 16271 5752
rect 2957 5747 3023 5750
rect 16205 5747 16271 5750
rect 17401 5674 17467 5677
rect 34605 5674 34671 5677
rect 17401 5672 34671 5674
rect 17401 5616 17406 5672
rect 17462 5616 34610 5672
rect 34666 5616 34671 5672
rect 17401 5614 34671 5616
rect 17401 5611 17467 5614
rect 34605 5611 34671 5614
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 16021 5130 16087 5133
rect 34973 5130 35039 5133
rect 16021 5128 35039 5130
rect 16021 5072 16026 5128
rect 16082 5072 34978 5128
rect 35034 5072 35039 5128
rect 16021 5070 35039 5072
rect 16021 5067 16087 5070
rect 34973 5067 35039 5070
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 34605 4042 34671 4045
rect 39520 4042 40000 4072
rect 34605 4040 40000 4042
rect 34605 3984 34610 4040
rect 34666 3984 40000 4040
rect 34605 3982 40000 3984
rect 34605 3979 34671 3982
rect 39520 3952 40000 3982
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 14917 2954 14983 2957
rect 20069 2954 20135 2957
rect 14917 2952 20135 2954
rect 14917 2896 14922 2952
rect 14978 2896 20074 2952
rect 20130 2896 20135 2952
rect 14917 2894 20135 2896
rect 14917 2891 14983 2894
rect 20069 2891 20135 2894
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 22185 2410 22251 2413
rect 33317 2410 33383 2413
rect 22185 2408 33383 2410
rect 22185 2352 22190 2408
rect 22246 2352 33322 2408
rect 33378 2352 33383 2408
rect 22185 2350 33383 2352
rect 22185 2347 22251 2350
rect 33317 2347 33383 2350
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 21725 1458 21791 1461
rect 24945 1458 25011 1461
rect 21725 1456 25011 1458
rect 21725 1400 21730 1456
rect 21786 1400 24950 1456
rect 25006 1400 25011 1456
rect 21725 1398 25011 1400
rect 21725 1395 21791 1398
rect 24945 1395 25011 1398
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_203 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__0__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _1_
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__1__A
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_323
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_330
timestamp 1586364061
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_342
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_354
timestamp 1586364061
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_288
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_300
timestamp 1586364061
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_312
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_scs8hd_dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_scs8hd_dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_293
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_dfxbp_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_scs8hd_dfxbp_1_mem.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_193
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_288
timestamp 1586364061
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_293
timestamp 1586364061
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_300
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_330
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_342
timestamp 1586364061
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_288
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_300
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_324
timestamp 1586364061
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_293
timestamp 1586364061
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_342
timestamp 1586364061
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_354
timestamp 1586364061
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_373
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_385
timestamp 1586364061
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_354
timestamp 1586364061
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_379
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_391
timestamp 1586364061
transform 1 0 37076 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_373
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_385
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _2_
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__2__A
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_176
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_373
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_379
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_391
timestamp 1586364061
transform 1 0 37076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_385
timestamp 1586364061
transform 1 0 36524 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_403
timestamp 1586364061
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_379
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_288
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_300
timestamp 1586364061
transform 1 0 28704 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_361
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_385
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _3_
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__3__A
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_154
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.ie_oe_inv tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.ie_oe_inv_A
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4986 0 5042 480 6 bottom_width_0_height_0__pin_0_
port 0 nsew default input
rlabel metal2 s 14922 0 14978 480 6 bottom_width_0_height_0__pin_1_lower
port 1 nsew default tristate
rlabel metal2 s 24950 0 25006 480 6 bottom_width_0_height_0__pin_1_upper
port 2 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 ccff_head
port 3 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 ccff_tail
port 4 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 gfpga_pad_GPIO_A
port 5 nsew default tristate
rlabel metal2 s 6642 15520 6698 16000 6 gfpga_pad_GPIO_IE
port 6 nsew default tristate
rlabel metal2 s 19982 15520 20038 16000 6 gfpga_pad_GPIO_OE
port 7 nsew default tristate
rlabel metal2 s 33322 15520 33378 16000 6 gfpga_pad_GPIO_Y
port 8 nsew default bidirectional
rlabel metal2 s 34978 0 35034 480 6 prog_clk
port 9 nsew default input
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 10 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 11 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
