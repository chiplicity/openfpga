magic
tech sky130A
magscale 1 2
timestamp 1608762085
<< checkpaint >>
rect -1260 -1260 24060 24060
<< locali >>
rect 16681 7395 16715 7497
rect 13277 7191 13311 7293
rect 11253 6783 11287 6953
rect 14565 5083 14599 5185
rect 11253 3587 11287 3689
<< viali >>
rect 20177 20009 20211 20043
rect 20729 20009 20763 20043
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 20729 19465 20763 19499
rect 6837 19261 6871 19295
rect 12817 19261 12851 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 7021 19125 7055 19159
rect 13001 19125 13035 19159
rect 20177 19125 20211 19159
rect 20453 18921 20487 18955
rect 20269 18785 20303 18819
rect 9873 18241 9907 18275
rect 12725 18241 12759 18275
rect 16129 18241 16163 18275
rect 18337 18241 18371 18275
rect 9597 18173 9631 18207
rect 12449 18173 12483 18207
rect 15853 18173 15887 18207
rect 18061 18173 18095 18207
rect 19533 18173 19567 18207
rect 19809 18173 19843 18207
rect 15485 17833 15519 17867
rect 7573 17697 7607 17731
rect 12173 17697 12207 17731
rect 15301 17697 15335 17731
rect 7849 17629 7883 17663
rect 12357 17561 12391 17595
rect 20177 17289 20211 17323
rect 20729 17289 20763 17323
rect 11621 17153 11655 17187
rect 14105 17153 14139 17187
rect 11345 17085 11379 17119
rect 13829 17085 13863 17119
rect 19993 17085 20027 17119
rect 20545 17085 20579 17119
rect 20453 16745 20487 16779
rect 19809 16677 19843 16711
rect 19533 16609 19567 16643
rect 20269 16609 20303 16643
rect 20729 16201 20763 16235
rect 19901 16065 19935 16099
rect 19625 15997 19659 16031
rect 20545 15997 20579 16031
rect 20453 15657 20487 15691
rect 14289 15589 14323 15623
rect 14013 15521 14047 15555
rect 20269 15521 20303 15555
rect 20177 15113 20211 15147
rect 12725 14977 12759 15011
rect 12449 14909 12483 14943
rect 19993 14909 20027 14943
rect 20545 14909 20579 14943
rect 20729 14773 20763 14807
rect 19901 14569 19935 14603
rect 8309 14433 8343 14467
rect 9689 14433 9723 14467
rect 9965 14433 9999 14467
rect 19717 14433 19751 14467
rect 20269 14433 20303 14467
rect 8585 14365 8619 14399
rect 20453 14297 20487 14331
rect 10701 13821 10735 13855
rect 10977 13821 11011 13855
rect 20085 13821 20119 13855
rect 20729 13753 20763 13787
rect 19257 13481 19291 13515
rect 19901 13413 19935 13447
rect 16396 13345 16430 13379
rect 19073 13345 19107 13379
rect 19625 13345 19659 13379
rect 16129 13277 16163 13311
rect 17509 13141 17543 13175
rect 18061 12937 18095 12971
rect 20913 12937 20947 12971
rect 18613 12801 18647 12835
rect 19441 12801 19475 12835
rect 20269 12801 20303 12835
rect 19257 12733 19291 12767
rect 19993 12733 20027 12767
rect 20729 12733 20763 12767
rect 18429 12597 18463 12631
rect 18521 12597 18555 12631
rect 17325 12393 17359 12427
rect 17868 12325 17902 12359
rect 16212 12257 16246 12291
rect 19257 12257 19291 12291
rect 19809 12257 19843 12291
rect 15485 12189 15519 12223
rect 15945 12189 15979 12223
rect 17601 12189 17635 12223
rect 20085 12189 20119 12223
rect 18981 12053 19015 12087
rect 19441 12053 19475 12087
rect 13185 11849 13219 11883
rect 17509 11849 17543 11883
rect 20729 11849 20763 11883
rect 13737 11713 13771 11747
rect 18061 11713 18095 11747
rect 18613 11713 18647 11747
rect 14473 11645 14507 11679
rect 16129 11645 16163 11679
rect 20545 11645 20579 11679
rect 13645 11577 13679 11611
rect 14740 11577 14774 11611
rect 16374 11577 16408 11611
rect 18880 11577 18914 11611
rect 13553 11509 13587 11543
rect 15853 11509 15887 11543
rect 19993 11509 20027 11543
rect 13001 11305 13035 11339
rect 15301 11305 15335 11339
rect 15669 11305 15703 11339
rect 16589 11305 16623 11339
rect 18889 11305 18923 11339
rect 19441 11305 19475 11339
rect 19901 11305 19935 11339
rect 13728 11237 13762 11271
rect 18797 11237 18831 11271
rect 20913 11237 20947 11271
rect 12173 11169 12207 11203
rect 16957 11169 16991 11203
rect 19809 11169 19843 11203
rect 12449 11101 12483 11135
rect 13461 11101 13495 11135
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 17049 11101 17083 11135
rect 17233 11101 17267 11135
rect 19073 11101 19107 11135
rect 19993 11101 20027 11135
rect 14841 11033 14875 11067
rect 18429 11033 18463 11067
rect 13921 10761 13955 10795
rect 14841 10761 14875 10795
rect 16129 10761 16163 10795
rect 15393 10625 15427 10659
rect 18981 10625 19015 10659
rect 12541 10557 12575 10591
rect 16313 10557 16347 10591
rect 19349 10557 19383 10591
rect 19605 10557 19639 10591
rect 12808 10489 12842 10523
rect 18705 10489 18739 10523
rect 14657 10421 14691 10455
rect 15209 10421 15243 10455
rect 15301 10421 15335 10455
rect 17509 10421 17543 10455
rect 18337 10421 18371 10455
rect 18797 10421 18831 10455
rect 20729 10421 20763 10455
rect 15669 10217 15703 10251
rect 17132 10149 17166 10183
rect 16037 10081 16071 10115
rect 18788 10081 18822 10115
rect 20269 10081 20303 10115
rect 16129 10013 16163 10047
rect 16313 10013 16347 10047
rect 16865 10013 16899 10047
rect 18521 10013 18555 10047
rect 20453 9945 20487 9979
rect 18245 9877 18279 9911
rect 19901 9877 19935 9911
rect 19441 9673 19475 9707
rect 17049 9537 17083 9571
rect 20269 9537 20303 9571
rect 20361 9537 20395 9571
rect 13001 9469 13035 9503
rect 13737 9469 13771 9503
rect 15393 9469 15427 9503
rect 18061 9469 18095 9503
rect 20821 9469 20855 9503
rect 13277 9401 13311 9435
rect 14004 9401 14038 9435
rect 15660 9401 15694 9435
rect 18328 9401 18362 9435
rect 15117 9333 15151 9367
rect 16773 9333 16807 9367
rect 19809 9333 19843 9367
rect 20177 9333 20211 9367
rect 21005 9333 21039 9367
rect 10425 9129 10459 9163
rect 17417 9129 17451 9163
rect 17785 9129 17819 9163
rect 17877 9129 17911 9163
rect 20545 9129 20579 9163
rect 15844 9061 15878 9095
rect 10609 8993 10643 9027
rect 11345 8993 11379 9027
rect 11612 8993 11646 9027
rect 13268 8993 13302 9027
rect 15577 8993 15611 9027
rect 19165 8993 19199 9027
rect 19432 8993 19466 9027
rect 13001 8925 13035 8959
rect 14657 8925 14691 8959
rect 18061 8925 18095 8959
rect 18705 8925 18739 8959
rect 12725 8857 12759 8891
rect 14381 8789 14415 8823
rect 16957 8789 16991 8823
rect 8861 8585 8895 8619
rect 14749 8585 14783 8619
rect 15577 8585 15611 8619
rect 20545 8585 20579 8619
rect 11621 8517 11655 8551
rect 16405 8517 16439 8551
rect 9413 8449 9447 8483
rect 15301 8449 15335 8483
rect 16129 8449 16163 8483
rect 16957 8449 16991 8483
rect 18613 8449 18647 8483
rect 18797 8449 18831 8483
rect 10241 8381 10275 8415
rect 12909 8381 12943 8415
rect 15117 8381 15151 8415
rect 16773 8381 16807 8415
rect 18521 8381 18555 8415
rect 19165 8381 19199 8415
rect 19432 8381 19466 8415
rect 9321 8313 9355 8347
rect 10508 8313 10542 8347
rect 11897 8313 11931 8347
rect 16037 8313 16071 8347
rect 16865 8313 16899 8347
rect 9229 8245 9263 8279
rect 14197 8245 14231 8279
rect 15209 8245 15243 8279
rect 15945 8245 15979 8279
rect 17233 8245 17267 8279
rect 18153 8245 18187 8279
rect 9321 8041 9355 8075
rect 11069 8041 11103 8075
rect 13553 8041 13587 8075
rect 15485 8041 15519 8075
rect 9934 7973 9968 8007
rect 13921 7973 13955 8007
rect 16212 7973 16246 8007
rect 7941 7905 7975 7939
rect 8208 7905 8242 7939
rect 9689 7905 9723 7939
rect 11897 7905 11931 7939
rect 12164 7905 12198 7939
rect 15669 7905 15703 7939
rect 15945 7905 15979 7939
rect 17601 7905 17635 7939
rect 18337 7905 18371 7939
rect 20177 7905 20211 7939
rect 14013 7837 14047 7871
rect 14105 7837 14139 7871
rect 17785 7837 17819 7871
rect 18613 7837 18647 7871
rect 19257 7837 19291 7871
rect 20269 7837 20303 7871
rect 20453 7837 20487 7871
rect 13277 7701 13311 7735
rect 17325 7701 17359 7735
rect 19809 7701 19843 7735
rect 12449 7497 12483 7531
rect 16681 7497 16715 7531
rect 18797 7497 18831 7531
rect 19809 7497 19843 7531
rect 10517 7429 10551 7463
rect 15761 7429 15795 7463
rect 9413 7361 9447 7395
rect 11069 7361 11103 7395
rect 12909 7361 12943 7395
rect 13001 7361 13035 7395
rect 16313 7361 16347 7395
rect 16681 7361 16715 7395
rect 17325 7361 17359 7395
rect 18337 7361 18371 7395
rect 19257 7361 19291 7395
rect 19349 7361 19383 7395
rect 20361 7361 20395 7395
rect 11713 7293 11747 7327
rect 12817 7293 12851 7327
rect 13277 7293 13311 7327
rect 13461 7293 13495 7327
rect 13728 7293 13762 7327
rect 17141 7293 17175 7327
rect 18061 7293 18095 7327
rect 19165 7293 19199 7327
rect 20269 7225 20303 7259
rect 10885 7157 10919 7191
rect 10977 7157 11011 7191
rect 11529 7157 11563 7191
rect 13277 7157 13311 7191
rect 14841 7157 14875 7191
rect 16129 7157 16163 7191
rect 16221 7157 16255 7191
rect 16773 7157 16807 7191
rect 17233 7157 17267 7191
rect 20177 7157 20211 7191
rect 11253 6953 11287 6987
rect 12725 6953 12759 6987
rect 15301 6953 15335 6987
rect 9689 6817 9723 6851
rect 9956 6817 9990 6851
rect 13185 6885 13219 6919
rect 13277 6885 13311 6919
rect 15669 6885 15703 6919
rect 11612 6817 11646 6851
rect 14013 6817 14047 6851
rect 16497 6817 16531 6851
rect 16948 6817 16982 6851
rect 18797 6817 18831 6851
rect 19064 6817 19098 6851
rect 9137 6749 9171 6783
rect 11253 6749 11287 6783
rect 11345 6749 11379 6783
rect 13369 6749 13403 6783
rect 14105 6749 14139 6783
rect 14197 6749 14231 6783
rect 15761 6749 15795 6783
rect 15945 6749 15979 6783
rect 16681 6749 16715 6783
rect 11069 6681 11103 6715
rect 12817 6681 12851 6715
rect 13645 6681 13679 6715
rect 16313 6613 16347 6647
rect 18061 6613 18095 6647
rect 20177 6613 20211 6647
rect 10241 6409 10275 6443
rect 10701 6409 10735 6443
rect 13185 6409 13219 6443
rect 17509 6409 17543 6443
rect 11345 6273 11379 6307
rect 13737 6273 13771 6307
rect 20361 6273 20395 6307
rect 7205 6205 7239 6239
rect 8861 6205 8895 6239
rect 12449 6205 12483 6239
rect 14473 6205 14507 6239
rect 16129 6205 16163 6239
rect 18061 6205 18095 6239
rect 18317 6205 18351 6239
rect 20729 6205 20763 6239
rect 7472 6137 7506 6171
rect 9106 6137 9140 6171
rect 13553 6137 13587 6171
rect 14740 6137 14774 6171
rect 16396 6137 16430 6171
rect 20177 6137 20211 6171
rect 8585 6069 8619 6103
rect 11069 6069 11103 6103
rect 11161 6069 11195 6103
rect 13645 6069 13679 6103
rect 15853 6069 15887 6103
rect 19441 6069 19475 6103
rect 19717 6069 19751 6103
rect 20085 6069 20119 6103
rect 20913 6069 20947 6103
rect 8033 5865 8067 5899
rect 10057 5865 10091 5899
rect 16221 5865 16255 5899
rect 17601 5865 17635 5899
rect 18705 5865 18739 5899
rect 20085 5865 20119 5899
rect 20913 5865 20947 5899
rect 14473 5797 14507 5831
rect 19073 5797 19107 5831
rect 6644 5729 6678 5763
rect 8401 5729 8435 5763
rect 9045 5729 9079 5763
rect 11049 5729 11083 5763
rect 12900 5729 12934 5763
rect 16589 5729 16623 5763
rect 16681 5729 16715 5763
rect 20177 5729 20211 5763
rect 6377 5661 6411 5695
rect 8493 5661 8527 5695
rect 8585 5661 8619 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 10793 5661 10827 5695
rect 12633 5661 12667 5695
rect 14565 5661 14599 5695
rect 14657 5661 14691 5695
rect 16773 5661 16807 5695
rect 17693 5661 17727 5695
rect 17785 5661 17819 5695
rect 19165 5661 19199 5695
rect 19349 5661 19383 5695
rect 20269 5661 20303 5695
rect 7757 5593 7791 5627
rect 9689 5593 9723 5627
rect 14013 5593 14047 5627
rect 12173 5525 12207 5559
rect 14105 5525 14139 5559
rect 17233 5525 17267 5559
rect 19717 5525 19751 5559
rect 8493 5321 8527 5355
rect 12633 5321 12667 5355
rect 13645 5321 13679 5355
rect 14657 5321 14691 5355
rect 16221 5321 16255 5355
rect 18337 5321 18371 5355
rect 19349 5321 19383 5355
rect 9965 5253 9999 5287
rect 9045 5185 9079 5219
rect 10241 5185 10275 5219
rect 13277 5185 13311 5219
rect 14197 5185 14231 5219
rect 14565 5185 14599 5219
rect 15117 5185 15151 5219
rect 15301 5185 15335 5219
rect 15669 5185 15703 5219
rect 16773 5185 16807 5219
rect 18889 5185 18923 5219
rect 19809 5185 19843 5219
rect 19901 5185 19935 5219
rect 6837 5117 6871 5151
rect 10149 5117 10183 5151
rect 14105 5117 14139 5151
rect 16681 5117 16715 5151
rect 19717 5117 19751 5151
rect 20545 5117 20579 5151
rect 7104 5049 7138 5083
rect 10508 5049 10542 5083
rect 13093 5049 13127 5083
rect 14013 5049 14047 5083
rect 14565 5049 14599 5083
rect 18705 5049 18739 5083
rect 8217 4981 8251 5015
rect 8861 4981 8895 5015
rect 8953 4981 8987 5015
rect 11621 4981 11655 5015
rect 13001 4981 13035 5015
rect 15025 4981 15059 5015
rect 16589 4981 16623 5015
rect 18797 4981 18831 5015
rect 20729 4981 20763 5015
rect 6653 4777 6687 4811
rect 7665 4777 7699 4811
rect 11621 4777 11655 4811
rect 13369 4777 13403 4811
rect 10977 4709 11011 4743
rect 19432 4709 19466 4743
rect 7021 4641 7055 4675
rect 7113 4641 7147 4675
rect 8033 4641 8067 4675
rect 17325 4641 17359 4675
rect 17592 4641 17626 4675
rect 19165 4641 19199 4675
rect 7205 4573 7239 4607
rect 8125 4573 8159 4607
rect 8217 4573 8251 4607
rect 11069 4573 11103 4607
rect 11253 4573 11287 4607
rect 10609 4505 10643 4539
rect 18705 4437 18739 4471
rect 20545 4437 20579 4471
rect 9137 4233 9171 4267
rect 7757 4097 7791 4131
rect 9873 4097 9907 4131
rect 9965 4097 9999 4131
rect 13001 4097 13035 4131
rect 14105 4097 14139 4131
rect 15761 4097 15795 4131
rect 18061 4097 18095 4131
rect 20361 4097 20395 4131
rect 17417 4029 17451 4063
rect 18328 4029 18362 4063
rect 20729 4029 20763 4063
rect 8024 3961 8058 3995
rect 9781 3961 9815 3995
rect 9413 3893 9447 3927
rect 10517 3893 10551 3927
rect 11621 3893 11655 3927
rect 12449 3893 12483 3927
rect 12817 3893 12851 3927
rect 12909 3893 12943 3927
rect 13553 3893 13587 3927
rect 13921 3893 13955 3927
rect 14013 3893 14047 3927
rect 15117 3893 15151 3927
rect 15485 3893 15519 3927
rect 15577 3893 15611 3927
rect 17601 3893 17635 3927
rect 19441 3893 19475 3927
rect 19717 3893 19751 3927
rect 20085 3893 20119 3927
rect 20177 3893 20211 3927
rect 20913 3893 20947 3927
rect 8493 3689 8527 3723
rect 11253 3689 11287 3723
rect 12725 3689 12759 3723
rect 17693 3689 17727 3723
rect 18061 3689 18095 3723
rect 18705 3689 18739 3723
rect 19073 3689 19107 3723
rect 19717 3689 19751 3723
rect 20085 3689 20119 3723
rect 15660 3621 15694 3655
rect 19165 3621 19199 3655
rect 20913 3621 20947 3655
rect 7113 3553 7147 3587
rect 7380 3553 7414 3587
rect 9689 3553 9723 3587
rect 9956 3553 9990 3587
rect 11253 3553 11287 3587
rect 11345 3553 11379 3587
rect 11612 3553 11646 3587
rect 13360 3553 13394 3587
rect 17141 3553 17175 3587
rect 20177 3553 20211 3587
rect 13093 3485 13127 3519
rect 14749 3485 14783 3519
rect 15393 3485 15427 3519
rect 18153 3485 18187 3519
rect 18245 3485 18279 3519
rect 19257 3485 19291 3519
rect 20361 3485 20395 3519
rect 14473 3417 14507 3451
rect 11069 3349 11103 3383
rect 16773 3349 16807 3383
rect 17325 3349 17359 3383
rect 8217 3145 8251 3179
rect 10701 3145 10735 3179
rect 10977 3145 11011 3179
rect 14381 3145 14415 3179
rect 16865 3145 16899 3179
rect 18061 3145 18095 3179
rect 20637 3145 20671 3179
rect 19533 3077 19567 3111
rect 6837 3009 6871 3043
rect 8493 3009 8527 3043
rect 11529 3009 11563 3043
rect 15209 3009 15243 3043
rect 17325 3009 17359 3043
rect 17417 3009 17451 3043
rect 18521 3009 18555 3043
rect 18705 3009 18739 3043
rect 9321 2941 9355 2975
rect 11345 2941 11379 2975
rect 12449 2941 12483 2975
rect 13001 2941 13035 2975
rect 13268 2941 13302 2975
rect 14657 2941 14691 2975
rect 15476 2941 15510 2975
rect 18429 2941 18463 2975
rect 19349 2941 19383 2975
rect 19901 2941 19935 2975
rect 20453 2941 20487 2975
rect 7104 2873 7138 2907
rect 9588 2873 9622 2907
rect 11437 2805 11471 2839
rect 12633 2805 12667 2839
rect 14841 2805 14875 2839
rect 16589 2805 16623 2839
rect 17233 2805 17267 2839
rect 20085 2805 20119 2839
rect 7389 2601 7423 2635
rect 10057 2601 10091 2635
rect 11713 2601 11747 2635
rect 13645 2601 13679 2635
rect 14289 2601 14323 2635
rect 14749 2601 14783 2635
rect 15669 2601 15703 2635
rect 16037 2601 16071 2635
rect 20085 2601 20119 2635
rect 10425 2533 10459 2567
rect 13737 2533 13771 2567
rect 7757 2465 7791 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 14657 2465 14691 2499
rect 16957 2465 16991 2499
rect 17509 2465 17543 2499
rect 18337 2465 18371 2499
rect 18889 2465 18923 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 7849 2397 7883 2431
rect 8033 2397 8067 2431
rect 10517 2397 10551 2431
rect 10701 2397 10735 2431
rect 11897 2397 11931 2431
rect 13829 2397 13863 2431
rect 14841 2397 14875 2431
rect 16129 2397 16163 2431
rect 16313 2397 16347 2431
rect 11345 2329 11379 2363
rect 13277 2329 13311 2363
rect 17693 2329 17727 2363
rect 19073 2329 19107 2363
rect 20637 2329 20671 2363
rect 12817 2261 12851 2295
rect 17141 2261 17175 2295
rect 18521 2261 18555 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 19978 19904 19984 19916
rect 19939 19876 19984 19904
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20070 19864 20076 19916
rect 20128 19904 20134 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 20128 19876 20545 19904
rect 20128 19864 20134 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 20714 19496 20720 19508
rect 20675 19468 20720 19496
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 5718 19252 5724 19304
rect 5776 19292 5782 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 5776 19264 6837 19292
rect 5776 19252 5782 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 12710 19252 12716 19304
rect 12768 19292 12774 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12768 19264 12817 19292
rect 12768 19252 12774 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 16172 19264 19993 19292
rect 16172 19252 16178 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 19981 19255 20039 19261
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 7006 19156 7012 19168
rect 6967 19128 7012 19156
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 12989 19159 13047 19165
rect 12989 19125 13001 19159
rect 13035 19156 13047 19159
rect 17954 19156 17960 19168
rect 13035 19128 17960 19156
rect 13035 19125 13047 19128
rect 12989 19119 13047 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 19300 19128 20177 19156
rect 19300 19116 19306 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 20165 19119 20223 19125
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 20438 18952 20444 18964
rect 20399 18924 20444 18952
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 20254 18816 20260 18828
rect 20215 18788 20260 18816
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 20530 18340 20536 18352
rect 9876 18312 20536 18340
rect 9876 18281 9904 18312
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18241 9919 18275
rect 12710 18272 12716 18284
rect 12671 18244 12716 18272
rect 9861 18235 9919 18241
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 16114 18272 16120 18284
rect 16075 18244 16120 18272
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 18325 18275 18383 18281
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 19978 18272 19984 18284
rect 18371 18244 19984 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18204 9643 18207
rect 9766 18204 9772 18216
rect 9631 18176 9772 18204
rect 9631 18173 9643 18176
rect 9585 18167 9643 18173
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 12437 18207 12495 18213
rect 12437 18173 12449 18207
rect 12483 18204 12495 18207
rect 13630 18204 13636 18216
rect 12483 18176 13636 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 13630 18164 13636 18176
rect 13688 18164 13694 18216
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15344 18176 15853 18204
rect 15344 18164 15350 18176
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 18012 18176 18061 18204
rect 18012 18164 18018 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18173 19579 18207
rect 19521 18167 19579 18173
rect 19797 18207 19855 18213
rect 19797 18173 19809 18207
rect 19843 18204 19855 18207
rect 20070 18204 20076 18216
rect 19843 18176 20076 18204
rect 19843 18173 19855 18176
rect 19797 18167 19855 18173
rect 19536 18136 19564 18167
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 19978 18136 19984 18148
rect 19536 18108 19984 18136
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 15473 17867 15531 17873
rect 15473 17833 15485 17867
rect 15519 17864 15531 17867
rect 17862 17864 17868 17876
rect 15519 17836 17868 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17728 7619 17731
rect 7650 17728 7656 17740
rect 7607 17700 7656 17728
rect 7607 17697 7619 17700
rect 7561 17691 7619 17697
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 12161 17731 12219 17737
rect 12161 17728 12173 17731
rect 11664 17700 12173 17728
rect 11664 17688 11670 17700
rect 12161 17697 12173 17700
rect 12207 17697 12219 17731
rect 12161 17691 12219 17697
rect 14090 17688 14096 17740
rect 14148 17728 14154 17740
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 14148 17700 15301 17728
rect 14148 17688 14154 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17660 7895 17663
rect 20254 17660 20260 17672
rect 7883 17632 20260 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 20254 17620 20260 17632
rect 20312 17620 20318 17672
rect 12345 17595 12403 17601
rect 12345 17561 12357 17595
rect 12391 17592 12403 17595
rect 18506 17592 18512 17604
rect 12391 17564 18512 17592
rect 12391 17561 12403 17564
rect 12345 17555 12403 17561
rect 18506 17552 18512 17564
rect 18564 17552 18570 17604
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 11606 17184 11612 17196
rect 11567 17156 11612 17184
rect 11606 17144 11612 17156
rect 11664 17144 11670 17196
rect 14090 17184 14096 17196
rect 14051 17156 14096 17184
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17116 11391 17119
rect 11790 17116 11796 17128
rect 11379 17088 11796 17116
rect 11379 17085 11391 17088
rect 11333 17079 11391 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 13814 17116 13820 17128
rect 13775 17088 13820 17116
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 19794 17076 19800 17128
rect 19852 17116 19858 17128
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 19852 17088 19993 17116
rect 19852 17076 19858 17088
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 20070 17076 20076 17128
rect 20128 17116 20134 17128
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 20128 17088 20545 17116
rect 20128 17076 20134 17088
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 20438 16776 20444 16788
rect 20399 16748 20444 16776
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 18506 16668 18512 16720
rect 18564 16708 18570 16720
rect 19794 16708 19800 16720
rect 18564 16680 19656 16708
rect 19755 16680 19800 16708
rect 18564 16668 18570 16680
rect 19518 16640 19524 16652
rect 19479 16612 19524 16640
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 19628 16640 19656 16680
rect 19794 16668 19800 16680
rect 19852 16668 19858 16720
rect 20257 16643 20315 16649
rect 20257 16640 20269 16643
rect 19628 16612 20269 16640
rect 20257 16609 20269 16612
rect 20303 16609 20315 16643
rect 20257 16603 20315 16609
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 19889 16099 19947 16105
rect 19889 16065 19901 16099
rect 19935 16096 19947 16099
rect 20070 16096 20076 16108
rect 19935 16068 20076 16096
rect 19935 16065 19947 16068
rect 19889 16059 19947 16065
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 19613 16031 19671 16037
rect 19613 16028 19625 16031
rect 17000 16000 19625 16028
rect 17000 15988 17006 16000
rect 19613 15997 19625 16000
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 16666 15920 16672 15972
rect 16724 15960 16730 15972
rect 20548 15960 20576 15991
rect 16724 15932 20576 15960
rect 16724 15920 16730 15932
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 14277 15623 14335 15629
rect 14277 15589 14289 15623
rect 14323 15620 14335 15623
rect 18506 15620 18512 15632
rect 14323 15592 18512 15620
rect 14323 15589 14335 15592
rect 14277 15583 14335 15589
rect 18506 15580 18512 15592
rect 18564 15580 18570 15632
rect 13998 15552 14004 15564
rect 13959 15524 14004 15552
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 19392 15524 20269 15552
rect 19392 15512 19398 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 20162 15144 20168 15156
rect 20123 15116 20168 15144
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 15008 12771 15011
rect 16666 15008 16672 15020
rect 12759 14980 16672 15008
rect 12759 14977 12771 14980
rect 12713 14971 12771 14977
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 19978 14940 19984 14952
rect 12492 14912 12537 14940
rect 19939 14912 19984 14940
rect 12492 14900 12498 14912
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20530 14940 20536 14952
rect 20491 14912 20536 14940
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 20714 14804 20720 14816
rect 20675 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 19886 14600 19892 14612
rect 19847 14572 19892 14600
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 9674 14464 9680 14476
rect 9635 14436 9680 14464
rect 9674 14424 9680 14436
rect 9732 14424 9738 14476
rect 9953 14467 10011 14473
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 19334 14464 19340 14476
rect 9999 14436 19340 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 19334 14424 19340 14436
rect 19392 14424 19398 14476
rect 19702 14464 19708 14476
rect 19663 14436 19708 14464
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 20254 14464 20260 14476
rect 20215 14436 20260 14464
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 19978 14396 19984 14408
rect 8619 14368 19984 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20438 14328 20444 14340
rect 20399 14300 20444 14328
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10870 13852 10876 13864
rect 10735 13824 10876 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 19702 13852 19708 13864
rect 11011 13824 19708 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13852 20131 13855
rect 20346 13852 20352 13864
rect 20119 13824 20352 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 18874 13744 18880 13796
rect 18932 13784 18938 13796
rect 20717 13787 20775 13793
rect 20717 13784 20729 13787
rect 18932 13756 20729 13784
rect 18932 13744 18938 13756
rect 20717 13753 20729 13756
rect 20763 13753 20775 13787
rect 20717 13747 20775 13753
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 19242 13512 19248 13524
rect 12584 13484 16804 13512
rect 19203 13484 19248 13512
rect 12584 13472 12590 13484
rect 16776 13444 16804 13484
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19889 13447 19947 13453
rect 16776 13416 19656 13444
rect 16384 13379 16442 13385
rect 16384 13345 16396 13379
rect 16430 13376 16442 13379
rect 17126 13376 17132 13388
rect 16430 13348 17132 13376
rect 16430 13345 16442 13348
rect 16384 13339 16442 13345
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 19061 13379 19119 13385
rect 19061 13345 19073 13379
rect 19107 13376 19119 13379
rect 19426 13376 19432 13388
rect 19107 13348 19432 13376
rect 19107 13345 19119 13348
rect 19061 13339 19119 13345
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 19628 13385 19656 13416
rect 19889 13413 19901 13447
rect 19935 13444 19947 13447
rect 20530 13444 20536 13456
rect 19935 13416 20536 13444
rect 19935 13413 19947 13416
rect 19889 13407 19947 13413
rect 20530 13404 20536 13416
rect 20588 13404 20594 13456
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13345 19671 13379
rect 19613 13339 19671 13345
rect 15930 13268 15936 13320
rect 15988 13308 15994 13320
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15988 13280 16129 13308
rect 15988 13268 15994 13280
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 17497 13175 17555 13181
rect 17497 13172 17509 13175
rect 16816 13144 17509 13172
rect 16816 13132 16822 13144
rect 17497 13141 17509 13144
rect 17543 13141 17555 13175
rect 17497 13135 17555 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18049 12971 18107 12977
rect 18049 12968 18061 12971
rect 18012 12940 18061 12968
rect 18012 12928 18018 12940
rect 18049 12937 18061 12940
rect 18095 12937 18107 12971
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 18049 12931 18107 12937
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 18598 12832 18604 12844
rect 18559 12804 18604 12832
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 19426 12832 19432 12844
rect 19387 12804 19432 12832
rect 19426 12792 19432 12804
rect 19484 12792 19490 12844
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 19058 12724 19064 12776
rect 19116 12764 19122 12776
rect 19245 12767 19303 12773
rect 19245 12764 19257 12767
rect 19116 12736 19257 12764
rect 19116 12724 19122 12736
rect 19245 12733 19257 12736
rect 19291 12733 19303 12767
rect 19245 12727 19303 12733
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12733 20039 12767
rect 19981 12727 20039 12733
rect 20717 12767 20775 12773
rect 20717 12733 20729 12767
rect 20763 12764 20775 12767
rect 20898 12764 20904 12776
rect 20763 12736 20904 12764
rect 20763 12733 20775 12736
rect 20717 12727 20775 12733
rect 14274 12656 14280 12708
rect 14332 12696 14338 12708
rect 19996 12696 20024 12727
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 14332 12668 20024 12696
rect 14332 12656 14338 12668
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18417 12631 18475 12637
rect 18417 12628 18429 12631
rect 18012 12600 18429 12628
rect 18012 12588 18018 12600
rect 18417 12597 18429 12600
rect 18463 12597 18475 12631
rect 18417 12591 18475 12597
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 18564 12600 18609 12628
rect 18564 12588 18570 12600
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 17313 12427 17371 12433
rect 17313 12393 17325 12427
rect 17359 12393 17371 12427
rect 17313 12387 17371 12393
rect 17328 12356 17356 12387
rect 17856 12359 17914 12365
rect 17856 12356 17868 12359
rect 17328 12328 17868 12356
rect 17856 12325 17868 12328
rect 17902 12356 17914 12359
rect 18598 12356 18604 12368
rect 17902 12328 18604 12356
rect 17902 12325 17914 12328
rect 17856 12319 17914 12325
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 16200 12291 16258 12297
rect 16200 12257 16212 12291
rect 16246 12288 16258 12291
rect 17494 12288 17500 12300
rect 16246 12260 17500 12288
rect 16246 12257 16258 12260
rect 16200 12251 16258 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 19242 12288 19248 12300
rect 19203 12260 19248 12288
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19794 12288 19800 12300
rect 19755 12260 19800 12288
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 15654 12220 15660 12232
rect 15519 12192 15660 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 15930 12220 15936 12232
rect 15891 12192 15936 12220
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12189 17647 12223
rect 17589 12183 17647 12189
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12220 20131 12223
rect 20530 12220 20536 12232
rect 20119 12192 20536 12220
rect 20119 12189 20131 12192
rect 20073 12183 20131 12189
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 17604 12084 17632 12183
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 18598 12084 18604 12096
rect 15988 12056 18604 12084
rect 15988 12044 15994 12056
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 18966 12084 18972 12096
rect 18927 12056 18972 12084
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 19429 12087 19487 12093
rect 19429 12053 19441 12087
rect 19475 12084 19487 12087
rect 20622 12084 20628 12096
rect 19475 12056 20628 12084
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 13173 11883 13231 11889
rect 13173 11849 13185 11883
rect 13219 11880 13231 11883
rect 17494 11880 17500 11892
rect 13219 11852 17080 11880
rect 17455 11852 17500 11880
rect 13219 11849 13231 11852
rect 13173 11843 13231 11849
rect 17052 11812 17080 11852
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 20070 11880 20076 11892
rect 17604 11852 20076 11880
rect 17604 11812 17632 11852
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20714 11880 20720 11892
rect 20675 11852 20720 11880
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 17052 11784 17632 11812
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 13906 11744 13912 11756
rect 13771 11716 13912 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 18012 11716 18061 11744
rect 18012 11704 18018 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 18049 11707 18107 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 13504 11648 14473 11676
rect 13504 11636 13510 11648
rect 14461 11645 14473 11648
rect 14507 11676 14519 11679
rect 15930 11676 15936 11688
rect 14507 11648 15936 11676
rect 14507 11645 14519 11648
rect 14461 11639 14519 11645
rect 15930 11636 15936 11648
rect 15988 11676 15994 11688
rect 16114 11676 16120 11688
rect 15988 11648 16120 11676
rect 15988 11636 15994 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 20530 11676 20536 11688
rect 20491 11648 20536 11676
rect 20530 11636 20536 11648
rect 20588 11636 20594 11688
rect 13354 11568 13360 11620
rect 13412 11608 13418 11620
rect 13633 11611 13691 11617
rect 13633 11608 13645 11611
rect 13412 11580 13645 11608
rect 13412 11568 13418 11580
rect 13633 11577 13645 11580
rect 13679 11577 13691 11611
rect 13633 11571 13691 11577
rect 14728 11611 14786 11617
rect 14728 11577 14740 11611
rect 14774 11608 14786 11611
rect 15378 11608 15384 11620
rect 14774 11580 15384 11608
rect 14774 11577 14786 11580
rect 14728 11571 14786 11577
rect 15378 11568 15384 11580
rect 15436 11568 15442 11620
rect 16362 11611 16420 11617
rect 16362 11608 16374 11611
rect 15856 11580 16374 11608
rect 15856 11552 15884 11580
rect 16362 11577 16374 11580
rect 16408 11577 16420 11611
rect 16362 11571 16420 11577
rect 18868 11611 18926 11617
rect 18868 11577 18880 11611
rect 18914 11608 18926 11611
rect 18966 11608 18972 11620
rect 18914 11580 18972 11608
rect 18914 11577 18926 11580
rect 18868 11571 18926 11577
rect 18966 11568 18972 11580
rect 19024 11608 19030 11620
rect 19426 11608 19432 11620
rect 19024 11580 19432 11608
rect 19024 11568 19030 11580
rect 19426 11568 19432 11580
rect 19484 11568 19490 11620
rect 13538 11540 13544 11552
rect 13499 11512 13544 11540
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 15838 11540 15844 11552
rect 15799 11512 15844 11540
rect 15838 11500 15844 11512
rect 15896 11500 15902 11552
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19981 11543 20039 11549
rect 19981 11540 19993 11543
rect 19392 11512 19993 11540
rect 19392 11500 19398 11512
rect 19981 11509 19993 11512
rect 20027 11509 20039 11543
rect 19981 11503 20039 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13538 11336 13544 11348
rect 13035 11308 13544 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 15286 11336 15292 11348
rect 13648 11308 15148 11336
rect 15247 11308 15292 11336
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 13648 11268 13676 11308
rect 4120 11240 13676 11268
rect 13716 11271 13774 11277
rect 4120 11228 4126 11240
rect 13716 11237 13728 11271
rect 13762 11268 13774 11271
rect 13906 11268 13912 11280
rect 13762 11240 13912 11268
rect 13762 11237 13774 11240
rect 13716 11231 13774 11237
rect 13906 11228 13912 11240
rect 13964 11228 13970 11280
rect 15120 11268 15148 11308
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15654 11336 15660 11348
rect 15615 11308 15660 11336
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16577 11339 16635 11345
rect 16577 11305 16589 11339
rect 16623 11336 16635 11339
rect 18506 11336 18512 11348
rect 16623 11308 18512 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 18923 11308 19441 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19886 11336 19892 11348
rect 19847 11308 19892 11336
rect 19429 11299 19487 11305
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 18785 11271 18843 11277
rect 15120 11240 18644 11268
rect 12161 11203 12219 11209
rect 12161 11169 12173 11203
rect 12207 11200 12219 11203
rect 16945 11203 17003 11209
rect 12207 11172 15516 11200
rect 12207 11169 12219 11172
rect 12161 11163 12219 11169
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 13170 11132 13176 11144
rect 12483 11104 13176 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 13446 11132 13452 11144
rect 13359 11104 13452 11132
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13078 11024 13084 11076
rect 13136 11064 13142 11076
rect 13464 11064 13492 11092
rect 13136 11036 13492 11064
rect 14829 11067 14887 11073
rect 13136 11024 13142 11036
rect 14829 11033 14841 11067
rect 14875 11064 14887 11067
rect 15378 11064 15384 11076
rect 14875 11036 15384 11064
rect 14875 11033 14887 11036
rect 14829 11027 14887 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 15488 11064 15516 11172
rect 16945 11169 16957 11203
rect 16991 11200 17003 11203
rect 17586 11200 17592 11212
rect 16991 11172 17592 11200
rect 16991 11169 17003 11172
rect 16945 11163 17003 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 18616 11200 18644 11240
rect 18785 11237 18797 11271
rect 18831 11268 18843 11271
rect 20901 11271 20959 11277
rect 20901 11268 20913 11271
rect 18831 11240 20913 11268
rect 18831 11237 18843 11240
rect 18785 11231 18843 11237
rect 20901 11237 20913 11240
rect 20947 11237 20959 11271
rect 20901 11231 20959 11237
rect 19150 11200 19156 11212
rect 18616 11172 19156 11200
rect 19150 11160 19156 11172
rect 19208 11160 19214 11212
rect 19797 11203 19855 11209
rect 19797 11169 19809 11203
rect 19843 11200 19855 11203
rect 20162 11200 20168 11212
rect 19843 11172 20168 11200
rect 19843 11169 19855 11172
rect 19797 11163 19855 11169
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 17034 11132 17040 11144
rect 15896 11104 15941 11132
rect 16995 11104 17040 11132
rect 15896 11092 15902 11104
rect 17034 11092 17040 11104
rect 17092 11092 17098 11144
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11132 17279 11135
rect 17494 11132 17500 11144
rect 17267 11104 17500 11132
rect 17267 11101 17279 11104
rect 17221 11095 17279 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 19061 11135 19119 11141
rect 19061 11101 19073 11135
rect 19107 11132 19119 11135
rect 19334 11132 19340 11144
rect 19107 11104 19340 11132
rect 19107 11101 19119 11104
rect 19061 11095 19119 11101
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 19981 11135 20039 11141
rect 19981 11132 19993 11135
rect 19484 11104 19993 11132
rect 19484 11092 19490 11104
rect 19981 11101 19993 11104
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 18417 11067 18475 11073
rect 18417 11064 18429 11067
rect 15488 11036 18429 11064
rect 18417 11033 18429 11036
rect 18463 11033 18475 11067
rect 18417 11027 18475 11033
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 13906 10792 13912 10804
rect 13867 10764 13912 10792
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 14829 10795 14887 10801
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15746 10792 15752 10804
rect 14875 10764 15752 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16114 10792 16120 10804
rect 16075 10764 16120 10792
rect 16114 10752 16120 10764
rect 16172 10792 16178 10804
rect 16574 10792 16580 10804
rect 16172 10764 16580 10792
rect 16172 10752 16178 10764
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 19334 10724 19340 10736
rect 18984 10696 19340 10724
rect 15378 10656 15384 10668
rect 15339 10628 15384 10656
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 18984 10665 19012 10696
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 11756 10560 12541 10588
rect 11756 10548 11762 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 16298 10588 16304 10600
rect 16259 10560 16304 10588
rect 12529 10551 12587 10557
rect 16298 10548 16304 10560
rect 16356 10548 16362 10600
rect 18506 10548 18512 10600
rect 18564 10588 18570 10600
rect 19337 10591 19395 10597
rect 19337 10588 19349 10591
rect 18564 10560 19349 10588
rect 18564 10548 18570 10560
rect 19337 10557 19349 10560
rect 19383 10557 19395 10591
rect 19337 10551 19395 10557
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19593 10591 19651 10597
rect 19593 10588 19605 10591
rect 19484 10560 19605 10588
rect 19484 10548 19490 10560
rect 19593 10557 19605 10560
rect 19639 10557 19651 10591
rect 19593 10551 19651 10557
rect 12796 10523 12854 10529
rect 12796 10489 12808 10523
rect 12842 10520 12854 10523
rect 13262 10520 13268 10532
rect 12842 10492 13268 10520
rect 12842 10489 12854 10492
rect 12796 10483 12854 10489
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 18693 10523 18751 10529
rect 18693 10489 18705 10523
rect 18739 10520 18751 10523
rect 20162 10520 20168 10532
rect 18739 10492 20168 10520
rect 18739 10489 18751 10492
rect 18693 10483 18751 10489
rect 20162 10480 20168 10492
rect 20220 10480 20226 10532
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14608 10424 14657 10452
rect 14608 10412 14614 10424
rect 14645 10421 14657 10424
rect 14691 10452 14703 10455
rect 15197 10455 15255 10461
rect 15197 10452 15209 10455
rect 14691 10424 15209 10452
rect 14691 10421 14703 10424
rect 14645 10415 14703 10421
rect 15197 10421 15209 10424
rect 15243 10421 15255 10455
rect 15197 10415 15255 10421
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 16022 10452 16028 10464
rect 15335 10424 16028 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 17494 10452 17500 10464
rect 17455 10424 17500 10452
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 18325 10455 18383 10461
rect 18325 10421 18337 10455
rect 18371 10452 18383 10455
rect 18598 10452 18604 10464
rect 18371 10424 18604 10452
rect 18371 10421 18383 10424
rect 18325 10415 18383 10421
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 18782 10412 18788 10464
rect 18840 10452 18846 10464
rect 18840 10424 18885 10452
rect 18840 10412 18846 10424
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 20404 10424 20729 10452
rect 20404 10412 20410 10424
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 20717 10415 20775 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 16942 10248 16948 10260
rect 15703 10220 16948 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 17120 10183 17178 10189
rect 17120 10149 17132 10183
rect 17166 10180 17178 10183
rect 20346 10180 20352 10192
rect 17166 10152 20352 10180
rect 17166 10149 17178 10152
rect 17120 10143 17178 10149
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 16025 10115 16083 10121
rect 16025 10081 16037 10115
rect 16071 10112 16083 10115
rect 16942 10112 16948 10124
rect 16071 10084 16948 10112
rect 16071 10081 16083 10084
rect 16025 10075 16083 10081
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 18776 10115 18834 10121
rect 18776 10081 18788 10115
rect 18822 10112 18834 10115
rect 19334 10112 19340 10124
rect 18822 10084 19340 10112
rect 18822 10081 18834 10084
rect 18776 10075 18834 10081
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 20254 10112 20260 10124
rect 20215 10084 20260 10112
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 15562 10004 15568 10056
rect 15620 10044 15626 10056
rect 16117 10047 16175 10053
rect 16117 10044 16129 10047
rect 15620 10016 16129 10044
rect 15620 10004 15626 10016
rect 16117 10013 16129 10016
rect 16163 10013 16175 10047
rect 16117 10007 16175 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10044 16359 10047
rect 16482 10044 16488 10056
rect 16347 10016 16488 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16632 10016 16865 10044
rect 16632 10004 16638 10016
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 17862 10004 17868 10056
rect 17920 10044 17926 10056
rect 18506 10044 18512 10056
rect 17920 10016 18512 10044
rect 17920 10004 17926 10016
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 20441 9979 20499 9985
rect 20441 9976 20453 9979
rect 19444 9948 20453 9976
rect 18233 9911 18291 9917
rect 18233 9877 18245 9911
rect 18279 9908 18291 9911
rect 18506 9908 18512 9920
rect 18279 9880 18512 9908
rect 18279 9877 18291 9880
rect 18233 9871 18291 9877
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 18690 9868 18696 9920
rect 18748 9908 18754 9920
rect 19444 9908 19472 9948
rect 20441 9945 20453 9948
rect 20487 9945 20499 9979
rect 20441 9939 20499 9945
rect 19886 9908 19892 9920
rect 18748 9880 19472 9908
rect 19847 9880 19892 9908
rect 18748 9868 18754 9880
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 12066 9664 12072 9716
rect 12124 9704 12130 9716
rect 18690 9704 18696 9716
rect 12124 9676 18696 9704
rect 12124 9664 12130 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 19334 9664 19340 9716
rect 19392 9704 19398 9716
rect 19429 9707 19487 9713
rect 19429 9704 19441 9707
rect 19392 9676 19441 9704
rect 19392 9664 19398 9676
rect 19429 9673 19441 9676
rect 19475 9673 19487 9707
rect 19429 9667 19487 9673
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 17000 9540 17049 9568
rect 17000 9528 17006 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19300 9540 20269 9568
rect 19300 9528 19306 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 20346 9528 20352 9580
rect 20404 9568 20410 9580
rect 20404 9540 20449 9568
rect 20404 9528 20410 9540
rect 12986 9500 12992 9512
rect 12947 9472 12992 9500
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13078 9460 13084 9512
rect 13136 9500 13142 9512
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13136 9472 13737 9500
rect 13136 9460 13142 9472
rect 13725 9469 13737 9472
rect 13771 9500 13783 9503
rect 15378 9500 15384 9512
rect 13771 9472 15384 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 17862 9500 17868 9512
rect 16632 9472 17868 9500
rect 16632 9460 16638 9472
rect 17862 9460 17868 9472
rect 17920 9500 17926 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17920 9472 18061 9500
rect 17920 9460 17926 9472
rect 18049 9469 18061 9472
rect 18095 9500 18107 9503
rect 18690 9500 18696 9512
rect 18095 9472 18696 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 20806 9500 20812 9512
rect 20767 9472 20812 9500
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 13265 9435 13323 9441
rect 13265 9432 13277 9435
rect 12952 9404 13277 9432
rect 12952 9392 12958 9404
rect 13265 9401 13277 9404
rect 13311 9401 13323 9435
rect 13265 9395 13323 9401
rect 13992 9435 14050 9441
rect 13992 9401 14004 9435
rect 14038 9432 14050 9435
rect 14366 9432 14372 9444
rect 14038 9404 14372 9432
rect 14038 9401 14050 9404
rect 13992 9395 14050 9401
rect 14366 9392 14372 9404
rect 14424 9392 14430 9444
rect 15648 9435 15706 9441
rect 15648 9432 15660 9435
rect 15120 9404 15660 9432
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 14550 9364 14556 9376
rect 10836 9336 14556 9364
rect 10836 9324 10842 9336
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 15120 9373 15148 9404
rect 15648 9401 15660 9404
rect 15694 9432 15706 9435
rect 16114 9432 16120 9444
rect 15694 9404 16120 9432
rect 15694 9401 15706 9404
rect 15648 9395 15706 9401
rect 16114 9392 16120 9404
rect 16172 9392 16178 9444
rect 18138 9392 18144 9444
rect 18196 9432 18202 9444
rect 18316 9435 18374 9441
rect 18316 9432 18328 9435
rect 18196 9404 18328 9432
rect 18196 9392 18202 9404
rect 18316 9401 18328 9404
rect 18362 9432 18374 9435
rect 18506 9432 18512 9444
rect 18362 9404 18512 9432
rect 18362 9401 18374 9404
rect 18316 9395 18374 9401
rect 18506 9392 18512 9404
rect 18564 9392 18570 9444
rect 15105 9367 15163 9373
rect 15105 9333 15117 9367
rect 15151 9333 15163 9367
rect 15105 9327 15163 9333
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 16540 9336 16773 9364
rect 16540 9324 16546 9336
rect 16761 9333 16773 9336
rect 16807 9333 16819 9367
rect 16761 9327 16819 9333
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 19797 9367 19855 9373
rect 19797 9364 19809 9367
rect 17920 9336 19809 9364
rect 17920 9324 17926 9336
rect 19797 9333 19809 9336
rect 19843 9333 19855 9367
rect 20162 9364 20168 9376
rect 20075 9336 20168 9364
rect 19797 9327 19855 9333
rect 20162 9324 20168 9336
rect 20220 9364 20226 9376
rect 20346 9364 20352 9376
rect 20220 9336 20352 9364
rect 20220 9324 20226 9336
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20990 9364 20996 9376
rect 20951 9336 20996 9364
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 10413 9163 10471 9169
rect 10413 9129 10425 9163
rect 10459 9129 10471 9163
rect 10413 9123 10471 9129
rect 10428 9092 10456 9123
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 17405 9163 17463 9169
rect 17405 9160 17417 9163
rect 13044 9132 17417 9160
rect 13044 9120 13050 9132
rect 17405 9129 17417 9132
rect 17451 9129 17463 9163
rect 17405 9123 17463 9129
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 17552 9132 17785 9160
rect 17552 9120 17558 9132
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 17773 9123 17831 9129
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 17920 9132 17965 9160
rect 17920 9120 17926 9132
rect 19150 9120 19156 9172
rect 19208 9160 19214 9172
rect 20533 9163 20591 9169
rect 20533 9160 20545 9163
rect 19208 9132 20545 9160
rect 19208 9120 19214 9132
rect 20533 9129 20545 9132
rect 20579 9129 20591 9163
rect 20533 9123 20591 9129
rect 11054 9092 11060 9104
rect 10428 9064 11060 9092
rect 11054 9052 11060 9064
rect 11112 9092 11118 9104
rect 11698 9092 11704 9104
rect 11112 9064 11704 9092
rect 11112 9052 11118 9064
rect 10594 9024 10600 9036
rect 10555 8996 10600 9024
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11348 9033 11376 9064
rect 11698 9052 11704 9064
rect 11756 9052 11762 9104
rect 15832 9095 15890 9101
rect 15832 9061 15844 9095
rect 15878 9092 15890 9095
rect 16482 9092 16488 9104
rect 15878 9064 16488 9092
rect 15878 9061 15890 9064
rect 15832 9055 15890 9061
rect 16482 9052 16488 9064
rect 16540 9052 16546 9104
rect 18690 9052 18696 9104
rect 18748 9092 18754 9104
rect 18748 9064 19196 9092
rect 18748 9052 18754 9064
rect 11606 9033 11612 9036
rect 11333 9027 11391 9033
rect 11333 8993 11345 9027
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11600 8987 11612 9033
rect 11664 9024 11670 9036
rect 13256 9027 13314 9033
rect 13256 9024 13268 9027
rect 11664 8996 11700 9024
rect 12728 8996 13268 9024
rect 11606 8984 11612 8987
rect 11664 8984 11670 8996
rect 12728 8897 12756 8996
rect 13256 8993 13268 8996
rect 13302 9024 13314 9027
rect 14090 9024 14096 9036
rect 13302 8996 14096 9024
rect 13302 8993 13314 8996
rect 13256 8987 13314 8993
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 15378 8984 15384 9036
rect 15436 9024 15442 9036
rect 19168 9033 19196 9064
rect 15565 9027 15623 9033
rect 15565 9024 15577 9027
rect 15436 8996 15577 9024
rect 15436 8984 15442 8996
rect 15565 8993 15577 8996
rect 15611 8993 15623 9027
rect 15565 8987 15623 8993
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 19420 9027 19478 9033
rect 19420 8993 19432 9027
rect 19466 9024 19478 9027
rect 20530 9024 20536 9036
rect 19466 8996 20536 9024
rect 19466 8993 19478 8996
rect 19420 8987 19478 8993
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 12986 8956 12992 8968
rect 12947 8928 12992 8956
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8956 14703 8959
rect 15102 8956 15108 8968
rect 14691 8928 15108 8956
rect 14691 8925 14703 8928
rect 14645 8919 14703 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 18049 8959 18107 8965
rect 18049 8925 18061 8959
rect 18095 8956 18107 8959
rect 18138 8956 18144 8968
rect 18095 8928 18144 8956
rect 18095 8925 18107 8928
rect 18049 8919 18107 8925
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 18693 8959 18751 8965
rect 18693 8956 18705 8959
rect 18564 8928 18705 8956
rect 18564 8916 18570 8928
rect 18693 8925 18705 8928
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 12713 8891 12771 8897
rect 12713 8857 12725 8891
rect 12759 8857 12771 8891
rect 18874 8888 18880 8900
rect 12713 8851 12771 8857
rect 16500 8860 18880 8888
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 13906 8820 13912 8832
rect 5132 8792 13912 8820
rect 5132 8780 5138 8792
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 14366 8820 14372 8832
rect 14327 8792 14372 8820
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 16500 8820 16528 8860
rect 18874 8848 18880 8860
rect 18932 8848 18938 8900
rect 16942 8820 16948 8832
rect 14516 8792 16528 8820
rect 16903 8792 16948 8820
rect 14516 8780 14522 8792
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 9674 8616 9680 8628
rect 8895 8588 9680 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9784 8588 13952 8616
rect 4890 8508 4896 8560
rect 4948 8548 4954 8560
rect 9784 8548 9812 8588
rect 11606 8548 11612 8560
rect 4948 8520 9812 8548
rect 11567 8520 11612 8548
rect 4948 8508 4954 8520
rect 11606 8508 11612 8520
rect 11664 8548 11670 8560
rect 12986 8548 12992 8560
rect 11664 8520 12992 8548
rect 11664 8508 11670 8520
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 13924 8548 13952 8588
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14737 8619 14795 8625
rect 14737 8616 14749 8619
rect 14056 8588 14749 8616
rect 14056 8576 14062 8588
rect 14737 8585 14749 8588
rect 14783 8585 14795 8619
rect 15562 8616 15568 8628
rect 15523 8588 15568 8616
rect 14737 8579 14795 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 20530 8616 20536 8628
rect 20491 8588 20536 8616
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 16393 8551 16451 8557
rect 13924 8520 15424 8548
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9364 8452 9413 8480
rect 9364 8440 9370 8452
rect 9401 8449 9413 8452
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 15289 8483 15347 8489
rect 15289 8480 15301 8483
rect 14424 8452 15301 8480
rect 14424 8440 14430 8452
rect 15289 8449 15301 8452
rect 15335 8449 15347 8483
rect 15289 8443 15347 8449
rect 10229 8415 10287 8421
rect 10229 8381 10241 8415
rect 10275 8412 10287 8415
rect 11054 8412 11060 8424
rect 10275 8384 11060 8412
rect 10275 8381 10287 8384
rect 10229 8375 10287 8381
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 14458 8412 14464 8424
rect 12943 8384 14464 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 15102 8412 15108 8424
rect 15063 8384 15108 8412
rect 15102 8372 15108 8384
rect 15160 8372 15166 8424
rect 15396 8412 15424 8520
rect 16393 8517 16405 8551
rect 16439 8548 16451 8551
rect 17126 8548 17132 8560
rect 16439 8520 17132 8548
rect 16439 8517 16451 8520
rect 16393 8511 16451 8517
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 16114 8480 16120 8492
rect 16075 8452 16120 8480
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16942 8480 16948 8492
rect 16903 8452 16948 8480
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 18598 8480 18604 8492
rect 18559 8452 18604 8480
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 18831 8452 19288 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 15396 8384 16773 8412
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 18506 8412 18512 8424
rect 18467 8384 18512 8412
rect 16761 8375 16819 8381
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 19153 8415 19211 8421
rect 19153 8412 19165 8415
rect 18748 8384 19165 8412
rect 18748 8372 18754 8384
rect 19153 8381 19165 8384
rect 19199 8381 19211 8415
rect 19260 8412 19288 8452
rect 19420 8415 19478 8421
rect 19420 8412 19432 8415
rect 19260 8384 19432 8412
rect 19153 8375 19211 8381
rect 19420 8381 19432 8384
rect 19466 8412 19478 8415
rect 19886 8412 19892 8424
rect 19466 8384 19892 8412
rect 19466 8381 19478 8384
rect 19420 8375 19478 8381
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 9309 8347 9367 8353
rect 9309 8313 9321 8347
rect 9355 8344 9367 8347
rect 9398 8344 9404 8356
rect 9355 8316 9404 8344
rect 9355 8313 9367 8316
rect 9309 8307 9367 8313
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 10496 8347 10554 8353
rect 10496 8313 10508 8347
rect 10542 8344 10554 8347
rect 10962 8344 10968 8356
rect 10542 8316 10968 8344
rect 10542 8313 10554 8316
rect 10496 8307 10554 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 11885 8347 11943 8353
rect 11885 8313 11897 8347
rect 11931 8344 11943 8347
rect 12802 8344 12808 8356
rect 11931 8316 12808 8344
rect 11931 8313 11943 8316
rect 11885 8307 11943 8313
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 13906 8304 13912 8356
rect 13964 8344 13970 8356
rect 16022 8344 16028 8356
rect 13964 8316 15884 8344
rect 15983 8316 16028 8344
rect 13964 8304 13970 8316
rect 9214 8276 9220 8288
rect 9175 8248 9220 8276
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 14182 8276 14188 8288
rect 14143 8248 14188 8276
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 15197 8279 15255 8285
rect 15197 8276 15209 8279
rect 15068 8248 15209 8276
rect 15068 8236 15074 8248
rect 15197 8245 15209 8248
rect 15243 8245 15255 8279
rect 15856 8276 15884 8316
rect 16022 8304 16028 8316
rect 16080 8344 16086 8356
rect 16482 8344 16488 8356
rect 16080 8316 16488 8344
rect 16080 8304 16086 8316
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 17034 8344 17040 8356
rect 16899 8316 17040 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 15933 8279 15991 8285
rect 15933 8276 15945 8279
rect 15856 8248 15945 8276
rect 15197 8239 15255 8245
rect 15933 8245 15945 8248
rect 15979 8245 15991 8279
rect 17218 8276 17224 8288
rect 17179 8248 17224 8276
rect 15933 8239 15991 8245
rect 17218 8236 17224 8248
rect 17276 8236 17282 8288
rect 18138 8276 18144 8288
rect 18099 8248 18144 8276
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 18782 8276 18788 8288
rect 18656 8248 18788 8276
rect 18656 8236 18662 8248
rect 18782 8236 18788 8248
rect 18840 8236 18846 8288
rect 19610 8236 19616 8288
rect 19668 8276 19674 8288
rect 19702 8276 19708 8288
rect 19668 8248 19708 8276
rect 19668 8236 19674 8248
rect 19702 8236 19708 8248
rect 19760 8236 19766 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 9306 8072 9312 8084
rect 9267 8044 9312 8072
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 10962 8032 10968 8084
rect 11020 8072 11026 8084
rect 11057 8075 11115 8081
rect 11057 8072 11069 8075
rect 11020 8044 11069 8072
rect 11020 8032 11026 8044
rect 11057 8041 11069 8044
rect 11103 8041 11115 8075
rect 11057 8035 11115 8041
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 15010 8072 15016 8084
rect 13587 8044 15016 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15473 8075 15531 8081
rect 15473 8041 15485 8075
rect 15519 8072 15531 8075
rect 16298 8072 16304 8084
rect 15519 8044 16304 8072
rect 15519 8041 15531 8044
rect 15473 8035 15531 8041
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 9324 8004 9352 8032
rect 9922 8007 9980 8013
rect 9922 8004 9934 8007
rect 7944 7976 9076 8004
rect 9324 7976 9934 8004
rect 7944 7945 7972 7976
rect 7929 7939 7987 7945
rect 7929 7905 7941 7939
rect 7975 7905 7987 7939
rect 7929 7899 7987 7905
rect 8196 7939 8254 7945
rect 8196 7905 8208 7939
rect 8242 7936 8254 7939
rect 8938 7936 8944 7948
rect 8242 7908 8944 7936
rect 8242 7905 8254 7908
rect 8196 7899 8254 7905
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 9048 7936 9076 7976
rect 9922 7973 9934 7976
rect 9968 7973 9980 8007
rect 9922 7967 9980 7973
rect 13909 8007 13967 8013
rect 13909 7973 13921 8007
rect 13955 8004 13967 8007
rect 13998 8004 14004 8016
rect 13955 7976 14004 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 13998 7964 14004 7976
rect 14056 7964 14062 8016
rect 16200 8007 16258 8013
rect 16200 7973 16212 8007
rect 16246 8004 16258 8007
rect 16942 8004 16948 8016
rect 16246 7976 16948 8004
rect 16246 7973 16258 7976
rect 16200 7967 16258 7973
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 9674 7936 9680 7948
rect 9048 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7936 9738 7948
rect 11054 7936 11060 7948
rect 9732 7908 11060 7936
rect 9732 7896 9738 7908
rect 11054 7896 11060 7908
rect 11112 7936 11118 7948
rect 11882 7936 11888 7948
rect 11112 7908 11888 7936
rect 11112 7896 11118 7908
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12152 7939 12210 7945
rect 12152 7905 12164 7939
rect 12198 7936 12210 7939
rect 12710 7936 12716 7948
rect 12198 7908 12716 7936
rect 12198 7905 12210 7908
rect 12152 7899 12210 7905
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 14240 7908 15669 7936
rect 14240 7896 14246 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15933 7939 15991 7945
rect 15933 7905 15945 7939
rect 15979 7936 15991 7939
rect 16022 7936 16028 7948
rect 15979 7908 16028 7936
rect 15979 7905 15991 7908
rect 15933 7899 15991 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 17589 7939 17647 7945
rect 17589 7905 17601 7939
rect 17635 7936 17647 7939
rect 18138 7936 18144 7948
rect 17635 7908 18144 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 18325 7939 18383 7945
rect 18325 7905 18337 7939
rect 18371 7936 18383 7939
rect 18782 7936 18788 7948
rect 18371 7908 18788 7936
rect 18371 7905 18383 7908
rect 18325 7899 18383 7905
rect 18782 7896 18788 7908
rect 18840 7896 18846 7948
rect 20165 7939 20223 7945
rect 20165 7905 20177 7939
rect 20211 7936 20223 7939
rect 20346 7936 20352 7948
rect 20211 7908 20352 7936
rect 20211 7905 20223 7908
rect 20165 7899 20223 7905
rect 20346 7896 20352 7908
rect 20404 7896 20410 7948
rect 14001 7871 14059 7877
rect 14001 7837 14013 7871
rect 14047 7837 14059 7871
rect 14001 7831 14059 7837
rect 14016 7800 14044 7831
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 14148 7840 14193 7868
rect 14148 7828 14154 7840
rect 16942 7828 16948 7880
rect 17000 7868 17006 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17000 7840 17785 7868
rect 17000 7828 17006 7840
rect 17773 7837 17785 7840
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 18601 7871 18659 7877
rect 18601 7837 18613 7871
rect 18647 7868 18659 7871
rect 18874 7868 18880 7880
rect 18647 7840 18880 7868
rect 18647 7837 18659 7840
rect 18601 7831 18659 7837
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19208 7840 19257 7868
rect 19208 7828 19214 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 20254 7868 20260 7880
rect 20215 7840 20260 7868
rect 19245 7831 19303 7837
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7868 20499 7871
rect 20530 7868 20536 7880
rect 20487 7840 20536 7868
rect 20487 7837 20499 7840
rect 20441 7831 20499 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 14458 7800 14464 7812
rect 14016 7772 14464 7800
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 13262 7732 13268 7744
rect 13223 7704 13268 7732
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 17310 7732 17316 7744
rect 17271 7704 17316 7732
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 19242 7692 19248 7744
rect 19300 7732 19306 7744
rect 19797 7735 19855 7741
rect 19797 7732 19809 7735
rect 19300 7704 19809 7732
rect 19300 7692 19306 7704
rect 19797 7701 19809 7704
rect 19843 7701 19855 7735
rect 19797 7695 19855 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 12492 7500 12537 7528
rect 15672 7500 16681 7528
rect 12492 7488 12498 7500
rect 10505 7463 10563 7469
rect 10505 7429 10517 7463
rect 10551 7460 10563 7463
rect 10551 7432 11468 7460
rect 10551 7429 10563 7432
rect 10505 7423 10563 7429
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9272 7364 9413 7392
rect 9272 7352 9278 7364
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 11020 7364 11069 7392
rect 11020 7352 11026 7364
rect 11057 7361 11069 7364
rect 11103 7361 11115 7395
rect 11440 7392 11468 7432
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 11440 7364 12909 7392
rect 11057 7355 11115 7361
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13044 7364 13089 7392
rect 13044 7352 13050 7364
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7293 11759 7327
rect 12802 7324 12808 7336
rect 12763 7296 12808 7324
rect 11701 7287 11759 7293
rect 10042 7216 10048 7268
rect 10100 7256 10106 7268
rect 10594 7256 10600 7268
rect 10100 7228 10600 7256
rect 10100 7216 10106 7228
rect 10594 7216 10600 7228
rect 10652 7256 10658 7268
rect 11716 7256 11744 7287
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7324 13323 7327
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 13311 7296 13461 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 13449 7293 13461 7296
rect 13495 7293 13507 7327
rect 13449 7287 13507 7293
rect 13716 7327 13774 7333
rect 13716 7293 13728 7327
rect 13762 7324 13774 7327
rect 15672 7324 15700 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 18782 7528 18788 7540
rect 18743 7500 18788 7528
rect 16669 7491 16727 7497
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 19794 7528 19800 7540
rect 19755 7500 19800 7528
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 15749 7463 15807 7469
rect 15749 7429 15761 7463
rect 15795 7460 15807 7463
rect 20898 7460 20904 7472
rect 15795 7432 18092 7460
rect 15795 7429 15807 7432
rect 15749 7423 15807 7429
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 17310 7392 17316 7404
rect 16715 7364 17316 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 13762 7296 15700 7324
rect 13762 7293 13774 7296
rect 13716 7287 13774 7293
rect 10652 7228 11560 7256
rect 11716 7228 13492 7256
rect 10652 7216 10658 7228
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 10873 7191 10931 7197
rect 10873 7188 10885 7191
rect 8628 7160 10885 7188
rect 8628 7148 8634 7160
rect 10873 7157 10885 7160
rect 10919 7157 10931 7191
rect 10873 7151 10931 7157
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11532 7197 11560 7228
rect 11517 7191 11575 7197
rect 11020 7160 11065 7188
rect 11020 7148 11026 7160
rect 11517 7157 11529 7191
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 11940 7160 13277 7188
rect 11940 7148 11946 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13464 7188 13492 7228
rect 13538 7216 13544 7268
rect 13596 7256 13602 7268
rect 16316 7256 16344 7355
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 17218 7324 17224 7336
rect 17175 7296 17224 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 17218 7284 17224 7296
rect 17276 7284 17282 7336
rect 18064 7333 18092 7432
rect 18340 7432 20904 7460
rect 18340 7401 18368 7432
rect 20898 7420 20904 7432
rect 20956 7420 20962 7472
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7361 18383 7395
rect 19242 7392 19248 7404
rect 19203 7364 19248 7392
rect 18325 7355 18383 7361
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 19334 7352 19340 7404
rect 19392 7392 19398 7404
rect 19392 7364 19437 7392
rect 19392 7352 19398 7364
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20349 7395 20407 7401
rect 20349 7392 20361 7395
rect 20220 7364 20361 7392
rect 20220 7352 20226 7364
rect 20349 7361 20361 7364
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 19150 7324 19156 7336
rect 19111 7296 19156 7324
rect 18049 7287 18107 7293
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19518 7324 19524 7336
rect 19260 7296 19524 7324
rect 16574 7256 16580 7268
rect 13596 7228 14872 7256
rect 16316 7228 16580 7256
rect 13596 7216 13602 7228
rect 14182 7188 14188 7200
rect 13464 7160 14188 7188
rect 13265 7151 13323 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14844 7197 14872 7228
rect 16574 7216 16580 7228
rect 16632 7216 16638 7268
rect 19260 7256 19288 7296
rect 19518 7284 19524 7296
rect 19576 7284 19582 7336
rect 16776 7228 19288 7256
rect 14829 7191 14887 7197
rect 14829 7157 14841 7191
rect 14875 7157 14887 7191
rect 16114 7188 16120 7200
rect 16075 7160 16120 7188
rect 14829 7151 14887 7157
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 16209 7191 16267 7197
rect 16209 7157 16221 7191
rect 16255 7188 16267 7191
rect 16666 7188 16672 7200
rect 16255 7160 16672 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 16776 7197 16804 7228
rect 19334 7216 19340 7268
rect 19392 7256 19398 7268
rect 20257 7259 20315 7265
rect 20257 7256 20269 7259
rect 19392 7228 20269 7256
rect 19392 7216 19398 7228
rect 20257 7225 20269 7228
rect 20303 7225 20315 7259
rect 20257 7219 20315 7225
rect 16761 7191 16819 7197
rect 16761 7157 16773 7191
rect 16807 7157 16819 7191
rect 16761 7151 16819 7157
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 17221 7191 17279 7197
rect 17221 7188 17233 7191
rect 17184 7160 17233 7188
rect 17184 7148 17190 7160
rect 17221 7157 17233 7160
rect 17267 7157 17279 7191
rect 17221 7151 17279 7157
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 18782 7188 18788 7200
rect 18656 7160 18788 7188
rect 18656 7148 18662 7160
rect 18782 7148 18788 7160
rect 18840 7148 18846 7200
rect 19518 7148 19524 7200
rect 19576 7188 19582 7200
rect 20165 7191 20223 7197
rect 20165 7188 20177 7191
rect 19576 7160 20177 7188
rect 19576 7148 19582 7160
rect 20165 7157 20177 7160
rect 20211 7157 20223 7191
rect 20165 7151 20223 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 11241 6987 11299 6993
rect 11241 6953 11253 6987
rect 11287 6984 11299 6987
rect 11882 6984 11888 6996
rect 11287 6956 11888 6984
rect 11287 6953 11299 6956
rect 11241 6947 11299 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12710 6984 12716 6996
rect 12671 6956 12716 6984
rect 12710 6944 12716 6956
rect 12768 6984 12774 6996
rect 15289 6987 15347 6993
rect 12768 6956 13768 6984
rect 12768 6944 12774 6956
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 2884 6888 13185 6916
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 2884 6848 2912 6888
rect 13173 6885 13185 6888
rect 13219 6885 13231 6919
rect 13173 6879 13231 6885
rect 13265 6919 13323 6925
rect 13265 6885 13277 6919
rect 13311 6916 13323 6919
rect 13446 6916 13452 6928
rect 13311 6888 13452 6916
rect 13311 6885 13323 6888
rect 13265 6879 13323 6885
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 13740 6916 13768 6956
rect 15289 6953 15301 6987
rect 15335 6984 15347 6987
rect 16114 6984 16120 6996
rect 15335 6956 16120 6984
rect 15335 6953 15347 6956
rect 15289 6947 15347 6953
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 15654 6916 15660 6928
rect 13740 6888 14136 6916
rect 15615 6888 15660 6916
rect 9674 6848 9680 6860
rect 2740 6820 2912 6848
rect 9635 6820 9680 6848
rect 2740 6808 2746 6820
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 9944 6851 10002 6857
rect 9944 6817 9956 6851
rect 9990 6848 10002 6851
rect 10226 6848 10232 6860
rect 9990 6820 10232 6848
rect 9990 6817 10002 6820
rect 9944 6811 10002 6817
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 11600 6851 11658 6857
rect 11600 6848 11612 6851
rect 11072 6820 11612 6848
rect 9122 6780 9128 6792
rect 9083 6752 9128 6780
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 11072 6721 11100 6820
rect 11600 6817 11612 6820
rect 11646 6848 11658 6851
rect 13998 6848 14004 6860
rect 11646 6820 13400 6848
rect 13959 6820 14004 6848
rect 11646 6817 11658 6820
rect 11600 6811 11658 6817
rect 13372 6789 13400 6820
rect 13998 6808 14004 6820
rect 14056 6808 14062 6860
rect 14108 6848 14136 6888
rect 15654 6876 15660 6888
rect 15712 6876 15718 6928
rect 14108 6820 14228 6848
rect 14200 6789 14228 6820
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 16356 6820 16497 6848
rect 16356 6808 16362 6820
rect 16485 6817 16497 6820
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16936 6851 16994 6857
rect 16936 6848 16948 6851
rect 16632 6820 16948 6848
rect 16632 6808 16638 6820
rect 16936 6817 16948 6820
rect 16982 6848 16994 6851
rect 17494 6848 17500 6860
rect 16982 6820 17500 6848
rect 16982 6817 16994 6820
rect 16936 6811 16994 6817
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 18785 6851 18843 6857
rect 18785 6848 18797 6851
rect 18748 6820 18797 6848
rect 18748 6808 18754 6820
rect 18785 6817 18797 6820
rect 18831 6817 18843 6851
rect 18785 6811 18843 6817
rect 19052 6851 19110 6857
rect 19052 6817 19064 6851
rect 19098 6848 19110 6851
rect 19426 6848 19432 6860
rect 19098 6820 19432 6848
rect 19098 6817 19110 6820
rect 19052 6811 19110 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 11287 6752 11345 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11333 6749 11345 6752
rect 11379 6749 11391 6783
rect 13357 6783 13415 6789
rect 11333 6743 11391 6749
rect 12820 6752 13308 6780
rect 12820 6721 12848 6752
rect 11057 6715 11115 6721
rect 11057 6681 11069 6715
rect 11103 6681 11115 6715
rect 11057 6675 11115 6681
rect 12805 6715 12863 6721
rect 12805 6681 12817 6715
rect 12851 6681 12863 6715
rect 13280 6712 13308 6752
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13357 6743 13415 6749
rect 13464 6752 14105 6780
rect 13464 6712 13492 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6749 14243 6783
rect 15746 6780 15752 6792
rect 15707 6752 15752 6780
rect 14185 6743 14243 6749
rect 15746 6740 15752 6752
rect 15804 6740 15810 6792
rect 15930 6780 15936 6792
rect 15891 6752 15936 6780
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16669 6783 16727 6789
rect 16669 6749 16681 6783
rect 16715 6749 16727 6783
rect 16669 6743 16727 6749
rect 13630 6712 13636 6724
rect 13280 6684 13492 6712
rect 13591 6684 13636 6712
rect 12805 6675 12863 6681
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 13446 6644 13452 6656
rect 11020 6616 13452 6644
rect 11020 6604 11026 6616
rect 13446 6604 13452 6616
rect 13504 6644 13510 6656
rect 15102 6644 15108 6656
rect 13504 6616 15108 6644
rect 13504 6604 13510 6616
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 16022 6604 16028 6656
rect 16080 6644 16086 6656
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 16080 6616 16313 6644
rect 16080 6604 16086 6616
rect 16301 6613 16313 6616
rect 16347 6644 16359 6647
rect 16684 6644 16712 6743
rect 16850 6644 16856 6656
rect 16347 6616 16856 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 18012 6616 18061 6644
rect 18012 6604 18018 6616
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 20162 6644 20168 6656
rect 20123 6616 20168 6644
rect 18049 6607 18107 6613
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 10226 6440 10232 6452
rect 10187 6412 10232 6440
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 10689 6443 10747 6449
rect 10689 6409 10701 6443
rect 10735 6440 10747 6443
rect 11790 6440 11796 6452
rect 10735 6412 11796 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13814 6440 13820 6452
rect 13219 6412 13820 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 16482 6400 16488 6452
rect 16540 6440 16546 6452
rect 17494 6440 17500 6452
rect 16540 6412 17356 6440
rect 17455 6412 17500 6440
rect 16540 6400 16546 6412
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 13906 6372 13912 6384
rect 13320 6344 13912 6372
rect 13320 6332 13326 6344
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 17328 6372 17356 6412
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 19242 6440 19248 6452
rect 18064 6412 19248 6440
rect 18064 6372 18092 6412
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 20254 6372 20260 6384
rect 17328 6344 18092 6372
rect 20167 6344 20260 6372
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11606 6304 11612 6316
rect 11379 6276 11612 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 13722 6304 13728 6316
rect 12360 6276 13728 6304
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6880 6208 7205 6236
rect 6880 6196 6886 6208
rect 7193 6205 7205 6208
rect 7239 6236 7251 6239
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 7239 6208 8861 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 8849 6205 8861 6208
rect 8895 6236 8907 6239
rect 9674 6236 9680 6248
rect 8895 6208 9680 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 12360 6236 12388 6276
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 17954 6264 17960 6316
rect 18012 6304 18018 6316
rect 18012 6276 18184 6304
rect 18012 6264 18018 6276
rect 10744 6208 12388 6236
rect 12437 6239 12495 6245
rect 10744 6196 10750 6208
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 13998 6236 14004 6248
rect 12483 6208 14004 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14461 6239 14519 6245
rect 14461 6205 14473 6239
rect 14507 6236 14519 6239
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 14507 6208 16129 6236
rect 14507 6205 14519 6208
rect 14461 6199 14519 6205
rect 16117 6205 16129 6208
rect 16163 6236 16175 6239
rect 16850 6236 16856 6248
rect 16163 6208 16856 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 17310 6236 17316 6248
rect 16908 6208 17316 6236
rect 16908 6196 16914 6208
rect 17310 6196 17316 6208
rect 17368 6236 17374 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17368 6208 18061 6236
rect 17368 6196 17374 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18156 6236 18184 6276
rect 18305 6239 18363 6245
rect 18305 6236 18317 6239
rect 18156 6208 18317 6236
rect 18049 6199 18107 6205
rect 18305 6205 18317 6208
rect 18351 6236 18363 6239
rect 20180 6236 20208 6344
rect 20254 6332 20260 6344
rect 20312 6372 20318 6384
rect 20312 6344 20392 6372
rect 20312 6332 20318 6344
rect 20364 6313 20392 6344
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6273 20407 6307
rect 20349 6267 20407 6273
rect 18351 6208 20208 6236
rect 18351 6205 18363 6208
rect 18305 6199 18363 6205
rect 7460 6171 7518 6177
rect 7460 6137 7472 6171
rect 7506 6168 7518 6171
rect 7742 6168 7748 6180
rect 7506 6140 7748 6168
rect 7506 6137 7518 6140
rect 7460 6131 7518 6137
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 9030 6168 9036 6180
rect 8588 6140 9036 6168
rect 8588 6109 8616 6140
rect 9030 6128 9036 6140
rect 9088 6177 9094 6180
rect 9088 6171 9152 6177
rect 9088 6137 9106 6171
rect 9140 6137 9152 6171
rect 9088 6131 9152 6137
rect 9088 6128 9094 6131
rect 12618 6128 12624 6180
rect 12676 6168 12682 6180
rect 13541 6171 13599 6177
rect 13541 6168 13553 6171
rect 12676 6140 13553 6168
rect 12676 6128 12682 6140
rect 13541 6137 13553 6140
rect 13587 6137 13599 6171
rect 13541 6131 13599 6137
rect 14728 6171 14786 6177
rect 14728 6137 14740 6171
rect 14774 6168 14786 6171
rect 15010 6168 15016 6180
rect 14774 6140 15016 6168
rect 14774 6137 14786 6140
rect 14728 6131 14786 6137
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 15930 6168 15936 6180
rect 15843 6140 15936 6168
rect 8573 6103 8631 6109
rect 8573 6069 8585 6103
rect 8619 6069 8631 6103
rect 11054 6100 11060 6112
rect 11015 6072 11060 6100
rect 8573 6063 8631 6069
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 13630 6100 13636 6112
rect 11204 6072 11249 6100
rect 13591 6072 13636 6100
rect 11204 6060 11210 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 15856 6109 15884 6140
rect 15930 6128 15936 6140
rect 15988 6168 15994 6180
rect 16384 6171 16442 6177
rect 16384 6168 16396 6171
rect 15988 6140 16396 6168
rect 15988 6128 15994 6140
rect 16384 6137 16396 6140
rect 16430 6168 16442 6171
rect 17770 6168 17776 6180
rect 16430 6140 17776 6168
rect 16430 6137 16442 6140
rect 16384 6131 16442 6137
rect 17770 6128 17776 6140
rect 17828 6128 17834 6180
rect 18064 6168 18092 6199
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 20717 6239 20775 6245
rect 20717 6236 20729 6239
rect 20680 6208 20729 6236
rect 20680 6196 20686 6208
rect 20717 6205 20729 6208
rect 20763 6205 20775 6239
rect 20717 6199 20775 6205
rect 18690 6168 18696 6180
rect 18064 6140 18696 6168
rect 18690 6128 18696 6140
rect 18748 6128 18754 6180
rect 20165 6171 20223 6177
rect 20165 6168 20177 6171
rect 18800 6140 20177 6168
rect 15841 6103 15899 6109
rect 15841 6069 15853 6103
rect 15887 6069 15899 6103
rect 15841 6063 15899 6069
rect 17126 6060 17132 6112
rect 17184 6100 17190 6112
rect 18800 6100 18828 6140
rect 20165 6137 20177 6140
rect 20211 6137 20223 6171
rect 20165 6131 20223 6137
rect 19426 6100 19432 6112
rect 17184 6072 18828 6100
rect 19387 6072 19432 6100
rect 17184 6060 17190 6072
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 19702 6100 19708 6112
rect 19663 6072 19708 6100
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 19852 6072 20085 6100
rect 19852 6060 19858 6072
rect 20073 6069 20085 6072
rect 20119 6069 20131 6103
rect 20898 6100 20904 6112
rect 20859 6072 20904 6100
rect 20073 6063 20131 6069
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7708 5868 8033 5896
rect 7708 5856 7714 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 9180 5868 10057 5896
rect 9180 5856 9186 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 10045 5859 10103 5865
rect 16209 5899 16267 5905
rect 16209 5865 16221 5899
rect 16255 5896 16267 5899
rect 17589 5899 17647 5905
rect 17589 5896 17601 5899
rect 16255 5868 17601 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 17589 5865 17601 5868
rect 17635 5865 17647 5899
rect 17589 5859 17647 5865
rect 18693 5899 18751 5905
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 19518 5896 19524 5908
rect 18739 5868 19524 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 19610 5856 19616 5908
rect 19668 5896 19674 5908
rect 20073 5899 20131 5905
rect 20073 5896 20085 5899
rect 19668 5868 20085 5896
rect 19668 5856 19674 5868
rect 20073 5865 20085 5868
rect 20119 5865 20131 5899
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20073 5859 20131 5865
rect 20180 5868 20913 5896
rect 1210 5788 1216 5840
rect 1268 5828 1274 5840
rect 12342 5828 12348 5840
rect 1268 5800 12348 5828
rect 1268 5788 1274 5800
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 12434 5788 12440 5840
rect 12492 5828 12498 5840
rect 14461 5831 14519 5837
rect 14461 5828 14473 5831
rect 12492 5800 14473 5828
rect 12492 5788 12498 5800
rect 14461 5797 14473 5800
rect 14507 5797 14519 5831
rect 14461 5791 14519 5797
rect 15102 5788 15108 5840
rect 15160 5828 15166 5840
rect 19061 5831 19119 5837
rect 15160 5800 16712 5828
rect 15160 5788 15166 5800
rect 6632 5763 6690 5769
rect 6632 5729 6644 5763
rect 6678 5760 6690 5763
rect 7190 5760 7196 5772
rect 6678 5732 7196 5760
rect 6678 5729 6690 5732
rect 6632 5723 6690 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 8389 5763 8447 5769
rect 8389 5729 8401 5763
rect 8435 5760 8447 5763
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8435 5732 9045 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9033 5723 9091 5729
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 11037 5763 11095 5769
rect 11037 5760 11049 5763
rect 10744 5732 11049 5760
rect 10744 5720 10750 5732
rect 11037 5729 11049 5732
rect 11083 5729 11095 5763
rect 11037 5723 11095 5729
rect 12888 5763 12946 5769
rect 12888 5729 12900 5763
rect 12934 5760 12946 5763
rect 13446 5760 13452 5772
rect 12934 5732 13452 5760
rect 12934 5729 12946 5732
rect 12888 5723 12946 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 13964 5732 14688 5760
rect 13964 5720 13970 5732
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6380 5556 6408 5655
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 7432 5664 8493 5692
rect 7432 5652 7438 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 8573 5655 8631 5661
rect 7742 5624 7748 5636
rect 7703 5596 7748 5624
rect 7742 5584 7748 5596
rect 7800 5624 7806 5636
rect 8588 5624 8616 5655
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10781 5695 10839 5701
rect 10284 5664 10329 5692
rect 10284 5652 10290 5664
rect 10781 5661 10793 5695
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 7800 5596 8616 5624
rect 9677 5627 9735 5633
rect 7800 5584 7806 5596
rect 9677 5593 9689 5627
rect 9723 5624 9735 5627
rect 9766 5624 9772 5636
rect 9723 5596 9772 5624
rect 9723 5593 9735 5596
rect 9677 5587 9735 5593
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 6730 5556 6736 5568
rect 6380 5528 6736 5556
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 10796 5556 10824 5655
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 11848 5664 12633 5692
rect 11848 5652 11854 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 14660 5701 14688 5732
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 16684 5769 16712 5800
rect 19061 5797 19073 5831
rect 19107 5828 19119 5831
rect 20180 5828 20208 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 19107 5800 20208 5828
rect 19107 5797 19119 5800
rect 19061 5791 19119 5797
rect 16577 5763 16635 5769
rect 16577 5760 16589 5763
rect 16540 5732 16589 5760
rect 16540 5720 16546 5732
rect 16577 5729 16589 5732
rect 16623 5729 16635 5763
rect 16577 5723 16635 5729
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5760 16727 5763
rect 16850 5760 16856 5772
rect 16715 5732 16856 5760
rect 16715 5729 16727 5732
rect 16669 5723 16727 5729
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 19794 5760 19800 5772
rect 19260 5732 19800 5760
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14516 5664 14565 5692
rect 14516 5652 14522 5664
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 16758 5692 16764 5704
rect 16719 5664 16764 5692
rect 14645 5655 14703 5661
rect 13722 5584 13728 5636
rect 13780 5624 13786 5636
rect 14001 5627 14059 5633
rect 14001 5624 14013 5627
rect 13780 5596 14013 5624
rect 13780 5584 13786 5596
rect 14001 5593 14013 5596
rect 14047 5593 14059 5627
rect 14568 5624 14596 5655
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 17218 5652 17224 5704
rect 17276 5652 17282 5704
rect 17678 5692 17684 5704
rect 17639 5664 17684 5692
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 17828 5664 17873 5692
rect 17828 5652 17834 5664
rect 18506 5652 18512 5704
rect 18564 5692 18570 5704
rect 19153 5695 19211 5701
rect 19153 5692 19165 5695
rect 18564 5664 19165 5692
rect 18564 5652 18570 5664
rect 19153 5661 19165 5664
rect 19199 5661 19211 5695
rect 19153 5655 19211 5661
rect 17126 5624 17132 5636
rect 14568 5596 17132 5624
rect 14001 5587 14059 5593
rect 17126 5584 17132 5596
rect 17184 5584 17190 5636
rect 17236 5624 17264 5652
rect 19260 5624 19288 5732
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 19996 5732 20177 5760
rect 19337 5695 19395 5701
rect 19337 5661 19349 5695
rect 19383 5692 19395 5695
rect 19426 5692 19432 5704
rect 19383 5664 19432 5692
rect 19383 5661 19395 5664
rect 19337 5655 19395 5661
rect 19426 5652 19432 5664
rect 19484 5692 19490 5704
rect 19886 5692 19892 5704
rect 19484 5664 19892 5692
rect 19484 5652 19490 5664
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 19996 5624 20024 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 20254 5692 20260 5704
rect 20215 5664 20260 5692
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 17236 5596 19288 5624
rect 19628 5596 20024 5624
rect 11882 5556 11888 5568
rect 10796 5528 11888 5556
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12158 5556 12164 5568
rect 12119 5528 12164 5556
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 13354 5516 13360 5568
rect 13412 5556 13418 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13412 5528 14105 5556
rect 13412 5516 13418 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 16724 5528 17233 5556
rect 16724 5516 16730 5528
rect 17221 5525 17233 5528
rect 17267 5525 17279 5559
rect 17221 5519 17279 5525
rect 18690 5516 18696 5568
rect 18748 5556 18754 5568
rect 19628 5556 19656 5596
rect 18748 5528 19656 5556
rect 19705 5559 19763 5565
rect 18748 5516 18754 5528
rect 19705 5525 19717 5559
rect 19751 5556 19763 5559
rect 19794 5556 19800 5568
rect 19751 5528 19800 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 8481 5355 8539 5361
rect 8481 5321 8493 5355
rect 8527 5352 8539 5355
rect 10134 5352 10140 5364
rect 8527 5324 10140 5352
rect 8527 5321 8539 5324
rect 8481 5315 8539 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 12618 5352 12624 5364
rect 12579 5324 12624 5352
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 13630 5352 13636 5364
rect 13591 5324 13636 5352
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 14645 5355 14703 5361
rect 14645 5321 14657 5355
rect 14691 5352 14703 5355
rect 15746 5352 15752 5364
rect 14691 5324 15752 5352
rect 14691 5321 14703 5324
rect 14645 5315 14703 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16209 5355 16267 5361
rect 16209 5321 16221 5355
rect 16255 5352 16267 5355
rect 17678 5352 17684 5364
rect 16255 5324 17684 5352
rect 16255 5321 16267 5324
rect 16209 5315 16267 5321
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 18325 5355 18383 5361
rect 18325 5321 18337 5355
rect 18371 5352 18383 5355
rect 19058 5352 19064 5364
rect 18371 5324 19064 5352
rect 18371 5321 18383 5324
rect 18325 5315 18383 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19334 5352 19340 5364
rect 19295 5324 19340 5352
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9953 5287 10011 5293
rect 9953 5284 9965 5287
rect 9732 5256 9965 5284
rect 9732 5244 9738 5256
rect 9953 5253 9965 5256
rect 9999 5253 10011 5287
rect 9953 5247 10011 5253
rect 9030 5216 9036 5228
rect 8991 5188 9036 5216
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9968 5216 9996 5247
rect 15010 5244 15016 5296
rect 15068 5284 15074 5296
rect 15068 5256 16804 5284
rect 15068 5244 15074 5256
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9968 5188 10241 5216
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5216 13323 5219
rect 13538 5216 13544 5228
rect 13311 5188 13544 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 13538 5176 13544 5188
rect 13596 5216 13602 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13596 5188 14197 5216
rect 13596 5176 13602 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5216 14611 5219
rect 15102 5216 15108 5228
rect 14599 5188 15108 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 15304 5225 15332 5256
rect 16776 5228 16804 5256
rect 15289 5219 15347 5225
rect 15289 5185 15301 5219
rect 15335 5185 15347 5219
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15289 5179 15347 5185
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 16758 5216 16764 5228
rect 16719 5188 16764 5216
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 17586 5176 17592 5228
rect 17644 5216 17650 5228
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 17644 5188 18889 5216
rect 17644 5176 17650 5188
rect 18877 5185 18889 5188
rect 18923 5185 18935 5219
rect 19794 5216 19800 5228
rect 19755 5188 19800 5216
rect 18877 5179 18935 5185
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 19944 5188 19989 5216
rect 19944 5176 19950 5188
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10100 5120 10149 5148
rect 10100 5108 10106 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 14093 5151 14151 5157
rect 14093 5117 14105 5151
rect 14139 5148 14151 5151
rect 14366 5148 14372 5160
rect 14139 5120 14372 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 14366 5108 14372 5120
rect 14424 5148 14430 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 14424 5120 16681 5148
rect 14424 5108 14430 5120
rect 16669 5117 16681 5120
rect 16715 5148 16727 5151
rect 18782 5148 18788 5160
rect 16715 5120 18788 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 18782 5108 18788 5120
rect 18840 5148 18846 5160
rect 19702 5148 19708 5160
rect 18840 5120 19012 5148
rect 19663 5120 19708 5148
rect 18840 5108 18846 5120
rect 7092 5083 7150 5089
rect 7092 5049 7104 5083
rect 7138 5080 7150 5083
rect 10496 5083 10554 5089
rect 7138 5052 10088 5080
rect 7138 5049 7150 5052
rect 7092 5043 7150 5049
rect 7190 4972 7196 5024
rect 7248 5012 7254 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 7248 4984 8217 5012
rect 7248 4972 7254 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8205 4975 8263 4981
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 8941 5015 8999 5021
rect 8941 4981 8953 5015
rect 8987 5012 8999 5015
rect 9858 5012 9864 5024
rect 8987 4984 9864 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10060 5012 10088 5052
rect 10496 5049 10508 5083
rect 10542 5080 10554 5083
rect 11238 5080 11244 5092
rect 10542 5052 11244 5080
rect 10542 5049 10554 5052
rect 10496 5043 10554 5049
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 11698 5040 11704 5092
rect 11756 5080 11762 5092
rect 13081 5083 13139 5089
rect 13081 5080 13093 5083
rect 11756 5052 13093 5080
rect 11756 5040 11762 5052
rect 13081 5049 13093 5052
rect 13127 5049 13139 5083
rect 13081 5043 13139 5049
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14001 5083 14059 5089
rect 14001 5080 14013 5083
rect 13872 5052 14013 5080
rect 13872 5040 13878 5052
rect 14001 5049 14013 5052
rect 14047 5080 14059 5083
rect 14553 5083 14611 5089
rect 14553 5080 14565 5083
rect 14047 5052 14565 5080
rect 14047 5049 14059 5052
rect 14001 5043 14059 5049
rect 14553 5049 14565 5052
rect 14599 5049 14611 5083
rect 14553 5043 14611 5049
rect 17678 5040 17684 5092
rect 17736 5080 17742 5092
rect 18693 5083 18751 5089
rect 18693 5080 18705 5083
rect 17736 5052 18705 5080
rect 17736 5040 17742 5052
rect 18693 5049 18705 5052
rect 18739 5049 18751 5083
rect 18984 5080 19012 5120
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 21082 5080 21088 5092
rect 18984 5052 21088 5080
rect 18693 5043 18751 5049
rect 21082 5040 21088 5052
rect 21140 5040 21146 5092
rect 11606 5012 11612 5024
rect 10060 4984 11612 5012
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 12986 5012 12992 5024
rect 12947 4984 12992 5012
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14240 4984 15025 5012
rect 14240 4972 14246 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 16574 5012 16580 5024
rect 16535 4984 16580 5012
rect 15013 4975 15071 4981
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 18840 4984 18885 5012
rect 18840 4972 18846 4984
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 20717 5015 20775 5021
rect 20717 5012 20729 5015
rect 19576 4984 20729 5012
rect 19576 4972 19582 4984
rect 20717 4981 20729 4984
rect 20763 4981 20775 5015
rect 20717 4975 20775 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 6641 4811 6699 4817
rect 6641 4777 6653 4811
rect 6687 4808 6699 4811
rect 7374 4808 7380 4820
rect 6687 4780 7380 4808
rect 6687 4777 6699 4780
rect 6641 4771 6699 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 8294 4808 8300 4820
rect 7699 4780 8300 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 11054 4768 11060 4820
rect 11112 4808 11118 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 11112 4780 11621 4808
rect 11112 4768 11118 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 12986 4768 12992 4820
rect 13044 4808 13050 4820
rect 13357 4811 13415 4817
rect 13357 4808 13369 4811
rect 13044 4780 13369 4808
rect 13044 4768 13050 4780
rect 13357 4777 13369 4780
rect 13403 4777 13415 4811
rect 19794 4808 19800 4820
rect 13357 4771 13415 4777
rect 16592 4780 19800 4808
rect 16592 4752 16620 4780
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 10965 4743 11023 4749
rect 10965 4740 10977 4743
rect 4764 4712 10977 4740
rect 4764 4700 4770 4712
rect 10965 4709 10977 4712
rect 11011 4709 11023 4743
rect 16574 4740 16580 4752
rect 10965 4703 11023 4709
rect 11072 4712 16580 4740
rect 4246 4632 4252 4684
rect 4304 4672 4310 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 4304 4644 7021 4672
rect 4304 4632 4310 4644
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7098 4632 7104 4684
rect 7156 4672 7162 4684
rect 8021 4675 8079 4681
rect 7156 4644 7328 4672
rect 7156 4632 7162 4644
rect 7190 4604 7196 4616
rect 7151 4576 7196 4604
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 7300 4536 7328 4644
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 8478 4672 8484 4684
rect 8067 4644 8484 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 11072 4672 11100 4712
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 19420 4743 19478 4749
rect 17328 4712 19196 4740
rect 17328 4684 17356 4712
rect 17310 4672 17316 4684
rect 8956 4644 11100 4672
rect 17271 4644 17316 4672
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 7432 4576 8125 4604
rect 7432 4564 7438 4576
rect 8113 4573 8125 4576
rect 8159 4573 8171 4607
rect 8113 4567 8171 4573
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8260 4576 8305 4604
rect 8260 4564 8266 4576
rect 8956 4536 8984 4644
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17580 4675 17638 4681
rect 17580 4641 17592 4675
rect 17626 4672 17638 4675
rect 17954 4672 17960 4684
rect 17626 4644 17960 4672
rect 17626 4641 17638 4644
rect 17580 4635 17638 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 19168 4681 19196 4712
rect 19420 4709 19432 4743
rect 19466 4740 19478 4743
rect 20162 4740 20168 4752
rect 19466 4712 20168 4740
rect 19466 4709 19478 4712
rect 19420 4703 19478 4709
rect 20162 4700 20168 4712
rect 20220 4700 20226 4752
rect 19153 4675 19211 4681
rect 19153 4641 19165 4675
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 10410 4564 10416 4616
rect 10468 4604 10474 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10468 4576 11069 4604
rect 10468 4564 10474 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11238 4604 11244 4616
rect 11151 4576 11244 4604
rect 11057 4567 11115 4573
rect 11238 4564 11244 4576
rect 11296 4604 11302 4616
rect 12158 4604 12164 4616
rect 11296 4576 12164 4604
rect 11296 4564 11302 4576
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 7300 4508 8984 4536
rect 10597 4539 10655 4545
rect 10597 4505 10609 4539
rect 10643 4536 10655 4539
rect 11146 4536 11152 4548
rect 10643 4508 11152 4536
rect 10643 4505 10655 4508
rect 10597 4499 10655 4505
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 17586 4428 17592 4480
rect 17644 4468 17650 4480
rect 18693 4471 18751 4477
rect 18693 4468 18705 4471
rect 17644 4440 18705 4468
rect 17644 4428 17650 4440
rect 18693 4437 18705 4440
rect 18739 4437 18751 4471
rect 20530 4468 20536 4480
rect 20491 4440 20536 4468
rect 18693 4431 18751 4437
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9125 4267 9183 4273
rect 9125 4264 9137 4267
rect 8996 4236 9137 4264
rect 8996 4224 9002 4236
rect 9125 4233 9137 4236
rect 9171 4233 9183 4267
rect 9125 4227 9183 4233
rect 9140 4196 9168 4227
rect 17034 4224 17040 4276
rect 17092 4264 17098 4276
rect 19058 4264 19064 4276
rect 17092 4236 19064 4264
rect 17092 4224 17098 4236
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 9140 4168 9996 4196
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 2682 4128 2688 4140
rect 1820 4100 2688 4128
rect 1820 4088 1826 4100
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 6880 4100 7757 4128
rect 6880 4088 6886 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 9858 4128 9864 4140
rect 9819 4100 9864 4128
rect 7745 4091 7803 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 9968 4137 9996 4168
rect 12820 4168 13124 4196
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 12820 4128 12848 4168
rect 12986 4128 12992 4140
rect 9953 4091 10011 4097
rect 10060 4100 12848 4128
rect 12947 4100 12992 4128
rect 10060 4060 10088 4100
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13096 4128 13124 4168
rect 13446 4156 13452 4208
rect 13504 4196 13510 4208
rect 13504 4168 14228 4196
rect 13504 4156 13510 4168
rect 13906 4128 13912 4140
rect 13096 4100 13912 4128
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 13998 4088 14004 4140
rect 14056 4128 14062 4140
rect 14093 4131 14151 4137
rect 14093 4128 14105 4131
rect 14056 4100 14105 4128
rect 14056 4088 14062 4100
rect 14093 4097 14105 4100
rect 14139 4097 14151 4131
rect 14200 4128 14228 4168
rect 15672 4168 16436 4196
rect 14200 4100 15148 4128
rect 14093 4091 14151 4097
rect 7852 4032 10088 4060
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 7852 3992 7880 4032
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 14182 4060 14188 4072
rect 10652 4032 14188 4060
rect 10652 4020 10658 4032
rect 14182 4020 14188 4032
rect 14240 4020 14246 4072
rect 15120 4060 15148 4100
rect 15378 4088 15384 4140
rect 15436 4128 15442 4140
rect 15672 4128 15700 4168
rect 15436 4100 15700 4128
rect 15436 4088 15442 4100
rect 15746 4088 15752 4140
rect 15804 4128 15810 4140
rect 16298 4128 16304 4140
rect 15804 4100 16304 4128
rect 15804 4088 15810 4100
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16408 4128 16436 4168
rect 19242 4156 19248 4208
rect 19300 4196 19306 4208
rect 19886 4196 19892 4208
rect 19300 4168 19892 4196
rect 19300 4156 19306 4168
rect 19886 4156 19892 4168
rect 19944 4156 19950 4208
rect 20272 4168 20668 4196
rect 17310 4128 17316 4140
rect 16408 4100 17316 4128
rect 17310 4088 17316 4100
rect 17368 4128 17374 4140
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17368 4100 18061 4128
rect 17368 4088 17374 4100
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18049 4091 18107 4097
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 20272 4128 20300 4168
rect 19208 4100 20300 4128
rect 20349 4131 20407 4137
rect 19208 4088 19214 4100
rect 20349 4097 20361 4131
rect 20395 4128 20407 4131
rect 20530 4128 20536 4140
rect 20395 4100 20536 4128
rect 20395 4097 20407 4100
rect 20349 4091 20407 4097
rect 17405 4063 17463 4069
rect 15120 4032 15884 4060
rect 5684 3964 7880 3992
rect 8012 3995 8070 4001
rect 5684 3952 5690 3964
rect 8012 3961 8024 3995
rect 8058 3992 8070 3995
rect 8202 3992 8208 4004
rect 8058 3964 8208 3992
rect 8058 3961 8070 3964
rect 8012 3955 8070 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 9769 3995 9827 4001
rect 9769 3992 9781 3995
rect 8312 3964 9781 3992
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 8312 3924 8340 3964
rect 9769 3961 9781 3964
rect 9815 3961 9827 3995
rect 9769 3955 9827 3961
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 13446 3992 13452 4004
rect 10008 3964 13452 3992
rect 10008 3952 10014 3964
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 15654 3992 15660 4004
rect 13688 3964 15660 3992
rect 13688 3952 13694 3964
rect 15654 3952 15660 3964
rect 15712 3952 15718 4004
rect 15856 3992 15884 4032
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17954 4060 17960 4072
rect 17451 4032 17960 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18316 4063 18374 4069
rect 18316 4029 18328 4063
rect 18362 4060 18374 4063
rect 19426 4060 19432 4072
rect 18362 4032 19432 4060
rect 18362 4029 18374 4032
rect 18316 4023 18374 4029
rect 19426 4020 19432 4032
rect 19484 4060 19490 4072
rect 20364 4060 20392 4091
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 20640 4128 20668 4168
rect 21358 4128 21364 4140
rect 20640 4100 21364 4128
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 19484 4032 20392 4060
rect 20717 4063 20775 4069
rect 19484 4020 19490 4032
rect 20717 4029 20729 4063
rect 20763 4060 20775 4063
rect 20806 4060 20812 4072
rect 20763 4032 20812 4060
rect 20763 4029 20775 4032
rect 20717 4023 20775 4029
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 18506 3992 18512 4004
rect 15856 3964 18512 3992
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 19058 3952 19064 4004
rect 19116 3992 19122 4004
rect 19116 3964 20944 3992
rect 19116 3952 19122 3964
rect 9398 3924 9404 3936
rect 6696 3896 8340 3924
rect 9359 3896 9404 3924
rect 6696 3884 6702 3896
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 10502 3924 10508 3936
rect 10463 3896 10508 3924
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 11606 3924 11612 3936
rect 11567 3896 11612 3924
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12526 3924 12532 3936
rect 12483 3896 12532 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 12768 3896 12817 3924
rect 12768 3884 12774 3896
rect 12805 3893 12817 3896
rect 12851 3893 12863 3927
rect 12805 3887 12863 3893
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 12943 3896 13553 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 13541 3887 13599 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 13909 3927 13967 3933
rect 13909 3924 13921 3927
rect 13872 3896 13921 3924
rect 13872 3884 13878 3896
rect 13909 3893 13921 3896
rect 13955 3893 13967 3927
rect 13909 3887 13967 3893
rect 14001 3927 14059 3933
rect 14001 3893 14013 3927
rect 14047 3924 14059 3927
rect 14366 3924 14372 3936
rect 14047 3896 14372 3924
rect 14047 3893 14059 3896
rect 14001 3887 14059 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 15102 3924 15108 3936
rect 15063 3896 15108 3924
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15470 3924 15476 3936
rect 15431 3896 15476 3924
rect 15470 3884 15476 3896
rect 15528 3884 15534 3936
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 15620 3896 15665 3924
rect 15620 3884 15626 3896
rect 15746 3884 15752 3936
rect 15804 3924 15810 3936
rect 17494 3924 17500 3936
rect 15804 3896 17500 3924
rect 15804 3884 15810 3896
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 17589 3927 17647 3933
rect 17589 3893 17601 3927
rect 17635 3924 17647 3927
rect 19150 3924 19156 3936
rect 17635 3896 19156 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 19242 3884 19248 3936
rect 19300 3924 19306 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 19300 3896 19441 3924
rect 19300 3884 19306 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 19702 3924 19708 3936
rect 19663 3896 19708 3924
rect 19429 3887 19487 3893
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 20073 3927 20131 3933
rect 20073 3924 20085 3927
rect 19944 3896 20085 3924
rect 19944 3884 19950 3896
rect 20073 3893 20085 3896
rect 20119 3893 20131 3927
rect 20073 3887 20131 3893
rect 20165 3927 20223 3933
rect 20165 3893 20177 3927
rect 20211 3924 20223 3927
rect 20346 3924 20352 3936
rect 20211 3896 20352 3924
rect 20211 3893 20223 3896
rect 20165 3887 20223 3893
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 20916 3933 20944 3964
rect 20901 3927 20959 3933
rect 20901 3893 20913 3927
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 4706 3720 4712 3732
rect 3476 3692 4712 3720
rect 3476 3680 3482 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8260 3692 8493 3720
rect 8260 3680 8266 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 9732 3692 11253 3720
rect 9732 3680 9738 3692
rect 11241 3689 11253 3692
rect 11287 3720 11299 3723
rect 11790 3720 11796 3732
rect 11287 3692 11796 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12713 3723 12771 3729
rect 12713 3689 12725 3723
rect 12759 3720 12771 3723
rect 12802 3720 12808 3732
rect 12759 3692 12808 3720
rect 12759 3689 12771 3692
rect 12713 3683 12771 3689
rect 12802 3680 12808 3692
rect 12860 3720 12866 3732
rect 12986 3720 12992 3732
rect 12860 3692 12992 3720
rect 12860 3680 12866 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 16942 3720 16948 3732
rect 14743 3692 16948 3720
rect 2314 3612 2320 3664
rect 2372 3652 2378 3664
rect 8846 3652 8852 3664
rect 2372 3624 8852 3652
rect 2372 3612 2378 3624
rect 8846 3612 8852 3624
rect 8904 3612 8910 3664
rect 8938 3612 8944 3664
rect 8996 3652 9002 3664
rect 11698 3652 11704 3664
rect 8996 3624 11704 3652
rect 8996 3612 9002 3624
rect 11698 3612 11704 3624
rect 11756 3612 11762 3664
rect 14642 3612 14648 3664
rect 14700 3652 14706 3664
rect 14743 3652 14771 3692
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17678 3720 17684 3732
rect 17639 3692 17684 3720
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3720 18107 3723
rect 18322 3720 18328 3732
rect 18095 3692 18328 3720
rect 18095 3689 18107 3692
rect 18049 3683 18107 3689
rect 18322 3680 18328 3692
rect 18380 3680 18386 3732
rect 18414 3680 18420 3732
rect 18472 3720 18478 3732
rect 18693 3723 18751 3729
rect 18472 3692 18644 3720
rect 18472 3680 18478 3692
rect 14700 3624 14771 3652
rect 15648 3655 15706 3661
rect 14700 3612 14706 3624
rect 15648 3621 15660 3655
rect 15694 3652 15706 3655
rect 17586 3652 17592 3664
rect 15694 3624 17592 3652
rect 15694 3621 15706 3624
rect 15648 3615 15706 3621
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 18506 3652 18512 3664
rect 17696 3624 18512 3652
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 4246 3584 4252 3596
rect 2924 3556 4252 3584
rect 2924 3544 2930 3556
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6880 3556 7113 3584
rect 6880 3544 6886 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 7368 3587 7426 3593
rect 7368 3553 7380 3587
rect 7414 3584 7426 3587
rect 8202 3584 8208 3596
rect 7414 3556 8208 3584
rect 7414 3553 7426 3556
rect 7368 3547 7426 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 9944 3587 10002 3593
rect 9944 3553 9956 3587
rect 9990 3584 10002 3587
rect 10686 3584 10692 3596
rect 9990 3556 10692 3584
rect 9990 3553 10002 3556
rect 9944 3547 10002 3553
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 11241 3587 11299 3593
rect 11241 3553 11253 3587
rect 11287 3584 11299 3587
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 11287 3556 11345 3584
rect 11287 3553 11299 3556
rect 11241 3547 11299 3553
rect 11333 3553 11345 3556
rect 11379 3553 11391 3587
rect 11333 3547 11391 3553
rect 11600 3587 11658 3593
rect 11600 3553 11612 3587
rect 11646 3584 11658 3587
rect 11882 3584 11888 3596
rect 11646 3556 11888 3584
rect 11646 3553 11658 3556
rect 11600 3547 11658 3553
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 13348 3587 13406 3593
rect 13348 3553 13360 3587
rect 13394 3584 13406 3587
rect 14366 3584 14372 3596
rect 13394 3556 14372 3584
rect 13394 3553 13406 3556
rect 13348 3547 13406 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 15068 3556 16436 3584
rect 15068 3544 15074 3556
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 13044 3488 13093 3516
rect 13044 3476 13050 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14737 3519 14795 3525
rect 14737 3516 14749 3519
rect 14148 3488 14749 3516
rect 14148 3476 14154 3488
rect 14737 3485 14749 3488
rect 14783 3485 14795 3519
rect 15378 3516 15384 3528
rect 15339 3488 15384 3516
rect 14737 3479 14795 3485
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 16408 3516 16436 3556
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 17092 3556 17141 3584
rect 17092 3544 17098 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 17696 3516 17724 3624
rect 18506 3612 18512 3624
rect 18564 3612 18570 3664
rect 18616 3652 18644 3692
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 18782 3720 18788 3732
rect 18739 3692 18788 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 19061 3723 19119 3729
rect 19061 3689 19073 3723
rect 19107 3689 19119 3723
rect 19705 3723 19763 3729
rect 19705 3720 19717 3723
rect 19061 3683 19119 3689
rect 19628 3692 19717 3720
rect 19076 3652 19104 3683
rect 18616 3624 19104 3652
rect 19153 3655 19211 3661
rect 19153 3621 19165 3655
rect 19199 3652 19211 3655
rect 19199 3624 19463 3652
rect 19199 3621 19211 3624
rect 19153 3615 19211 3621
rect 18046 3544 18052 3596
rect 18104 3584 18110 3596
rect 19435 3584 19463 3624
rect 19628 3584 19656 3692
rect 19705 3689 19717 3692
rect 19751 3689 19763 3723
rect 19705 3683 19763 3689
rect 19794 3680 19800 3732
rect 19852 3720 19858 3732
rect 20073 3723 20131 3729
rect 20073 3720 20085 3723
rect 19852 3692 20085 3720
rect 19852 3680 19858 3692
rect 20073 3689 20085 3692
rect 20119 3720 20131 3723
rect 20162 3720 20168 3732
rect 20119 3692 20168 3720
rect 20119 3689 20131 3692
rect 20073 3683 20131 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 21910 3720 21916 3732
rect 20680 3692 21916 3720
rect 20680 3680 20686 3692
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 20901 3655 20959 3661
rect 20901 3652 20913 3655
rect 20772 3624 20913 3652
rect 20772 3612 20778 3624
rect 20901 3621 20913 3624
rect 20947 3621 20959 3655
rect 20901 3615 20959 3621
rect 18104 3556 18276 3584
rect 19435 3556 19656 3584
rect 20165 3587 20223 3593
rect 18104 3544 18110 3556
rect 16408 3488 17724 3516
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18248 3525 18276 3556
rect 20165 3553 20177 3587
rect 20211 3584 20223 3587
rect 21082 3584 21088 3596
rect 20211 3556 21088 3584
rect 20211 3553 20223 3556
rect 20165 3547 20223 3553
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 18012 3488 18153 3516
rect 18012 3476 18018 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 20349 3519 20407 3525
rect 20349 3485 20361 3519
rect 20395 3516 20407 3519
rect 20530 3516 20536 3528
rect 20395 3488 20536 3516
rect 20395 3485 20407 3488
rect 20349 3479 20407 3485
rect 14458 3448 14464 3460
rect 14419 3420 14464 3448
rect 14458 3408 14464 3420
rect 14516 3408 14522 3460
rect 17494 3448 17500 3460
rect 16316 3420 17500 3448
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 10778 3380 10784 3392
rect 6972 3352 10784 3380
rect 6972 3340 6978 3352
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 11054 3380 11060 3392
rect 11015 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 12342 3340 12348 3392
rect 12400 3380 12406 3392
rect 16316 3380 16344 3420
rect 17494 3408 17500 3420
rect 17552 3408 17558 3460
rect 18248 3448 18276 3479
rect 19150 3448 19156 3460
rect 18248 3420 19156 3448
rect 19150 3408 19156 3420
rect 19208 3448 19214 3460
rect 19260 3448 19288 3479
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 19208 3420 19288 3448
rect 19208 3408 19214 3420
rect 19702 3408 19708 3460
rect 19760 3448 19766 3460
rect 20898 3448 20904 3460
rect 19760 3420 20904 3448
rect 19760 3408 19766 3420
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 12400 3352 16344 3380
rect 12400 3340 12406 3352
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 16761 3383 16819 3389
rect 16761 3380 16773 3383
rect 16540 3352 16773 3380
rect 16540 3340 16546 3352
rect 16761 3349 16773 3352
rect 16807 3349 16819 3383
rect 16761 3343 16819 3349
rect 17313 3383 17371 3389
rect 17313 3349 17325 3383
rect 17359 3380 17371 3383
rect 20806 3380 20812 3392
rect 17359 3352 20812 3380
rect 17359 3349 17371 3352
rect 17313 3343 17371 3349
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 3970 3136 3976 3188
rect 4028 3176 4034 3188
rect 8202 3176 8208 3188
rect 4028 3148 7788 3176
rect 8163 3148 8208 3176
rect 4028 3136 4034 3148
rect 7760 3108 7788 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 10686 3176 10692 3188
rect 9548 3148 10272 3176
rect 10647 3148 10692 3176
rect 9548 3136 9554 3148
rect 8938 3108 8944 3120
rect 7760 3080 8944 3108
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 10244 3108 10272 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10870 3136 10876 3188
rect 10928 3176 10934 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10928 3148 10977 3176
rect 10928 3136 10934 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 14366 3176 14372 3188
rect 11204 3148 14228 3176
rect 14327 3148 14372 3176
rect 11204 3136 11210 3148
rect 12250 3108 12256 3120
rect 10244 3080 12256 3108
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 12986 3108 12992 3120
rect 12360 3080 12992 3108
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 8478 3040 8484 3052
rect 8439 3012 8484 3040
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 11054 3040 11060 3052
rect 10428 3012 11060 3040
rect 9309 2975 9367 2981
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 9398 2972 9404 2984
rect 9355 2944 9404 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10428 2972 10456 3012
rect 11054 3000 11060 3012
rect 11112 3040 11118 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11112 3012 11529 3040
rect 11112 3000 11118 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 12360 3040 12388 3080
rect 12986 3068 12992 3080
rect 13044 3068 13050 3120
rect 14200 3108 14228 3148
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 15378 3176 15384 3188
rect 15212 3148 15384 3176
rect 14200 3080 15148 3108
rect 11848 3012 12388 3040
rect 11848 3000 11854 3012
rect 9508 2944 10456 2972
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 6914 2904 6920 2916
rect 716 2876 6920 2904
rect 716 2864 722 2876
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 7092 2907 7150 2913
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 9508 2904 9536 2944
rect 10502 2932 10508 2984
rect 10560 2972 10566 2984
rect 11333 2975 11391 2981
rect 11333 2972 11345 2975
rect 10560 2944 11345 2972
rect 10560 2932 10566 2944
rect 11333 2941 11345 2944
rect 11379 2941 11391 2975
rect 11333 2935 11391 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12894 2972 12900 2984
rect 12483 2944 12900 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13256 2975 13314 2981
rect 13044 2944 13089 2972
rect 13044 2932 13050 2944
rect 13256 2941 13268 2975
rect 13302 2972 13314 2975
rect 13630 2972 13636 2984
rect 13302 2944 13636 2972
rect 13302 2941 13314 2944
rect 13256 2935 13314 2941
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 7138 2876 9536 2904
rect 9576 2907 9634 2913
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 9576 2873 9588 2907
rect 9622 2904 9634 2907
rect 12802 2904 12808 2916
rect 9622 2876 12808 2904
rect 9622 2873 9634 2876
rect 9576 2867 9634 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 13722 2864 13728 2916
rect 13780 2904 13786 2916
rect 15120 2904 15148 3080
rect 15212 3049 15240 3148
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15470 3136 15476 3188
rect 15528 3176 15534 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 15528 3148 16865 3176
rect 15528 3136 15534 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 17126 3136 17132 3188
rect 17184 3176 17190 3188
rect 17586 3176 17592 3188
rect 17184 3148 17592 3176
rect 17184 3136 17190 3148
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 18012 3148 18061 3176
rect 18012 3136 18018 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 18049 3139 18107 3145
rect 18156 3148 20637 3176
rect 16206 3068 16212 3120
rect 16264 3108 16270 3120
rect 18156 3108 18184 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 20625 3139 20683 3145
rect 16264 3080 18184 3108
rect 19521 3111 19579 3117
rect 16264 3068 16270 3080
rect 19521 3077 19533 3111
rect 19567 3108 19579 3111
rect 20254 3108 20260 3120
rect 19567 3080 20260 3108
rect 19567 3077 19579 3080
rect 19521 3071 19579 3077
rect 20254 3068 20260 3080
rect 20312 3068 20318 3120
rect 15197 3043 15255 3049
rect 15197 3009 15209 3043
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 17184 3012 17325 3040
rect 17184 3000 17190 3012
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 17313 3003 17371 3009
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 18506 3040 18512 3052
rect 18467 3012 18512 3040
rect 17405 3003 17463 3009
rect 15464 2975 15522 2981
rect 15464 2941 15476 2975
rect 15510 2972 15522 2975
rect 16482 2972 16488 2984
rect 15510 2944 16488 2972
rect 15510 2941 15522 2944
rect 15464 2935 15522 2941
rect 16482 2932 16488 2944
rect 16540 2972 16546 2984
rect 17420 2972 17448 3003
rect 18506 3000 18512 3012
rect 18564 3000 18570 3052
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 19426 3040 19432 3052
rect 18739 3012 19432 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 16540 2944 17448 2972
rect 16540 2932 16546 2944
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17552 2944 18429 2972
rect 17552 2932 17558 2944
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 19334 2972 19340 2984
rect 19295 2944 19340 2972
rect 18417 2935 18475 2941
rect 19334 2932 19340 2944
rect 19392 2932 19398 2984
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2972 19947 2975
rect 19978 2972 19984 2984
rect 19935 2944 19984 2972
rect 19935 2941 19947 2944
rect 19889 2935 19947 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20070 2932 20076 2984
rect 20128 2972 20134 2984
rect 20441 2975 20499 2981
rect 20441 2972 20453 2975
rect 20128 2944 20453 2972
rect 20128 2932 20134 2944
rect 20441 2941 20453 2944
rect 20487 2941 20499 2975
rect 20441 2935 20499 2941
rect 15746 2904 15752 2916
rect 13780 2876 14872 2904
rect 15120 2876 15752 2904
rect 13780 2864 13786 2876
rect 6086 2796 6092 2848
rect 6144 2836 6150 2848
rect 8570 2836 8576 2848
rect 6144 2808 8576 2836
rect 6144 2796 6150 2808
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 10502 2836 10508 2848
rect 8904 2808 10508 2836
rect 8904 2796 8910 2808
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 12618 2836 12624 2848
rect 12579 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 14844 2845 14872 2876
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 15838 2864 15844 2916
rect 15896 2904 15902 2916
rect 15896 2876 20116 2904
rect 15896 2864 15902 2876
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 15010 2796 15016 2848
rect 15068 2836 15074 2848
rect 16206 2836 16212 2848
rect 15068 2808 16212 2836
rect 15068 2796 15074 2808
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 16298 2796 16304 2848
rect 16356 2836 16362 2848
rect 16577 2839 16635 2845
rect 16577 2836 16589 2839
rect 16356 2808 16589 2836
rect 16356 2796 16362 2808
rect 16577 2805 16589 2808
rect 16623 2805 16635 2839
rect 17218 2836 17224 2848
rect 17131 2808 17224 2836
rect 16577 2799 16635 2805
rect 17218 2796 17224 2808
rect 17276 2836 17282 2848
rect 17954 2836 17960 2848
rect 17276 2808 17960 2836
rect 17276 2796 17282 2808
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 19426 2836 19432 2848
rect 18656 2808 19432 2836
rect 18656 2796 18662 2808
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 20088 2845 20116 2876
rect 20073 2839 20131 2845
rect 20073 2805 20085 2839
rect 20119 2805 20131 2839
rect 20073 2799 20131 2805
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 10045 2635 10103 2641
rect 10045 2601 10057 2635
rect 10091 2632 10103 2635
rect 11422 2632 11428 2644
rect 10091 2604 11428 2632
rect 10091 2601 10103 2604
rect 10045 2595 10103 2601
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 11606 2592 11612 2644
rect 11664 2632 11670 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11664 2604 11713 2632
rect 11664 2592 11670 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 13633 2635 13691 2641
rect 13633 2601 13645 2635
rect 13679 2632 13691 2635
rect 14090 2632 14096 2644
rect 13679 2604 14096 2632
rect 13679 2601 13691 2604
rect 13633 2595 13691 2601
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 14274 2632 14280 2644
rect 14235 2604 14280 2632
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 14737 2635 14795 2641
rect 14737 2601 14749 2635
rect 14783 2632 14795 2635
rect 15102 2632 15108 2644
rect 14783 2604 15108 2632
rect 14783 2601 14795 2604
rect 14737 2595 14795 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 15562 2592 15568 2644
rect 15620 2632 15626 2644
rect 15657 2635 15715 2641
rect 15657 2632 15669 2635
rect 15620 2604 15669 2632
rect 15620 2592 15626 2604
rect 15657 2601 15669 2604
rect 15703 2601 15715 2635
rect 16022 2632 16028 2644
rect 15935 2604 16028 2632
rect 15657 2595 15715 2601
rect 16022 2592 16028 2604
rect 16080 2632 16086 2644
rect 19610 2632 19616 2644
rect 16080 2604 19616 2632
rect 16080 2592 16086 2604
rect 19610 2592 19616 2604
rect 19668 2632 19674 2644
rect 19978 2632 19984 2644
rect 19668 2604 19984 2632
rect 19668 2592 19674 2604
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20073 2635 20131 2641
rect 20073 2601 20085 2635
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 7834 2524 7840 2576
rect 7892 2564 7898 2576
rect 10413 2567 10471 2573
rect 10413 2564 10425 2567
rect 7892 2536 10425 2564
rect 7892 2524 7898 2536
rect 10413 2533 10425 2536
rect 10459 2533 10471 2567
rect 10413 2527 10471 2533
rect 10502 2524 10508 2576
rect 10560 2564 10566 2576
rect 13725 2567 13783 2573
rect 13725 2564 13737 2567
rect 10560 2536 13737 2564
rect 10560 2524 10566 2536
rect 13725 2533 13737 2536
rect 13771 2533 13783 2567
rect 13725 2527 13783 2533
rect 15378 2524 15384 2576
rect 15436 2564 15442 2576
rect 20088 2564 20116 2595
rect 15436 2536 20116 2564
rect 15436 2524 15442 2536
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 7248 2468 7757 2496
rect 7248 2456 7254 2468
rect 7745 2465 7757 2468
rect 7791 2465 7803 2499
rect 7745 2459 7803 2465
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 8352 2468 11805 2496
rect 8352 2456 8358 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13354 2496 13360 2508
rect 12667 2468 13360 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 13924 2468 14657 2496
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7156 2400 7849 2428
rect 7156 2388 7162 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8202 2428 8208 2440
rect 8067 2400 8208 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 10468 2400 10517 2428
rect 10468 2388 10474 2400
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 10686 2428 10692 2440
rect 10647 2400 10692 2428
rect 10505 2391 10563 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 11882 2428 11888 2440
rect 11843 2400 11888 2428
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 13630 2388 13636 2440
rect 13688 2428 13694 2440
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 13688 2400 13829 2428
rect 13688 2388 13694 2400
rect 13817 2397 13829 2400
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 11333 2363 11391 2369
rect 11333 2329 11345 2363
rect 11379 2360 11391 2363
rect 12710 2360 12716 2372
rect 11379 2332 12716 2360
rect 11379 2329 11391 2332
rect 11333 2323 11391 2329
rect 12710 2320 12716 2332
rect 12768 2320 12774 2372
rect 13265 2363 13323 2369
rect 13265 2329 13277 2363
rect 13311 2360 13323 2363
rect 13924 2360 13952 2468
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17402 2496 17408 2508
rect 16991 2468 17408 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17402 2456 17408 2468
rect 17460 2456 17466 2508
rect 17497 2499 17555 2505
rect 17497 2465 17509 2499
rect 17543 2496 17555 2499
rect 17770 2496 17776 2508
rect 17543 2468 17776 2496
rect 17543 2465 17555 2468
rect 17497 2459 17555 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18690 2496 18696 2508
rect 18371 2468 18696 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 18874 2496 18880 2508
rect 18835 2468 18880 2496
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19794 2456 19800 2508
rect 19852 2496 19858 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19852 2468 19901 2496
rect 19852 2456 19858 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 20438 2496 20444 2508
rect 20399 2468 20444 2496
rect 19889 2459 19947 2465
rect 20438 2456 20444 2468
rect 20496 2456 20502 2508
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14424 2400 14841 2428
rect 14424 2388 14430 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 14829 2391 14887 2397
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16482 2428 16488 2440
rect 16347 2400 16488 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 16592 2400 20668 2428
rect 13311 2332 13952 2360
rect 13311 2329 13323 2332
rect 13265 2323 13323 2329
rect 14274 2320 14280 2372
rect 14332 2360 14338 2372
rect 16592 2360 16620 2400
rect 14332 2332 16620 2360
rect 14332 2320 14338 2332
rect 17034 2320 17040 2372
rect 17092 2360 17098 2372
rect 17681 2363 17739 2369
rect 17681 2360 17693 2363
rect 17092 2332 17693 2360
rect 17092 2320 17098 2332
rect 17681 2329 17693 2332
rect 17727 2329 17739 2363
rect 17681 2323 17739 2329
rect 17954 2320 17960 2372
rect 18012 2360 18018 2372
rect 20640 2369 20668 2400
rect 19061 2363 19119 2369
rect 19061 2360 19073 2363
rect 18012 2332 19073 2360
rect 18012 2320 18018 2332
rect 19061 2329 19073 2332
rect 19107 2329 19119 2363
rect 19061 2323 19119 2329
rect 20625 2363 20683 2369
rect 20625 2329 20637 2363
rect 20671 2329 20683 2363
rect 20625 2323 20683 2329
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 11664 2264 12817 2292
rect 11664 2252 11670 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 16482 2252 16488 2304
rect 16540 2292 16546 2304
rect 17129 2295 17187 2301
rect 17129 2292 17141 2295
rect 16540 2264 17141 2292
rect 16540 2252 16546 2264
rect 17129 2261 17141 2264
rect 17175 2261 17187 2295
rect 17129 2255 17187 2261
rect 17494 2252 17500 2304
rect 17552 2292 17558 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 17552 2264 18521 2292
rect 17552 2252 17558 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 10410 2048 10416 2100
rect 10468 2088 10474 2100
rect 16114 2088 16120 2100
rect 10468 2060 16120 2088
rect 10468 2048 10474 2060
rect 16114 2048 16120 2060
rect 16172 2088 16178 2100
rect 18782 2088 18788 2100
rect 16172 2060 18788 2088
rect 16172 2048 16178 2060
rect 18782 2048 18788 2060
rect 18840 2088 18846 2100
rect 20070 2088 20076 2100
rect 18840 2060 20076 2088
rect 18840 2048 18846 2060
rect 20070 2048 20076 2060
rect 20128 2048 20134 2100
rect 9858 1980 9864 2032
rect 9916 2020 9922 2032
rect 16022 2020 16028 2032
rect 9916 1992 16028 2020
rect 9916 1980 9922 1992
rect 16022 1980 16028 1992
rect 16080 1980 16086 2032
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20628 20000 20680 20052
rect 19984 19907 20036 19916
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 20076 19864 20128 19916
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 20720 19499 20772 19508
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 5724 19252 5776 19304
rect 12716 19252 12768 19304
rect 16120 19252 16172 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 17960 19116 18012 19168
rect 19248 19116 19300 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 20444 18955 20496 18964
rect 20444 18921 20453 18955
rect 20453 18921 20487 18955
rect 20487 18921 20496 18955
rect 20444 18912 20496 18921
rect 20260 18819 20312 18828
rect 20260 18785 20269 18819
rect 20269 18785 20303 18819
rect 20303 18785 20312 18819
rect 20260 18776 20312 18785
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 20536 18300 20588 18352
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 19984 18232 20036 18284
rect 9772 18164 9824 18216
rect 13636 18164 13688 18216
rect 15292 18164 15344 18216
rect 17960 18164 18012 18216
rect 20076 18164 20128 18216
rect 19984 18096 20036 18148
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 17868 17824 17920 17876
rect 7656 17688 7708 17740
rect 11612 17688 11664 17740
rect 14096 17688 14148 17740
rect 20260 17620 20312 17672
rect 18512 17552 18564 17604
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 11612 17187 11664 17196
rect 11612 17153 11621 17187
rect 11621 17153 11655 17187
rect 11655 17153 11664 17187
rect 11612 17144 11664 17153
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 11796 17076 11848 17128
rect 13820 17119 13872 17128
rect 13820 17085 13829 17119
rect 13829 17085 13863 17119
rect 13863 17085 13872 17119
rect 13820 17076 13872 17085
rect 19800 17076 19852 17128
rect 20076 17076 20128 17128
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 18512 16668 18564 16720
rect 19800 16711 19852 16720
rect 19524 16643 19576 16652
rect 19524 16609 19533 16643
rect 19533 16609 19567 16643
rect 19567 16609 19576 16643
rect 19524 16600 19576 16609
rect 19800 16677 19809 16711
rect 19809 16677 19843 16711
rect 19843 16677 19852 16711
rect 19800 16668 19852 16677
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 20076 16056 20128 16108
rect 16948 15988 17000 16040
rect 16672 15920 16724 15972
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 18512 15580 18564 15632
rect 14004 15555 14056 15564
rect 14004 15521 14013 15555
rect 14013 15521 14047 15555
rect 14047 15521 14056 15555
rect 14004 15512 14056 15521
rect 19340 15512 19392 15564
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 20168 15147 20220 15156
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 16672 14968 16724 15020
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 19984 14943 20036 14952
rect 12440 14900 12492 14909
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 20536 14943 20588 14952
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 20720 14807 20772 14816
rect 20720 14773 20729 14807
rect 20729 14773 20763 14807
rect 20763 14773 20772 14807
rect 20720 14764 20772 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 19892 14603 19944 14612
rect 19892 14569 19901 14603
rect 19901 14569 19935 14603
rect 19935 14569 19944 14603
rect 19892 14560 19944 14569
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 9680 14467 9732 14476
rect 9680 14433 9689 14467
rect 9689 14433 9723 14467
rect 9723 14433 9732 14467
rect 9680 14424 9732 14433
rect 19340 14424 19392 14476
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 20260 14467 20312 14476
rect 20260 14433 20269 14467
rect 20269 14433 20303 14467
rect 20303 14433 20312 14467
rect 20260 14424 20312 14433
rect 19984 14356 20036 14408
rect 20444 14331 20496 14340
rect 20444 14297 20453 14331
rect 20453 14297 20487 14331
rect 20487 14297 20496 14331
rect 20444 14288 20496 14297
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 10876 13812 10928 13864
rect 19708 13812 19760 13864
rect 20352 13812 20404 13864
rect 18880 13744 18932 13796
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 12532 13472 12584 13524
rect 19248 13515 19300 13524
rect 19248 13481 19257 13515
rect 19257 13481 19291 13515
rect 19291 13481 19300 13515
rect 19248 13472 19300 13481
rect 17132 13336 17184 13388
rect 19432 13336 19484 13388
rect 20536 13404 20588 13456
rect 15936 13268 15988 13320
rect 16764 13132 16816 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 17960 12928 18012 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 19432 12835 19484 12844
rect 19432 12801 19441 12835
rect 19441 12801 19475 12835
rect 19475 12801 19484 12835
rect 19432 12792 19484 12801
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 19064 12724 19116 12776
rect 14280 12656 14332 12708
rect 20904 12724 20956 12776
rect 17960 12588 18012 12640
rect 18512 12631 18564 12640
rect 18512 12597 18521 12631
rect 18521 12597 18555 12631
rect 18555 12597 18564 12631
rect 18512 12588 18564 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 18604 12316 18656 12368
rect 17500 12248 17552 12300
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 15660 12180 15712 12232
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 15936 12044 15988 12096
rect 20536 12180 20588 12232
rect 18604 12044 18656 12096
rect 18972 12087 19024 12096
rect 18972 12053 18981 12087
rect 18981 12053 19015 12087
rect 19015 12053 19024 12087
rect 18972 12044 19024 12053
rect 20628 12044 20680 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 20076 11840 20128 11892
rect 20720 11883 20772 11892
rect 20720 11849 20729 11883
rect 20729 11849 20763 11883
rect 20763 11849 20772 11883
rect 20720 11840 20772 11849
rect 13912 11704 13964 11756
rect 17960 11704 18012 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 13452 11636 13504 11688
rect 15936 11636 15988 11688
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 20536 11679 20588 11688
rect 20536 11645 20545 11679
rect 20545 11645 20579 11679
rect 20579 11645 20588 11679
rect 20536 11636 20588 11645
rect 13360 11568 13412 11620
rect 15384 11568 15436 11620
rect 18972 11568 19024 11620
rect 19432 11568 19484 11620
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 19340 11500 19392 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 13544 11296 13596 11348
rect 15292 11339 15344 11348
rect 4068 11228 4120 11280
rect 13912 11228 13964 11280
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 18512 11296 18564 11348
rect 19892 11339 19944 11348
rect 19892 11305 19901 11339
rect 19901 11305 19935 11339
rect 19935 11305 19944 11339
rect 19892 11296 19944 11305
rect 13176 11092 13228 11144
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 13084 11024 13136 11076
rect 15384 11024 15436 11076
rect 17592 11160 17644 11212
rect 19156 11160 19208 11212
rect 20168 11160 20220 11212
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 17040 11135 17092 11144
rect 15844 11092 15896 11101
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 17500 11092 17552 11144
rect 19340 11092 19392 11144
rect 19432 11092 19484 11144
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 13912 10795 13964 10804
rect 13912 10761 13921 10795
rect 13921 10761 13955 10795
rect 13955 10761 13964 10795
rect 13912 10752 13964 10761
rect 15752 10752 15804 10804
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 16580 10752 16632 10804
rect 15384 10659 15436 10668
rect 15384 10625 15393 10659
rect 15393 10625 15427 10659
rect 15427 10625 15436 10659
rect 15384 10616 15436 10625
rect 19340 10684 19392 10736
rect 11704 10548 11756 10600
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 18512 10548 18564 10600
rect 19432 10548 19484 10600
rect 13268 10480 13320 10532
rect 20168 10480 20220 10532
rect 14556 10412 14608 10464
rect 16028 10412 16080 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 18604 10412 18656 10464
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 20352 10412 20404 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 16948 10208 17000 10260
rect 20352 10140 20404 10192
rect 16948 10072 17000 10124
rect 19340 10072 19392 10124
rect 20260 10115 20312 10124
rect 20260 10081 20269 10115
rect 20269 10081 20303 10115
rect 20303 10081 20312 10115
rect 20260 10072 20312 10081
rect 15568 10004 15620 10056
rect 16488 10004 16540 10056
rect 16580 10004 16632 10056
rect 17868 10004 17920 10056
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 18512 9868 18564 9920
rect 18696 9868 18748 9920
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 12072 9664 12124 9716
rect 18696 9664 18748 9716
rect 19340 9664 19392 9716
rect 16948 9528 17000 9580
rect 19248 9528 19300 9580
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 12992 9503 13044 9512
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 13084 9460 13136 9512
rect 15384 9503 15436 9512
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 16580 9460 16632 9512
rect 17868 9460 17920 9512
rect 18696 9460 18748 9512
rect 20812 9503 20864 9512
rect 20812 9469 20821 9503
rect 20821 9469 20855 9503
rect 20855 9469 20864 9503
rect 20812 9460 20864 9469
rect 12900 9392 12952 9444
rect 14372 9392 14424 9444
rect 10784 9324 10836 9376
rect 14556 9324 14608 9376
rect 16120 9392 16172 9444
rect 18144 9392 18196 9444
rect 18512 9392 18564 9444
rect 16488 9324 16540 9376
rect 17868 9324 17920 9376
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 20352 9324 20404 9376
rect 20996 9367 21048 9376
rect 20996 9333 21005 9367
rect 21005 9333 21039 9367
rect 21039 9333 21048 9367
rect 20996 9324 21048 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 12992 9120 13044 9172
rect 17500 9120 17552 9172
rect 17868 9163 17920 9172
rect 17868 9129 17877 9163
rect 17877 9129 17911 9163
rect 17911 9129 17920 9163
rect 17868 9120 17920 9129
rect 19156 9120 19208 9172
rect 11060 9052 11112 9104
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 11704 9052 11756 9104
rect 16488 9052 16540 9104
rect 18696 9052 18748 9104
rect 11612 9027 11664 9036
rect 11612 8993 11646 9027
rect 11646 8993 11664 9027
rect 11612 8984 11664 8993
rect 14096 8984 14148 9036
rect 15384 8984 15436 9036
rect 20536 8984 20588 9036
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 15108 8916 15160 8968
rect 18144 8916 18196 8968
rect 18512 8916 18564 8968
rect 5080 8780 5132 8832
rect 13912 8780 13964 8832
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 14464 8780 14516 8832
rect 18880 8848 18932 8900
rect 16948 8823 17000 8832
rect 16948 8789 16957 8823
rect 16957 8789 16991 8823
rect 16991 8789 17000 8823
rect 16948 8780 17000 8789
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 9680 8576 9732 8628
rect 4896 8508 4948 8560
rect 11612 8551 11664 8560
rect 11612 8517 11621 8551
rect 11621 8517 11655 8551
rect 11655 8517 11664 8551
rect 11612 8508 11664 8517
rect 12992 8508 13044 8560
rect 14004 8576 14056 8628
rect 15568 8619 15620 8628
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 9312 8440 9364 8492
rect 14372 8440 14424 8492
rect 11060 8372 11112 8424
rect 14464 8372 14516 8424
rect 15108 8415 15160 8424
rect 15108 8381 15117 8415
rect 15117 8381 15151 8415
rect 15151 8381 15160 8415
rect 15108 8372 15160 8381
rect 17132 8508 17184 8560
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 18696 8372 18748 8424
rect 19892 8372 19944 8424
rect 9404 8304 9456 8356
rect 10968 8304 11020 8356
rect 12808 8304 12860 8356
rect 13912 8304 13964 8356
rect 16028 8347 16080 8356
rect 9220 8279 9272 8288
rect 9220 8245 9229 8279
rect 9229 8245 9263 8279
rect 9263 8245 9272 8279
rect 9220 8236 9272 8245
rect 14188 8279 14240 8288
rect 14188 8245 14197 8279
rect 14197 8245 14231 8279
rect 14231 8245 14240 8279
rect 14188 8236 14240 8245
rect 15016 8236 15068 8288
rect 16028 8313 16037 8347
rect 16037 8313 16071 8347
rect 16071 8313 16080 8347
rect 16028 8304 16080 8313
rect 16488 8304 16540 8356
rect 17040 8304 17092 8356
rect 17224 8279 17276 8288
rect 17224 8245 17233 8279
rect 17233 8245 17267 8279
rect 17267 8245 17276 8279
rect 17224 8236 17276 8245
rect 18144 8279 18196 8288
rect 18144 8245 18153 8279
rect 18153 8245 18187 8279
rect 18187 8245 18196 8279
rect 18144 8236 18196 8245
rect 18604 8236 18656 8288
rect 18788 8236 18840 8288
rect 19616 8236 19668 8288
rect 19708 8236 19760 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 10968 8032 11020 8084
rect 15016 8032 15068 8084
rect 16304 8032 16356 8084
rect 8944 7896 8996 7948
rect 14004 7964 14056 8016
rect 16948 7964 17000 8016
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 11060 7896 11112 7948
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 11888 7896 11940 7905
rect 12716 7896 12768 7948
rect 14188 7896 14240 7948
rect 16028 7896 16080 7948
rect 18144 7896 18196 7948
rect 18788 7896 18840 7948
rect 20352 7896 20404 7948
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 16948 7828 17000 7880
rect 18880 7828 18932 7880
rect 19156 7828 19208 7880
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 20260 7828 20312 7837
rect 20536 7828 20588 7880
rect 14464 7760 14516 7812
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 19248 7692 19300 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 9220 7352 9272 7404
rect 10968 7352 11020 7404
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 12808 7327 12860 7336
rect 10048 7216 10100 7268
rect 10600 7216 10652 7268
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 19800 7531 19852 7540
rect 19800 7497 19809 7531
rect 19809 7497 19843 7531
rect 19843 7497 19852 7531
rect 19800 7488 19852 7497
rect 17316 7395 17368 7404
rect 8576 7148 8628 7200
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 11888 7148 11940 7200
rect 13544 7216 13596 7268
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 17316 7352 17368 7361
rect 17224 7284 17276 7336
rect 20904 7420 20956 7472
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 20168 7352 20220 7404
rect 19156 7327 19208 7336
rect 19156 7293 19165 7327
rect 19165 7293 19199 7327
rect 19199 7293 19208 7327
rect 19156 7284 19208 7293
rect 14188 7148 14240 7200
rect 16580 7216 16632 7268
rect 19524 7284 19576 7336
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 16672 7148 16724 7200
rect 19340 7216 19392 7268
rect 17132 7148 17184 7200
rect 18604 7148 18656 7200
rect 18788 7148 18840 7200
rect 19524 7148 19576 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 11888 6944 11940 6996
rect 12716 6987 12768 6996
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 2688 6808 2740 6860
rect 13452 6876 13504 6928
rect 16120 6944 16172 6996
rect 15660 6919 15712 6928
rect 9680 6851 9732 6860
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 9680 6808 9732 6817
rect 10232 6808 10284 6860
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 14004 6851 14056 6860
rect 14004 6817 14013 6851
rect 14013 6817 14047 6851
rect 14047 6817 14056 6851
rect 14004 6808 14056 6817
rect 15660 6885 15669 6919
rect 15669 6885 15703 6919
rect 15703 6885 15712 6919
rect 15660 6876 15712 6885
rect 16304 6808 16356 6860
rect 16580 6808 16632 6860
rect 17500 6808 17552 6860
rect 18696 6808 18748 6860
rect 19432 6808 19484 6860
rect 15752 6783 15804 6792
rect 15752 6749 15761 6783
rect 15761 6749 15795 6783
rect 15795 6749 15804 6783
rect 15752 6740 15804 6749
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 13636 6715 13688 6724
rect 13636 6681 13645 6715
rect 13645 6681 13679 6715
rect 13679 6681 13688 6715
rect 13636 6672 13688 6681
rect 10968 6604 11020 6656
rect 13452 6604 13504 6656
rect 15108 6604 15160 6656
rect 16028 6604 16080 6656
rect 16856 6604 16908 6656
rect 17960 6604 18012 6656
rect 20168 6647 20220 6656
rect 20168 6613 20177 6647
rect 20177 6613 20211 6647
rect 20211 6613 20220 6647
rect 20168 6604 20220 6613
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 10232 6443 10284 6452
rect 10232 6409 10241 6443
rect 10241 6409 10275 6443
rect 10275 6409 10284 6443
rect 10232 6400 10284 6409
rect 11796 6400 11848 6452
rect 13820 6400 13872 6452
rect 16488 6400 16540 6452
rect 17500 6443 17552 6452
rect 13268 6332 13320 6384
rect 13912 6332 13964 6384
rect 17500 6409 17509 6443
rect 17509 6409 17543 6443
rect 17543 6409 17552 6443
rect 17500 6400 17552 6409
rect 19248 6400 19300 6452
rect 11612 6264 11664 6316
rect 13728 6307 13780 6316
rect 6828 6196 6880 6248
rect 9680 6196 9732 6248
rect 10692 6196 10744 6248
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 17960 6264 18012 6316
rect 14004 6196 14056 6248
rect 16856 6196 16908 6248
rect 17316 6196 17368 6248
rect 20260 6332 20312 6384
rect 7748 6128 7800 6180
rect 9036 6128 9088 6180
rect 12624 6128 12676 6180
rect 15016 6128 15068 6180
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 13636 6103 13688 6112
rect 11152 6060 11204 6069
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 15936 6128 15988 6180
rect 17776 6128 17828 6180
rect 20628 6196 20680 6248
rect 18696 6128 18748 6180
rect 17132 6060 17184 6112
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 19708 6103 19760 6112
rect 19708 6069 19717 6103
rect 19717 6069 19751 6103
rect 19751 6069 19760 6103
rect 19708 6060 19760 6069
rect 19800 6060 19852 6112
rect 20904 6103 20956 6112
rect 20904 6069 20913 6103
rect 20913 6069 20947 6103
rect 20947 6069 20956 6103
rect 20904 6060 20956 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 7656 5856 7708 5908
rect 9128 5856 9180 5908
rect 19524 5856 19576 5908
rect 19616 5856 19668 5908
rect 1216 5788 1268 5840
rect 12348 5788 12400 5840
rect 12440 5788 12492 5840
rect 15108 5788 15160 5840
rect 7196 5720 7248 5772
rect 10692 5720 10744 5772
rect 13452 5720 13504 5772
rect 13912 5720 13964 5772
rect 7380 5652 7432 5704
rect 10140 5695 10192 5704
rect 7748 5627 7800 5636
rect 7748 5593 7757 5627
rect 7757 5593 7791 5627
rect 7791 5593 7800 5627
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 7748 5584 7800 5593
rect 9772 5584 9824 5636
rect 6736 5516 6788 5568
rect 11796 5652 11848 5704
rect 14464 5652 14516 5704
rect 16488 5720 16540 5772
rect 16856 5720 16908 5772
rect 16764 5695 16816 5704
rect 13728 5584 13780 5636
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 17224 5652 17276 5704
rect 17684 5695 17736 5704
rect 17684 5661 17693 5695
rect 17693 5661 17727 5695
rect 17727 5661 17736 5695
rect 17684 5652 17736 5661
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 18512 5652 18564 5704
rect 17132 5584 17184 5636
rect 19800 5720 19852 5772
rect 19432 5652 19484 5704
rect 19892 5652 19944 5704
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 11888 5516 11940 5568
rect 12164 5559 12216 5568
rect 12164 5525 12173 5559
rect 12173 5525 12207 5559
rect 12207 5525 12216 5559
rect 12164 5516 12216 5525
rect 13360 5516 13412 5568
rect 16672 5516 16724 5568
rect 18696 5516 18748 5568
rect 19800 5516 19852 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 10140 5312 10192 5364
rect 12624 5355 12676 5364
rect 12624 5321 12633 5355
rect 12633 5321 12667 5355
rect 12667 5321 12676 5355
rect 12624 5312 12676 5321
rect 13636 5355 13688 5364
rect 13636 5321 13645 5355
rect 13645 5321 13679 5355
rect 13679 5321 13688 5355
rect 13636 5312 13688 5321
rect 15752 5312 15804 5364
rect 17684 5312 17736 5364
rect 19064 5312 19116 5364
rect 19340 5355 19392 5364
rect 19340 5321 19349 5355
rect 19349 5321 19383 5355
rect 19383 5321 19392 5355
rect 19340 5312 19392 5321
rect 9680 5244 9732 5296
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 15016 5244 15068 5296
rect 13544 5176 13596 5228
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 17592 5176 17644 5228
rect 19800 5219 19852 5228
rect 19800 5185 19809 5219
rect 19809 5185 19843 5219
rect 19843 5185 19852 5219
rect 19800 5176 19852 5185
rect 19892 5219 19944 5228
rect 19892 5185 19901 5219
rect 19901 5185 19935 5219
rect 19935 5185 19944 5219
rect 19892 5176 19944 5185
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 10048 5108 10100 5160
rect 14372 5108 14424 5160
rect 18788 5108 18840 5160
rect 19708 5151 19760 5160
rect 7196 4972 7248 5024
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 9864 4972 9916 5024
rect 11244 5040 11296 5092
rect 11704 5040 11756 5092
rect 13820 5040 13872 5092
rect 17684 5040 17736 5092
rect 19708 5117 19717 5151
rect 19717 5117 19751 5151
rect 19751 5117 19760 5151
rect 19708 5108 19760 5117
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 21088 5040 21140 5092
rect 11612 5015 11664 5024
rect 11612 4981 11621 5015
rect 11621 4981 11655 5015
rect 11655 4981 11664 5015
rect 11612 4972 11664 4981
rect 12992 5015 13044 5024
rect 12992 4981 13001 5015
rect 13001 4981 13035 5015
rect 13035 4981 13044 5015
rect 12992 4972 13044 4981
rect 14188 4972 14240 5024
rect 16580 5015 16632 5024
rect 16580 4981 16589 5015
rect 16589 4981 16623 5015
rect 16623 4981 16632 5015
rect 16580 4972 16632 4981
rect 18788 5015 18840 5024
rect 18788 4981 18797 5015
rect 18797 4981 18831 5015
rect 18831 4981 18840 5015
rect 18788 4972 18840 4981
rect 19524 4972 19576 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 7380 4768 7432 4820
rect 8300 4768 8352 4820
rect 11060 4768 11112 4820
rect 12992 4768 13044 4820
rect 19800 4768 19852 4820
rect 4712 4700 4764 4752
rect 4252 4632 4304 4684
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 8484 4632 8536 4684
rect 16580 4700 16632 4752
rect 17316 4675 17368 4684
rect 7380 4564 7432 4616
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 17960 4632 18012 4684
rect 20168 4700 20220 4752
rect 10416 4564 10468 4616
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 12164 4564 12216 4616
rect 11152 4496 11204 4548
rect 17592 4428 17644 4480
rect 20536 4471 20588 4480
rect 20536 4437 20545 4471
rect 20545 4437 20579 4471
rect 20579 4437 20588 4471
rect 20536 4428 20588 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 8944 4224 8996 4276
rect 17040 4224 17092 4276
rect 19064 4224 19116 4276
rect 1768 4088 1820 4140
rect 2688 4088 2740 4140
rect 6828 4088 6880 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 13452 4156 13504 4208
rect 13912 4088 13964 4140
rect 14004 4088 14056 4140
rect 5632 3952 5684 4004
rect 10600 4020 10652 4072
rect 14188 4020 14240 4072
rect 15384 4088 15436 4140
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 16304 4088 16356 4140
rect 19248 4156 19300 4208
rect 19892 4156 19944 4208
rect 17316 4088 17368 4140
rect 19156 4088 19208 4140
rect 8208 3952 8260 4004
rect 6644 3884 6696 3936
rect 9956 3952 10008 4004
rect 13452 3952 13504 4004
rect 13636 3952 13688 4004
rect 15660 3952 15712 4004
rect 17960 4020 18012 4072
rect 19432 4020 19484 4072
rect 20536 4088 20588 4140
rect 21364 4088 21416 4140
rect 20812 4020 20864 4072
rect 18512 3952 18564 4004
rect 19064 3952 19116 4004
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 12532 3884 12584 3936
rect 12716 3884 12768 3936
rect 13820 3884 13872 3936
rect 14372 3884 14424 3936
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 15476 3884 15528 3893
rect 15568 3927 15620 3936
rect 15568 3893 15577 3927
rect 15577 3893 15611 3927
rect 15611 3893 15620 3927
rect 15568 3884 15620 3893
rect 15752 3884 15804 3936
rect 17500 3884 17552 3936
rect 19156 3884 19208 3936
rect 19248 3884 19300 3936
rect 19708 3927 19760 3936
rect 19708 3893 19717 3927
rect 19717 3893 19751 3927
rect 19751 3893 19760 3927
rect 19708 3884 19760 3893
rect 19892 3884 19944 3936
rect 20352 3884 20404 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3424 3680 3476 3732
rect 4712 3680 4764 3732
rect 8208 3680 8260 3732
rect 9680 3680 9732 3732
rect 11796 3680 11848 3732
rect 12808 3680 12860 3732
rect 12992 3680 13044 3732
rect 2320 3612 2372 3664
rect 8852 3612 8904 3664
rect 8944 3612 8996 3664
rect 11704 3612 11756 3664
rect 14648 3612 14700 3664
rect 16948 3680 17000 3732
rect 17684 3723 17736 3732
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 18328 3680 18380 3732
rect 18420 3680 18472 3732
rect 17592 3612 17644 3664
rect 2872 3544 2924 3596
rect 4252 3544 4304 3596
rect 6828 3544 6880 3596
rect 8208 3544 8260 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10692 3544 10744 3596
rect 11888 3544 11940 3596
rect 14372 3544 14424 3596
rect 15016 3544 15068 3596
rect 12992 3476 13044 3528
rect 14096 3476 14148 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 17040 3544 17092 3596
rect 18512 3612 18564 3664
rect 18788 3680 18840 3732
rect 18052 3544 18104 3596
rect 19800 3680 19852 3732
rect 20168 3680 20220 3732
rect 20628 3680 20680 3732
rect 21916 3680 21968 3732
rect 20720 3612 20772 3664
rect 17960 3476 18012 3528
rect 21088 3544 21140 3596
rect 14464 3451 14516 3460
rect 14464 3417 14473 3451
rect 14473 3417 14507 3451
rect 14507 3417 14516 3451
rect 14464 3408 14516 3417
rect 6920 3340 6972 3392
rect 10784 3340 10836 3392
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 12348 3340 12400 3392
rect 17500 3408 17552 3460
rect 19156 3408 19208 3460
rect 20536 3476 20588 3528
rect 19708 3408 19760 3460
rect 20904 3408 20956 3460
rect 16488 3340 16540 3392
rect 20812 3340 20864 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 3976 3136 4028 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 9496 3136 9548 3188
rect 10692 3179 10744 3188
rect 8944 3068 8996 3120
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 10876 3136 10928 3188
rect 11152 3136 11204 3188
rect 14372 3179 14424 3188
rect 12256 3068 12308 3120
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8484 3043 8536 3052
rect 8484 3009 8493 3043
rect 8493 3009 8527 3043
rect 8527 3009 8536 3043
rect 8484 3000 8536 3009
rect 9404 2932 9456 2984
rect 11060 3000 11112 3052
rect 11796 3000 11848 3052
rect 12992 3068 13044 3120
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 664 2864 716 2916
rect 6920 2864 6972 2916
rect 10508 2932 10560 2984
rect 12900 2932 12952 2984
rect 12992 2975 13044 2984
rect 12992 2941 13001 2975
rect 13001 2941 13035 2975
rect 13035 2941 13044 2975
rect 12992 2932 13044 2941
rect 13636 2932 13688 2984
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 12808 2864 12860 2916
rect 13728 2864 13780 2916
rect 15384 3136 15436 3188
rect 15476 3136 15528 3188
rect 17132 3136 17184 3188
rect 17592 3136 17644 3188
rect 17960 3136 18012 3188
rect 16212 3068 16264 3120
rect 20260 3068 20312 3120
rect 17132 3000 17184 3052
rect 18512 3043 18564 3052
rect 16488 2932 16540 2984
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 19432 3000 19484 3052
rect 17500 2932 17552 2984
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 19340 2932 19392 2941
rect 19984 2932 20036 2984
rect 20076 2932 20128 2984
rect 6092 2796 6144 2848
rect 8576 2796 8628 2848
rect 8852 2796 8904 2848
rect 10508 2796 10560 2848
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 15752 2864 15804 2916
rect 15844 2864 15896 2916
rect 15016 2796 15068 2848
rect 16212 2796 16264 2848
rect 16304 2796 16356 2848
rect 17224 2839 17276 2848
rect 17224 2805 17233 2839
rect 17233 2805 17267 2839
rect 17267 2805 17276 2839
rect 17224 2796 17276 2805
rect 17960 2796 18012 2848
rect 18604 2796 18656 2848
rect 19432 2796 19484 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 11428 2592 11480 2644
rect 11612 2592 11664 2644
rect 14096 2592 14148 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 14280 2592 14332 2601
rect 15108 2592 15160 2644
rect 15568 2592 15620 2644
rect 16028 2635 16080 2644
rect 16028 2601 16037 2635
rect 16037 2601 16071 2635
rect 16071 2601 16080 2635
rect 16028 2592 16080 2601
rect 19616 2592 19668 2644
rect 19984 2592 20036 2644
rect 7840 2524 7892 2576
rect 10508 2524 10560 2576
rect 15384 2524 15436 2576
rect 7196 2456 7248 2508
rect 8300 2456 8352 2508
rect 13360 2456 13412 2508
rect 7104 2388 7156 2440
rect 8208 2388 8260 2440
rect 10416 2388 10468 2440
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 13636 2388 13688 2440
rect 12716 2320 12768 2372
rect 17408 2456 17460 2508
rect 17776 2456 17828 2508
rect 18696 2456 18748 2508
rect 18880 2499 18932 2508
rect 18880 2465 18889 2499
rect 18889 2465 18923 2499
rect 18923 2465 18932 2499
rect 18880 2456 18932 2465
rect 19800 2456 19852 2508
rect 20444 2499 20496 2508
rect 20444 2465 20453 2499
rect 20453 2465 20487 2499
rect 20487 2465 20496 2499
rect 20444 2456 20496 2465
rect 14372 2388 14424 2440
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 16488 2388 16540 2440
rect 14280 2320 14332 2372
rect 17040 2320 17092 2372
rect 17960 2320 18012 2372
rect 11612 2252 11664 2304
rect 16488 2252 16540 2304
rect 17500 2252 17552 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 10416 2048 10468 2100
rect 16120 2048 16172 2100
rect 18788 2048 18840 2100
rect 20076 2048 20128 2100
rect 9864 1980 9916 2032
rect 16028 1980 16080 2032
<< metal2 >>
rect 5722 22000 5778 22800
rect 17130 22000 17186 22800
rect 18786 22536 18842 22545
rect 18786 22471 18842 22480
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 5736 19310 5764 22000
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4066 11520 4122 11529
rect 4066 11455 4122 11464
rect 4080 11286 4108 11455
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 1216 5840 1268 5846
rect 1216 5782 1268 5788
rect 202 3496 258 3505
rect 202 3431 258 3440
rect 216 800 244 3431
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 676 800 704 2858
rect 1228 800 1256 5782
rect 2700 4146 2728 6802
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 1780 800 1808 4082
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2332 800 2360 3606
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2884 800 2912 3538
rect 3436 800 3464 3674
rect 4264 3602 4292 4626
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4724 3738 4752 4694
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3988 800 4016 3130
rect 4908 2802 4936 8502
rect 4724 2774 4936 2802
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 1986 4752 2774
rect 4540 1958 4752 1986
rect 4540 800 4568 1958
rect 5092 800 5120 8774
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6736 5568 6788 5574
rect 6840 5522 6868 6190
rect 6788 5516 6868 5522
rect 6736 5510 6868 5516
rect 6748 5494 6868 5510
rect 6840 5166 6868 5494
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4146 6868 5102
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5644 800 5672 3946
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 6104 800 6132 2790
rect 6656 800 6684 3878
rect 6840 3602 6868 4082
rect 7024 3641 7052 19110
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 12728 18290 12756 19246
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 16132 18290 16160 19246
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7668 5914 7696 17682
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 5030 7236 5714
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7010 3632 7066 3641
rect 6828 3596 6880 3602
rect 7010 3567 7066 3576
rect 6828 3538 6880 3544
rect 6840 3058 6868 3538
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6932 2922 6960 3334
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 7116 2446 7144 4626
rect 7208 4622 7236 4966
rect 7392 4826 7420 5646
rect 7760 5642 7788 6122
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8312 4826 8340 14418
rect 9692 8634 9720 14418
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 7392 2650 7420 4558
rect 8220 4010 8248 4558
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3738 8248 3946
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8220 3194 8248 3538
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7208 800 7236 2450
rect 7852 1306 7880 2518
rect 8220 2446 8248 3130
rect 8496 3058 8524 4626
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8588 2854 8616 7142
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8864 3670 8892 4966
rect 8956 4282 8984 7890
rect 9232 7410 9260 8230
rect 9324 8090 9352 8434
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 9048 5234 9076 6122
rect 9140 5914 9168 6734
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9416 3942 9444 8298
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9692 6866 9720 7890
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9692 5302 9720 6190
rect 9784 5642 9812 18158
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 17202 11652 17682
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10612 7274 10640 8978
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9692 3738 9720 5238
rect 10060 5166 10088 7210
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10244 6458 10272 6802
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10244 5710 10272 6394
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10704 5778 10732 6190
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10152 5370 10180 5646
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4146 9904 4966
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8956 3126 8984 3606
rect 9692 3602 9720 3674
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9692 3346 9720 3538
rect 9416 3318 9720 3346
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 9416 2990 9444 3318
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8852 2848 8904 2854
rect 9508 2836 9536 3130
rect 8852 2790 8904 2796
rect 9416 2808 9536 2836
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 7760 1278 7880 1306
rect 7760 800 7788 1278
rect 8312 800 8340 2450
rect 8864 800 8892 2790
rect 9416 800 9444 2808
rect 9876 2038 9904 4082
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9864 2032 9916 2038
rect 9864 1974 9916 1980
rect 9968 800 9996 3946
rect 10428 2446 10456 4558
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 2990 10548 3878
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10520 2582 10548 2790
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10416 2440 10468 2446
rect 10612 2394 10640 4014
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10704 3194 10732 3538
rect 10796 3398 10824 9318
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10888 3194 10916 13806
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11716 9110 11744 10542
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11072 8430 11100 9046
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8566 11652 8978
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10980 8090 11008 8298
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10980 7410 11008 8026
rect 11072 7954 11100 8366
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6662 11008 7142
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11808 6458 11836 17070
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7206 11928 7890
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 7002 11928 7142
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11072 4826 11100 6054
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 11164 4554 11192 6054
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11256 4622 11284 5034
rect 11624 5030 11652 6258
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10704 2446 10732 3130
rect 11072 3058 11100 3334
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10416 2382 10468 2388
rect 10428 2106 10456 2382
rect 10520 2366 10640 2394
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10416 2100 10468 2106
rect 10416 2042 10468 2048
rect 10520 800 10548 2366
rect 11164 1442 11192 3130
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11440 2650 11468 2790
rect 11624 2650 11652 3878
rect 11716 3670 11744 5034
rect 11808 3738 11836 5646
rect 11900 5574 11928 6938
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11808 3058 11836 3674
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11900 3369 11928 3538
rect 11886 3360 11942 3369
rect 11886 3295 11942 3304
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11900 2446 11928 3295
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11072 1414 11192 1442
rect 11072 800 11100 1414
rect 11624 800 11652 2246
rect 12084 800 12112 9658
rect 12452 7546 12480 14894
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 5840 12400 5846
rect 12440 5840 12492 5846
rect 12400 5800 12440 5828
rect 12348 5782 12400 5788
rect 12440 5782 12492 5788
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 4622 12204 5510
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12544 3942 12572 13466
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13360 11620 13412 11626
rect 13360 11562 13412 11568
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 13096 9518 13124 11018
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12728 7002 12756 7890
rect 12820 7342 12848 8298
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12636 5370 12664 6122
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12360 3210 12388 3334
rect 12268 3182 12388 3210
rect 12268 3126 12296 3182
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12636 800 12664 2790
rect 12728 2378 12756 3878
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12820 2922 12848 3674
rect 12912 2990 12940 9386
rect 13004 9178 13032 9454
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12992 8968 13044 8974
rect 13096 8956 13124 9454
rect 13044 8928 13124 8956
rect 12992 8910 13044 8916
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 13004 7410 13032 8502
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13188 5386 13216 11086
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13280 7750 13308 10474
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 6390 13308 7686
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13372 5574 13400 11562
rect 13464 11150 13492 11630
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 11354 13584 11494
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13544 7268 13596 7274
rect 13544 7210 13596 7216
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13464 6662 13492 6870
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13556 5794 13584 7210
rect 13648 6730 13676 18158
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14108 17202 14136 17682
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13832 6458 13860 17070
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13924 11286 13952 11698
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13924 10810 13952 11222
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 8362 13952 8774
rect 14016 8634 14044 15506
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 14016 7018 14044 7958
rect 14108 7886 14136 8978
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 7954 14228 8230
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14200 7206 14228 7890
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14016 6990 14136 7018
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13464 5778 13584 5794
rect 13452 5772 13584 5778
rect 13504 5766 13584 5772
rect 13452 5714 13504 5720
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13188 5358 13400 5386
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13004 4826 13032 4966
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13004 3738 13032 4082
rect 13174 4040 13230 4049
rect 13174 3975 13230 3984
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3126 13032 3470
rect 12992 3120 13044 3126
rect 12992 3062 13044 3068
rect 13004 2990 13032 3062
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 13188 800 13216 3975
rect 13372 2514 13400 5358
rect 13556 5234 13584 5766
rect 13648 5370 13676 6054
rect 13740 5642 13768 6258
rect 13924 5778 13952 6326
rect 14016 6254 14044 6802
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13464 4010 13492 4150
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13648 2990 13676 3946
rect 13832 3942 13860 5034
rect 14108 4298 14136 6990
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 13924 4270 14136 4298
rect 13924 4146 13952 4270
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 14016 3369 14044 4082
rect 14200 4078 14228 4966
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14002 3360 14058 3369
rect 14002 3295 14058 3304
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13648 2446 13676 2926
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13740 800 13768 2858
rect 14108 2650 14136 3470
rect 14292 2650 14320 12650
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15304 11354 15332 18158
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16672 15972 16724 15978
rect 16672 15914 16724 15920
rect 16684 15026 16712 15914
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12238 15976 13262
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15396 11082 15424 11562
rect 15672 11354 15700 12174
rect 15948 12102 15976 12174
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15948 11694 15976 12038
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15856 11150 15884 11494
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15396 10674 15424 11018
rect 15764 10810 15792 11086
rect 16132 10810 16160 11630
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 14384 8838 14412 9386
rect 14568 9382 14596 10406
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15396 9042 15424 9454
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14384 8498 14412 8774
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14476 8430 14504 8774
rect 15120 8430 15148 8910
rect 15580 8634 15608 9998
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 16040 8362 16068 10406
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16132 8498 16160 9386
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15028 8090 15056 8230
rect 16316 8090 16344 10542
rect 16592 10062 16620 10746
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16500 9382 16528 9998
rect 16592 9518 16620 9998
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16500 9110 16528 9318
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14476 5710 14504 7754
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 15028 5302 15056 6122
rect 15120 5846 15148 6598
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 15672 5234 15700 6870
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15764 5370 15792 6734
rect 15948 6186 15976 6734
rect 16040 6662 16068 7890
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16132 7002 16160 7142
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16316 6866 16344 8026
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16500 6458 16528 8298
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16592 6866 16620 7210
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16500 5778 16528 6394
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16684 5574 16712 7142
rect 16776 5710 16804 13126
rect 16960 10266 16988 15982
rect 17144 13394 17172 22000
rect 17958 20224 18014 20233
rect 17958 20159 18014 20168
rect 17972 19174 18000 20159
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18800 19292 18828 22471
rect 20350 22128 20406 22137
rect 20350 22063 20406 22072
rect 20166 21584 20222 21593
rect 20166 21519 20222 21528
rect 19246 21176 19302 21185
rect 19246 21111 19302 21120
rect 18800 19264 18911 19292
rect 17960 19168 18012 19174
rect 18883 19145 18911 19264
rect 19260 19174 19288 21111
rect 20180 20058 20208 21519
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19248 19168 19300 19174
rect 17960 19110 18012 19116
rect 18878 19136 18934 19145
rect 19248 19110 19300 19116
rect 18878 19071 18934 19080
rect 18510 18864 18566 18873
rect 18510 18799 18566 18808
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17866 18320 17922 18329
rect 17866 18255 17922 18264
rect 17880 17882 17908 18255
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17972 12986 18000 18158
rect 18524 17610 18552 18799
rect 19996 18290 20024 19858
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 20088 18222 20116 19858
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 19800 17128 19852 17134
rect 19800 17070 19852 17076
rect 19812 16726 19840 17070
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 19800 16720 19852 16726
rect 19800 16662 19852 16668
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18524 15638 18552 16662
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 18512 15632 18564 15638
rect 18512 15574 18564 15580
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 19352 14482 19380 15506
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 19246 13832 19302 13841
rect 18880 13796 18932 13802
rect 19246 13767 19302 13776
rect 18880 13738 18932 13744
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17512 11898 17540 12242
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17512 11150 17540 11834
rect 17972 11762 18000 12582
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18524 11354 18552 12582
rect 18616 12374 18644 12786
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18616 11762 18644 12038
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16960 9586 16988 10066
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16960 8498 16988 8774
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16960 8022 16988 8434
rect 17052 8362 17080 11086
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 9178 17540 10406
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 6254 16896 6598
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 16776 5234 16804 5646
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14384 3942 14412 5102
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15120 4026 15148 5170
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4758 16620 4966
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 15028 3998 15148 4026
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14384 3194 14412 3538
rect 14464 3460 14516 3466
rect 14464 3402 14516 3408
rect 14476 3369 14504 3402
rect 14462 3360 14518 3369
rect 14462 3295 14518 3304
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14384 2446 14412 3130
rect 14660 2990 14688 3606
rect 15028 3602 15056 3998
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14292 800 14320 2314
rect 15028 1442 15056 2790
rect 15120 2650 15148 3878
rect 15396 3534 15424 4082
rect 15764 4026 15792 4082
rect 15672 4010 15792 4026
rect 15660 4004 15792 4010
rect 15712 3998 15792 4004
rect 15660 3946 15712 3952
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 3194 15424 3470
rect 15488 3194 15516 3878
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15580 2650 15608 3878
rect 15764 2922 15792 3878
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 14844 1414 15056 1442
rect 14844 800 14872 1414
rect 15396 800 15424 2518
rect 15856 898 15884 2858
rect 16224 2854 16252 3062
rect 16316 2854 16344 4082
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16500 2990 16528 3334
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16040 2038 16068 2586
rect 16500 2446 16528 2926
rect 16868 2689 16896 5714
rect 16960 3738 16988 7822
rect 17052 7018 17080 8298
rect 17144 7206 17172 8502
rect 17224 8288 17276 8294
rect 17224 8230 17276 8236
rect 17236 7342 17264 8230
rect 17406 7984 17462 7993
rect 17406 7919 17462 7928
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 7410 17356 7686
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17052 6990 17264 7018
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17144 5642 17172 6054
rect 17236 5710 17264 6990
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17052 3602 17080 4218
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17144 3194 17172 5578
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17144 3058 17172 3130
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17236 2854 17264 5646
rect 17328 4690 17356 6190
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17328 4146 17356 4626
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 16854 2680 16910 2689
rect 16854 2615 16910 2624
rect 17420 2514 17448 7919
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17512 6458 17540 6802
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17604 5386 17632 11154
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18524 10062 18552 10542
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 17880 9518 17908 9998
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 18524 9450 18552 9862
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17880 9178 17908 9318
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 18156 8974 18184 9386
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18524 8430 18552 8910
rect 18616 8498 18644 10406
rect 18800 10169 18828 10406
rect 18786 10160 18842 10169
rect 18786 10095 18842 10104
rect 18786 10024 18842 10033
rect 18786 9959 18842 9968
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18708 9722 18736 9862
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18708 9110 18736 9454
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18156 7954 18184 8230
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17866 7440 17922 7449
rect 17866 7375 17922 7384
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5710 17816 6122
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17512 5358 17632 5386
rect 17696 5370 17724 5646
rect 17684 5364 17736 5370
rect 17512 3942 17540 5358
rect 17684 5306 17736 5312
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17604 4486 17632 5170
rect 17880 5114 17908 7375
rect 18616 7206 18644 8230
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18602 7032 18658 7041
rect 18602 6967 18658 6976
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6322 18000 6598
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17684 5092 17736 5098
rect 17684 5034 17736 5040
rect 17788 5086 17908 5114
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17604 3670 17632 4422
rect 17696 3738 17724 5034
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 17512 2990 17540 3402
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16132 2106 16160 2382
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16120 2100 16172 2106
rect 16120 2042 16172 2048
rect 16028 2032 16080 2038
rect 16028 1974 16080 1980
rect 15856 870 15976 898
rect 15948 800 15976 870
rect 16500 800 16528 2246
rect 17052 800 17080 2314
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17512 800 17540 2246
rect 17604 2009 17632 3130
rect 17788 2514 17816 5086
rect 17960 4684 18012 4690
rect 17960 4626 18012 4632
rect 17972 4162 18000 4626
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18326 4176 18382 4185
rect 17972 4134 18092 4162
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17972 3777 18000 4014
rect 17958 3768 18014 3777
rect 17958 3703 18014 3712
rect 18064 3602 18092 4134
rect 18326 4111 18382 4120
rect 18340 3738 18368 4111
rect 18524 4010 18552 5646
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18418 3904 18474 3913
rect 18418 3839 18474 3848
rect 18432 3738 18460 3839
rect 18328 3732 18380 3738
rect 18328 3674 18380 3680
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18512 3664 18564 3670
rect 18512 3606 18564 3612
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17972 3194 18000 3470
rect 18524 3369 18552 3606
rect 18616 3516 18644 6967
rect 18708 6866 18736 8366
rect 18800 8294 18828 9959
rect 18892 8906 18920 13738
rect 19260 13530 19288 13767
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19444 12850 19472 13330
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11626 19012 12038
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18800 7546 18828 7890
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18708 6186 18736 6802
rect 18696 6180 18748 6186
rect 18696 6122 18748 6128
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18708 3618 18736 5510
rect 18800 5166 18828 7142
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18800 3738 18828 4966
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18708 3590 18828 3618
rect 18616 3488 18736 3516
rect 18510 3360 18566 3369
rect 18116 3292 18412 3312
rect 18510 3295 18566 3304
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18524 3058 18552 3295
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 17958 2952 18014 2961
rect 17958 2887 18014 2896
rect 17972 2854 18000 2887
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17590 2000 17646 2009
rect 17590 1935 17646 1944
rect 17972 1170 18000 2314
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18092 1170
rect 18064 800 18092 1142
rect 18616 800 18644 2790
rect 18708 2514 18736 3488
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18800 2106 18828 3590
rect 18892 2514 18920 7822
rect 19076 5370 19104 12718
rect 19246 12472 19302 12481
rect 19246 12407 19302 12416
rect 19260 12306 19288 12407
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19432 11620 19484 11626
rect 19432 11562 19484 11568
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19168 9178 19196 11154
rect 19352 11150 19380 11494
rect 19444 11150 19472 11562
rect 19340 11144 19392 11150
rect 19246 11112 19302 11121
rect 19340 11086 19392 11092
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19246 11047 19302 11056
rect 19260 9586 19288 11047
rect 19352 10826 19380 11086
rect 19352 10798 19472 10826
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19352 10130 19380 10678
rect 19444 10606 19472 10798
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19352 9722 19380 10066
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19168 7970 19196 9114
rect 19168 7942 19288 7970
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19260 7834 19288 7942
rect 19168 7342 19196 7822
rect 19260 7806 19380 7834
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 7410 19288 7686
rect 19352 7410 19380 7806
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19536 7342 19564 16594
rect 19996 15314 20024 18090
rect 20166 18048 20222 18057
rect 20166 17983 20222 17992
rect 20180 17338 20208 17983
rect 20272 17678 20300 18770
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20088 16114 20116 17070
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20166 15736 20222 15745
rect 20166 15671 20222 15680
rect 19996 15286 20116 15314
rect 19890 15192 19946 15201
rect 19890 15127 19946 15136
rect 19904 14618 19932 15127
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19720 13870 19748 14418
rect 19996 14414 20024 14894
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19614 8800 19670 8809
rect 19614 8735 19670 8744
rect 19628 8294 19656 8735
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19062 4312 19118 4321
rect 19062 4247 19064 4256
rect 19116 4247 19118 4256
rect 19064 4218 19116 4224
rect 19260 4214 19288 6394
rect 19352 5370 19380 7210
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6118 19472 6802
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19444 5710 19472 6054
rect 19536 5914 19564 7142
rect 19720 6225 19748 8230
rect 19812 7546 19840 12242
rect 19890 12064 19946 12073
rect 19890 11999 19946 12008
rect 19904 11354 19932 11999
rect 20088 11898 20116 15286
rect 20180 15162 20208 15671
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20272 12850 20300 14418
rect 20364 13870 20392 22063
rect 20626 20768 20682 20777
rect 20626 20703 20682 20712
rect 20640 20058 20668 20703
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20732 19514 20760 19751
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20442 19408 20498 19417
rect 20442 19343 20498 19352
rect 20456 18970 20484 19343
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20548 18358 20576 19246
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20718 17504 20774 17513
rect 20718 17439 20774 17448
rect 20732 17338 20760 17439
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20442 17096 20498 17105
rect 20442 17031 20498 17040
rect 20456 16794 20484 17031
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20718 16552 20774 16561
rect 20718 16487 20774 16496
rect 20732 16250 20760 16487
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20442 16144 20498 16153
rect 20442 16079 20498 16088
rect 20456 15706 20484 16079
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20442 14376 20498 14385
rect 20442 14311 20444 14320
rect 20496 14311 20498 14320
rect 20444 14282 20496 14288
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20548 13462 20576 14894
rect 20720 14816 20772 14822
rect 20718 14784 20720 14793
rect 20772 14784 20774 14793
rect 20718 14719 20774 14728
rect 20536 13456 20588 13462
rect 20536 13398 20588 13404
rect 20718 13424 20774 13433
rect 20718 13359 20774 13368
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20548 11694 20576 12174
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20536 11688 20588 11694
rect 20258 11656 20314 11665
rect 20536 11630 20588 11636
rect 20258 11591 20314 11600
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20180 10538 20208 11154
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 8430 19932 9862
rect 20180 9382 20208 10474
rect 20272 10130 20300 11591
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10198 20392 10406
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20364 9586 20392 10134
rect 20442 9752 20498 9761
rect 20442 9687 20498 9696
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20168 9376 20220 9382
rect 20074 9344 20130 9353
rect 20168 9318 20220 9324
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20074 9279 20130 9288
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19982 8392 20038 8401
rect 19982 8327 20038 8336
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19706 6216 19762 6225
rect 19706 6151 19762 6160
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19338 4720 19394 4729
rect 19338 4655 19394 4664
rect 19248 4208 19300 4214
rect 19248 4150 19300 4156
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 19076 1442 19104 3946
rect 19168 3942 19196 4082
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19156 3460 19208 3466
rect 19260 3448 19288 3878
rect 19208 3420 19288 3448
rect 19156 3402 19208 3408
rect 19352 2990 19380 4655
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19444 3058 19472 4014
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19340 2984 19392 2990
rect 19536 2938 19564 4966
rect 19340 2926 19392 2932
rect 19444 2910 19564 2938
rect 19444 2854 19472 2910
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19628 2650 19656 5850
rect 19720 5166 19748 6054
rect 19812 5778 19840 6054
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19812 5234 19840 5510
rect 19904 5234 19932 5646
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19708 3936 19760 3942
rect 19706 3904 19708 3913
rect 19760 3904 19762 3913
rect 19706 3839 19762 3848
rect 19812 3738 19840 4762
rect 19892 4208 19944 4214
rect 19892 4150 19944 4156
rect 19904 3942 19932 4150
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19076 1414 19196 1442
rect 19168 800 19196 1414
rect 19720 800 19748 3402
rect 19798 3224 19854 3233
rect 19798 3159 19854 3168
rect 19812 2514 19840 3159
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19904 2417 19932 3878
rect 19996 2990 20024 8327
rect 20088 2990 20116 9279
rect 20364 7954 20392 9318
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 20180 6662 20208 7346
rect 20168 6656 20220 6662
rect 20272 6633 20300 7822
rect 20168 6598 20220 6604
rect 20258 6624 20314 6633
rect 20180 4758 20208 6598
rect 20258 6559 20314 6568
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20272 5710 20300 6326
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20364 5556 20392 7890
rect 20272 5528 20392 5556
rect 20168 4752 20220 4758
rect 20168 4694 20220 4700
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19890 2408 19946 2417
rect 19890 2343 19946 2352
rect 19996 1057 20024 2586
rect 20076 2100 20128 2106
rect 20076 2042 20128 2048
rect 19982 1048 20038 1057
rect 19982 983 20038 992
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6090 0 6146 800
rect 6642 0 6698 800
rect 7194 0 7250 800
rect 7746 0 7802 800
rect 8298 0 8354 800
rect 8850 0 8906 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10506 0 10562 800
rect 11058 0 11114 800
rect 11610 0 11666 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20088 241 20116 2042
rect 20180 649 20208 3674
rect 20272 3505 20300 5528
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20258 3496 20314 3505
rect 20258 3431 20314 3440
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 20272 800 20300 3062
rect 20364 2689 20392 3878
rect 20350 2680 20406 2689
rect 20350 2615 20406 2624
rect 20364 1601 20392 2615
rect 20456 2514 20484 9687
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20548 8634 20576 8978
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20548 7886 20576 8570
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20640 6338 20668 12038
rect 20732 11898 20760 13359
rect 20902 13016 20958 13025
rect 20902 12951 20904 12960
rect 20956 12951 20958 12960
rect 20904 12922 20956 12928
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20810 10704 20866 10713
rect 20810 10639 20866 10648
rect 20824 9518 20852 10639
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20916 7478 20944 12718
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20640 6310 20760 6338
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20534 6080 20590 6089
rect 20534 6015 20590 6024
rect 20548 5166 20576 6015
rect 20536 5160 20588 5166
rect 20640 5137 20668 6190
rect 20536 5102 20588 5108
rect 20626 5128 20682 5137
rect 20626 5063 20682 5072
rect 20732 4978 20760 6310
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20810 5672 20866 5681
rect 20810 5607 20866 5616
rect 20640 4950 20760 4978
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 4146 20576 4422
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20548 3534 20576 4082
rect 20640 3738 20668 4950
rect 20718 4176 20774 4185
rect 20718 4111 20774 4120
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20732 3670 20760 4111
rect 20824 4078 20852 5607
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20916 3466 20944 6054
rect 21008 4049 21036 9318
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 20994 4040 21050 4049
rect 20994 3975 21050 3984
rect 21100 3602 21128 5034
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 20350 1592 20406 1601
rect 20350 1527 20406 1536
rect 20824 800 20852 3334
rect 21376 800 21404 4082
rect 21836 3862 22048 3890
rect 21836 3641 21864 3862
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21822 3632 21878 3641
rect 21822 3567 21878 3576
rect 21928 800 21956 3674
rect 22020 898 22048 3862
rect 22020 870 22508 898
rect 22480 800 22508 870
rect 20166 640 20222 649
rect 20166 575 20222 584
rect 20074 232 20130 241
rect 20074 167 20130 176
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
<< via2 >>
rect 18786 22480 18842 22536
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4066 11464 4122 11520
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 202 3440 258 3496
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7010 3576 7066 3632
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11886 3304 11942 3360
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 13174 3984 13230 4040
rect 14002 3304 14058 3360
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 17958 20168 18014 20224
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 20350 22072 20406 22128
rect 20166 21528 20222 21584
rect 19246 21120 19302 21176
rect 18878 19080 18934 19136
rect 18510 18808 18566 18864
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 17866 18264 17922 18320
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 19246 13776 19302 13832
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14462 3304 14518 3360
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 17406 7928 17462 7984
rect 16854 2624 16910 2680
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18786 10104 18842 10160
rect 18786 9968 18842 10024
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 17866 7384 17922 7440
rect 18602 6976 18658 7032
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17958 3712 18014 3768
rect 18326 4120 18382 4176
rect 18418 3848 18474 3904
rect 18510 3304 18566 3360
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 17958 2896 18014 2952
rect 17590 1944 17646 2000
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 19246 12416 19302 12472
rect 19246 11056 19302 11112
rect 20166 17992 20222 18048
rect 20166 15680 20222 15736
rect 19890 15136 19946 15192
rect 19614 8744 19670 8800
rect 19062 4276 19118 4312
rect 19062 4256 19064 4276
rect 19064 4256 19116 4276
rect 19116 4256 19118 4276
rect 19890 12008 19946 12064
rect 20626 20712 20682 20768
rect 20718 19760 20774 19816
rect 20442 19352 20498 19408
rect 20718 17448 20774 17504
rect 20442 17040 20498 17096
rect 20718 16496 20774 16552
rect 20442 16088 20498 16144
rect 20442 14340 20498 14376
rect 20442 14320 20444 14340
rect 20444 14320 20496 14340
rect 20496 14320 20498 14340
rect 20718 14764 20720 14784
rect 20720 14764 20772 14784
rect 20772 14764 20774 14784
rect 20718 14728 20774 14764
rect 20718 13368 20774 13424
rect 20258 11600 20314 11656
rect 20442 9696 20498 9752
rect 20074 9288 20130 9344
rect 19982 8336 20038 8392
rect 19706 6160 19762 6216
rect 19338 4664 19394 4720
rect 19706 3884 19708 3904
rect 19708 3884 19760 3904
rect 19760 3884 19762 3904
rect 19706 3848 19762 3884
rect 19798 3168 19854 3224
rect 20258 6568 20314 6624
rect 19890 2352 19946 2408
rect 19982 992 20038 1048
rect 20258 3440 20314 3496
rect 20350 2624 20406 2680
rect 20902 12980 20958 13016
rect 20902 12960 20904 12980
rect 20904 12960 20956 12980
rect 20956 12960 20958 12980
rect 20810 10648 20866 10704
rect 20534 6024 20590 6080
rect 20626 5072 20682 5128
rect 20810 5616 20866 5672
rect 20718 4120 20774 4176
rect 20994 3984 21050 4040
rect 20350 1536 20406 1592
rect 21822 3576 21878 3632
rect 20166 584 20222 640
rect 20074 176 20130 232
<< metal3 >>
rect 18781 22538 18847 22541
rect 22000 22538 22800 22568
rect 18781 22536 22800 22538
rect 18781 22480 18786 22536
rect 18842 22480 22800 22536
rect 18781 22478 22800 22480
rect 18781 22475 18847 22478
rect 22000 22448 22800 22478
rect 20345 22130 20411 22133
rect 22000 22130 22800 22160
rect 20345 22128 22800 22130
rect 20345 22072 20350 22128
rect 20406 22072 22800 22128
rect 20345 22070 22800 22072
rect 20345 22067 20411 22070
rect 22000 22040 22800 22070
rect 20161 21586 20227 21589
rect 22000 21586 22800 21616
rect 20161 21584 22800 21586
rect 20161 21528 20166 21584
rect 20222 21528 22800 21584
rect 20161 21526 22800 21528
rect 20161 21523 20227 21526
rect 22000 21496 22800 21526
rect 19241 21178 19307 21181
rect 22000 21178 22800 21208
rect 19241 21176 22800 21178
rect 19241 21120 19246 21176
rect 19302 21120 22800 21176
rect 19241 21118 22800 21120
rect 19241 21115 19307 21118
rect 22000 21088 22800 21118
rect 20621 20770 20687 20773
rect 22000 20770 22800 20800
rect 20621 20768 22800 20770
rect 20621 20712 20626 20768
rect 20682 20712 22800 20768
rect 20621 20710 22800 20712
rect 20621 20707 20687 20710
rect 22000 20680 22800 20710
rect 17953 20226 18019 20229
rect 22000 20226 22800 20256
rect 17953 20224 22800 20226
rect 17953 20168 17958 20224
rect 18014 20168 22800 20224
rect 17953 20166 22800 20168
rect 17953 20163 18019 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22000 20136 22800 20166
rect 14672 20095 14992 20096
rect 20713 19818 20779 19821
rect 22000 19818 22800 19848
rect 20713 19816 22800 19818
rect 20713 19760 20718 19816
rect 20774 19760 22800 19816
rect 20713 19758 22800 19760
rect 20713 19755 20779 19758
rect 22000 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 20437 19410 20503 19413
rect 22000 19410 22800 19440
rect 20437 19408 22800 19410
rect 20437 19352 20442 19408
rect 20498 19352 22800 19408
rect 20437 19350 22800 19352
rect 20437 19347 20503 19350
rect 22000 19320 22800 19350
rect 18873 19140 18939 19141
rect 18822 19138 18828 19140
rect 18782 19078 18828 19138
rect 18892 19136 18939 19140
rect 18934 19080 18939 19136
rect 18822 19076 18828 19078
rect 18892 19076 18939 19080
rect 18873 19075 18939 19076
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 18505 18866 18571 18869
rect 22000 18866 22800 18896
rect 18505 18864 22800 18866
rect 18505 18808 18510 18864
rect 18566 18808 22800 18864
rect 18505 18806 22800 18808
rect 18505 18803 18571 18806
rect 22000 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 22000 18458 22800 18488
rect 18830 18398 22800 18458
rect 17861 18322 17927 18325
rect 18830 18322 18890 18398
rect 22000 18368 22800 18398
rect 17861 18320 18890 18322
rect 17861 18264 17866 18320
rect 17922 18264 18890 18320
rect 17861 18262 18890 18264
rect 17861 18259 17927 18262
rect 20161 18050 20227 18053
rect 22000 18050 22800 18080
rect 20161 18048 22800 18050
rect 20161 17992 20166 18048
rect 20222 17992 22800 18048
rect 20161 17990 22800 17992
rect 20161 17987 20227 17990
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 22000 17960 22800 17990
rect 14672 17919 14992 17920
rect 20713 17506 20779 17509
rect 22000 17506 22800 17536
rect 20713 17504 22800 17506
rect 20713 17448 20718 17504
rect 20774 17448 22800 17504
rect 20713 17446 22800 17448
rect 20713 17443 20779 17446
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 22000 17416 22800 17446
rect 18104 17375 18424 17376
rect 20437 17098 20503 17101
rect 22000 17098 22800 17128
rect 20437 17096 22800 17098
rect 20437 17040 20442 17096
rect 20498 17040 22800 17096
rect 20437 17038 22800 17040
rect 20437 17035 20503 17038
rect 22000 17008 22800 17038
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 20713 16554 20779 16557
rect 22000 16554 22800 16584
rect 20713 16552 22800 16554
rect 20713 16496 20718 16552
rect 20774 16496 22800 16552
rect 20713 16494 22800 16496
rect 20713 16491 20779 16494
rect 22000 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 20437 16146 20503 16149
rect 22000 16146 22800 16176
rect 20437 16144 22800 16146
rect 20437 16088 20442 16144
rect 20498 16088 22800 16144
rect 20437 16086 22800 16088
rect 20437 16083 20503 16086
rect 22000 16056 22800 16086
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 20161 15738 20227 15741
rect 22000 15738 22800 15768
rect 20161 15736 22800 15738
rect 20161 15680 20166 15736
rect 20222 15680 22800 15736
rect 20161 15678 22800 15680
rect 20161 15675 20227 15678
rect 22000 15648 22800 15678
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 19885 15194 19951 15197
rect 22000 15194 22800 15224
rect 19885 15192 22800 15194
rect 19885 15136 19890 15192
rect 19946 15136 22800 15192
rect 19885 15134 22800 15136
rect 19885 15131 19951 15134
rect 22000 15104 22800 15134
rect 20713 14786 20779 14789
rect 22000 14786 22800 14816
rect 20713 14784 22800 14786
rect 20713 14728 20718 14784
rect 20774 14728 22800 14784
rect 20713 14726 22800 14728
rect 20713 14723 20779 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 22000 14696 22800 14726
rect 14672 14655 14992 14656
rect 20437 14378 20503 14381
rect 22000 14378 22800 14408
rect 20437 14376 22800 14378
rect 20437 14320 20442 14376
rect 20498 14320 22800 14376
rect 20437 14318 22800 14320
rect 20437 14315 20503 14318
rect 22000 14288 22800 14318
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 19241 13834 19307 13837
rect 22000 13834 22800 13864
rect 19241 13832 22800 13834
rect 19241 13776 19246 13832
rect 19302 13776 22800 13832
rect 19241 13774 22800 13776
rect 19241 13771 19307 13774
rect 22000 13744 22800 13774
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 20713 13426 20779 13429
rect 22000 13426 22800 13456
rect 20713 13424 22800 13426
rect 20713 13368 20718 13424
rect 20774 13368 22800 13424
rect 20713 13366 22800 13368
rect 20713 13363 20779 13366
rect 22000 13336 22800 13366
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 20897 13018 20963 13021
rect 22000 13018 22800 13048
rect 20897 13016 22800 13018
rect 20897 12960 20902 13016
rect 20958 12960 22800 13016
rect 20897 12958 22800 12960
rect 20897 12955 20963 12958
rect 22000 12928 22800 12958
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 19241 12474 19307 12477
rect 22000 12474 22800 12504
rect 19241 12472 22800 12474
rect 19241 12416 19246 12472
rect 19302 12416 22800 12472
rect 19241 12414 22800 12416
rect 19241 12411 19307 12414
rect 22000 12384 22800 12414
rect 19885 12066 19951 12069
rect 22000 12066 22800 12096
rect 19885 12064 22800 12066
rect 19885 12008 19890 12064
rect 19946 12008 22800 12064
rect 19885 12006 22800 12008
rect 19885 12003 19951 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 22000 11976 22800 12006
rect 18104 11935 18424 11936
rect 20253 11658 20319 11661
rect 22000 11658 22800 11688
rect 20253 11656 22800 11658
rect 20253 11600 20258 11656
rect 20314 11600 22800 11656
rect 20253 11598 22800 11600
rect 20253 11595 20319 11598
rect 22000 11568 22800 11598
rect 0 11522 800 11552
rect 4061 11522 4127 11525
rect 0 11520 4127 11522
rect 0 11464 4066 11520
rect 4122 11464 4127 11520
rect 0 11462 4127 11464
rect 0 11432 800 11462
rect 4061 11459 4127 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 19241 11114 19307 11117
rect 22000 11114 22800 11144
rect 19241 11112 22800 11114
rect 19241 11056 19246 11112
rect 19302 11056 22800 11112
rect 19241 11054 22800 11056
rect 19241 11051 19307 11054
rect 22000 11024 22800 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 20805 10706 20871 10709
rect 22000 10706 22800 10736
rect 20805 10704 22800 10706
rect 20805 10648 20810 10704
rect 20866 10648 22800 10704
rect 20805 10646 22800 10648
rect 20805 10643 20871 10646
rect 22000 10616 22800 10646
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 18781 10162 18847 10165
rect 22000 10162 22800 10192
rect 18781 10160 22800 10162
rect 18781 10104 18786 10160
rect 18842 10104 22800 10160
rect 18781 10102 22800 10104
rect 18781 10099 18847 10102
rect 22000 10072 22800 10102
rect 18781 10028 18847 10029
rect 18781 10026 18828 10028
rect 18736 10024 18828 10026
rect 18736 9968 18786 10024
rect 18736 9966 18828 9968
rect 18781 9964 18828 9966
rect 18892 9964 18898 10028
rect 18781 9963 18847 9964
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 20437 9754 20503 9757
rect 22000 9754 22800 9784
rect 20437 9752 22800 9754
rect 20437 9696 20442 9752
rect 20498 9696 22800 9752
rect 20437 9694 22800 9696
rect 20437 9691 20503 9694
rect 22000 9664 22800 9694
rect 20069 9346 20135 9349
rect 22000 9346 22800 9376
rect 20069 9344 22800 9346
rect 20069 9288 20074 9344
rect 20130 9288 22800 9344
rect 20069 9286 22800 9288
rect 20069 9283 20135 9286
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 22000 9256 22800 9286
rect 14672 9215 14992 9216
rect 19609 8802 19675 8805
rect 22000 8802 22800 8832
rect 19609 8800 22800 8802
rect 19609 8744 19614 8800
rect 19670 8744 22800 8800
rect 19609 8742 22800 8744
rect 19609 8739 19675 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 22000 8712 22800 8742
rect 18104 8671 18424 8672
rect 19977 8394 20043 8397
rect 22000 8394 22800 8424
rect 19977 8392 22800 8394
rect 19977 8336 19982 8392
rect 20038 8336 22800 8392
rect 19977 8334 22800 8336
rect 19977 8331 20043 8334
rect 22000 8304 22800 8334
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 17401 7986 17467 7989
rect 22000 7986 22800 8016
rect 17401 7984 22800 7986
rect 17401 7928 17406 7984
rect 17462 7928 22800 7984
rect 17401 7926 22800 7928
rect 17401 7923 17467 7926
rect 22000 7896 22800 7926
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 17861 7442 17927 7445
rect 22000 7442 22800 7472
rect 17861 7440 22800 7442
rect 17861 7384 17866 7440
rect 17922 7384 22800 7440
rect 17861 7382 22800 7384
rect 17861 7379 17927 7382
rect 22000 7352 22800 7382
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 18597 7034 18663 7037
rect 22000 7034 22800 7064
rect 18597 7032 22800 7034
rect 18597 6976 18602 7032
rect 18658 6976 22800 7032
rect 18597 6974 22800 6976
rect 18597 6971 18663 6974
rect 22000 6944 22800 6974
rect 20253 6626 20319 6629
rect 22000 6626 22800 6656
rect 20253 6624 22800 6626
rect 20253 6568 20258 6624
rect 20314 6568 22800 6624
rect 20253 6566 22800 6568
rect 20253 6563 20319 6566
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 22000 6536 22800 6566
rect 18104 6495 18424 6496
rect 19701 6220 19767 6221
rect 19701 6218 19748 6220
rect 19656 6216 19748 6218
rect 19656 6160 19706 6216
rect 19656 6158 19748 6160
rect 19701 6156 19748 6158
rect 19812 6156 19818 6220
rect 19701 6155 19767 6156
rect 20529 6082 20595 6085
rect 22000 6082 22800 6112
rect 20529 6080 22800 6082
rect 20529 6024 20534 6080
rect 20590 6024 22800 6080
rect 20529 6022 22800 6024
rect 20529 6019 20595 6022
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 22000 5992 22800 6022
rect 14672 5951 14992 5952
rect 20805 5674 20871 5677
rect 22000 5674 22800 5704
rect 20805 5672 22800 5674
rect 20805 5616 20810 5672
rect 20866 5616 22800 5672
rect 20805 5614 22800 5616
rect 20805 5611 20871 5614
rect 22000 5584 22800 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 20621 5130 20687 5133
rect 22000 5130 22800 5160
rect 20621 5128 22800 5130
rect 20621 5072 20626 5128
rect 20682 5072 22800 5128
rect 20621 5070 22800 5072
rect 20621 5067 20687 5070
rect 22000 5040 22800 5070
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 19333 4722 19399 4725
rect 22000 4722 22800 4752
rect 19333 4720 22800 4722
rect 19333 4664 19338 4720
rect 19394 4664 22800 4720
rect 19333 4662 22800 4664
rect 19333 4659 19399 4662
rect 22000 4632 22800 4662
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 19057 4314 19123 4317
rect 22000 4314 22800 4344
rect 19057 4312 22800 4314
rect 19057 4256 19062 4312
rect 19118 4256 22800 4312
rect 19057 4254 22800 4256
rect 19057 4251 19123 4254
rect 22000 4224 22800 4254
rect 18321 4178 18387 4181
rect 20713 4178 20779 4181
rect 18321 4176 20779 4178
rect 18321 4120 18326 4176
rect 18382 4120 20718 4176
rect 20774 4120 20779 4176
rect 18321 4118 20779 4120
rect 18321 4115 18387 4118
rect 20713 4115 20779 4118
rect 13169 4042 13235 4045
rect 20989 4042 21055 4045
rect 13169 4040 21055 4042
rect 13169 3984 13174 4040
rect 13230 3984 20994 4040
rect 21050 3984 21055 4040
rect 13169 3982 21055 3984
rect 13169 3979 13235 3982
rect 20989 3979 21055 3982
rect 18413 3906 18479 3909
rect 19701 3906 19767 3909
rect 18413 3904 19767 3906
rect 18413 3848 18418 3904
rect 18474 3848 19706 3904
rect 19762 3848 19767 3904
rect 18413 3846 19767 3848
rect 18413 3843 18479 3846
rect 19701 3843 19767 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 17953 3770 18019 3773
rect 22000 3770 22800 3800
rect 17953 3768 22800 3770
rect 17953 3712 17958 3768
rect 18014 3712 22800 3768
rect 17953 3710 22800 3712
rect 17953 3707 18019 3710
rect 22000 3680 22800 3710
rect 7005 3634 7071 3637
rect 21817 3634 21883 3637
rect 7005 3632 21883 3634
rect 7005 3576 7010 3632
rect 7066 3576 21822 3632
rect 21878 3576 21883 3632
rect 7005 3574 21883 3576
rect 7005 3571 7071 3574
rect 21817 3571 21883 3574
rect 197 3498 263 3501
rect 20253 3498 20319 3501
rect 197 3496 20319 3498
rect 197 3440 202 3496
rect 258 3440 20258 3496
rect 20314 3440 20319 3496
rect 197 3438 20319 3440
rect 197 3435 263 3438
rect 20253 3435 20319 3438
rect 11881 3362 11947 3365
rect 13997 3362 14063 3365
rect 14457 3362 14523 3365
rect 11881 3360 14523 3362
rect 11881 3304 11886 3360
rect 11942 3304 14002 3360
rect 14058 3304 14462 3360
rect 14518 3304 14523 3360
rect 11881 3302 14523 3304
rect 11881 3299 11947 3302
rect 13997 3299 14063 3302
rect 14457 3299 14523 3302
rect 18505 3362 18571 3365
rect 22000 3362 22800 3392
rect 18505 3360 22800 3362
rect 18505 3304 18510 3360
rect 18566 3304 22800 3360
rect 18505 3302 22800 3304
rect 18505 3299 18571 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 22000 3272 22800 3302
rect 18104 3231 18424 3232
rect 19793 3228 19859 3229
rect 19742 3226 19748 3228
rect 19702 3166 19748 3226
rect 19812 3224 19859 3228
rect 19854 3168 19859 3224
rect 19742 3164 19748 3166
rect 19812 3164 19859 3168
rect 19793 3163 19859 3164
rect 17953 2954 18019 2957
rect 22000 2954 22800 2984
rect 17953 2952 22800 2954
rect 17953 2896 17958 2952
rect 18014 2896 22800 2952
rect 17953 2894 22800 2896
rect 17953 2891 18019 2894
rect 22000 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 16849 2682 16915 2685
rect 20345 2682 20411 2685
rect 16849 2680 20411 2682
rect 16849 2624 16854 2680
rect 16910 2624 20350 2680
rect 20406 2624 20411 2680
rect 16849 2622 20411 2624
rect 16849 2619 16915 2622
rect 20345 2619 20411 2622
rect 19885 2410 19951 2413
rect 22000 2410 22800 2440
rect 19885 2408 22800 2410
rect 19885 2352 19890 2408
rect 19946 2352 22800 2408
rect 19885 2350 22800 2352
rect 19885 2347 19951 2350
rect 22000 2320 22800 2350
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 17585 2002 17651 2005
rect 22000 2002 22800 2032
rect 17585 2000 22800 2002
rect 17585 1944 17590 2000
rect 17646 1944 22800 2000
rect 17585 1942 22800 1944
rect 17585 1939 17651 1942
rect 22000 1912 22800 1942
rect 20345 1594 20411 1597
rect 22000 1594 22800 1624
rect 20345 1592 22800 1594
rect 20345 1536 20350 1592
rect 20406 1536 22800 1592
rect 20345 1534 22800 1536
rect 20345 1531 20411 1534
rect 22000 1504 22800 1534
rect 19977 1050 20043 1053
rect 22000 1050 22800 1080
rect 19977 1048 22800 1050
rect 19977 992 19982 1048
rect 20038 992 22800 1048
rect 19977 990 22800 992
rect 19977 987 20043 990
rect 22000 960 22800 990
rect 20161 642 20227 645
rect 22000 642 22800 672
rect 20161 640 22800 642
rect 20161 584 20166 640
rect 20222 584 22800 640
rect 20161 582 22800 584
rect 20161 579 20227 582
rect 22000 552 22800 582
rect 20069 234 20135 237
rect 22000 234 22800 264
rect 20069 232 22800 234
rect 20069 176 20074 232
rect 20130 176 22800 232
rect 20069 174 22800 176
rect 20069 171 20135 174
rect 22000 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 18828 19136 18892 19140
rect 18828 19080 18878 19136
rect 18878 19080 18892 19136
rect 18828 19076 18892 19080
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 18828 10024 18892 10028
rect 18828 9968 18842 10024
rect 18842 9968 18892 10024
rect 18828 9964 18892 9968
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 19748 6216 19812 6220
rect 19748 6160 19762 6216
rect 19762 6160 19812 6216
rect 19748 6156 19812 6160
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 19748 3224 19812 3228
rect 19748 3168 19798 3224
rect 19798 3168 19812 3224
rect 19748 3164 19812 3168
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18827 19140 18893 19141
rect 18827 19076 18828 19140
rect 18892 19076 18893 19140
rect 18827 19075 18893 19076
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18830 10029 18890 19075
rect 18827 10028 18893 10029
rect 18827 9964 18828 10028
rect 18892 9964 18893 10028
rect 18827 9963 18893 9964
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 19747 6220 19813 6221
rect 19747 6156 19748 6220
rect 19812 6156 19813 6220
rect 19747 6155 19813 6156
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 19750 3229 19810 6155
rect 19747 3228 19813 3229
rect 19747 3164 19748 3228
rect 19812 3164 19813 3228
rect 19747 3163 19813 3164
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608762085
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608762085
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608762085
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1608762085
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1608762085
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608762085
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608762085
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_199
timestamp 1608762085
transform 1 0 19412 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608762085
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1608762085
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1608762085
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1608762085
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608762085
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1608762085
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1608762085
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1608762085
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608762085
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1608762085
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1608762085
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1608762085
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608762085
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1608762085
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1608762085
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1608762085
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1608762085
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608762085
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608762085
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1608762085
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608762085
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608762085
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608762085
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608762085
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608762085
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608762085
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608762085
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608762085
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1608762085
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1608762085
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1608762085
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608762085
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_196
timestamp 1608762085
transform 1 0 19136 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_204
timestamp 1608762085
transform 1 0 19872 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608762085
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_167
timestamp 1608762085
transform 1 0 16468 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1608762085
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1608762085
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_155
timestamp 1608762085
transform 1 0 15364 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608762085
transform 1 0 12788 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_131
timestamp 1608762085
transform 1 0 13156 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_143
timestamp 1608762085
transform 1 0 14260 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608762085
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_114
timestamp 1608762085
transform 1 0 11592 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1608762085
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_90
timestamp 1608762085
transform 1 0 9384 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_102
timestamp 1608762085
transform 1 0 10488 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_66
timestamp 1608762085
transform 1 0 7176 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_78
timestamp 1608762085
transform 1 0 8280 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608762085
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608762085
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1608762085
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608762085
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1608762085
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1608762085
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608762085
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1608762085
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1608762085
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608762085
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608762085
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1608762085
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608762085
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608762085
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608762085
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1608762085
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_202
timestamp 1608762085
transform 1 0 19688 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1608762085
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608762085
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1608762085
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1608762085
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1608762085
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1608762085
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1608762085
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1608762085
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608762085
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1608762085
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1608762085
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1608762085
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1608762085
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1608762085
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608762085
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608762085
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1608762085
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608762085
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1608762085
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1608762085
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608762085
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_218
timestamp 1608762085
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 19504 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_190
timestamp 1608762085
transform 1 0 18584 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_198
timestamp 1608762085
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_206
timestamp 1608762085
transform 1 0 20056 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608762085
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1608762085
transform 1 0 17480 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1608762085
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 15824 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_153
timestamp 1608762085
transform 1 0 15180 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_159
timestamp 1608762085
transform 1 0 15732 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_166
timestamp 1608762085
transform 1 0 16376 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_129
timestamp 1608762085
transform 1 0 12972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_141
timestamp 1608762085
transform 1 0 14076 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608762085
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1608762085
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 9568 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_86
timestamp 1608762085
transform 1 0 9016 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1608762085
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1608762085
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608762085
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1608762085
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608762085
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1608762085
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1608762085
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1608762085
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608762085
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608762085
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1608762085
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608762085
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608762085
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1608762085
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608762085
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_194
timestamp 1608762085
transform 1 0 18952 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1608762085
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_170
timestamp 1608762085
transform 1 0 16744 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_182
timestamp 1608762085
transform 1 0 17848 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608762085
transform 1 0 15272 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608762085
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_148
timestamp 1608762085
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1608762085
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_158
timestamp 1608762085
transform 1 0 15640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_136
timestamp 1608762085
transform 1 0 13616 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608762085
transform 1 0 12144 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1608762085
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_117
timestamp 1608762085
transform 1 0 11868 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_124
timestamp 1608762085
transform 1 0 12512 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608762085
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1608762085
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1608762085
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 7544 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1608762085
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_76
timestamp 1608762085
transform 1 0 8096 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1608762085
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1608762085
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608762085
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1608762085
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1608762085
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608762085
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1608762085
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1608762085
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608762085
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608762085
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608762085
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1608762085
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608762085
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1608762085
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1608762085
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608762085
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1608762085
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1608762085
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608762085
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608762085
transform 1 0 19964 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 19504 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_190
timestamp 1608762085
transform 1 0 18584 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_198
timestamp 1608762085
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1608762085
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1608762085
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1608762085
transform 1 0 19872 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608762085
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1608762085
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1608762085
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1608762085
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608762085
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608762085
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1608762085
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1608762085
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1608762085
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 13800 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1608762085
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1608762085
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_135
timestamp 1608762085
transform 1 0 13524 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_144
timestamp 1608762085
transform 1 0 14352 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 11316 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608762085
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1608762085
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1608762085
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_110
timestamp 1608762085
transform 1 0 11224 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_117
timestamp 1608762085
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1608762085
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1608762085
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608762085
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1608762085
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1608762085
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1608762085
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1608762085
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1608762085
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1608762085
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608762085
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1608762085
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1608762085
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1608762085
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1608762085
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1608762085
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608762085
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608762085
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1608762085
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1608762085
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1608762085
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608762085
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608762085
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608762085
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1608762085
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1608762085
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1608762085
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608762085
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608762085
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1608762085
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1608762085
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 19596 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1608762085
transform 1 0 19136 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_200
timestamp 1608762085
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1608762085
transform 1 0 20148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608762085
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1608762085
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608762085
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1608762085
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1608762085
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1608762085
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608762085
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1608762085
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1608762085
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1608762085
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1608762085
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1608762085
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608762085
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1608762085
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608762085
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1608762085
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1608762085
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1608762085
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608762085
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608762085
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1608762085
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608762085
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608762085
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1608762085
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608762085
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608762085
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608762085
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1608762085
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_202
timestamp 1608762085
transform 1 0 19688 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1608762085
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608762085
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1608762085
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1608762085
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1608762085
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1608762085
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 13984 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_129
timestamp 1608762085
transform 1 0 12972 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1608762085
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1608762085
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1608762085
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608762085
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1608762085
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1608762085
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1608762085
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1608762085
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1608762085
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608762085
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1608762085
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1608762085
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608762085
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1608762085
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1608762085
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608762085
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608762085
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1608762085
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1608762085
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1608762085
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608762085
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1608762085
transform 1 0 19136 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_204
timestamp 1608762085
transform 1 0 19872 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608762085
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_177
timestamp 1608762085
transform 1 0 17388 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1608762085
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_153
timestamp 1608762085
transform 1 0 15180 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_165
timestamp 1608762085
transform 1 0 16284 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_129
timestamp 1608762085
transform 1 0 12972 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_141
timestamp 1608762085
transform 1 0 14076 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608762085
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1608762085
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1608762085
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1608762085
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1608762085
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608762085
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1608762085
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1608762085
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1608762085
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1608762085
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1608762085
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608762085
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1608762085
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1608762085
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608762085
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608762085
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608762085
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1608762085
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1608762085
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608762085
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608762085
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1608762085
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1608762085
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1608762085
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608762085
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1608762085
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1608762085
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1608762085
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_135
timestamp 1608762085
transform 1 0 13524 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1608762085
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1608762085
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608762085
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1608762085
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1608762085
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 8280 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_68
timestamp 1608762085
transform 1 0 7360 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1608762085
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608762085
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1608762085
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608762085
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608762085
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608762085
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608762085
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608762085
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608762085
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608762085
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_216
timestamp 1608762085
transform 1 0 20976 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608762085
transform 1 0 19872 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_196
timestamp 1608762085
transform 1 0 19136 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608762085
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1608762085
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1608762085
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1608762085
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1608762085
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1608762085
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608762085
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1608762085
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608762085
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 10672 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1608762085
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_98
timestamp 1608762085
transform 1 0 10120 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1608762085
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608762085
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1608762085
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608762085
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1608762085
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1608762085
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1608762085
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608762085
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608762085
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608762085
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608762085
transform 1 0 20700 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608762085
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608762085
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608762085
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1608762085
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1608762085
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1608762085
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608762085
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608762085
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608762085
transform 1 0 19044 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 19228 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 19964 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 19596 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1608762085
transform 1 0 18860 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1608762085
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1608762085
transform 1 0 18676 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1608762085
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1608762085
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1608762085
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608762085
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1608762085
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_179
timestamp 1608762085
transform 1 0 17572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 16100 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608762085
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608762085
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1608762085
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1608762085
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1608762085
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608762085
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1608762085
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608762085
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608762085
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1608762085
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608762085
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608762085
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608762085
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608762085
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1608762085
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1608762085
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608762085
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608762085
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608762085
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1608762085
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608762085
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608762085
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608762085
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1608762085
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608762085
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608762085
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608762085
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1608762085
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608762085
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608762085
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608762085
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608762085
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608762085
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608762085
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608762085
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608762085
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608762085
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608762085
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608762085
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1608762085
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1608762085
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1608762085
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1608762085
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1608762085
transform 1 0 19228 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 19780 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_195
timestamp 1608762085
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1608762085
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 17572 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1608762085
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608762085
transform 1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 15916 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608762085
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1608762085
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_159
timestamp 1608762085
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1608762085
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1608762085
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1608762085
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1608762085
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608762085
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1608762085
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1608762085
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1608762085
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1608762085
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1608762085
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608762085
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608762085
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608762085
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608762085
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608762085
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608762085
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608762085
transform 1 0 20516 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608762085
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_210
timestamp 1608762085
transform 1 0 20424 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1608762085
transform 1 0 20884 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1608762085
transform 1 0 21252 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 18584 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1608762085
transform 1 0 20056 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1608762085
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608762085
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1608762085
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_187
timestamp 1608762085
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 16100 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1608762085
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 14444 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1608762085
transform 1 0 13156 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 1608762085
transform 1 0 13984 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_144
timestamp 1608762085
transform 1 0 14352 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608762085
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1608762085
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1608762085
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1608762085
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1608762085
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1608762085
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608762085
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1608762085
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608762085
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1608762085
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1608762085
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1608762085
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608762085
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608762085
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608762085
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1608762085
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608762085
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608762085
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1608762085
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608762085
transform 1 0 19412 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608762085
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1608762085
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_208
timestamp 1608762085
transform 1 0 20240 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1608762085
transform 1 0 16560 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_167
timestamp 1608762085
transform 1 0 16468 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 1608762085
transform 1 0 17388 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_185
timestamp 1608762085
transform 1 0 18124 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1608762085
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608762085
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1608762085
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1608762085
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608762085
transform 1 0 12972 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 13432 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_126
timestamp 1608762085
transform 1 0 12696 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1608762085
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 12144 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1608762085
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_117
timestamp 1608762085
transform 1 0 11868 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608762085
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1608762085
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1608762085
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1608762085
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608762085
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1608762085
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608762085
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608762085
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608762085
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608762085
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608762085
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608762085
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608762085
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_214
timestamp 1608762085
transform 1 0 20792 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 19320 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1608762085
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1608762085
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608762085
transform 1 0 18308 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608762085
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608762085
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1608762085
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1608762085
transform 1 0 14812 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608762085
transform 1 0 16100 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1608762085
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_146
timestamp 1608762085
transform 1 0 14536 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_158
timestamp 1608762085
transform 1 0 15640 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_162
timestamp 1608762085
transform 1 0 16008 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_166
timestamp 1608762085
transform 1 0 16376 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_140
timestamp 1608762085
transform 1 0 13984 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 12512 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608762085
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1608762085
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_123
timestamp 1608762085
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1608762085
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1608762085
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1608762085
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608762085
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1608762085
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608762085
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1608762085
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1608762085
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1608762085
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608762085
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608762085
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608762085
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608762085
transform 1 0 20792 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608762085
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608762085
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608762085
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1608762085
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1608762085
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1608762085
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608762085
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608762085
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608762085
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 18492 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608762085
transform 1 0 19780 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_200
timestamp 1608762085
transform 1 0 19504 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_205
timestamp 1608762085
transform 1 0 19964 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1608762085
transform 1 0 17020 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 16836 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608762085
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1608762085
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1608762085
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1608762085
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_167
timestamp 1608762085
transform 1 0 16468 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1608762085
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 15364 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1608762085
transform 1 0 15640 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608762085
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1608762085
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1608762085
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 13708 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 12972 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1608762085
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1608762085
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1608762085
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608762085
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1608762085
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1608762085
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1608762085
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1608762085
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608762085
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1608762085
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1608762085
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1608762085
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1608762085
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1608762085
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1608762085
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608762085
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1608762085
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608762085
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1608762085
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1608762085
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1608762085
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608762085
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1608762085
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1608762085
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608762085
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608762085
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608762085
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608762085
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608762085
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608762085
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608762085
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608762085
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608762085
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608762085
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1608762085
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608762085
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608762085
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1608762085
transform 1 0 18676 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 19136 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1608762085
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1608762085
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608762085
transform 1 0 17388 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_173
timestamp 1608762085
transform 1 0 17020 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1608762085
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1608762085
transform 1 0 14628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 15548 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608762085
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1608762085
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1608762085
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 12972 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1608762085
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1608762085
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 11316 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 1608762085
transform 1 0 11224 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608762085
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762085
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1608762085
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_104
timestamp 1608762085
transform 1 0 10672 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1608762085
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1608762085
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608762085
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1608762085
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608762085
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608762085
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608762085
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608762085
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608762085
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608762085
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608762085
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_212
timestamp 1608762085
transform 1 0 20608 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 19136 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1608762085
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608762085
transform 1 0 17204 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608762085
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608762085
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1608762085
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1608762085
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_184
timestamp 1608762085
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1608762085
transform 1 0 14720 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1608762085
transform 1 0 15548 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1608762085
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk
timestamp 1608762085
transform 1 0 12880 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1608762085
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1608762085
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608762085
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1608762085
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1608762085
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1608762085
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 10212 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1608762085
transform 1 0 8832 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_93
timestamp 1608762085
transform 1 0 9660 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_74
timestamp 1608762085
transform 1 0 7912 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1608762085
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608762085
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608762085
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608762085
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1608762085
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608762085
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608762085
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608762085
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608762085
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608762085
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608762085
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608762085
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1608762085
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1608762085
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1608762085
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1608762085
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608762085
transform 1 0 19780 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_193
timestamp 1608762085
transform 1 0 18860 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp 1608762085
transform 1 0 19504 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 18308 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 17572 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1608762085
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_185
timestamp 1608762085
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 15916 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608762085
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608762085
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1608762085
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1608762085
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_159
timestamp 1608762085
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1608762085
transform 1 0 13524 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1608762085
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_144
timestamp 1608762085
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 11868 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_109
timestamp 1608762085
transform 1 0 11132 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608762085
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608762085
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_68
timestamp 1608762085
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608762085
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608762085
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608762085
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608762085
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608762085
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608762085
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608762085
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608762085
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608762085
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_212
timestamp 1608762085
transform 1 0 20608 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608762085
transform 1 0 18768 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608762085
transform 1 0 19780 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_190
timestamp 1608762085
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1608762085
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608762085
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1608762085
transform 1 0 16744 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608762085
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_168
timestamp 1608762085
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_179
timestamp 1608762085
transform 1 0 17572 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608762085
transform 1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_150
timestamp 1608762085
transform 1 0 14904 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_158
timestamp 1608762085
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 13432 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1608762085
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608762085
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608762085
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762085
transform 1 0 11500 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_111
timestamp 1608762085
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1608762085
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1608762085
transform 1 0 9384 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608762085
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 1608762085
transform 1 0 9016 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1608762085
transform 1 0 9660 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1608762085
transform 1 0 10396 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1608762085
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608762085
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1608762085
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608762085
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608762085
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1608762085
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1608762085
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608762085
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608762085
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608762085
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608762085
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608762085
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608762085
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608762085
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762085
transform 1 0 18768 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_191
timestamp 1608762085
transform 1 0 18676 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_208
timestamp 1608762085
transform 1 0 20240 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 16652 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_168
timestamp 1608762085
transform 1 0 16560 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_185
timestamp 1608762085
transform 1 0 18124 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608762085
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608762085
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608762085
transform 1 0 16284 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1608762085
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608762085
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608762085
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1608762085
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 11316 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1608762085
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608762085
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608762085
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_86
timestamp 1608762085
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608762085
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1608762085
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_80
timestamp 1608762085
transform 1 0 8464 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608762085
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608762085
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608762085
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608762085
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608762085
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608762085
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608762085
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608762085
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1608762085
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1608762085
transform 1 0 20700 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608762085
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608762085
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608762085
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1608762085
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_218
timestamp 1608762085
transform 1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_211
timestamp 1608762085
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 1608762085
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608762085
transform 1 0 19688 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608762085
transform 1 0 19688 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608762085
transform 1 0 18676 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_190
timestamp 1608762085
transform 1 0 18584 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_200
timestamp 1608762085
transform 1 0 19504 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_200
timestamp 1608762085
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 18032 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608762085
transform 1 0 17204 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608762085
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_173
timestamp 1608762085
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_184
timestamp 1608762085
transform 1 0 18032 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1608762085
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762085
transform 1 0 16100 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608762085
transform 1 0 16192 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608762085
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 1608762085
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_154
timestamp 1608762085
transform 1 0 15272 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_162
timestamp 1608762085
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_161
timestamp 1608762085
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 14444 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608762085
transform 1 0 13156 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1608762085
transform 1 0 14076 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_126
timestamp 1608762085
transform 1 0 12696 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_130
timestamp 1608762085
transform 1 0 13064 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_140
timestamp 1608762085
transform 1 0 13984 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_144
timestamp 1608762085
transform 1 0 14352 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608762085
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 10764 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608762085
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1608762085
transform 1 0 12236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1608762085
transform 1 0 11500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1608762085
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608762085
transform 1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 8832 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1608762085
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1608762085
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608762085
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1608762085
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1608762085
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_102
timestamp 1608762085
transform 1 0 10488 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_100
timestamp 1608762085
transform 1 0 10304 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 7176 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1608762085
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_73
timestamp 1608762085
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1608762085
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 6348 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608762085
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608762085
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1608762085
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608762085
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608762085
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1608762085
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608762085
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608762085
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608762085
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608762085
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608762085
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608762085
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608762085
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608762085
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608762085
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608762085
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608762085
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1608762085
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608762085
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1608762085
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1608762085
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608762085
transform 1 0 19320 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1608762085
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_207
timestamp 1608762085
transform 1 0 20148 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608762085
transform 1 0 18308 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608762085
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_173
timestamp 1608762085
transform 1 0 17020 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1608762085
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 1608762085
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1608762085
transform 1 0 15640 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608762085
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608762085
transform 1 0 14628 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1608762085
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_161
timestamp 1608762085
transform 1 0 15916 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608762085
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_134
timestamp 1608762085
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_145
timestamp 1608762085
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1608762085
transform 1 0 12604 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608762085
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1608762085
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608762085
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1608762085
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 10212 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608762085
transform 1 0 9936 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_89
timestamp 1608762085
transform 1 0 9292 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1608762085
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1608762085
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1608762085
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608762085
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608762085
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608762085
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608762085
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608762085
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608762085
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608762085
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608762085
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608762085
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608762085
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1608762085
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1608762085
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1608762085
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 19136 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1608762085
transform 1 0 18768 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762085
transform 1 0 17296 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1608762085
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608762085
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1608762085
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1608762085
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1608762085
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_166
timestamp 1608762085
transform 1 0 16376 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608762085
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1608762085
transform 1 0 12972 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_136
timestamp 1608762085
transform 1 0 13616 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608762085
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1608762085
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1608762085
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1608762085
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608762085
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1608762085
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1608762085
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1608762085
transform 1 0 7636 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_69
timestamp 1608762085
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608762085
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1608762085
transform 1 0 6624 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608762085
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1608762085
transform 1 0 6256 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608762085
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608762085
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608762085
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608762085
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608762085
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608762085
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1608762085
transform 1 0 20700 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608762085
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_211
timestamp 1608762085
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 1608762085
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608762085
transform 1 0 19688 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1608762085
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1608762085
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608762085
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_173
timestamp 1608762085
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1608762085
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1608762085
transform 1 0 15088 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_161
timestamp 1608762085
transform 1 0 15916 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608762085
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_132
timestamp 1608762085
transform 1 0 13248 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_144
timestamp 1608762085
transform 1 0 14352 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1608762085
transform 1 0 11592 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608762085
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608762085
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_105
timestamp 1608762085
transform 1 0 10764 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1608762085
transform 1 0 11500 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1608762085
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1608762085
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1608762085
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1608762085
transform 1 0 9384 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1608762085
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_99
timestamp 1608762085
transform 1 0 10212 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 7728 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1608762085
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608762085
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608762085
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608762085
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1608762085
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608762085
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608762085
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608762085
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608762085
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608762085
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1608762085
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608762085
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608762085
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_211
timestamp 1608762085
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1608762085
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608762085
transform 1 0 19688 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608762085
transform 1 0 18676 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_189
timestamp 1608762085
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_200
timestamp 1608762085
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1608762085
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608762085
transform 1 0 17664 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_171
timestamp 1608762085
transform 1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_178
timestamp 1608762085
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1608762085
transform 1 0 14720 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 15364 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608762085
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_146
timestamp 1608762085
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1608762085
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_154
timestamp 1608762085
transform 1 0 15272 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 13064 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_127
timestamp 1608762085
transform 1 0 12788 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 11316 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_109
timestamp 1608762085
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608762085
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1608762085
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 7084 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1608762085
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_81
timestamp 1608762085
transform 1 0 8556 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608762085
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_56
timestamp 1608762085
transform 1 0 6256 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608762085
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608762085
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608762085
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608762085
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608762085
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608762085
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608762085
transform 1 0 20424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1608762085
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608762085
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608762085
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608762085
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_214
timestamp 1608762085
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608762085
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_214
timestamp 1608762085
transform 1 0 20792 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1608762085
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1608762085
transform 1 0 19872 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1608762085
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1608762085
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_202
timestamp 1608762085
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_208
timestamp 1608762085
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1608762085
transform 1 0 19320 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1608762085
transform 1 0 19228 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_197
timestamp 1608762085
transform 1 0 19228 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1608762085
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1608762085
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1608762085
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1608762085
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1608762085
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608762085
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608762085
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608762085
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1608762085
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_180
timestamp 1608762085
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1608762085
transform 1 0 16928 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1608762085
transform 1 0 16836 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_167
timestamp 1608762085
transform 1 0 16468 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_171
timestamp 1608762085
transform 1 0 16836 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1608762085
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1608762085
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608762085
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608762085
transform 1 0 15180 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1608762085
transform 1 0 15640 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608762085
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1608762085
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1608762085
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1608762085
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608762085
transform 1 0 12972 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1608762085
transform 1 0 13248 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1608762085
transform 1 0 14260 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_129
timestamp 1608762085
transform 1 0 12972 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1608762085
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1608762085
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_145
timestamp 1608762085
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608762085
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608762085
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608762085
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608762085
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1608762085
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116
timestamp 1608762085
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1608762085
transform 1 0 10948 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1608762085
transform 1 0 11316 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_106
timestamp 1608762085
transform 1 0 10856 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_110
timestamp 1608762085
transform 1 0 11224 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_105
timestamp 1608762085
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 9292 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1608762085
transform 1 0 10028 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608762085
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1608762085
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1608762085
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1608762085
transform 1 0 8464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1608762085
transform 1 0 7360 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1608762085
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1608762085
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_77
timestamp 1608762085
transform 1 0 8188 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1608762085
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_83
timestamp 1608762085
transform 1 0 8740 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608762085
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608762085
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608762085
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608762085
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608762085
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51
timestamp 1608762085
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608762085
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608762085
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608762085
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608762085
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608762085
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608762085
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608762085
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608762085
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608762085
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608762085
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608762085
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1608762085
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 5722 22000 5778 22800 4 SC_IN_TOP
port 1 nsew
rlabel metal2 s 22466 0 22522 800 4 SC_OUT_BOT
port 2 nsew
rlabel metal2 s 202 0 258 800 4 bottom_left_grid_pin_1_
port 3 nsew
rlabel metal2 s 17130 22000 17186 22800 4 ccff_head
port 4 nsew
rlabel metal3 s 0 11432 800 11552 4 ccff_tail
port 5 nsew
rlabel metal3 s 22000 3680 22800 3800 4 chanx_right_in[0]
port 6 nsew
rlabel metal3 s 22000 8304 22800 8424 4 chanx_right_in[10]
port 7 nsew
rlabel metal3 s 22000 8712 22800 8832 4 chanx_right_in[11]
port 8 nsew
rlabel metal3 s 22000 9256 22800 9376 4 chanx_right_in[12]
port 9 nsew
rlabel metal3 s 22000 9664 22800 9784 4 chanx_right_in[13]
port 10 nsew
rlabel metal3 s 22000 10072 22800 10192 4 chanx_right_in[14]
port 11 nsew
rlabel metal3 s 22000 10616 22800 10736 4 chanx_right_in[15]
port 12 nsew
rlabel metal3 s 22000 11024 22800 11144 4 chanx_right_in[16]
port 13 nsew
rlabel metal3 s 22000 11568 22800 11688 4 chanx_right_in[17]
port 14 nsew
rlabel metal3 s 22000 11976 22800 12096 4 chanx_right_in[18]
port 15 nsew
rlabel metal3 s 22000 12384 22800 12504 4 chanx_right_in[19]
port 16 nsew
rlabel metal3 s 22000 4224 22800 4344 4 chanx_right_in[1]
port 17 nsew
rlabel metal3 s 22000 4632 22800 4752 4 chanx_right_in[2]
port 18 nsew
rlabel metal3 s 22000 5040 22800 5160 4 chanx_right_in[3]
port 19 nsew
rlabel metal3 s 22000 5584 22800 5704 4 chanx_right_in[4]
port 20 nsew
rlabel metal3 s 22000 5992 22800 6112 4 chanx_right_in[5]
port 21 nsew
rlabel metal3 s 22000 6536 22800 6656 4 chanx_right_in[6]
port 22 nsew
rlabel metal3 s 22000 6944 22800 7064 4 chanx_right_in[7]
port 23 nsew
rlabel metal3 s 22000 7352 22800 7472 4 chanx_right_in[8]
port 24 nsew
rlabel metal3 s 22000 7896 22800 8016 4 chanx_right_in[9]
port 25 nsew
rlabel metal3 s 22000 12928 22800 13048 4 chanx_right_out[0]
port 26 nsew
rlabel metal3 s 22000 17416 22800 17536 4 chanx_right_out[10]
port 27 nsew
rlabel metal3 s 22000 17960 22800 18080 4 chanx_right_out[11]
port 28 nsew
rlabel metal3 s 22000 18368 22800 18488 4 chanx_right_out[12]
port 29 nsew
rlabel metal3 s 22000 18776 22800 18896 4 chanx_right_out[13]
port 30 nsew
rlabel metal3 s 22000 19320 22800 19440 4 chanx_right_out[14]
port 31 nsew
rlabel metal3 s 22000 19728 22800 19848 4 chanx_right_out[15]
port 32 nsew
rlabel metal3 s 22000 20136 22800 20256 4 chanx_right_out[16]
port 33 nsew
rlabel metal3 s 22000 20680 22800 20800 4 chanx_right_out[17]
port 34 nsew
rlabel metal3 s 22000 21088 22800 21208 4 chanx_right_out[18]
port 35 nsew
rlabel metal3 s 22000 21496 22800 21616 4 chanx_right_out[19]
port 36 nsew
rlabel metal3 s 22000 13336 22800 13456 4 chanx_right_out[1]
port 37 nsew
rlabel metal3 s 22000 13744 22800 13864 4 chanx_right_out[2]
port 38 nsew
rlabel metal3 s 22000 14288 22800 14408 4 chanx_right_out[3]
port 39 nsew
rlabel metal3 s 22000 14696 22800 14816 4 chanx_right_out[4]
port 40 nsew
rlabel metal3 s 22000 15104 22800 15224 4 chanx_right_out[5]
port 41 nsew
rlabel metal3 s 22000 15648 22800 15768 4 chanx_right_out[6]
port 42 nsew
rlabel metal3 s 22000 16056 22800 16176 4 chanx_right_out[7]
port 43 nsew
rlabel metal3 s 22000 16464 22800 16584 4 chanx_right_out[8]
port 44 nsew
rlabel metal3 s 22000 17008 22800 17128 4 chanx_right_out[9]
port 45 nsew
rlabel metal2 s 662 0 718 800 4 chany_bottom_in[0]
port 46 nsew
rlabel metal2 s 6090 0 6146 800 4 chany_bottom_in[10]
port 47 nsew
rlabel metal2 s 6642 0 6698 800 4 chany_bottom_in[11]
port 48 nsew
rlabel metal2 s 7194 0 7250 800 4 chany_bottom_in[12]
port 49 nsew
rlabel metal2 s 7746 0 7802 800 4 chany_bottom_in[13]
port 50 nsew
rlabel metal2 s 8298 0 8354 800 4 chany_bottom_in[14]
port 51 nsew
rlabel metal2 s 8850 0 8906 800 4 chany_bottom_in[15]
port 52 nsew
rlabel metal2 s 9402 0 9458 800 4 chany_bottom_in[16]
port 53 nsew
rlabel metal2 s 9954 0 10010 800 4 chany_bottom_in[17]
port 54 nsew
rlabel metal2 s 10506 0 10562 800 4 chany_bottom_in[18]
port 55 nsew
rlabel metal2 s 11058 0 11114 800 4 chany_bottom_in[19]
port 56 nsew
rlabel metal2 s 1214 0 1270 800 4 chany_bottom_in[1]
port 57 nsew
rlabel metal2 s 1766 0 1822 800 4 chany_bottom_in[2]
port 58 nsew
rlabel metal2 s 2318 0 2374 800 4 chany_bottom_in[3]
port 59 nsew
rlabel metal2 s 2870 0 2926 800 4 chany_bottom_in[4]
port 60 nsew
rlabel metal2 s 3422 0 3478 800 4 chany_bottom_in[5]
port 61 nsew
rlabel metal2 s 3974 0 4030 800 4 chany_bottom_in[6]
port 62 nsew
rlabel metal2 s 4526 0 4582 800 4 chany_bottom_in[7]
port 63 nsew
rlabel metal2 s 5078 0 5134 800 4 chany_bottom_in[8]
port 64 nsew
rlabel metal2 s 5630 0 5686 800 4 chany_bottom_in[9]
port 65 nsew
rlabel metal2 s 11610 0 11666 800 4 chany_bottom_out[0]
port 66 nsew
rlabel metal2 s 17038 0 17094 800 4 chany_bottom_out[10]
port 67 nsew
rlabel metal2 s 17498 0 17554 800 4 chany_bottom_out[11]
port 68 nsew
rlabel metal2 s 18050 0 18106 800 4 chany_bottom_out[12]
port 69 nsew
rlabel metal2 s 18602 0 18658 800 4 chany_bottom_out[13]
port 70 nsew
rlabel metal2 s 19154 0 19210 800 4 chany_bottom_out[14]
port 71 nsew
rlabel metal2 s 19706 0 19762 800 4 chany_bottom_out[15]
port 72 nsew
rlabel metal2 s 20258 0 20314 800 4 chany_bottom_out[16]
port 73 nsew
rlabel metal2 s 20810 0 20866 800 4 chany_bottom_out[17]
port 74 nsew
rlabel metal2 s 21362 0 21418 800 4 chany_bottom_out[18]
port 75 nsew
rlabel metal2 s 21914 0 21970 800 4 chany_bottom_out[19]
port 76 nsew
rlabel metal2 s 12070 0 12126 800 4 chany_bottom_out[1]
port 77 nsew
rlabel metal2 s 12622 0 12678 800 4 chany_bottom_out[2]
port 78 nsew
rlabel metal2 s 13174 0 13230 800 4 chany_bottom_out[3]
port 79 nsew
rlabel metal2 s 13726 0 13782 800 4 chany_bottom_out[4]
port 80 nsew
rlabel metal2 s 14278 0 14334 800 4 chany_bottom_out[5]
port 81 nsew
rlabel metal2 s 14830 0 14886 800 4 chany_bottom_out[6]
port 82 nsew
rlabel metal2 s 15382 0 15438 800 4 chany_bottom_out[7]
port 83 nsew
rlabel metal2 s 15934 0 15990 800 4 chany_bottom_out[8]
port 84 nsew
rlabel metal2 s 16486 0 16542 800 4 chany_bottom_out[9]
port 85 nsew
rlabel metal3 s 22000 22040 22800 22160 4 prog_clk_0_E_in
port 86 nsew
rlabel metal3 s 22000 144 22800 264 4 right_bottom_grid_pin_34_
port 87 nsew
rlabel metal3 s 22000 552 22800 672 4 right_bottom_grid_pin_35_
port 88 nsew
rlabel metal3 s 22000 960 22800 1080 4 right_bottom_grid_pin_36_
port 89 nsew
rlabel metal3 s 22000 1504 22800 1624 4 right_bottom_grid_pin_37_
port 90 nsew
rlabel metal3 s 22000 1912 22800 2032 4 right_bottom_grid_pin_38_
port 91 nsew
rlabel metal3 s 22000 2320 22800 2440 4 right_bottom_grid_pin_39_
port 92 nsew
rlabel metal3 s 22000 2864 22800 2984 4 right_bottom_grid_pin_40_
port 93 nsew
rlabel metal3 s 22000 3272 22800 3392 4 right_bottom_grid_pin_41_
port 94 nsew
rlabel metal3 s 22000 22448 22800 22568 4 right_top_grid_pin_1_
port 95 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 96 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 97 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22800
string GDS_FILE /ef/openfpga/openlane/runs/sb_0__2_/results/magic/sb_0__2_.gds
string GDS_END 669778
string GDS_START 81916
<< end >>
