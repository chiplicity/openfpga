VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 5378.840 BY 5966.160 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 142.080 51.880 142.680 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 588.160 5329.480 588.760 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 76.800 51.880 77.400 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 207.360 51.880 207.960 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.430 5921.720 91.710 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2330.320 5329.480 2330.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[100]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2403.080 5329.480 2403.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[101]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1971.280 51.880 1971.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[102]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2475.160 5329.480 2475.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[103]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 2036.560 51.880 2037.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[104]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2437.890 5921.720 2438.170 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[105]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3070.390 44.120 3070.670 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[106]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2547.920 5329.480 2548.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[107]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1056.050 44.120 1056.330 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1110.790 44.120 1111.070 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1165.070 44.120 1165.350 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1219.350 44.120 1219.630 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1274.090 44.120 1274.370 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1328.370 44.120 1328.650 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 272.640 51.880 273.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 468.480 51.880 469.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 729.600 51.880 730.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[18]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 594.210 5921.720 594.490 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[19]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.150 5921.720 175.430 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2035.850 44.120 2036.130 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[20]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2090.590 44.120 2090.870 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[21]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.930 5921.720 678.210 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[22]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 761.650 5921.720 761.930 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[23]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 794.880 51.880 795.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[24]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 860.160 51.880 860.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[25]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.370 5921.720 845.650 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[26]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 926.120 51.880 926.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[27]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 991.400 51.880 992.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[28]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2144.870 44.120 2145.150 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[29]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 152.280 5329.480 152.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2199.150 44.120 2199.430 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[30]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1056.680 51.880 1057.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[31]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 929.090 5921.720 929.370 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[32]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1121.960 51.880 1122.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[33]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.270 5921.720 1013.550 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[34]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 733.000 5329.480 733.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[35]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 805.760 5329.480 806.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[36]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 878.520 5329.480 879.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[37]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2253.890 44.120 2254.170 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[38]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2308.170 44.120 2308.450 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[39]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 370.560 5329.480 371.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2362.450 44.120 2362.730 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[40]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2417.190 44.120 2417.470 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[41]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 951.280 5329.480 951.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[42]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2471.470 44.120 2471.750 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[43]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1023.360 5329.480 1023.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[44]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1096.990 5921.720 1097.270 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[45]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1096.120 5329.480 1096.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[46]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1187.240 51.880 1187.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[47]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1180.710 5921.720 1180.990 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[48]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1168.880 5329.480 1169.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[49]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.710 44.120 76.990 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2525.750 44.120 2526.030 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[50]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1241.640 5329.480 1242.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[51]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1313.720 5329.480 1314.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[52]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1264.430 5921.720 1264.710 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[53]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1252.520 51.880 1253.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[54]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1348.150 5921.720 1348.430 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[55]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1386.480 5329.480 1387.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[56]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2580.490 44.120 2580.770 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[57]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2634.770 44.120 2635.050 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[58]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2689.050 44.120 2689.330 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[59]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.990 44.120 131.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1459.240 5329.480 1459.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[60]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1317.800 51.880 1318.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[61]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1532.000 5329.480 1532.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[62]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2743.790 44.120 2744.070 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[63]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1604.080 5329.480 1604.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[64]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1383.080 51.880 1383.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[65]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1432.330 5921.720 1432.610 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[66]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1448.360 51.880 1448.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[67]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1516.050 5921.720 1516.330 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[68]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1513.640 51.880 1514.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[69]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.270 44.120 185.550 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1578.920 51.880 1579.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[70]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1599.770 5921.720 1600.050 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[71]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1644.200 51.880 1644.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[72]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1709.480 51.880 1710.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[73]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1683.490 5921.720 1683.770 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[74]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1767.210 5921.720 1767.490 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[75]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1676.840 5329.480 1677.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[76]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.390 5921.720 1851.670 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[77]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2798.070 44.120 2798.350 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[78]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1935.110 5921.720 1935.390 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[79]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.550 44.120 239.830 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1775.440 51.880 1776.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[80]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1749.600 5329.480 1750.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[81]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2852.350 44.120 2852.630 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[82]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2907.090 44.120 2907.370 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[83]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2961.370 44.120 2961.650 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[84]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1822.360 5329.480 1822.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[85]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1894.440 5329.480 1895.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[86]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2018.830 5921.720 2019.110 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[87]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 1967.200 5329.480 1967.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[88]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1840.720 51.880 1841.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[89]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.290 44.120 294.570 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2102.550 5921.720 2102.830 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[90]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2039.960 5329.480 2040.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[91]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3015.650 44.120 3015.930 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[92]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2112.720 5329.480 2113.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[93]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1906.000 51.880 1906.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[94]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2186.270 5921.720 2186.550 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[95]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2269.990 5921.720 2270.270 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[96]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2184.800 5329.480 2185.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[97]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2257.560 5329.480 2258.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[98]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2354.170 5921.720 2354.450 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[99]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.570 44.120 348.850 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.870 5921.720 259.150 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3999.720 5329.480 4000.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[100]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[101]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 4126.880 51.880 4127.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[101]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3611.350 5921.720 3611.630 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[102]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4158.750 44.120 4159.030 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[103]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4213.490 44.120 4213.770 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[104]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[105]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4072.480 5329.480 4073.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[105]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4267.770 44.120 4268.050 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[106]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4322.050 44.120 4322.330 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[107]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.650 44.120 1382.930 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1437.390 44.120 1437.670 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1491.670 44.120 1491.950 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1545.950 44.120 1546.230 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1600.690 44.120 1600.970 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1654.970 44.120 1655.250 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 337.920 51.880 338.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 533.760 51.880 534.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2101.840 51.880 2102.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[18]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2620.680 5329.480 2621.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[19]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 342.590 5921.720 342.870 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3124.670 44.120 3124.950 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[20]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2521.610 5921.720 2521.890 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[21]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2605.330 5921.720 2605.610 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[22]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2689.050 5921.720 2689.330 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[23]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2167.120 51.880 2167.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[24]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2232.400 51.880 2233.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[25]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2297.680 51.880 2298.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[26]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3178.950 44.120 3179.230 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[27]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2362.960 51.880 2363.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[28]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2693.440 5329.480 2694.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[29]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 225.040 5329.480 225.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2428.240 51.880 2428.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[30]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2765.520 5329.480 2766.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[31]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2493.520 51.880 2494.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[32]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2558.800 51.880 2559.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[33]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2838.280 5329.480 2838.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[34]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2911.040 5329.480 2911.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[35]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3233.690 44.120 3233.970 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[36]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2624.760 51.880 2625.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[37]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3287.970 44.120 3288.250 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[38]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3342.250 44.120 3342.530 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[39]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 442.640 5329.480 443.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 2983.800 5329.480 2984.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[40]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2690.040 51.880 2690.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[41]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[42]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2755.320 51.880 2755.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[42]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[43]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3055.880 5329.480 3056.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[43]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3396.990 44.120 3397.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[44]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3451.270 44.120 3451.550 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[45]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.230 5921.720 2773.510 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[46]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2856.950 5921.720 2857.230 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[47]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[48]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2820.600 51.880 2821.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[48]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[49]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2885.880 51.880 2886.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[49]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 402.850 44.120 403.130 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[50]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2951.160 51.880 2951.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[50]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3505.550 44.120 3505.830 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[51]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3560.290 44.120 3560.570 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[52]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3614.570 44.120 3614.850 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[53]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3016.440 51.880 3017.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[54]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3668.850 44.120 3669.130 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[55]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3128.640 5329.480 3129.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[56]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2940.670 5921.720 2940.950 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[57]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[58]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3081.720 51.880 3082.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[58]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[59]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3147.000 51.880 3147.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[59]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.590 44.120 457.870 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3024.390 5921.720 3024.670 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[60]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3201.400 5329.480 3202.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[61]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[62]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3212.280 51.880 3212.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[62]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3723.590 44.120 3723.870 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[63]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[64]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3274.160 5329.480 3274.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[64]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3277.560 51.880 3278.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[65]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[66]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3346.240 5329.480 3346.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[66]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3777.870 44.120 3778.150 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[67]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3832.150 44.120 3832.430 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[68]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[69]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3342.840 51.880 3343.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[69]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.870 44.120 512.150 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3108.110 5921.720 3108.390 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[70]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[71]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3419.000 5329.480 3419.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[71]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3886.890 44.120 3887.170 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[72]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[73]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3491.760 5329.480 3492.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[73]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3408.120 51.880 3408.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[74]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[75]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3474.080 51.880 3474.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[75]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[76]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3539.360 51.880 3539.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[76]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[77]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3564.520 5329.480 3565.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[77]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3192.290 5921.720 3192.570 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[78]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[79]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3636.600 5329.480 3637.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[79]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.150 44.120 566.430 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3941.170 44.120 3941.450 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[80]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[81]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3604.640 51.880 3605.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[81]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[82]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3669.920 51.880 3670.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[82]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3276.010 5921.720 3276.290 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[83]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3709.360 5329.480 3709.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[84]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3995.450 44.120 3995.730 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[85]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3782.120 5329.480 3782.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[86]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[87]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3735.200 51.880 3735.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[87]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[88]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3854.880 5329.480 3855.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[88]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[89]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3800.480 51.880 3801.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[89]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.890 44.120 621.170 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4050.190 44.120 4050.470 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[90]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[91]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3865.760 51.880 3866.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[91]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4104.470 44.120 4104.750 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[92]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[93]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3931.040 51.880 3931.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[93]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3996.320 51.880 3996.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[94]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3359.730 5921.720 3360.010 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[95]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 3926.960 5329.480 3927.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[96]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3443.450 5921.720 3443.730 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[97]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 4061.600 51.880 4062.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[98]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3527.170 5921.720 3527.450 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[99]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.170 44.120 675.450 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 426.310 5921.720 426.590 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5890.800 51.880 5891.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[100]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5247.570 44.120 5247.850 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[101]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5597.040 5329.480 5597.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[102]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5669.120 5329.480 5669.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[103]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5741.880 5329.480 5742.480 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[104]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5814.640 5329.480 5815.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[105]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5301.850 44.120 5302.130 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[106]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5887.400 5329.480 5888.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[107]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.250 44.120 1709.530 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1763.990 44.120 1764.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1818.270 44.120 1818.550 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1872.550 44.120 1872.830 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1927.290 44.120 1927.570 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1981.570 44.120 1981.850 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 403.200 51.880 403.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 599.040 51.880 599.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4145.240 5329.480 4145.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[18]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4192.160 51.880 4192.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[19]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 510.030 5921.720 510.310 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3695.070 5921.720 3695.350 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[20]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4217.320 5329.480 4217.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[21]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3778.790 5921.720 3779.070 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[22]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4376.790 44.120 4377.070 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[23]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4431.070 44.120 4431.350 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[24]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4257.440 51.880 4258.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[25]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4323.400 51.880 4324.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[26]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4388.680 51.880 4389.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[27]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3862.510 5921.720 3862.790 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[28]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4453.960 51.880 4454.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[29]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 297.800 5329.480 298.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4519.240 51.880 4519.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[30]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4584.520 51.880 4585.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[31]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3946.230 5921.720 3946.510 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[32]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4029.950 5921.720 4030.230 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[33]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4114.130 5921.720 4114.410 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[34]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4290.080 5329.480 4290.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[35]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4649.800 51.880 4650.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[36]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4715.080 51.880 4715.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[37]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4485.350 44.120 4485.630 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[38]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4197.850 5921.720 4198.130 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[39]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 515.400 5329.480 516.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4540.090 44.120 4540.370 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[40]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4780.360 51.880 4780.960 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[41]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4281.570 5921.720 4281.850 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[42]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4365.290 5921.720 4365.570 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[43]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4449.010 5921.720 4449.290 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[44]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4533.190 5921.720 4533.470 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[45]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4362.840 5329.480 4363.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[46]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4435.600 5329.480 4436.200 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[47]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4845.640 51.880 4846.240 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[48]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4507.680 5329.480 4508.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[49]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 729.450 44.120 729.730 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4910.920 51.880 4911.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[50]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4580.440 5329.480 4581.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[51]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4594.370 44.120 4594.650 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[52]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4648.650 44.120 4648.930 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[53]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4653.200 5329.480 4653.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[54]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 4976.200 51.880 4976.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[55]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4725.960 5329.480 4726.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[56]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4703.390 44.120 4703.670 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[57]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4798.040 5329.480 4798.640 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[58]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4616.910 5921.720 4617.190 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[59]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 784.190 44.120 784.470 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4870.800 5329.480 4871.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[60]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 4943.560 5329.480 4944.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[61]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4700.630 5921.720 4700.910 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[62]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4757.670 44.120 4757.950 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[63]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5041.480 51.880 5042.080 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[64]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4784.350 5921.720 4784.630 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[65]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4811.950 44.120 4812.230 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[66]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5106.760 51.880 5107.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[67]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5016.320 5329.480 5016.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[68]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5172.720 51.880 5173.320 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[69]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 838.470 44.120 838.750 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5088.400 5329.480 5089.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[70]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5161.160 5329.480 5161.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[71]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4866.690 44.120 4866.970 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[72]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4920.970 44.120 4921.250 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[73]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4868.070 5921.720 4868.350 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[74]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5238.000 51.880 5238.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[75]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4975.250 44.120 4975.530 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[76]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4952.250 5921.720 4952.530 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[77]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5029.990 44.120 5030.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[78]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5233.920 5329.480 5234.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[79]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 892.750 44.120 893.030 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5035.970 5921.720 5036.250 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[80]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5303.280 51.880 5303.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[81]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5306.680 5329.480 5307.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[82]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5378.760 5329.480 5379.360 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[83]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5451.520 5329.480 5452.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[84]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5368.560 51.880 5369.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[85]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5433.840 51.880 5434.440 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[86]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5119.690 5921.720 5119.970 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[87]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5499.120 51.880 5499.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[88]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5084.270 44.120 5084.550 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[89]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 947.490 44.120 947.770 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5564.400 51.880 5565.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[90]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 5524.280 5329.480 5524.880 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[91]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5138.550 44.120 5138.830 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[92]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5629.680 51.880 5630.280 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[93]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5694.960 51.880 5695.560 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[94]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5760.240 51.880 5760.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[95]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5193.290 44.120 5193.570 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[96]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5203.410 5921.720 5203.690 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[97]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 5825.520 51.880 5826.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[98]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5287.130 5921.720 5287.410 5924.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[99]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1001.770 44.120 1002.050 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 5327.080 80.200 5329.480 80.800 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 664.320 51.880 664.920 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 5327.080 660.920 5329.480 661.520 ;
    END
  END sc_tail
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 5353.840 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 5378.840 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 105.000 81.945 5288.275 5906.655 ;
      LAYER met1 ;
        RECT 63.350 46.880 5314.110 5908.060 ;
      LAYER met2 ;
        RECT 63.370 5921.440 91.150 5921.770 ;
        RECT 91.990 5921.440 174.870 5921.770 ;
        RECT 175.710 5921.440 258.590 5921.770 ;
        RECT 259.430 5921.440 342.310 5921.770 ;
        RECT 343.150 5921.440 426.030 5921.770 ;
        RECT 426.870 5921.440 509.750 5921.770 ;
        RECT 510.590 5921.440 593.930 5921.770 ;
        RECT 594.770 5921.440 677.650 5921.770 ;
        RECT 678.490 5921.440 761.370 5921.770 ;
        RECT 762.210 5921.440 845.090 5921.770 ;
        RECT 845.930 5921.440 928.810 5921.770 ;
        RECT 929.650 5921.440 1012.990 5921.770 ;
        RECT 1013.830 5921.440 1096.710 5921.770 ;
        RECT 1097.550 5921.440 1180.430 5921.770 ;
        RECT 1181.270 5921.440 1264.150 5921.770 ;
        RECT 1264.990 5921.440 1347.870 5921.770 ;
        RECT 1348.710 5921.440 1432.050 5921.770 ;
        RECT 1432.890 5921.440 1515.770 5921.770 ;
        RECT 1516.610 5921.440 1599.490 5921.770 ;
        RECT 1600.330 5921.440 1683.210 5921.770 ;
        RECT 1684.050 5921.440 1766.930 5921.770 ;
        RECT 1767.770 5921.440 1851.110 5921.770 ;
        RECT 1851.950 5921.440 1934.830 5921.770 ;
        RECT 1935.670 5921.440 2018.550 5921.770 ;
        RECT 2019.390 5921.440 2102.270 5921.770 ;
        RECT 2103.110 5921.440 2185.990 5921.770 ;
        RECT 2186.830 5921.440 2269.710 5921.770 ;
        RECT 2270.550 5921.440 2353.890 5921.770 ;
        RECT 2354.730 5921.440 2437.610 5921.770 ;
        RECT 2438.450 5921.440 2521.330 5921.770 ;
        RECT 2522.170 5921.440 2605.050 5921.770 ;
        RECT 2605.890 5921.440 2688.770 5921.770 ;
        RECT 2689.610 5921.440 2772.950 5921.770 ;
        RECT 2773.790 5921.440 2856.670 5921.770 ;
        RECT 2857.510 5921.440 2940.390 5921.770 ;
        RECT 2941.230 5921.440 3024.110 5921.770 ;
        RECT 3024.950 5921.440 3107.830 5921.770 ;
        RECT 3108.670 5921.440 3192.010 5921.770 ;
        RECT 3192.850 5921.440 3275.730 5921.770 ;
        RECT 3276.570 5921.440 3359.450 5921.770 ;
        RECT 3360.290 5921.440 3443.170 5921.770 ;
        RECT 3444.010 5921.440 3526.890 5921.770 ;
        RECT 3527.730 5921.440 3611.070 5921.770 ;
        RECT 3611.910 5921.440 3694.790 5921.770 ;
        RECT 3695.630 5921.440 3778.510 5921.770 ;
        RECT 3779.350 5921.440 3862.230 5921.770 ;
        RECT 3863.070 5921.440 3945.950 5921.770 ;
        RECT 3946.790 5921.440 4029.670 5921.770 ;
        RECT 4030.510 5921.440 4113.850 5921.770 ;
        RECT 4114.690 5921.440 4197.570 5921.770 ;
        RECT 4198.410 5921.440 4281.290 5921.770 ;
        RECT 4282.130 5921.440 4365.010 5921.770 ;
        RECT 4365.850 5921.440 4448.730 5921.770 ;
        RECT 4449.570 5921.440 4532.910 5921.770 ;
        RECT 4533.750 5921.440 4616.630 5921.770 ;
        RECT 4617.470 5921.440 4700.350 5921.770 ;
        RECT 4701.190 5921.440 4784.070 5921.770 ;
        RECT 4784.910 5921.440 4867.790 5921.770 ;
        RECT 4868.630 5921.440 4951.970 5921.770 ;
        RECT 4952.810 5921.440 5035.690 5921.770 ;
        RECT 5036.530 5921.440 5119.410 5921.770 ;
        RECT 5120.250 5921.440 5203.130 5921.770 ;
        RECT 5203.970 5921.440 5286.850 5921.770 ;
        RECT 5287.690 5921.440 5314.090 5921.770 ;
        RECT 63.370 46.800 5314.090 5921.440 ;
        RECT 63.370 46.520 76.430 46.800 ;
        RECT 77.270 46.520 130.710 46.800 ;
        RECT 131.550 46.520 184.990 46.800 ;
        RECT 185.830 46.520 239.270 46.800 ;
        RECT 240.110 46.520 294.010 46.800 ;
        RECT 294.850 46.520 348.290 46.800 ;
        RECT 349.130 46.520 402.570 46.800 ;
        RECT 403.410 46.520 457.310 46.800 ;
        RECT 458.150 46.520 511.590 46.800 ;
        RECT 512.430 46.520 565.870 46.800 ;
        RECT 566.710 46.520 620.610 46.800 ;
        RECT 621.450 46.520 674.890 46.800 ;
        RECT 675.730 46.520 729.170 46.800 ;
        RECT 730.010 46.520 783.910 46.800 ;
        RECT 784.750 46.520 838.190 46.800 ;
        RECT 839.030 46.520 892.470 46.800 ;
        RECT 893.310 46.520 947.210 46.800 ;
        RECT 948.050 46.520 1001.490 46.800 ;
        RECT 1002.330 46.520 1055.770 46.800 ;
        RECT 1056.610 46.520 1110.510 46.800 ;
        RECT 1111.350 46.520 1164.790 46.800 ;
        RECT 1165.630 46.520 1219.070 46.800 ;
        RECT 1219.910 46.520 1273.810 46.800 ;
        RECT 1274.650 46.520 1328.090 46.800 ;
        RECT 1328.930 46.520 1382.370 46.800 ;
        RECT 1383.210 46.520 1437.110 46.800 ;
        RECT 1437.950 46.520 1491.390 46.800 ;
        RECT 1492.230 46.520 1545.670 46.800 ;
        RECT 1546.510 46.520 1600.410 46.800 ;
        RECT 1601.250 46.520 1654.690 46.800 ;
        RECT 1655.530 46.520 1708.970 46.800 ;
        RECT 1709.810 46.520 1763.710 46.800 ;
        RECT 1764.550 46.520 1817.990 46.800 ;
        RECT 1818.830 46.520 1872.270 46.800 ;
        RECT 1873.110 46.520 1927.010 46.800 ;
        RECT 1927.850 46.520 1981.290 46.800 ;
        RECT 1982.130 46.520 2035.570 46.800 ;
        RECT 2036.410 46.520 2090.310 46.800 ;
        RECT 2091.150 46.520 2144.590 46.800 ;
        RECT 2145.430 46.520 2198.870 46.800 ;
        RECT 2199.710 46.520 2253.610 46.800 ;
        RECT 2254.450 46.520 2307.890 46.800 ;
        RECT 2308.730 46.520 2362.170 46.800 ;
        RECT 2363.010 46.520 2416.910 46.800 ;
        RECT 2417.750 46.520 2471.190 46.800 ;
        RECT 2472.030 46.520 2525.470 46.800 ;
        RECT 2526.310 46.520 2580.210 46.800 ;
        RECT 2581.050 46.520 2634.490 46.800 ;
        RECT 2635.330 46.520 2688.770 46.800 ;
        RECT 2689.610 46.520 2743.510 46.800 ;
        RECT 2744.350 46.520 2797.790 46.800 ;
        RECT 2798.630 46.520 2852.070 46.800 ;
        RECT 2852.910 46.520 2906.810 46.800 ;
        RECT 2907.650 46.520 2961.090 46.800 ;
        RECT 2961.930 46.520 3015.370 46.800 ;
        RECT 3016.210 46.520 3070.110 46.800 ;
        RECT 3070.950 46.520 3124.390 46.800 ;
        RECT 3125.230 46.520 3178.670 46.800 ;
        RECT 3179.510 46.520 3233.410 46.800 ;
        RECT 3234.250 46.520 3287.690 46.800 ;
        RECT 3288.530 46.520 3341.970 46.800 ;
        RECT 3342.810 46.520 3396.710 46.800 ;
        RECT 3397.550 46.520 3450.990 46.800 ;
        RECT 3451.830 46.520 3505.270 46.800 ;
        RECT 3506.110 46.520 3560.010 46.800 ;
        RECT 3560.850 46.520 3614.290 46.800 ;
        RECT 3615.130 46.520 3668.570 46.800 ;
        RECT 3669.410 46.520 3723.310 46.800 ;
        RECT 3724.150 46.520 3777.590 46.800 ;
        RECT 3778.430 46.520 3831.870 46.800 ;
        RECT 3832.710 46.520 3886.610 46.800 ;
        RECT 3887.450 46.520 3940.890 46.800 ;
        RECT 3941.730 46.520 3995.170 46.800 ;
        RECT 3996.010 46.520 4049.910 46.800 ;
        RECT 4050.750 46.520 4104.190 46.800 ;
        RECT 4105.030 46.520 4158.470 46.800 ;
        RECT 4159.310 46.520 4213.210 46.800 ;
        RECT 4214.050 46.520 4267.490 46.800 ;
        RECT 4268.330 46.520 4321.770 46.800 ;
        RECT 4322.610 46.520 4376.510 46.800 ;
        RECT 4377.350 46.520 4430.790 46.800 ;
        RECT 4431.630 46.520 4485.070 46.800 ;
        RECT 4485.910 46.520 4539.810 46.800 ;
        RECT 4540.650 46.520 4594.090 46.800 ;
        RECT 4594.930 46.520 4648.370 46.800 ;
        RECT 4649.210 46.520 4703.110 46.800 ;
        RECT 4703.950 46.520 4757.390 46.800 ;
        RECT 4758.230 46.520 4811.670 46.800 ;
        RECT 4812.510 46.520 4866.410 46.800 ;
        RECT 4867.250 46.520 4920.690 46.800 ;
        RECT 4921.530 46.520 4974.970 46.800 ;
        RECT 4975.810 46.520 5029.710 46.800 ;
        RECT 5030.550 46.520 5083.990 46.800 ;
        RECT 5084.830 46.520 5138.270 46.800 ;
        RECT 5139.110 46.520 5193.010 46.800 ;
        RECT 5193.850 46.520 5247.290 46.800 ;
        RECT 5248.130 46.520 5301.570 46.800 ;
        RECT 5302.410 46.520 5314.090 46.800 ;
      LAYER met3 ;
        RECT 51.880 5891.800 5327.210 5908.945 ;
        RECT 52.280 5890.400 5327.210 5891.800 ;
        RECT 51.880 5888.400 5327.210 5890.400 ;
        RECT 51.880 5887.000 5326.680 5888.400 ;
        RECT 51.880 5826.520 5327.210 5887.000 ;
        RECT 52.280 5825.120 5327.210 5826.520 ;
        RECT 51.880 5815.640 5327.210 5825.120 ;
        RECT 51.880 5814.240 5326.680 5815.640 ;
        RECT 51.880 5761.240 5327.210 5814.240 ;
        RECT 52.280 5759.840 5327.210 5761.240 ;
        RECT 51.880 5742.880 5327.210 5759.840 ;
        RECT 51.880 5741.480 5326.680 5742.880 ;
        RECT 51.880 5695.960 5327.210 5741.480 ;
        RECT 52.280 5694.560 5327.210 5695.960 ;
        RECT 51.880 5670.120 5327.210 5694.560 ;
        RECT 51.880 5668.720 5326.680 5670.120 ;
        RECT 51.880 5630.680 5327.210 5668.720 ;
        RECT 52.280 5629.280 5327.210 5630.680 ;
        RECT 51.880 5598.040 5327.210 5629.280 ;
        RECT 51.880 5596.640 5326.680 5598.040 ;
        RECT 51.880 5565.400 5327.210 5596.640 ;
        RECT 52.280 5564.000 5327.210 5565.400 ;
        RECT 51.880 5525.280 5327.210 5564.000 ;
        RECT 51.880 5523.880 5326.680 5525.280 ;
        RECT 51.880 5500.120 5327.210 5523.880 ;
        RECT 52.280 5498.720 5327.210 5500.120 ;
        RECT 51.880 5452.520 5327.210 5498.720 ;
        RECT 51.880 5451.120 5326.680 5452.520 ;
        RECT 51.880 5434.840 5327.210 5451.120 ;
        RECT 52.280 5433.440 5327.210 5434.840 ;
        RECT 51.880 5379.760 5327.210 5433.440 ;
        RECT 51.880 5378.360 5326.680 5379.760 ;
        RECT 51.880 5369.560 5327.210 5378.360 ;
        RECT 52.280 5368.160 5327.210 5369.560 ;
        RECT 51.880 5307.680 5327.210 5368.160 ;
        RECT 51.880 5306.280 5326.680 5307.680 ;
        RECT 51.880 5304.280 5327.210 5306.280 ;
        RECT 52.280 5302.880 5327.210 5304.280 ;
        RECT 51.880 5239.000 5327.210 5302.880 ;
        RECT 52.280 5237.600 5327.210 5239.000 ;
        RECT 51.880 5234.920 5327.210 5237.600 ;
        RECT 51.880 5233.520 5326.680 5234.920 ;
        RECT 51.880 5173.720 5327.210 5233.520 ;
        RECT 52.280 5172.320 5327.210 5173.720 ;
        RECT 51.880 5162.160 5327.210 5172.320 ;
        RECT 51.880 5160.760 5326.680 5162.160 ;
        RECT 51.880 5107.760 5327.210 5160.760 ;
        RECT 52.280 5106.360 5327.210 5107.760 ;
        RECT 51.880 5089.400 5327.210 5106.360 ;
        RECT 51.880 5088.000 5326.680 5089.400 ;
        RECT 51.880 5042.480 5327.210 5088.000 ;
        RECT 52.280 5041.080 5327.210 5042.480 ;
        RECT 51.880 5017.320 5327.210 5041.080 ;
        RECT 51.880 5015.920 5326.680 5017.320 ;
        RECT 51.880 4977.200 5327.210 5015.920 ;
        RECT 52.280 4975.800 5327.210 4977.200 ;
        RECT 51.880 4944.560 5327.210 4975.800 ;
        RECT 51.880 4943.160 5326.680 4944.560 ;
        RECT 51.880 4911.920 5327.210 4943.160 ;
        RECT 52.280 4910.520 5327.210 4911.920 ;
        RECT 51.880 4871.800 5327.210 4910.520 ;
        RECT 51.880 4870.400 5326.680 4871.800 ;
        RECT 51.880 4846.640 5327.210 4870.400 ;
        RECT 52.280 4845.240 5327.210 4846.640 ;
        RECT 51.880 4799.040 5327.210 4845.240 ;
        RECT 51.880 4797.640 5326.680 4799.040 ;
        RECT 51.880 4781.360 5327.210 4797.640 ;
        RECT 52.280 4779.960 5327.210 4781.360 ;
        RECT 51.880 4726.960 5327.210 4779.960 ;
        RECT 51.880 4725.560 5326.680 4726.960 ;
        RECT 51.880 4716.080 5327.210 4725.560 ;
        RECT 52.280 4714.680 5327.210 4716.080 ;
        RECT 51.880 4654.200 5327.210 4714.680 ;
        RECT 51.880 4652.800 5326.680 4654.200 ;
        RECT 51.880 4650.800 5327.210 4652.800 ;
        RECT 52.280 4649.400 5327.210 4650.800 ;
        RECT 51.880 4585.520 5327.210 4649.400 ;
        RECT 52.280 4584.120 5327.210 4585.520 ;
        RECT 51.880 4581.440 5327.210 4584.120 ;
        RECT 51.880 4580.040 5326.680 4581.440 ;
        RECT 51.880 4520.240 5327.210 4580.040 ;
        RECT 52.280 4518.840 5327.210 4520.240 ;
        RECT 51.880 4508.680 5327.210 4518.840 ;
        RECT 51.880 4507.280 5326.680 4508.680 ;
        RECT 51.880 4454.960 5327.210 4507.280 ;
        RECT 52.280 4453.560 5327.210 4454.960 ;
        RECT 51.880 4436.600 5327.210 4453.560 ;
        RECT 51.880 4435.200 5326.680 4436.600 ;
        RECT 51.880 4389.680 5327.210 4435.200 ;
        RECT 52.280 4388.280 5327.210 4389.680 ;
        RECT 51.880 4363.840 5327.210 4388.280 ;
        RECT 51.880 4362.440 5326.680 4363.840 ;
        RECT 51.880 4324.400 5327.210 4362.440 ;
        RECT 52.280 4323.000 5327.210 4324.400 ;
        RECT 51.880 4291.080 5327.210 4323.000 ;
        RECT 51.880 4289.680 5326.680 4291.080 ;
        RECT 51.880 4258.440 5327.210 4289.680 ;
        RECT 52.280 4257.040 5327.210 4258.440 ;
        RECT 51.880 4218.320 5327.210 4257.040 ;
        RECT 51.880 4216.920 5326.680 4218.320 ;
        RECT 51.880 4193.160 5327.210 4216.920 ;
        RECT 52.280 4191.760 5327.210 4193.160 ;
        RECT 51.880 4146.240 5327.210 4191.760 ;
        RECT 51.880 4144.840 5326.680 4146.240 ;
        RECT 51.880 4127.880 5327.210 4144.840 ;
        RECT 52.280 4126.480 5327.210 4127.880 ;
        RECT 51.880 4073.480 5327.210 4126.480 ;
        RECT 51.880 4072.080 5326.680 4073.480 ;
        RECT 51.880 4062.600 5327.210 4072.080 ;
        RECT 52.280 4061.200 5327.210 4062.600 ;
        RECT 51.880 4000.720 5327.210 4061.200 ;
        RECT 51.880 3999.320 5326.680 4000.720 ;
        RECT 51.880 3997.320 5327.210 3999.320 ;
        RECT 52.280 3995.920 5327.210 3997.320 ;
        RECT 51.880 3932.040 5327.210 3995.920 ;
        RECT 52.280 3930.640 5327.210 3932.040 ;
        RECT 51.880 3927.960 5327.210 3930.640 ;
        RECT 51.880 3926.560 5326.680 3927.960 ;
        RECT 51.880 3866.760 5327.210 3926.560 ;
        RECT 52.280 3865.360 5327.210 3866.760 ;
        RECT 51.880 3855.880 5327.210 3865.360 ;
        RECT 51.880 3854.480 5326.680 3855.880 ;
        RECT 51.880 3801.480 5327.210 3854.480 ;
        RECT 52.280 3800.080 5327.210 3801.480 ;
        RECT 51.880 3783.120 5327.210 3800.080 ;
        RECT 51.880 3781.720 5326.680 3783.120 ;
        RECT 51.880 3736.200 5327.210 3781.720 ;
        RECT 52.280 3734.800 5327.210 3736.200 ;
        RECT 51.880 3710.360 5327.210 3734.800 ;
        RECT 51.880 3708.960 5326.680 3710.360 ;
        RECT 51.880 3670.920 5327.210 3708.960 ;
        RECT 52.280 3669.520 5327.210 3670.920 ;
        RECT 51.880 3637.600 5327.210 3669.520 ;
        RECT 51.880 3636.200 5326.680 3637.600 ;
        RECT 51.880 3605.640 5327.210 3636.200 ;
        RECT 52.280 3604.240 5327.210 3605.640 ;
        RECT 51.880 3565.520 5327.210 3604.240 ;
        RECT 51.880 3564.120 5326.680 3565.520 ;
        RECT 51.880 3540.360 5327.210 3564.120 ;
        RECT 52.280 3538.960 5327.210 3540.360 ;
        RECT 51.880 3492.760 5327.210 3538.960 ;
        RECT 51.880 3491.360 5326.680 3492.760 ;
        RECT 51.880 3475.080 5327.210 3491.360 ;
        RECT 52.280 3473.680 5327.210 3475.080 ;
        RECT 51.880 3420.000 5327.210 3473.680 ;
        RECT 51.880 3418.600 5326.680 3420.000 ;
        RECT 51.880 3409.120 5327.210 3418.600 ;
        RECT 52.280 3407.720 5327.210 3409.120 ;
        RECT 51.880 3347.240 5327.210 3407.720 ;
        RECT 51.880 3345.840 5326.680 3347.240 ;
        RECT 51.880 3343.840 5327.210 3345.840 ;
        RECT 52.280 3342.440 5327.210 3343.840 ;
        RECT 51.880 3278.560 5327.210 3342.440 ;
        RECT 52.280 3277.160 5327.210 3278.560 ;
        RECT 51.880 3275.160 5327.210 3277.160 ;
        RECT 51.880 3273.760 5326.680 3275.160 ;
        RECT 51.880 3213.280 5327.210 3273.760 ;
        RECT 52.280 3211.880 5327.210 3213.280 ;
        RECT 51.880 3202.400 5327.210 3211.880 ;
        RECT 51.880 3201.000 5326.680 3202.400 ;
        RECT 51.880 3148.000 5327.210 3201.000 ;
        RECT 52.280 3146.600 5327.210 3148.000 ;
        RECT 51.880 3129.640 5327.210 3146.600 ;
        RECT 51.880 3128.240 5326.680 3129.640 ;
        RECT 51.880 3082.720 5327.210 3128.240 ;
        RECT 52.280 3081.320 5327.210 3082.720 ;
        RECT 51.880 3056.880 5327.210 3081.320 ;
        RECT 51.880 3055.480 5326.680 3056.880 ;
        RECT 51.880 3017.440 5327.210 3055.480 ;
        RECT 52.280 3016.040 5327.210 3017.440 ;
        RECT 51.880 2984.800 5327.210 3016.040 ;
        RECT 51.880 2983.400 5326.680 2984.800 ;
        RECT 51.880 2952.160 5327.210 2983.400 ;
        RECT 52.280 2950.760 5327.210 2952.160 ;
        RECT 51.880 2912.040 5327.210 2950.760 ;
        RECT 51.880 2910.640 5326.680 2912.040 ;
        RECT 51.880 2886.880 5327.210 2910.640 ;
        RECT 52.280 2885.480 5327.210 2886.880 ;
        RECT 51.880 2839.280 5327.210 2885.480 ;
        RECT 51.880 2837.880 5326.680 2839.280 ;
        RECT 51.880 2821.600 5327.210 2837.880 ;
        RECT 52.280 2820.200 5327.210 2821.600 ;
        RECT 51.880 2766.520 5327.210 2820.200 ;
        RECT 51.880 2765.120 5326.680 2766.520 ;
        RECT 51.880 2756.320 5327.210 2765.120 ;
        RECT 52.280 2754.920 5327.210 2756.320 ;
        RECT 51.880 2694.440 5327.210 2754.920 ;
        RECT 51.880 2693.040 5326.680 2694.440 ;
        RECT 51.880 2691.040 5327.210 2693.040 ;
        RECT 52.280 2689.640 5327.210 2691.040 ;
        RECT 51.880 2625.760 5327.210 2689.640 ;
        RECT 52.280 2624.360 5327.210 2625.760 ;
        RECT 51.880 2621.680 5327.210 2624.360 ;
        RECT 51.880 2620.280 5326.680 2621.680 ;
        RECT 51.880 2559.800 5327.210 2620.280 ;
        RECT 52.280 2558.400 5327.210 2559.800 ;
        RECT 51.880 2548.920 5327.210 2558.400 ;
        RECT 51.880 2547.520 5326.680 2548.920 ;
        RECT 51.880 2494.520 5327.210 2547.520 ;
        RECT 52.280 2493.120 5327.210 2494.520 ;
        RECT 51.880 2476.160 5327.210 2493.120 ;
        RECT 51.880 2474.760 5326.680 2476.160 ;
        RECT 51.880 2429.240 5327.210 2474.760 ;
        RECT 52.280 2427.840 5327.210 2429.240 ;
        RECT 51.880 2404.080 5327.210 2427.840 ;
        RECT 51.880 2402.680 5326.680 2404.080 ;
        RECT 51.880 2363.960 5327.210 2402.680 ;
        RECT 52.280 2362.560 5327.210 2363.960 ;
        RECT 51.880 2331.320 5327.210 2362.560 ;
        RECT 51.880 2329.920 5326.680 2331.320 ;
        RECT 51.880 2298.680 5327.210 2329.920 ;
        RECT 52.280 2297.280 5327.210 2298.680 ;
        RECT 51.880 2258.560 5327.210 2297.280 ;
        RECT 51.880 2257.160 5326.680 2258.560 ;
        RECT 51.880 2233.400 5327.210 2257.160 ;
        RECT 52.280 2232.000 5327.210 2233.400 ;
        RECT 51.880 2185.800 5327.210 2232.000 ;
        RECT 51.880 2184.400 5326.680 2185.800 ;
        RECT 51.880 2168.120 5327.210 2184.400 ;
        RECT 52.280 2166.720 5327.210 2168.120 ;
        RECT 51.880 2113.720 5327.210 2166.720 ;
        RECT 51.880 2112.320 5326.680 2113.720 ;
        RECT 51.880 2102.840 5327.210 2112.320 ;
        RECT 52.280 2101.440 5327.210 2102.840 ;
        RECT 51.880 2040.960 5327.210 2101.440 ;
        RECT 51.880 2039.560 5326.680 2040.960 ;
        RECT 51.880 2037.560 5327.210 2039.560 ;
        RECT 52.280 2036.160 5327.210 2037.560 ;
        RECT 51.880 1972.280 5327.210 2036.160 ;
        RECT 52.280 1970.880 5327.210 1972.280 ;
        RECT 51.880 1968.200 5327.210 1970.880 ;
        RECT 51.880 1966.800 5326.680 1968.200 ;
        RECT 51.880 1907.000 5327.210 1966.800 ;
        RECT 52.280 1905.600 5327.210 1907.000 ;
        RECT 51.880 1895.440 5327.210 1905.600 ;
        RECT 51.880 1894.040 5326.680 1895.440 ;
        RECT 51.880 1841.720 5327.210 1894.040 ;
        RECT 52.280 1840.320 5327.210 1841.720 ;
        RECT 51.880 1823.360 5327.210 1840.320 ;
        RECT 51.880 1821.960 5326.680 1823.360 ;
        RECT 51.880 1776.440 5327.210 1821.960 ;
        RECT 52.280 1775.040 5327.210 1776.440 ;
        RECT 51.880 1750.600 5327.210 1775.040 ;
        RECT 51.880 1749.200 5326.680 1750.600 ;
        RECT 51.880 1710.480 5327.210 1749.200 ;
        RECT 52.280 1709.080 5327.210 1710.480 ;
        RECT 51.880 1677.840 5327.210 1709.080 ;
        RECT 51.880 1676.440 5326.680 1677.840 ;
        RECT 51.880 1645.200 5327.210 1676.440 ;
        RECT 52.280 1643.800 5327.210 1645.200 ;
        RECT 51.880 1605.080 5327.210 1643.800 ;
        RECT 51.880 1603.680 5326.680 1605.080 ;
        RECT 51.880 1579.920 5327.210 1603.680 ;
        RECT 52.280 1578.520 5327.210 1579.920 ;
        RECT 51.880 1533.000 5327.210 1578.520 ;
        RECT 51.880 1531.600 5326.680 1533.000 ;
        RECT 51.880 1514.640 5327.210 1531.600 ;
        RECT 52.280 1513.240 5327.210 1514.640 ;
        RECT 51.880 1460.240 5327.210 1513.240 ;
        RECT 51.880 1458.840 5326.680 1460.240 ;
        RECT 51.880 1449.360 5327.210 1458.840 ;
        RECT 52.280 1447.960 5327.210 1449.360 ;
        RECT 51.880 1387.480 5327.210 1447.960 ;
        RECT 51.880 1386.080 5326.680 1387.480 ;
        RECT 51.880 1384.080 5327.210 1386.080 ;
        RECT 52.280 1382.680 5327.210 1384.080 ;
        RECT 51.880 1318.800 5327.210 1382.680 ;
        RECT 52.280 1317.400 5327.210 1318.800 ;
        RECT 51.880 1314.720 5327.210 1317.400 ;
        RECT 51.880 1313.320 5326.680 1314.720 ;
        RECT 51.880 1253.520 5327.210 1313.320 ;
        RECT 52.280 1252.120 5327.210 1253.520 ;
        RECT 51.880 1242.640 5327.210 1252.120 ;
        RECT 51.880 1241.240 5326.680 1242.640 ;
        RECT 51.880 1188.240 5327.210 1241.240 ;
        RECT 52.280 1186.840 5327.210 1188.240 ;
        RECT 51.880 1169.880 5327.210 1186.840 ;
        RECT 51.880 1168.480 5326.680 1169.880 ;
        RECT 51.880 1122.960 5327.210 1168.480 ;
        RECT 52.280 1121.560 5327.210 1122.960 ;
        RECT 51.880 1097.120 5327.210 1121.560 ;
        RECT 51.880 1095.720 5326.680 1097.120 ;
        RECT 51.880 1057.680 5327.210 1095.720 ;
        RECT 52.280 1056.280 5327.210 1057.680 ;
        RECT 51.880 1024.360 5327.210 1056.280 ;
        RECT 51.880 1022.960 5326.680 1024.360 ;
        RECT 51.880 992.400 5327.210 1022.960 ;
        RECT 52.280 991.000 5327.210 992.400 ;
        RECT 51.880 952.280 5327.210 991.000 ;
        RECT 51.880 950.880 5326.680 952.280 ;
        RECT 51.880 927.120 5327.210 950.880 ;
        RECT 52.280 925.720 5327.210 927.120 ;
        RECT 51.880 879.520 5327.210 925.720 ;
        RECT 51.880 878.120 5326.680 879.520 ;
        RECT 51.880 861.160 5327.210 878.120 ;
        RECT 52.280 859.760 5327.210 861.160 ;
        RECT 51.880 806.760 5327.210 859.760 ;
        RECT 51.880 805.360 5326.680 806.760 ;
        RECT 51.880 795.880 5327.210 805.360 ;
        RECT 52.280 794.480 5327.210 795.880 ;
        RECT 51.880 734.000 5327.210 794.480 ;
        RECT 51.880 732.600 5326.680 734.000 ;
        RECT 51.880 730.600 5327.210 732.600 ;
        RECT 52.280 729.200 5327.210 730.600 ;
        RECT 51.880 665.320 5327.210 729.200 ;
        RECT 52.280 663.920 5327.210 665.320 ;
        RECT 51.880 661.920 5327.210 663.920 ;
        RECT 51.880 660.520 5326.680 661.920 ;
        RECT 51.880 600.040 5327.210 660.520 ;
        RECT 52.280 598.640 5327.210 600.040 ;
        RECT 51.880 589.160 5327.210 598.640 ;
        RECT 51.880 587.760 5326.680 589.160 ;
        RECT 51.880 534.760 5327.210 587.760 ;
        RECT 52.280 533.360 5327.210 534.760 ;
        RECT 51.880 516.400 5327.210 533.360 ;
        RECT 51.880 515.000 5326.680 516.400 ;
        RECT 51.880 469.480 5327.210 515.000 ;
        RECT 52.280 468.080 5327.210 469.480 ;
        RECT 51.880 443.640 5327.210 468.080 ;
        RECT 51.880 442.240 5326.680 443.640 ;
        RECT 51.880 404.200 5327.210 442.240 ;
        RECT 52.280 402.800 5327.210 404.200 ;
        RECT 51.880 371.560 5327.210 402.800 ;
        RECT 51.880 370.160 5326.680 371.560 ;
        RECT 51.880 338.920 5327.210 370.160 ;
        RECT 52.280 337.520 5327.210 338.920 ;
        RECT 51.880 298.800 5327.210 337.520 ;
        RECT 51.880 297.400 5326.680 298.800 ;
        RECT 51.880 273.640 5327.210 297.400 ;
        RECT 52.280 272.240 5327.210 273.640 ;
        RECT 51.880 226.040 5327.210 272.240 ;
        RECT 51.880 224.640 5326.680 226.040 ;
        RECT 51.880 208.360 5327.210 224.640 ;
        RECT 52.280 206.960 5327.210 208.360 ;
        RECT 51.880 153.280 5327.210 206.960 ;
        RECT 51.880 151.880 5326.680 153.280 ;
        RECT 51.880 143.080 5327.210 151.880 ;
        RECT 52.280 141.680 5327.210 143.080 ;
        RECT 51.880 81.200 5327.210 141.680 ;
        RECT 51.880 79.800 5326.680 81.200 ;
        RECT 51.880 77.800 5327.210 79.800 ;
        RECT 52.280 76.400 5327.210 77.800 ;
        RECT 51.880 59.935 5327.210 76.400 ;
      LAYER met4 ;
        RECT 0.000 0.000 5378.840 5966.160 ;
      LAYER met5 ;
        RECT 0.000 79.200 5378.840 5966.160 ;
  END
END fpga_core
END LIBRARY

