* NGSPICE file created from sb_1__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt sb_1__1_ Test_en_N_out Test_en_S_in bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] clk_1_E_out clk_1_N_in clk_1_S_in clk_1_W_out clk_2_E_in clk_2_E_out
+ clk_2_N_in clk_2_N_out clk_2_S_in clk_2_S_out clk_2_W_in clk_2_W_out clk_3_E_in
+ clk_3_E_out clk_3_N_in clk_3_N_out clk_3_S_in clk_3_S_out clk_3_W_in clk_3_W_out
+ left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_ left_bottom_grid_pin_37_
+ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_ left_bottom_grid_pin_41_
+ prog_clk_0_N_in prog_clk_1_E_out prog_clk_1_N_in prog_clk_1_S_in prog_clk_1_W_out
+ prog_clk_2_E_in prog_clk_2_E_out prog_clk_2_N_in prog_clk_2_N_out prog_clk_2_S_in
+ prog_clk_2_S_out prog_clk_2_W_in prog_clk_2_W_out prog_clk_3_E_in prog_clk_3_E_out
+ prog_clk_3_N_in prog_clk_3_N_out prog_clk_3_S_in prog_clk_3_S_out prog_clk_3_W_in
+ prog_clk_3_W_out right_bottom_grid_pin_34_ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_
+ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_
+ right_bottom_grid_pin_41_ top_left_grid_pin_42_ top_left_grid_pin_43_ top_left_grid_pin_44_
+ top_left_grid_pin_45_ top_left_grid_pin_46_ top_left_grid_pin_47_ top_left_grid_pin_48_
+ top_left_grid_pin_49_ VPWR VGND
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[4] mux_bottom_track_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_131_ _131_/A VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
X_062_ chanx_right_in[12] VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_045_ VGND VGND VPWR VPWR _045_/HI _045_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_114_ _114_/A VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_028_ VGND VGND VPWR VPWR _028_/HI _028_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_5 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _114_/A sky130_fd_sc_hd__buf_4
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_130_ chany_bottom_in[4] VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_2_W_FTB01 prog_clk_2_E_in VGND VGND VPWR VPWR prog_clk_2_W_out sky130_fd_sc_hd__buf_4
X_061_ chanx_right_in[13] VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _071_/A sky130_fd_sc_hd__buf_4
X_113_ _113_/A VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
X_044_ VGND VGND VPWR VPWR _044_/HI _044_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_6 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_3_ _036_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_3_ _037_/HI chanx_left_in[12] mux_top_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _063_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_mem_bottom_track_1.prog_clk clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l1_in_4_ chanx_left_in[0] chany_bottom_in[12] mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_060_ chanx_right_in[14] VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_043_ VGND VGND VPWR VPWR _043_/HI _043_/LO sky130_fd_sc_hd__conb_1
X_112_ chany_top_in[2] VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclk_2_E_FTB01 clk_2_E_in VGND VGND VPWR VPWR clk_2_E_out sky130_fd_sc_hd__buf_4
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_7 chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[16] mux_right_track_8.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[2] mux_top_track_0.mux_l1_in_4_/X mux_top_track_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_0.mux_l1_in_3_ chany_bottom_in[2] chanx_right_in[12] mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_042_ VGND VGND VPWR VPWR _042_/HI _042_/LO sky130_fd_sc_hd__conb_1
X_111_ _111_/A VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xprog_clk_3_N_FTB01 prog_clk_3_E_in VGND VGND VPWR VPWR prog_clk_3_N_out sky130_fd_sc_hd__buf_4
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ mux_top_track_0.mux_l1_in_3_/X mux_top_track_0.mux_l1_in_2_/X
+ mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ chany_bottom_in[6] mux_right_track_8.mux_l1_in_2_/X
+ mux_right_track_8.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l1_in_2_ chany_bottom_in[3] right_bottom_grid_pin_38_ mux_right_track_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_2_ chanx_right_in[2] chanx_right_in[1] mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _127_/A sky130_fd_sc_hd__buf_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_3_ _046_/HI chanx_left_in[19] mux_bottom_track_25.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_041_ VGND VGND VPWR VPWR _041_/HI _041_/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_110_ chany_top_in[4] VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xmux_right_track_4.mux_l2_in_7_ _035_/HI chanx_left_in[14] mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_9 chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_3_ _050_/HI chanx_left_in[16] mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _135_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l4_in_0_ mux_bottom_track_25.mux_l3_in_1_/X mux_bottom_track_25.mux_l3_in_0_/X
+ mux_bottom_track_25.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ mux_right_track_8.mux_l1_in_1_/X mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l3_in_1_ mux_bottom_track_25.mux_l2_in_3_/X mux_bottom_track_25.mux_l2_in_2_/X
+ mux_bottom_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l1_in_1_ right_bottom_grid_pin_34_ chany_top_in[16] mux_right_track_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l4_in_0_ mux_bottom_track_9.mux_l3_in_1_/X mux_bottom_track_9.mux_l3_in_0_/X
+ mux_bottom_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_2_ chanx_left_in[18] chanx_left_in[9] mux_bottom_track_25.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l3_in_1_ mux_bottom_track_9.mux_l2_in_3_/X mux_bottom_track_9.mux_l2_in_2_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_040_ VGND VGND VPWR VPWR _040_/HI _040_/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_6_ chanx_left_in[5] chany_bottom_in[14] mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_6_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[6] mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__buf_4
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[6] chany_top_in[3] mux_right_track_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_0.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclk_3_W_FTB01 clk_3_E_in VGND VGND VPWR VPWR clk_3_W_out sky130_fd_sc_hd__buf_4
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _091_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_25.mux_l2_in_1_ bottom_left_grid_pin_48_ mux_bottom_track_25.mux_l1_in_2_/X
+ mux_bottom_track_25.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_2_S_FTB01 prog_clk_2_E_in VGND VGND VPWR VPWR prog_clk_2_S_out sky130_fd_sc_hd__buf_4
Xmux_right_track_4.mux_l2_in_5_ chany_bottom_in[7] chany_bottom_in[5] mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_5_/X sky130_fd_sc_hd__mux2_1
X_099_ _099_/A VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xmux_top_track_16.mux_l2_in_3_ _038_/HI chanx_left_in[17] mux_top_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l5_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_3_0_mem_bottom_track_1.prog_clk clkbuf_3_2_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l1_in_2_ bottom_left_grid_pin_44_ chanx_right_in[18] mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l2_in_1_ bottom_left_grid_pin_46_ mux_bottom_track_9.mux_l1_in_2_/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__buf_4
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l1_in_2_ bottom_left_grid_pin_42_ chanx_right_in[16] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l4_in_0_ mux_top_track_16.mux_l3_in_1_/X mux_top_track_16.mux_l3_in_0_/X
+ mux_top_track_16.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_3_ _054_/HI left_bottom_grid_pin_41_ mux_left_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_4.mux_l3_in_3_ mux_right_track_4.mux_l2_in_7_/X mux_right_track_4.mux_l2_in_6_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l3_in_1_ mux_top_track_16.mux_l2_in_3_/X mux_top_track_16.mux_l2_in_2_/X
+ mux_top_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_7_ _049_/HI chanx_left_in[14] mux_bottom_track_5.mux_l2_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l1_in_4_ left_bottom_grid_pin_37_ left_bottom_grid_pin_35_ mux_left_track_3.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_4.mux_l2_in_4_ right_bottom_grid_pin_41_ right_bottom_grid_pin_40_
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_4_/X
+ sky130_fd_sc_hd__mux2_1
X_098_ chany_top_in[16] VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xmux_top_track_16.mux_l2_in_2_ chanx_left_in[8] chanx_left_in[7] mux_top_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l5_in_0_ mux_right_track_4.mux_l4_in_1_/X mux_right_track_4.mux_l4_in_0_/X
+ mux_right_track_4.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l1_in_1_ chanx_right_in[9] chanx_right_in[0] mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l4_in_1_ mux_right_track_4.mux_l3_in_3_/X mux_right_track_4.mux_l3_in_2_/X
+ mux_right_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l5_in_0_/X VGND VGND
+ VPWR VPWR _073_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_9.mux_l1_in_1_ chanx_right_in[6] chanx_right_in[3] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_2_ left_bottom_grid_pin_39_ mux_left_track_3.mux_l1_in_4_/X
+ mux_left_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l3_in_2_ mux_right_track_4.mux_l2_in_5_/X mux_right_track_4.mux_l2_in_4_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_6_ chanx_left_in[7] chanx_left_in[5] mux_bottom_track_5.mux_l2_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_6_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l1_in_3_ chany_bottom_in[13] chany_bottom_in[4] mux_left_track_3.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l5_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_4.mux_l2_in_3_ right_bottom_grid_pin_39_ right_bottom_grid_pin_38_
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_16.mux_l2_in_3_ _031_/HI chanx_left_in[17] mux_right_track_16.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l2_in_1_ chany_bottom_in[17] mux_top_track_16.mux_l1_in_2_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ chany_top_in[17] VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_149_ prog_clk_3_E_in VGND VGND VPWR VPWR prog_clk_3_W_in sky130_fd_sc_hd__buf_2
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_ chany_bottom_in[8] chanx_right_in[17] mux_top_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.mux_l4_in_0_ mux_right_track_16.mux_l3_in_1_/X mux_right_track_16.mux_l3_in_0_/X
+ mux_right_track_16.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _111_/A sky130_fd_sc_hd__buf_4
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l3_in_1_ mux_right_track_16.mux_l2_in_3_/X mux_right_track_16.mux_l2_in_2_/X
+ mux_right_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ mux_left_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l4_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_5_ bottom_left_grid_pin_49_ bottom_left_grid_pin_48_
+ mux_bottom_track_5.mux_l2_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_5_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_2_ chanx_left_in[8] chany_bottom_in[17] mux_right_track_16.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l1_in_2_ chany_bottom_in[0] chanx_right_in[13] mux_left_track_3.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_2_ right_bottom_grid_pin_37_ right_bottom_grid_pin_36_
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_096_ chany_top_in[18] VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_148_ prog_clk_3_E_in VGND VGND VPWR VPWR prog_clk_3_S_in sky130_fd_sc_hd__buf_2
X_079_ _079_/A VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l1_in_1_ chanx_right_in[15] chanx_right_in[8] mux_top_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l3_in_3_ mux_bottom_track_5.mux_l2_in_7_/X mux_bottom_track_5.mux_l2_in_6_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_4_ bottom_left_grid_pin_47_ bottom_left_grid_pin_46_
+ mux_bottom_track_5.mux_l2_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_4_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_1_ chany_bottom_in[8] mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l1_in_1_ chanx_right_in[4] chany_top_in[19] mux_left_track_3.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xprog_clk_1_W_FTB01 prog_clk_1_N_in VGND VGND VPWR VPWR prog_clk_1_W_out sky130_fd_sc_hd__buf_4
Xmux_right_track_4.mux_l2_in_1_ right_bottom_grid_pin_35_ right_bottom_grid_pin_34_
+ mux_right_track_4.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_095_ _095_/A VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_5.mux_l5_in_0_ mux_bottom_track_5.mux_l4_in_1_/X mux_bottom_track_5.mux_l4_in_0_/X
+ mux_bottom_track_5.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_078_ chanx_left_in[16] VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_2_ chany_bottom_in[1] right_bottom_grid_pin_39_ mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_147_ prog_clk_3_E_in VGND VGND VPWR VPWR prog_clk_3_N_in sky130_fd_sc_hd__buf_2
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l4_in_1_ mux_bottom_track_5.mux_l3_in_3_/X mux_bottom_track_5.mux_l3_in_2_/X
+ mux_bottom_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l1_in_0_ top_left_grid_pin_47_ top_left_grid_pin_43_ mux_top_track_16.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l3_in_2_ mux_bottom_track_5.mux_l2_in_5_/X mux_bottom_track_5.mux_l2_in_4_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_mem_bottom_track_1.prog_clk clkbuf_3_2_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_4.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_3_ bottom_left_grid_pin_45_ bottom_left_grid_pin_44_
+ mux_bottom_track_5.mux_l2_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xclk_3_S_FTB01 clk_3_E_in VGND VGND VPWR VPWR clk_3_S_out sky130_fd_sc_hd__buf_4
Xmux_left_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_left_track_3.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ chany_top_in[14] ANTENNA_18/DIODE mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_4.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_094_ _094_/A VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_1_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_077_ chanx_left_in[17] VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
X_146_ prog_clk_2_E_in VGND VGND VPWR VPWR prog_clk_2_W_in sky130_fd_sc_hd__buf_2
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclk_1_E_FTB01 clk_1_N_in VGND VGND VPWR VPWR clk_1_E_out sky130_fd_sc_hd__buf_4
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_1_ right_bottom_grid_pin_35_ chany_top_in[17] mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l4_in_0_ mux_bottom_track_5.mux_l3_in_1_/X mux_bottom_track_5.mux_l3_in_0_/X
+ mux_bottom_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_129_ chany_bottom_in[5] VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l3_in_1_ mux_bottom_track_5.mux_l2_in_3_/X mux_bottom_track_5.mux_l2_in_2_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_2_ bottom_left_grid_pin_43_ bottom_left_grid_pin_42_
+ mux_bottom_track_5.mux_l2_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l5_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_4.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_093_ _093_/A VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_076_ chanx_left_in[18] VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_145_ prog_clk_2_E_in VGND VGND VPWR VPWR prog_clk_2_S_in sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_right_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[5] chany_top_in[1] mux_right_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR ANTENNA_18/DIODE sky130_fd_sc_hd__mux2_1
Xprog_clk_2_N_FTB01 prog_clk_2_E_in VGND VGND VPWR VPWR prog_clk_2_N_out sky130_fd_sc_hd__buf_4
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l5_in_0_/X VGND
+ VGND VPWR VPWR _093_/A sky130_fd_sc_hd__buf_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ chany_bottom_in[6] VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
X_059_ _059_/A VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_1_ chanx_right_in[14] chanx_right_in[7] mux_bottom_track_5.mux_l2_in_6_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l3_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ chanx_left_in[2] VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
X_144_ prog_clk_2_E_in VGND VGND VPWR VPWR prog_clk_2_N_in sky130_fd_sc_hd__buf_2
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_075_ _075_/A VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_33.mux_l1_in_3_ _048_/HI chanx_left_in[10] mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__buf_4
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_127_ _127_/A VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
X_058_ chanx_right_in[16] VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l3_in_0_ mux_bottom_track_33.mux_l2_in_1_/X mux_bottom_track_33.mux_l2_in_0_/X
+ mux_bottom_track_33.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l2_in_1_ mux_bottom_track_33.mux_l1_in_3_/X mux_bottom_track_33.mux_l1_in_2_/X
+ mux_bottom_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_5.mux_l2_in_0_ chanx_right_in[5] mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_6_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _075_/A sky130_fd_sc_hd__buf_4
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_091_ _091_/A VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l2_in_3_ _040_/HI chanx_left_in[18] mux_top_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_143_ prog_clk_1_N_in VGND VGND VPWR VPWR prog_clk_1_S_in sky130_fd_sc_hd__buf_2
X_074_ _074_/A VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_33.mux_l1_in_2_ chanx_left_in[0] bottom_left_grid_pin_49_ mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l2_in_3_ _052_/HI left_bottom_grid_pin_39_ mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_057_ chanx_right_in[17] VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xclkbuf_2_3_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
X_126_ chany_bottom_in[8] VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l4_in_0_ mux_top_track_24.mux_l3_in_1_/X mux_top_track_24.mux_l3_in_0_/X
+ mux_top_track_24.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_3_ _029_/HI left_bottom_grid_pin_38_ mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_109_ chany_top_in[5] VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xprog_clk_3_E_FTB01 prog_clk_3_E_in VGND VGND VPWR VPWR prog_clk_3_E_out sky130_fd_sc_hd__buf_4
XFILLER_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l4_in_0_ mux_left_track_17.mux_l3_in_1_/X mux_left_track_17.mux_l3_in_0_/X
+ mux_left_track_17.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_3_ _030_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l3_in_1_ mux_top_track_24.mux_l2_in_3_/X mux_top_track_24.mux_l2_in_2_/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ mux_bottom_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_6_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclk_2_W_FTB01 clk_2_E_in VGND VGND VPWR VPWR clk_2_W_out sky130_fd_sc_hd__buf_4
Xmux_left_track_17.mux_l3_in_1_ mux_left_track_17.mux_l2_in_3_/X mux_left_track_17.mux_l2_in_2_/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_090_ chanx_left_in[4] VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
Xmux_right_track_0.mux_l1_in_4_ chany_bottom_in[15] chany_bottom_in[12] mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l5_in_0_/X VGND
+ VGND VPWR VPWR _113_/A sky130_fd_sc_hd__buf_4
X_142_ clk_3_E_in VGND VGND VPWR VPWR clk_3_W_in sky130_fd_sc_hd__buf_2
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l2_in_2_ chanx_left_in[9] chanx_left_in[3] mux_top_track_24.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l1_in_1_ bottom_left_grid_pin_45_ chanx_right_in[19] mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_073_ _073_/A VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l2_in_2_ left_bottom_grid_pin_35_ chany_bottom_in[17] mux_left_track_17.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_056_ chanx_right_in[18] VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_125_ chany_bottom_in[9] VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_039_ VGND VGND VPWR VPWR _039_/HI _039_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_108_ chany_top_in[6] VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XFILLER_7_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_9.mux_l2_in_2_ left_bottom_grid_pin_34_ chany_bottom_in[16] mux_left_track_9.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] mux_right_track_0.mux_l1_in_4_/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _059_/A sky130_fd_sc_hd__buf_4
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_2.mux_l2_in_3_ _039_/HI chanx_left_in[19] mux_top_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_3_ _033_/HI chanx_left_in[18] mux_right_track_24.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l1_in_3_ chany_bottom_in[2] right_bottom_grid_pin_40_ mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l2_in_1_ chany_bottom_in[18] mux_top_track_24.mux_l1_in_2_/X
+ mux_top_track_24.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_0_ chanx_right_in[10] chany_top_in[10] mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ chanx_right_in[2] VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
X_141_ clk_3_E_in VGND VGND VPWR VPWR clk_3_S_in sky130_fd_sc_hd__buf_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_4_ chanx_left_in[4] chany_bottom_in[13] mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_17.mux_l2_in_1_ chany_bottom_in[8] mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_10 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ chany_bottom_in[10] VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
X_055_ VGND VGND VPWR VPWR _055_/HI _055_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_2.mux_l4_in_0_ mux_top_track_2.mux_l3_in_1_/X mux_top_track_2.mux_l3_in_0_/X
+ mux_top_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l1_in_2_ chany_bottom_in[9] chanx_right_in[19] mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l4_in_0_ mux_right_track_24.mux_l3_in_1_/X mux_right_track_24.mux_l3_in_0_/X
+ mux_right_track_24.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_038_ VGND VGND VPWR VPWR _038_/HI _038_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_2_ chany_bottom_in[7] chanx_right_in[17] mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ _107_/A VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_9.mux_l2_in_1_ chany_bottom_in[6] mux_left_track_9.mux_l1_in_2_/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_1_ mux_top_track_2.mux_l2_in_3_/X mux_top_track_2.mux_l2_in_2_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l2_in_1_ mux_right_track_0.mux_l1_in_3_/X mux_right_track_0.mux_l1_in_2_/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_1_ mux_right_track_24.mux_l2_in_3_/X mux_right_track_24.mux_l2_in_2_/X
+ mux_right_track_24.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_2_ chany_bottom_in[3] chanx_right_in[16] mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_2_ chanx_left_in[13] mux_top_track_2.mux_l1_in_4_/X mux_top_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l1_in_2_ right_bottom_grid_pin_38_ right_bottom_grid_pin_36_
+ mux_right_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l2_in_2_ chanx_left_in[9] chany_bottom_in[18] mux_right_track_24.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_140_ clk_3_E_in VGND VGND VPWR VPWR clk_3_N_in sky130_fd_sc_hd__buf_2
X_071_ _071_/A VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_2.mux_l1_in_3_ chany_bottom_in[4] chanx_right_in[13] mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclk_3_N_FTB01 clk_3_E_in VGND VGND VPWR VPWR clk_3_N_out sky130_fd_sc_hd__buf_4
Xmux_left_track_5.mux_l2_in_7_ _028_/HI left_bottom_grid_pin_41_ mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
XANTENNA_11 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_1_ chanx_right_in[18] chanx_right_in[9] mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_123_ _123_/A VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
X_054_ VGND VGND VPWR VPWR _054_/HI _054_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_037_ VGND VGND VPWR VPWR _037_/HI _037_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_1_ chanx_right_in[8] chany_top_in[17] mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l2_in_3_ _044_/HI chanx_left_in[12] mux_bottom_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_106_ chany_top_in[8] VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l1_in_4_ chanx_left_in[1] bottom_left_grid_pin_48_ mux_bottom_track_1.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_1_ chanx_right_in[6] chany_top_in[16] mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l4_in_0_ mux_bottom_track_1.mux_l3_in_1_/X mux_bottom_track_1.mux_l3_in_0_/X
+ mux_bottom_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_34_ chany_top_in[19] mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ chany_bottom_in[9] mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_070_ chanx_right_in[4] VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _123_/A sky130_fd_sc_hd__buf_4
XFILLER_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l3_in_1_ mux_bottom_track_1.mux_l2_in_3_/X mux_bottom_track_1.mux_l2_in_2_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_2.mux_l1_in_2_ chanx_right_in[4] chanx_right_in[3] mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_2_ chany_bottom_in[0] right_bottom_grid_pin_40_ mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l2_in_6_ left_bottom_grid_pin_40_ left_bottom_grid_pin_39_ mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_6_/X sky130_fd_sc_hd__mux2_1
XANTENNA_12 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_0_ top_left_grid_pin_48_ top_left_grid_pin_44_ mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_053_ VGND VGND VPWR VPWR _053_/HI _053_/LO sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_122_ chany_bottom_in[12] VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l2_in_2_ chanx_left_in[2] mux_bottom_track_1.mux_l1_in_4_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
X_105_ chany_top_in[9] VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_036_ VGND VGND VPWR VPWR _036_/HI _036_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _095_/A sky130_fd_sc_hd__buf_4
Xmux_bottom_track_1.mux_l1_in_3_ bottom_left_grid_pin_46_ bottom_left_grid_pin_44_
+ mux_bottom_track_1.mux_l1_in_4_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_9.mux_l1_in_0_ chany_top_in[11] chany_top_in[6] mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_right_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _134_/A sky130_fd_sc_hd__buf_4
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_mem_bottom_track_1.prog_clk clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_24.mux_l1_in_1_ right_bottom_grid_pin_36_ chany_top_in[18] mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l2_in_5_ left_bottom_grid_pin_38_ left_bottom_grid_pin_37_ mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_5_/X sky130_fd_sc_hd__mux2_1
XANTENNA_13 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_052_ VGND VGND VPWR VPWR _052_/HI _052_/LO sky130_fd_sc_hd__conb_1
X_121_ chany_bottom_in[13] VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l1_in_3_/X mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_035_ VGND VGND VPWR VPWR _035_/HI _035_/LO sky130_fd_sc_hd__conb_1
X_104_ chany_top_in[10] VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_42_ chanx_right_in[15] mux_bottom_track_1.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l3_in_3_ mux_left_track_5.mux_l2_in_7_/X mux_left_track_5.mux_l2_in_6_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xclk_2_S_FTB01 clk_2_E_in VGND VGND VPWR VPWR clk_2_S_out sky130_fd_sc_hd__buf_4
Xclkbuf_3_0_0_mem_bottom_track_1.prog_clk clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_0_ chany_top_in[11] chany_top_in[9] mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_4_ left_bottom_grid_pin_36_ left_bottom_grid_pin_35_ mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_4_/X sky130_fd_sc_hd__mux2_1
XANTENNA_14 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_120_ chany_bottom_in[14] VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
X_051_ VGND VGND VPWR VPWR _051_/HI _051_/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_5.mux_l5_in_0_ mux_left_track_5.mux_l4_in_1_/X mux_left_track_5.mux_l4_in_0_/X
+ mux_left_track_5.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_034_ VGND VGND VPWR VPWR _034_/HI _034_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ _103_/A VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l4_in_1_ mux_left_track_5.mux_l3_in_3_/X mux_left_track_5.mux_l3_in_2_/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l1_in_1_ chanx_right_in[12] chanx_right_in[2] mux_bottom_track_1.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_2_ mux_left_track_5.mux_l2_in_5_/X mux_left_track_5.mux_l2_in_4_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_4_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ ccff_head VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_3_ left_bottom_grid_pin_34_ chany_bottom_in[14] mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_050_ VGND VGND VPWR VPWR _050_/HI _050_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_033_ VGND VGND VPWR VPWR _033_/HI _033_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _115_/A sky130_fd_sc_hd__buf_4
X_102_ chany_top_in[12] VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
XFILLER_8_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_4_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_4_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_16 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_25.mux_l2_in_3_ _053_/HI left_bottom_grid_pin_40_ mux_left_track_25.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
Xmux_left_track_5.mux_l2_in_2_ chany_bottom_in[5] chany_bottom_in[1] mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_101_ chany_top_in[13] VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
X_032_ VGND VGND VPWR VPWR _032_/HI _032_/LO sky130_fd_sc_hd__conb_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l4_in_0_ mux_left_track_25.mux_l3_in_1_/X mux_left_track_25.mux_l3_in_0_/X
+ mux_left_track_25.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _067_/A sky130_fd_sc_hd__buf_4
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_0.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l3_in_1_ mux_left_track_25.mux_l2_in_3_/X mux_left_track_25.mux_l2_in_2_/X
+ mux_left_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_17 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_25.mux_l2_in_2_ left_bottom_grid_pin_36_ chany_bottom_in[18] mux_left_track_25.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l2_in_1_ chanx_right_in[14] chanx_right_in[5] mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l1_in_3_ _041_/HI chanx_left_in[10] mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
X_031_ VGND VGND VPWR VPWR _031_/HI _031_/LO sky130_fd_sc_hd__conb_1
Xclkbuf_3_7_0_mem_bottom_track_1.prog_clk clkbuf_3_6_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_100_ chany_top_in[14] VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_2_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__dfxtp_1
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_2_E_FTB01 prog_clk_2_E_in VGND VGND VPWR VPWR prog_clk_2_E_out sky130_fd_sc_hd__buf_4
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l2_in_3_ _043_/HI chanx_left_in[16] mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.mux_l2_in_1_ mux_top_track_32.mux_l1_in_3_/X mux_top_track_32.mux_l1_in_2_/X
+ mux_top_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclk_1_W_FTB01 clk_1_N_in VGND VGND VPWR VPWR clk_1_W_out sky130_fd_sc_hd__buf_4
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_18 ANTENNA_18/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_0_ chany_top_in[15] mux_left_track_5.mux_l1_in_0_/X mux_left_track_5.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_8.mux_l4_in_0_ mux_top_track_8.mux_l3_in_1_/X mux_top_track_8.mux_l3_in_0_/X
+ mux_top_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l2_in_1_ chany_bottom_in[11] mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.mux_l1_in_2_ chanx_left_in[1] chany_bottom_in[10] mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_030_ VGND VGND VPWR VPWR _030_/HI _030_/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_8.mux_l3_in_1_ mux_top_track_8.mux_l2_in_3_/X mux_top_track_8.mux_l2_in_2_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l1_in_2_ chany_bottom_in[9] chanx_right_in[18] mux_left_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_33.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[6] mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_32.mux_l2_in_0_ mux_top_track_32.mux_l1_in_1_/X mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_32.mux_l1_in_3_ _034_/HI chanx_left_in[10] mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l1_in_1_ chanx_right_in[10] chanx_right_in[0] mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_left_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_089_ chanx_left_in[5] VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l1_in_1_ chanx_right_in[9] chany_top_in[18] mux_left_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_4_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l2_in_1_ chany_bottom_in[16] mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_32.mux_l2_in_1_ mux_right_track_32.mux_l1_in_3_/X mux_right_track_32.mux_l1_in_2_/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l1_in_2_ chany_bottom_in[6] chanx_right_in[16] mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_32.mux_l1_in_2_ chany_bottom_in[19] chany_bottom_in[10] mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.mux_l1_in_0_ top_left_grid_pin_49_ top_left_grid_pin_45_ mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclk_2_N_FTB01 clk_2_E_in VGND VGND VPWR VPWR clk_2_N_out sky130_fd_sc_hd__buf_4
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_0_ chany_top_in[9] chany_top_in[3] mux_left_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_088_ chanx_left_in[6] VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XFILLER_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.mux_l2_in_7_ _042_/HI chanx_left_in[15] mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_7_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_32.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_4_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__buf_4
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _131_/A sky130_fd_sc_hd__buf_4
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[6] mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_32.mux_l1_in_1_ right_bottom_grid_pin_41_ right_bottom_grid_pin_37_
+ mux_right_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_3_W_FTB01 prog_clk_3_E_in VGND VGND VPWR VPWR prog_clk_3_W_out sky130_fd_sc_hd__buf_4
X_087_ _087_/A VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.mux_l2_in_6_ chanx_left_in[14] chanx_left_in[5] mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_139_ clk_2_E_in VGND VGND VPWR VPWR clk_2_W_in sky130_fd_sc_hd__buf_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__buf_4
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_1.mux_l2_in_3_ _051_/HI left_bottom_grid_pin_40_ mux_left_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_mem_bottom_track_1.prog_clk clkbuf_3_6_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l1_in_0_ top_left_grid_pin_46_ top_left_grid_pin_42_ mux_top_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_4_ left_bottom_grid_pin_36_ left_bottom_grid_pin_34_ mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l1_in_0_ chany_top_in[15] chany_top_in[10] mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_right_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_0_0_mem_bottom_track_1.prog_clk clkbuf_2_1_0_mem_bottom_track_1.prog_clk/A
+ VGND VGND VPWR VPWR clkbuf_2_0_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_086_ chanx_left_in[8] VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XFILLER_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l2_in_5_ chany_bottom_in[14] chany_bottom_in[5] mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_5_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _074_/A sky130_fd_sc_hd__buf_4
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_069_ chanx_right_in[5] VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
X_138_ clk_2_E_in VGND VGND VPWR VPWR clk_2_S_in sky130_fd_sc_hd__buf_2
Xclk_3_E_FTB01 clk_3_E_in VGND VGND VPWR VPWR clk_3_E_out sky130_fd_sc_hd__buf_4
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_2_ left_bottom_grid_pin_38_ mux_left_track_1.mux_l1_in_4_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_16.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_3_ chany_bottom_in[19] chany_bottom_in[12] mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_3_ mux_top_track_4.mux_l2_in_7_/X mux_top_track_4.mux_l2_in_6_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_2.mux_l2_in_3_ _032_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l2_in_4_ chanx_right_in[14] chanx_right_in[7] mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_4_/X sky130_fd_sc_hd__mux2_1
X_085_ chanx_left_in[9] VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_4_ chany_bottom_in[13] chany_bottom_in[11] mux_right_track_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_137_ clk_2_E_in VGND VGND VPWR VPWR clk_2_N_in sky130_fd_sc_hd__buf_2
Xmux_top_track_4.mux_l5_in_0_ mux_top_track_4.mux_l4_in_1_/X mux_top_track_4.mux_l4_in_0_/X
+ mux_top_track_4.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l5_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_068_ chanx_right_in[6] VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l1_in_3_/X mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.mux_l4_in_1_ mux_top_track_4.mux_l3_in_3_/X mux_top_track_4.mux_l3_in_2_/X
+ mux_top_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_right_track_16.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l1_in_2_ chany_bottom_in[2] chanx_right_in[12] mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_2_ mux_top_track_4.mux_l2_in_5_/X mux_top_track_4.mux_l2_in_4_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] mux_right_track_2.mux_l1_in_4_/X
+ mux_right_track_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l5_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
X_084_ chanx_left_in[10] VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_2.mux_l1_in_3_ chany_bottom_in[4] right_bottom_grid_pin_41_ mux_right_track_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l2_in_3_ chanx_right_in[5] top_left_grid_pin_49_ mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_136_ clk_1_N_in VGND VGND VPWR VPWR clk_1_S_in sky130_fd_sc_hd__buf_2
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_067_ _067_/A VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_2_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_119_ _119_/A VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l4_in_0_ mux_top_track_4.mux_l3_in_1_/X mux_top_track_4.mux_l3_in_0_/X
+ mux_top_track_4.mux_l4_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_0 Test_en_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_1_ chanx_right_in[2] chany_top_in[12] mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_1_ mux_top_track_4.mux_l2_in_3_/X mux_top_track_4.mux_l2_in_2_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_083_ _083_/A VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_2.mux_l1_in_2_ right_bottom_grid_pin_39_ right_bottom_grid_pin_37_
+ mux_right_track_2.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l2_in_2_ top_left_grid_pin_48_ top_left_grid_pin_47_ mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.mux_l1_in_3_ _055_/HI left_bottom_grid_pin_41_ mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_135_ _135_/A VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l2_in_3_ _045_/HI chanx_left_in[17] mux_bottom_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_066_ chanx_right_in[8] VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_2_3_0_mem_bottom_track_1.prog_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_049_ VGND VGND VPWR VPWR _049_/HI _049_/LO sky130_fd_sc_hd__conb_1
X_118_ chany_bottom_in[16] VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail VGND VGND VPWR VPWR mux_left_track_33.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_17.mux_l4_in_0_ mux_bottom_track_17.mux_l3_in_1_/X mux_bottom_track_17.mux_l3_in_0_/X
+ mux_bottom_track_17.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l2_in_3_ _047_/HI chanx_left_in[13] mux_bottom_track_3.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[2] chany_top_in[0] mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ mux_left_track_33.mux_l1_in_3_/X mux_left_track_33.mux_l1_in_2_/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l3_in_1_ mux_bottom_track_17.mux_l2_in_3_/X mux_bottom_track_17.mux_l2_in_2_/X
+ mux_bottom_track_17.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_4_ chanx_left_in[3] bottom_left_grid_pin_49_ mux_bottom_track_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
X_082_ chanx_left_in[12] VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _119_/A sky130_fd_sc_hd__buf_4
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ top_left_grid_pin_46_ top_left_grid_pin_45_ mux_top_track_4.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_35_ chany_top_in[13] mux_right_track_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l4_in_0_ mux_bottom_track_3.mux_l3_in_1_/X mux_bottom_track_3.mux_l3_in_0_/X
+ mux_bottom_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_2_ left_bottom_grid_pin_37_ chany_bottom_in[15] mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xprog_clk_3_S_FTB01 prog_clk_3_E_in VGND VGND VPWR VPWR prog_clk_3_S_out sky130_fd_sc_hd__buf_4
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_134_ _134_/A VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_17.mux_l2_in_2_ chanx_left_in[15] chanx_left_in[8] mux_bottom_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_065_ chanx_right_in[9] VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xclkbuf_3_5_0_mem_bottom_track_1.prog_clk clkbuf_2_2_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l3_in_1_ mux_bottom_track_3.mux_l2_in_3_/X mux_bottom_track_3.mux_l2_in_2_/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_117_ chany_bottom_in[17] VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_048_ VGND VGND VPWR VPWR _048_/HI _048_/LO sky130_fd_sc_hd__conb_1
Xprog_clk_1_E_FTB01 prog_clk_1_N_in VGND VGND VPWR VPWR prog_clk_1_E_out sky130_fd_sc_hd__buf_4
XANTENNA_2 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l2_in_2_ chanx_left_in[4] mux_bottom_track_3.mux_l1_in_4_/X
+ mux_bottom_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l3_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l1_in_3_ bottom_left_grid_pin_47_ bottom_left_grid_pin_45_
+ mux_bottom_track_3.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_3_/X
+ sky130_fd_sc_hd__mux2_1
X_081_ chanx_left_in[13] VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _094_/A sky130_fd_sc_hd__buf_4
Xmux_top_track_4.mux_l2_in_0_ top_left_grid_pin_44_ mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTest_en_N_FTB01 Test_en_S_in VGND VGND VPWR VPWR Test_en_N_out sky130_fd_sc_hd__buf_4
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[4] chany_top_in[0] mux_right_track_2.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_right_track_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_1_ chany_bottom_in[10] chanx_right_in[10] mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l5_in_0_/X VGND VGND
+ VPWR VPWR _133_/A sky130_fd_sc_hd__buf_4
X_133_ _133_/A VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_17.mux_l2_in_1_ bottom_left_grid_pin_47_ mux_bottom_track_17.mux_l1_in_2_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_064_ chanx_right_in[10] VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_047_ VGND VGND VPWR VPWR _047_/HI _047_/LO sky130_fd_sc_hd__conb_1
X_116_ chany_bottom_in[18] VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_2_ bottom_left_grid_pin_43_ chanx_right_in[17] mux_bottom_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_3 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l1_in_3_/X mux_bottom_track_3.mux_l1_in_2_/X
+ mux_bottom_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_2.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_track_2.mux_l2_in_2_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l1_in_2_ bottom_left_grid_pin_43_ chanx_right_in[13] mux_bottom_track_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
X_080_ chanx_left_in[14] VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0_0_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l1_in_0_ chany_top_in[10] chany_top_in[1] mux_left_track_33.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_132_ chany_bottom_in[2] VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
X_063_ _063_/A VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_right_track_8.mux_l2_in_2_/S VGND VGND VPWR VPWR mux_right_track_8.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_43_ top_left_grid_pin_42_ mux_top_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_046_ VGND VGND VPWR VPWR _046_/HI _046_/LO sky130_fd_sc_hd__conb_1
X_115_ _115_/A VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l5_in_0_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4_0_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l4_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ chanx_right_in[8] chanx_right_in[1] mux_bottom_track_17.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_029_ VGND VGND VPWR VPWR _029_/HI _029_/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6_0_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

