magic
tech EFS8A
magscale 1 2
timestamp 1603804930
<< locali >>
rect 395129 385595 395163 395149
rect 395313 364991 395347 366317
rect 76257 353907 76291 357545
rect 104961 354927 104995 355097
rect 122165 354995 122199 355165
rect 216465 354995 216499 355165
rect 96773 350371 96807 351493
rect 191257 350371 191291 351833
rect 284545 350371 284579 351561
rect 75429 331603 75463 334765
rect 75429 330107 75463 331569
rect 75521 331671 75555 334697
rect 75981 334527 76015 349657
rect 395313 345611 395347 363461
rect 212785 334459 212819 334561
rect 221065 334255 221099 334561
rect 201745 331739 201779 331841
rect 75521 330175 75555 331637
rect 211313 331603 211347 331841
rect 154825 329087 154859 329189
rect 147775 329053 148017 329087
rect 174145 328883 174179 329189
rect 176847 329053 176905 329087
rect 182425 328883 182459 329257
rect 191993 329155 192027 329257
rect 186507 329053 186657 329087
rect 163381 327319 163415 327489
rect 168257 327251 168291 327421
rect 168349 327319 168383 327489
rect 174053 327251 174087 327421
rect 181045 327387 181079 327489
rect 183805 326979 183839 327421
rect 196225 327047 196259 327421
rect 248113 326979 248147 327217
rect 32039 326469 32097 326503
rect 19585 326299 19619 326401
rect 29153 326299 29187 326469
rect 58225 326163 58259 326401
rect 73865 326299 73899 326673
rect 162369 326639 162403 326945
rect 253023 326741 253173 326775
rect 258233 326503 258267 327353
rect 345909 326911 345943 327285
rect 348025 326571 348059 327285
rect 338365 326435 338399 326537
rect 347933 326435 347967 326537
rect 67793 326163 67827 326265
rect 137713 316643 137747 326197
rect 352809 325211 352843 326809
rect 354465 326367 354499 326877
rect 352717 291007 352751 291721
rect 367345 291075 367379 291177
rect 352993 279379 353027 290973
rect 357685 290871 357719 290973
rect 362469 290871 362503 291041
rect 376913 291007 376947 291177
rect 386665 291143 386699 291245
rect 379673 291109 379857 291143
rect 379673 291007 379707 291109
rect 396233 291075 396267 291245
rect 399027 291041 399085 291075
rect 395129 282099 395163 288865
rect 154733 274415 154767 274721
rect 154825 274279 154859 274857
rect 51417 269723 51451 272477
rect 253633 266459 253667 266765
rect 252989 266255 253023 266357
rect 154825 263603 154859 263705
rect 164393 263535 164427 263705
rect 203125 263671 203159 263773
rect 174145 263535 174179 263637
rect 167153 263501 167245 263535
rect 183713 263535 183747 263637
rect 212693 263603 212727 263773
rect 186507 263501 186565 263535
rect 167153 263467 167187 263501
rect 215545 263467 215579 263569
rect 241673 263535 241707 263637
rect 321747 263637 321805 263671
rect 241765 263467 241799 263569
rect 73865 262515 73899 263433
rect 250597 263331 250631 263569
rect 312145 263467 312179 263637
rect 272769 263331 272803 263433
rect 277645 263263 277679 263433
rect 287213 263263 287247 263433
rect 296965 263263 296999 263433
rect 331373 263467 331407 263637
rect 336893 263467 336927 263569
rect 336985 263467 337019 263569
rect 341159 263501 341309 263535
rect 302669 263263 302703 263433
rect 237809 262311 237843 262753
rect 263845 262311 263879 262753
rect 156849 232935 156883 233309
rect 341343 225285 341493 225319
rect 335605 224435 335639 224809
rect 341217 224775 341251 225217
rect 343149 224367 343183 230317
rect 345909 224571 345943 225217
rect 348025 223075 348059 224333
rect 34857 213895 34891 220457
rect 369093 216887 369127 219437
rect 369369 216751 369403 219369
rect 369001 214439 369035 214541
rect 34857 204715 34891 206857
rect 369829 192407 369863 199445
rect 369829 182751 369863 192237
rect 345357 180779 345391 181153
rect 345265 180575 345299 180745
rect 254921 172211 254955 172925
rect 73497 168879 73531 169389
rect 369829 153715 369863 156469
rect 173685 150655 173719 151641
rect 186749 142223 186783 142325
rect 193465 142223 193499 142801
rect 203033 142291 203067 142801
rect 85825 140659 85859 140761
rect 157953 139639 157987 139877
rect 253265 138959 253299 139469
rect 253357 138891 253391 139401
rect 254921 139299 254955 139537
rect 255933 139503 255967 139877
rect 254829 139163 254863 139265
rect 341769 138687 341803 138789
rect 236245 124815 236279 134369
rect 340021 130867 340055 131037
rect 345265 130799 345299 130901
rect 357685 130323 357719 134369
rect 357685 124815 357719 130289
rect 369553 124883 369587 132873
rect 74049 117743 74083 124713
rect 369645 124679 369679 132941
rect 51693 108019 51727 115057
rect 360295 115057 360445 115091
rect 369863 115057 370047 115091
rect 236245 105503 236279 115057
rect 370013 115023 370047 115057
rect 236245 95031 236279 95745
rect 340389 86735 340423 86905
rect 340757 86667 340791 86973
rect 65401 78371 65435 78745
rect 369921 76467 369955 81329
rect 155377 73747 155411 75481
rect 249217 73747 249251 75413
rect 129433 57155 129467 66709
rect 134033 54911 134067 55013
rect 96773 48519 96807 50933
rect 357317 48927 357351 49505
rect 357317 48179 357351 48893
rect 109377 47635 109411 47669
rect 109227 47601 109411 47635
rect 124465 47635 124499 47737
rect 134033 47635 134067 47737
rect 95117 47227 95151 47533
rect 95485 47431 95519 47533
rect 105053 47431 105087 47601
rect 86101 46139 86135 46785
<< viali >>
rect 395129 395149 395163 395183
rect 395129 385561 395163 385595
rect 395313 366317 395347 366351
rect 395313 364957 395347 364991
rect 395313 363461 395347 363495
rect 76257 357545 76291 357579
rect 122165 355165 122199 355199
rect 104961 355097 104995 355131
rect 122165 354961 122199 354995
rect 216465 355165 216499 355199
rect 216465 354961 216499 354995
rect 104961 354893 104995 354927
rect 76257 353873 76291 353907
rect 191257 351833 191291 351867
rect 96773 351493 96807 351527
rect 96773 350337 96807 350371
rect 191257 350337 191291 350371
rect 284545 351561 284579 351595
rect 284545 350337 284579 350371
rect 75981 349657 76015 349691
rect 75429 334765 75463 334799
rect 75429 331569 75463 331603
rect 75521 334697 75555 334731
rect 395313 345577 395347 345611
rect 75981 334493 76015 334527
rect 212785 334561 212819 334595
rect 212785 334425 212819 334459
rect 221065 334561 221099 334595
rect 221065 334221 221099 334255
rect 201745 331841 201779 331875
rect 201745 331705 201779 331739
rect 211313 331841 211347 331875
rect 75521 331637 75555 331671
rect 211313 331569 211347 331603
rect 75521 330141 75555 330175
rect 75429 330073 75463 330107
rect 182425 329257 182459 329291
rect 154825 329189 154859 329223
rect 147741 329053 147775 329087
rect 148017 329053 148051 329087
rect 154825 329053 154859 329087
rect 174145 329189 174179 329223
rect 176813 329053 176847 329087
rect 176905 329053 176939 329087
rect 174145 328849 174179 328883
rect 191993 329257 192027 329291
rect 191993 329121 192027 329155
rect 186473 329053 186507 329087
rect 186657 329053 186691 329087
rect 182425 328849 182459 328883
rect 163381 327489 163415 327523
rect 168349 327489 168383 327523
rect 163381 327285 163415 327319
rect 168257 327421 168291 327455
rect 181045 327489 181079 327523
rect 168349 327285 168383 327319
rect 174053 327421 174087 327455
rect 168257 327217 168291 327251
rect 181045 327353 181079 327387
rect 183805 327421 183839 327455
rect 174053 327217 174087 327251
rect 196225 327421 196259 327455
rect 258233 327353 258267 327387
rect 196225 327013 196259 327047
rect 248113 327217 248147 327251
rect 162369 326945 162403 326979
rect 183805 326945 183839 326979
rect 248113 326945 248147 326979
rect 73865 326673 73899 326707
rect 29153 326469 29187 326503
rect 32005 326469 32039 326503
rect 32097 326469 32131 326503
rect 19585 326401 19619 326435
rect 19585 326265 19619 326299
rect 29153 326265 29187 326299
rect 58225 326401 58259 326435
rect 252989 326741 253023 326775
rect 253173 326741 253207 326775
rect 162369 326605 162403 326639
rect 345909 327285 345943 327319
rect 345909 326877 345943 326911
rect 348025 327285 348059 327319
rect 354465 326877 354499 326911
rect 258233 326469 258267 326503
rect 338365 326537 338399 326571
rect 338365 326401 338399 326435
rect 347933 326537 347967 326571
rect 348025 326537 348059 326571
rect 352809 326809 352843 326843
rect 347933 326401 347967 326435
rect 58225 326129 58259 326163
rect 67793 326265 67827 326299
rect 73865 326265 73899 326299
rect 67793 326129 67827 326163
rect 137713 326197 137747 326231
rect 354465 326333 354499 326367
rect 352809 325177 352843 325211
rect 137713 316609 137747 316643
rect 352717 291721 352751 291755
rect 386665 291245 386699 291279
rect 367345 291177 367379 291211
rect 362469 291041 362503 291075
rect 367345 291041 367379 291075
rect 376913 291177 376947 291211
rect 352717 290973 352751 291007
rect 352993 290973 353027 291007
rect 357685 290973 357719 291007
rect 357685 290837 357719 290871
rect 376913 290973 376947 291007
rect 379857 291109 379891 291143
rect 386665 291109 386699 291143
rect 396233 291245 396267 291279
rect 396233 291041 396267 291075
rect 398993 291041 399027 291075
rect 399085 291041 399119 291075
rect 379673 290973 379707 291007
rect 362469 290837 362503 290871
rect 395129 288865 395163 288899
rect 395129 282065 395163 282099
rect 352993 279345 353027 279379
rect 154825 274857 154859 274891
rect 154733 274721 154767 274755
rect 154733 274381 154767 274415
rect 154825 274245 154859 274279
rect 51417 272477 51451 272511
rect 51417 269689 51451 269723
rect 253633 266765 253667 266799
rect 253633 266425 253667 266459
rect 252989 266357 253023 266391
rect 252989 266221 253023 266255
rect 203125 263773 203159 263807
rect 154825 263705 154859 263739
rect 154825 263569 154859 263603
rect 164393 263705 164427 263739
rect 174145 263637 174179 263671
rect 164393 263501 164427 263535
rect 167245 263501 167279 263535
rect 174145 263501 174179 263535
rect 183713 263637 183747 263671
rect 203125 263637 203159 263671
rect 212693 263773 212727 263807
rect 241673 263637 241707 263671
rect 212693 263569 212727 263603
rect 215545 263569 215579 263603
rect 183713 263501 183747 263535
rect 186473 263501 186507 263535
rect 186565 263501 186599 263535
rect 73865 263433 73899 263467
rect 167153 263433 167187 263467
rect 312145 263637 312179 263671
rect 321713 263637 321747 263671
rect 321805 263637 321839 263671
rect 331373 263637 331407 263671
rect 241673 263501 241707 263535
rect 241765 263569 241799 263603
rect 215545 263433 215579 263467
rect 241765 263433 241799 263467
rect 250597 263569 250631 263603
rect 250597 263297 250631 263331
rect 272769 263433 272803 263467
rect 272769 263297 272803 263331
rect 277645 263433 277679 263467
rect 277645 263229 277679 263263
rect 287213 263433 287247 263467
rect 287213 263229 287247 263263
rect 296965 263433 296999 263467
rect 296965 263229 296999 263263
rect 302669 263433 302703 263467
rect 312145 263433 312179 263467
rect 331373 263433 331407 263467
rect 336893 263569 336927 263603
rect 336893 263433 336927 263467
rect 336985 263569 337019 263603
rect 341125 263501 341159 263535
rect 341309 263501 341343 263535
rect 336985 263433 337019 263467
rect 302669 263229 302703 263263
rect 73865 262481 73899 262515
rect 237809 262753 237843 262787
rect 237809 262277 237843 262311
rect 263845 262753 263879 262787
rect 263845 262277 263879 262311
rect 156849 233309 156883 233343
rect 156849 232901 156883 232935
rect 343149 230317 343183 230351
rect 341309 225285 341343 225319
rect 341493 225285 341527 225319
rect 341217 225217 341251 225251
rect 335605 224809 335639 224843
rect 341217 224741 341251 224775
rect 335605 224401 335639 224435
rect 345909 225217 345943 225251
rect 345909 224537 345943 224571
rect 343149 224333 343183 224367
rect 348025 224333 348059 224367
rect 348025 223041 348059 223075
rect 34857 220457 34891 220491
rect 369093 219437 369127 219471
rect 369093 216853 369127 216887
rect 369369 219369 369403 219403
rect 369369 216717 369403 216751
rect 369001 214541 369035 214575
rect 369001 214405 369035 214439
rect 34857 213861 34891 213895
rect 34857 206857 34891 206891
rect 34857 204681 34891 204715
rect 369829 199445 369863 199479
rect 369829 192373 369863 192407
rect 369829 192237 369863 192271
rect 369829 182717 369863 182751
rect 345357 181153 345391 181187
rect 345265 180745 345299 180779
rect 345357 180745 345391 180779
rect 345265 180541 345299 180575
rect 254921 172925 254955 172959
rect 254921 172177 254955 172211
rect 73497 169389 73531 169423
rect 73497 168845 73531 168879
rect 369829 156469 369863 156503
rect 369829 153681 369863 153715
rect 173685 151641 173719 151675
rect 173685 150621 173719 150655
rect 193465 142801 193499 142835
rect 186749 142325 186783 142359
rect 186749 142189 186783 142223
rect 203033 142801 203067 142835
rect 203033 142257 203067 142291
rect 193465 142189 193499 142223
rect 85825 140761 85859 140795
rect 85825 140625 85859 140659
rect 157953 139877 157987 139911
rect 157953 139605 157987 139639
rect 255933 139877 255967 139911
rect 254921 139537 254955 139571
rect 253265 139469 253299 139503
rect 253265 138925 253299 138959
rect 253357 139401 253391 139435
rect 255933 139469 255967 139503
rect 254829 139265 254863 139299
rect 254921 139265 254955 139299
rect 254829 139129 254863 139163
rect 253357 138857 253391 138891
rect 341769 138789 341803 138823
rect 341769 138653 341803 138687
rect 236245 134369 236279 134403
rect 357685 134369 357719 134403
rect 340021 131037 340055 131071
rect 340021 130833 340055 130867
rect 345265 130901 345299 130935
rect 345265 130765 345299 130799
rect 236245 124781 236279 124815
rect 369645 132941 369679 132975
rect 357685 130289 357719 130323
rect 369553 132873 369587 132907
rect 369553 124849 369587 124883
rect 357685 124781 357719 124815
rect 74049 124713 74083 124747
rect 369645 124645 369679 124679
rect 74049 117709 74083 117743
rect 51693 115057 51727 115091
rect 51693 107985 51727 108019
rect 236245 115057 236279 115091
rect 360261 115057 360295 115091
rect 360445 115057 360479 115091
rect 369829 115057 369863 115091
rect 370013 114989 370047 115023
rect 236245 105469 236279 105503
rect 236245 95745 236279 95779
rect 236245 94997 236279 95031
rect 340757 86973 340791 87007
rect 340389 86905 340423 86939
rect 340389 86701 340423 86735
rect 340757 86633 340791 86667
rect 369921 81329 369955 81363
rect 65401 78745 65435 78779
rect 65401 78337 65435 78371
rect 369921 76433 369955 76467
rect 155377 75481 155411 75515
rect 155377 73713 155411 73747
rect 249217 75413 249251 75447
rect 249217 73713 249251 73747
rect 129433 66709 129467 66743
rect 129433 57121 129467 57155
rect 134033 55013 134067 55047
rect 134033 54877 134067 54911
rect 96773 50933 96807 50967
rect 96773 48485 96807 48519
rect 357317 49505 357351 49539
rect 357317 48893 357351 48927
rect 357317 48145 357351 48179
rect 124465 47737 124499 47771
rect 109377 47669 109411 47703
rect 105053 47601 105087 47635
rect 109193 47601 109227 47635
rect 124465 47601 124499 47635
rect 134033 47737 134067 47771
rect 134033 47601 134067 47635
rect 95117 47533 95151 47567
rect 95485 47533 95519 47567
rect 95485 47397 95519 47431
rect 105053 47397 105087 47431
rect 95117 47193 95151 47227
rect 86101 46785 86135 46819
rect 86101 46105 86135 46139
<< metal1 >>
rect 395114 395180 395120 395192
rect 395075 395152 395120 395180
rect 395114 395140 395120 395152
rect 395172 395140 395178 395192
rect 22330 393780 22336 393832
rect 22388 393820 22394 393832
rect 23158 393820 23164 393832
rect 22388 393792 23164 393820
rect 22388 393780 22394 393792
rect 23158 393780 23164 393792
rect 23216 393780 23222 393832
rect 48550 393780 48556 393832
rect 48608 393820 48614 393832
rect 49654 393820 49660 393832
rect 48608 393792 49660 393820
rect 48608 393780 48614 393792
rect 49654 393780 49660 393792
rect 49712 393780 49718 393832
rect 128590 393780 128596 393832
rect 128648 393820 128654 393832
rect 129418 393820 129424 393832
rect 128648 393792 129424 393820
rect 128648 393780 128654 393792
rect 129418 393780 129424 393792
rect 129476 393780 129482 393832
rect 154810 393780 154816 393832
rect 154868 393820 154874 393832
rect 155914 393820 155920 393832
rect 154868 393792 155920 393820
rect 154868 393780 154874 393792
rect 155914 393780 155920 393792
rect 155972 393780 155978 393832
rect 234850 393780 234856 393832
rect 234908 393820 234914 393832
rect 235678 393820 235684 393832
rect 234908 393792 235684 393820
rect 234908 393780 234914 393792
rect 235678 393780 235684 393792
rect 235736 393780 235742 393832
rect 261070 393780 261076 393832
rect 261128 393820 261134 393832
rect 262174 393820 262180 393832
rect 261128 393792 262180 393820
rect 261128 393780 261134 393792
rect 262174 393780 262180 393792
rect 262232 393780 262238 393832
rect 279654 393168 279660 393220
rect 279712 393208 279718 393220
rect 315350 393208 315356 393220
rect 279712 393180 315356 393208
rect 279712 393168 279718 393180
rect 315350 393168 315356 393180
rect 315408 393168 315414 393220
rect 102830 393100 102836 393152
rect 102888 393140 102894 393152
rect 108902 393140 108908 393152
rect 102888 393112 108908 393140
rect 102888 393100 102894 393112
rect 108902 393100 108908 393112
rect 108960 393100 108966 393152
rect 314614 393100 314620 393152
rect 314672 393140 314678 393152
rect 421610 393140 421616 393152
rect 314672 393112 421616 393140
rect 314672 393100 314678 393112
rect 421610 393100 421616 393112
rect 421668 393100 421674 393152
rect 284438 392488 284444 392540
rect 284496 392528 284502 392540
rect 288762 392528 288768 392540
rect 284496 392500 288768 392528
rect 284496 392488 284502 392500
rect 288762 392488 288768 392500
rect 288820 392488 288826 392540
rect 13130 391060 13136 391112
rect 13188 391100 13194 391112
rect 87190 391100 87196 391112
rect 13188 391072 87196 391100
rect 13188 391060 13194 391072
rect 87190 391060 87196 391072
rect 87248 391060 87254 391112
rect 299618 389700 299624 389752
rect 299676 389740 299682 389752
rect 429430 389740 429436 389752
rect 299676 389712 429436 389740
rect 299676 389700 299682 389712
rect 429430 389700 429436 389712
rect 429488 389700 429494 389752
rect 108902 389428 108908 389480
rect 108960 389468 108966 389480
rect 111294 389468 111300 389480
rect 108960 389440 111300 389468
rect 108960 389428 108966 389440
rect 111294 389428 111300 389440
rect 111352 389428 111358 389480
rect 195290 389156 195296 389208
rect 195348 389196 195354 389208
rect 208630 389196 208636 389208
rect 195348 389168 208636 389196
rect 195348 389156 195354 389168
rect 208630 389156 208636 389168
rect 208688 389156 208694 389208
rect 76150 389088 76156 389140
rect 76208 389128 76214 389140
rect 116262 389128 116268 389140
rect 76208 389100 116268 389128
rect 76208 389088 76214 389100
rect 116262 389088 116268 389100
rect 116320 389088 116326 389140
rect 182410 389088 182416 389140
rect 182468 389128 182474 389140
rect 200350 389128 200356 389140
rect 182468 389100 200356 389128
rect 182468 389088 182474 389100
rect 200350 389088 200356 389100
rect 200408 389088 200414 389140
rect 48550 389020 48556 389072
rect 48608 389060 48614 389072
rect 121322 389060 121328 389072
rect 48608 389032 121328 389060
rect 48608 389020 48614 389032
rect 121322 389020 121328 389032
rect 121380 389020 121386 389072
rect 154810 389020 154816 389072
rect 154868 389060 154874 389072
rect 205318 389060 205324 389072
rect 154868 389032 205324 389060
rect 154868 389020 154874 389032
rect 205318 389020 205324 389032
rect 205376 389020 205382 389072
rect 261070 389020 261076 389072
rect 261128 389060 261134 389072
rect 288946 389060 288952 389072
rect 261128 389032 288952 389060
rect 261128 389020 261134 389032
rect 288946 389020 288952 389032
rect 289004 389020 289010 389072
rect 22330 388952 22336 389004
rect 22388 388992 22394 389004
rect 126290 388992 126296 389004
rect 22388 388964 126296 388992
rect 22388 388952 22394 388964
rect 126290 388952 126296 388964
rect 126348 388952 126354 389004
rect 128590 388952 128596 389004
rect 128648 388992 128654 389004
rect 210286 388992 210292 389004
rect 128648 388964 210292 388992
rect 128648 388952 128654 388964
rect 210286 388952 210292 388964
rect 210344 388952 210350 389004
rect 234850 388952 234856 389004
rect 234908 388992 234914 389004
rect 294190 388992 294196 389004
rect 234908 388964 294196 388992
rect 234908 388952 234914 388964
rect 294190 388952 294196 388964
rect 294248 388952 294254 389004
rect 91330 388680 91336 388732
rect 91388 388720 91394 388732
rect 358498 388720 358504 388732
rect 91388 388692 358504 388720
rect 91388 388680 91394 388692
rect 358498 388680 358504 388692
rect 358556 388680 358562 388732
rect 13498 388612 13504 388664
rect 13556 388652 13562 388664
rect 96298 388652 96304 388664
rect 13556 388624 96304 388652
rect 13556 388612 13562 388624
rect 96298 388612 96304 388624
rect 96356 388612 96362 388664
rect 13314 388544 13320 388596
rect 13372 388584 13378 388596
rect 106326 388584 106332 388596
rect 13372 388556 106332 388584
rect 13372 388544 13378 388556
rect 106326 388544 106332 388556
rect 106384 388544 106390 388596
rect 13682 388476 13688 388528
rect 13740 388516 13746 388528
rect 185354 388516 185360 388528
rect 13740 388488 185360 388516
rect 13740 388476 13746 388488
rect 185354 388476 185360 388488
rect 185412 388476 185418 388528
rect 190322 388476 190328 388528
rect 190380 388516 190386 388528
rect 223074 388516 223080 388528
rect 190380 388488 223080 388516
rect 190380 388476 190386 388488
rect 223074 388476 223080 388488
rect 223132 388476 223138 388528
rect 304586 388476 304592 388528
rect 304644 388516 304650 388528
rect 322526 388516 322532 388528
rect 304644 388488 322532 388516
rect 304644 388476 304650 388488
rect 322526 388476 322532 388488
rect 322584 388476 322590 388528
rect 13590 388408 13596 388460
rect 13648 388448 13654 388460
rect 215346 388448 215352 388460
rect 13648 388420 215352 388448
rect 13648 388408 13654 388420
rect 215346 388408 215352 388420
rect 215404 388408 215410 388460
rect 220314 388408 220320 388460
rect 220372 388448 220378 388460
rect 362454 388448 362460 388460
rect 220372 388420 362460 388448
rect 220372 388408 220378 388420
rect 362454 388408 362460 388420
rect 362512 388408 362518 388460
rect 13406 388340 13412 388392
rect 13464 388380 13470 388392
rect 101266 388380 101272 388392
rect 13464 388352 101272 388380
rect 13464 388340 13470 388352
rect 101266 388340 101272 388352
rect 101324 388340 101330 388392
rect 309278 388340 309284 388392
rect 309336 388380 309342 388392
rect 315626 388380 315632 388392
rect 309336 388352 315632 388380
rect 309336 388340 309342 388352
rect 315626 388340 315632 388352
rect 315684 388340 315690 388392
rect 395117 385595 395175 385601
rect 395117 385561 395129 385595
rect 395163 385592 395175 385595
rect 395206 385592 395212 385604
rect 395163 385564 395212 385592
rect 395163 385561 395175 385564
rect 395117 385555 395175 385561
rect 395206 385552 395212 385564
rect 395264 385552 395270 385604
rect 315810 378616 315816 378668
rect 315868 378656 315874 378668
rect 429430 378656 429436 378668
rect 315868 378628 429436 378656
rect 315868 378616 315874 378628
rect 429430 378616 429436 378628
rect 429488 378616 429494 378668
rect 131810 371748 131816 371800
rect 131868 371788 131874 371800
rect 134754 371788 134760 371800
rect 131868 371760 134760 371788
rect 131868 371748 131874 371760
rect 134754 371748 134760 371760
rect 134812 371748 134818 371800
rect 225834 371748 225840 371800
rect 225892 371788 225898 371800
rect 265854 371788 265860 371800
rect 225892 371760 265860 371788
rect 225892 371748 225898 371760
rect 265854 371748 265860 371760
rect 265912 371748 265918 371800
rect 320134 371748 320140 371800
rect 320192 371788 320198 371800
rect 323814 371788 323820 371800
rect 320192 371760 323820 371788
rect 320192 371748 320198 371760
rect 323814 371748 323820 371760
rect 323872 371748 323878 371800
rect 189034 368552 189040 368604
rect 189092 368592 189098 368604
rect 190690 368592 190696 368604
rect 189092 368564 190696 368592
rect 189092 368552 189098 368564
rect 190690 368552 190696 368564
rect 190748 368552 190754 368604
rect 208998 368552 209004 368604
rect 209056 368592 209062 368604
rect 210010 368592 210016 368604
rect 209056 368564 210016 368592
rect 209056 368552 209062 368564
rect 210010 368552 210016 368564
rect 210068 368552 210074 368604
rect 219026 368552 219032 368604
rect 219084 368592 219090 368604
rect 220314 368592 220320 368604
rect 219084 368564 220320 368592
rect 219084 368552 219090 368564
rect 220314 368552 220320 368564
rect 220372 368552 220378 368604
rect 277538 368280 277544 368332
rect 277596 368320 277602 368332
rect 280390 368320 280396 368332
rect 277596 368292 280396 368320
rect 277596 368280 277602 368292
rect 280390 368280 280396 368292
rect 280448 368280 280454 368332
rect 89858 367668 89864 367720
rect 89916 367708 89922 367720
rect 92526 367708 92532 367720
rect 89916 367680 92532 367708
rect 89916 367668 89922 367680
rect 92526 367668 92532 367680
rect 92584 367668 92590 367720
rect 90042 367600 90048 367652
rect 90100 367640 90106 367652
rect 91330 367640 91336 367652
rect 90100 367612 91336 367640
rect 90100 367600 90106 367612
rect 91330 367600 91336 367612
rect 91388 367600 91394 367652
rect 99978 367600 99984 367652
rect 100036 367640 100042 367652
rect 100898 367640 100904 367652
rect 100036 367612 100904 367640
rect 100036 367600 100042 367612
rect 100898 367600 100904 367612
rect 100956 367600 100962 367652
rect 110006 367600 110012 367652
rect 110064 367640 110070 367652
rect 112030 367640 112036 367652
rect 110064 367612 112036 367640
rect 110064 367600 110070 367612
rect 112030 367600 112036 367612
rect 112088 367600 112094 367652
rect 114974 367600 114980 367652
rect 115032 367640 115038 367652
rect 116170 367640 116176 367652
rect 115032 367612 116176 367640
rect 115032 367600 115038 367612
rect 116170 367600 116176 367612
rect 116228 367600 116234 367652
rect 125002 367600 125008 367652
rect 125060 367640 125066 367652
rect 126474 367640 126480 367652
rect 125060 367612 126480 367640
rect 125060 367600 125066 367612
rect 126474 367600 126480 367612
rect 126532 367600 126538 367652
rect 184066 367600 184072 367652
rect 184124 367640 184130 367652
rect 185078 367640 185084 367652
rect 184124 367612 185084 367640
rect 184124 367600 184130 367612
rect 185078 367600 185084 367612
rect 185136 367600 185142 367652
rect 185262 367600 185268 367652
rect 185320 367640 185326 367652
rect 186550 367640 186556 367652
rect 185320 367612 186556 367640
rect 185320 367600 185326 367612
rect 186550 367600 186556 367612
rect 186608 367600 186614 367652
rect 199062 367600 199068 367652
rect 199120 367640 199126 367652
rect 200258 367640 200264 367652
rect 199120 367612 200264 367640
rect 199120 367600 199126 367612
rect 200258 367600 200264 367612
rect 200316 367600 200322 367652
rect 204030 367600 204036 367652
rect 204088 367640 204094 367652
rect 205870 367640 205876 367652
rect 204088 367612 205876 367640
rect 204088 367600 204094 367612
rect 205870 367600 205876 367612
rect 205928 367600 205934 367652
rect 278366 367600 278372 367652
rect 278424 367640 278430 367652
rect 280482 367640 280488 367652
rect 278424 367612 280488 367640
rect 278424 367600 278430 367612
rect 280482 367600 280488 367612
rect 280540 367600 280546 367652
rect 293362 367600 293368 367652
rect 293420 367640 293426 367652
rect 294282 367640 294288 367652
rect 293420 367612 294288 367640
rect 293420 367600 293426 367612
rect 294282 367600 294288 367612
rect 294340 367600 294346 367652
rect 298238 367600 298244 367652
rect 298296 367640 298302 367652
rect 299710 367640 299716 367652
rect 298296 367612 299716 367640
rect 298296 367600 298302 367612
rect 299710 367600 299716 367612
rect 299768 367600 299774 367652
rect 303298 367600 303304 367652
rect 303356 367640 303362 367652
rect 305230 367640 305236 367652
rect 303356 367612 305236 367640
rect 303356 367600 303362 367612
rect 305230 367600 305236 367612
rect 305288 367600 305294 367652
rect 308358 367600 308364 367652
rect 308416 367640 308422 367652
rect 309278 367640 309284 367652
rect 308416 367612 309284 367640
rect 308416 367600 308422 367612
rect 309278 367600 309284 367612
rect 309336 367600 309342 367652
rect 223074 367532 223080 367584
rect 223132 367572 223138 367584
rect 429430 367572 429436 367584
rect 223132 367544 429436 367572
rect 223132 367532 223138 367544
rect 429430 367532 429436 367544
rect 429488 367532 429494 367584
rect 395298 366348 395304 366360
rect 395259 366320 395304 366348
rect 395298 366308 395304 366320
rect 395356 366308 395362 366360
rect 395206 364948 395212 365000
rect 395264 364988 395270 365000
rect 395301 364991 395359 364997
rect 395301 364988 395313 364991
rect 395264 364960 395313 364988
rect 395264 364948 395270 364960
rect 395301 364957 395313 364960
rect 395347 364957 395359 364991
rect 395301 364951 395359 364957
rect 91330 363452 91336 363504
rect 91388 363492 91394 363504
rect 92066 363492 92072 363504
rect 91388 363464 92072 363492
rect 91388 363452 91394 363464
rect 92066 363452 92072 363464
rect 92124 363452 92130 363504
rect 116170 363452 116176 363504
rect 116228 363492 116234 363504
rect 116814 363492 116820 363504
rect 116228 363464 116820 363492
rect 116228 363452 116234 363464
rect 116814 363452 116820 363464
rect 116872 363452 116878 363504
rect 210010 363452 210016 363504
rect 210068 363492 210074 363504
rect 210838 363492 210844 363504
rect 210068 363464 210844 363492
rect 210068 363452 210074 363464
rect 210838 363452 210844 363464
rect 210896 363452 210902 363504
rect 395298 363492 395304 363504
rect 395259 363464 395304 363492
rect 395298 363452 395304 363464
rect 395356 363452 395362 363504
rect 53702 359780 53708 359832
rect 53760 359820 53766 359832
rect 76978 359820 76984 359832
rect 53760 359792 76984 359820
rect 53760 359780 53766 359792
rect 76978 359780 76984 359792
rect 77036 359780 77042 359832
rect 50206 359712 50212 359764
rect 50264 359752 50270 359764
rect 76794 359752 76800 359764
rect 50264 359724 76800 359752
rect 50264 359712 50270 359724
rect 76794 359712 76800 359724
rect 76852 359712 76858 359764
rect 64190 359644 64196 359696
rect 64248 359684 64254 359696
rect 76058 359684 76064 359696
rect 64248 359656 76064 359684
rect 64248 359644 64254 359656
rect 76058 359644 76064 359656
rect 76116 359644 76122 359696
rect 60694 359576 60700 359628
rect 60752 359616 60758 359628
rect 75874 359616 75880 359628
rect 60752 359588 75880 359616
rect 60752 359576 60758 359588
rect 75874 359576 75880 359588
rect 75932 359576 75938 359628
rect 57198 359508 57204 359560
rect 57256 359548 57262 359560
rect 75782 359548 75788 359560
rect 57256 359520 75788 359548
rect 57256 359508 57262 359520
rect 75782 359508 75788 359520
rect 75840 359508 75846 359560
rect 67686 359372 67692 359424
rect 67744 359412 67750 359424
rect 75966 359412 75972 359424
rect 67744 359384 75972 359412
rect 67744 359372 67750 359384
rect 75966 359372 75972 359384
rect 76024 359372 76030 359424
rect 80198 357876 80204 357928
rect 80256 357916 80262 357928
rect 127210 357916 127216 357928
rect 80256 357888 127216 357916
rect 80256 357876 80262 357888
rect 127210 357876 127216 357888
rect 127268 357916 127274 357928
rect 139630 357916 139636 357928
rect 127268 357888 139636 357916
rect 127268 357876 127274 357888
rect 139630 357876 139636 357888
rect 139688 357876 139694 357928
rect 174038 357876 174044 357928
rect 174096 357916 174102 357928
rect 221050 357916 221056 357928
rect 174096 357888 221056 357916
rect 174096 357876 174102 357888
rect 221050 357876 221056 357888
rect 221108 357916 221114 357928
rect 233470 357916 233476 357928
rect 221108 357888 233476 357916
rect 221108 357876 221114 357888
rect 233470 357876 233476 357888
rect 233528 357876 233534 357928
rect 266590 357876 266596 357928
rect 266648 357916 266654 357928
rect 314890 357916 314896 357928
rect 266648 357888 314896 357916
rect 266648 357876 266654 357888
rect 314890 357876 314896 357888
rect 314948 357916 314954 357928
rect 328414 357916 328420 357928
rect 314948 357888 328420 357916
rect 314948 357876 314954 357888
rect 328414 357876 328420 357888
rect 328472 357876 328478 357928
rect 75874 357604 75880 357656
rect 75932 357644 75938 357656
rect 76150 357644 76156 357656
rect 75932 357616 76156 357644
rect 75932 357604 75938 357616
rect 76150 357604 76156 357616
rect 76208 357604 76214 357656
rect 75782 357536 75788 357588
rect 75840 357576 75846 357588
rect 76245 357579 76303 357585
rect 76245 357576 76257 357579
rect 75840 357548 76257 357576
rect 75840 357536 75846 357548
rect 76245 357545 76257 357548
rect 76291 357545 76303 357579
rect 76245 357539 76303 357545
rect 71458 357468 71464 357520
rect 71516 357508 71522 357520
rect 75874 357508 75880 357520
rect 71516 357480 75880 357508
rect 71516 357468 71522 357480
rect 75874 357468 75880 357480
rect 75932 357468 75938 357520
rect 74770 357400 74776 357452
rect 74828 357440 74834 357452
rect 76886 357440 76892 357452
rect 74828 357412 76892 357440
rect 74828 357400 74834 357412
rect 76886 357400 76892 357412
rect 76944 357400 76950 357452
rect 80198 356516 80204 356568
rect 80256 356556 80262 356568
rect 121690 356556 121696 356568
rect 80256 356528 121696 356556
rect 80256 356516 80262 356528
rect 121690 356516 121696 356528
rect 121748 356556 121754 356568
rect 139630 356556 139636 356568
rect 121748 356528 139636 356556
rect 121748 356516 121754 356528
rect 139630 356516 139636 356528
rect 139688 356516 139694 356568
rect 173486 356516 173492 356568
rect 173544 356556 173550 356568
rect 215530 356556 215536 356568
rect 173544 356528 215536 356556
rect 173544 356516 173550 356528
rect 215530 356516 215536 356528
rect 215588 356556 215594 356568
rect 233470 356556 233476 356568
rect 215588 356528 233476 356556
rect 215588 356516 215594 356528
rect 233470 356516 233476 356528
rect 233528 356516 233534 356568
rect 266590 356516 266596 356568
rect 266648 356556 266654 356568
rect 309370 356556 309376 356568
rect 266648 356528 309376 356556
rect 266648 356516 266654 356528
rect 309370 356516 309376 356528
rect 309428 356556 309434 356568
rect 328322 356556 328328 356568
rect 309428 356528 328328 356556
rect 309428 356516 309434 356528
rect 328322 356516 328328 356528
rect 328380 356516 328386 356568
rect 80198 355156 80204 355208
rect 80256 355196 80262 355208
rect 117550 355196 117556 355208
rect 80256 355168 117556 355196
rect 80256 355156 80262 355168
rect 117550 355156 117556 355168
rect 117608 355196 117614 355208
rect 118010 355196 118016 355208
rect 117608 355168 118016 355196
rect 117608 355156 117614 355168
rect 118010 355156 118016 355168
rect 118068 355156 118074 355208
rect 120218 355156 120224 355208
rect 120276 355196 120282 355208
rect 122058 355196 122064 355208
rect 120276 355168 122064 355196
rect 120276 355156 120282 355168
rect 122058 355156 122064 355168
rect 122116 355156 122122 355208
rect 122153 355199 122211 355205
rect 122153 355165 122165 355199
rect 122199 355196 122211 355199
rect 139630 355196 139636 355208
rect 122199 355168 139636 355196
rect 122199 355165 122211 355168
rect 122153 355159 122211 355165
rect 139630 355156 139636 355168
rect 139688 355156 139694 355208
rect 174038 355156 174044 355208
rect 174096 355196 174102 355208
rect 211390 355196 211396 355208
rect 174096 355168 211396 355196
rect 174096 355156 174102 355168
rect 211390 355156 211396 355168
rect 211448 355196 211454 355208
rect 212678 355196 212684 355208
rect 211448 355168 212684 355196
rect 211448 355156 211454 355168
rect 212678 355156 212684 355168
rect 212736 355156 212742 355208
rect 214058 355156 214064 355208
rect 214116 355196 214122 355208
rect 216358 355196 216364 355208
rect 214116 355168 216364 355196
rect 214116 355156 214122 355168
rect 216358 355156 216364 355168
rect 216416 355156 216422 355208
rect 216453 355199 216511 355205
rect 216453 355165 216465 355199
rect 216499 355196 216511 355199
rect 233470 355196 233476 355208
rect 216499 355168 233476 355196
rect 216499 355165 216511 355168
rect 216453 355159 216511 355165
rect 233470 355156 233476 355168
rect 233528 355156 233534 355208
rect 266590 355156 266596 355208
rect 266648 355196 266654 355208
rect 305322 355196 305328 355208
rect 266648 355168 305328 355196
rect 266648 355156 266654 355168
rect 305322 355156 305328 355168
rect 305380 355196 305386 355208
rect 328414 355196 328420 355208
rect 305380 355168 328420 355196
rect 305380 355156 305386 355168
rect 328414 355156 328420 355168
rect 328472 355156 328478 355208
rect 79278 355088 79284 355140
rect 79336 355128 79342 355140
rect 104949 355131 105007 355137
rect 104949 355128 104961 355131
rect 79336 355100 104961 355128
rect 79336 355088 79342 355100
rect 104949 355097 104961 355100
rect 104995 355097 105007 355131
rect 104949 355091 105007 355097
rect 105038 355088 105044 355140
rect 105096 355128 105102 355140
rect 107062 355128 107068 355140
rect 105096 355100 107068 355128
rect 105096 355088 105102 355100
rect 107062 355088 107068 355100
rect 107120 355088 107126 355140
rect 139722 355128 139728 355140
rect 112324 355100 139728 355128
rect 95378 355020 95384 355072
rect 95436 355060 95442 355072
rect 97034 355060 97040 355072
rect 95436 355032 97040 355060
rect 95436 355020 95442 355032
rect 97034 355020 97040 355032
rect 97092 355020 97098 355072
rect 100898 355020 100904 355072
rect 100956 355060 100962 355072
rect 102370 355060 102376 355072
rect 100956 355032 102376 355060
rect 100956 355020 100962 355032
rect 102370 355020 102376 355032
rect 102428 355020 102434 355072
rect 104949 354927 105007 354933
rect 104949 354893 104961 354927
rect 104995 354924 105007 354927
rect 112122 354924 112128 354936
rect 104995 354896 112128 354924
rect 104995 354893 105007 354896
rect 104949 354887 105007 354893
rect 112122 354884 112128 354896
rect 112180 354924 112186 354936
rect 112324 354924 112352 355100
rect 139722 355088 139728 355100
rect 139780 355088 139786 355140
rect 173762 355088 173768 355140
rect 173820 355128 173826 355140
rect 205962 355128 205968 355140
rect 173820 355100 205968 355128
rect 173820 355088 173826 355100
rect 205962 355088 205968 355100
rect 206020 355128 206026 355140
rect 233562 355128 233568 355140
rect 206020 355100 233568 355128
rect 206020 355088 206026 355100
rect 233562 355088 233568 355100
rect 233620 355088 233626 355140
rect 266682 355088 266688 355140
rect 266740 355128 266746 355140
rect 299802 355128 299808 355140
rect 266740 355100 299808 355128
rect 266740 355088 266746 355100
rect 299802 355088 299808 355100
rect 299860 355128 299866 355140
rect 328506 355128 328512 355140
rect 299860 355100 328512 355128
rect 299860 355088 299866 355100
rect 328506 355088 328512 355100
rect 328564 355088 328570 355140
rect 126474 355020 126480 355072
rect 126532 355060 126538 355072
rect 127210 355060 127216 355072
rect 126532 355032 127216 355060
rect 126532 355020 126538 355032
rect 127210 355020 127216 355032
rect 127268 355020 127274 355072
rect 185078 355020 185084 355072
rect 185136 355060 185142 355072
rect 186366 355060 186372 355072
rect 185136 355032 186372 355060
rect 185136 355020 185142 355032
rect 186366 355020 186372 355032
rect 186424 355020 186430 355072
rect 194738 355020 194744 355072
rect 194796 355060 194802 355072
rect 196302 355060 196308 355072
rect 194796 355032 196308 355060
rect 194796 355020 194802 355032
rect 196302 355020 196308 355032
rect 196360 355020 196366 355072
rect 220314 355020 220320 355072
rect 220372 355060 220378 355072
rect 221326 355060 221332 355072
rect 220372 355032 221332 355060
rect 220372 355020 220378 355032
rect 221326 355020 221332 355032
rect 221384 355020 221390 355072
rect 283058 355020 283064 355072
rect 283116 355060 283122 355072
rect 285358 355060 285364 355072
rect 283116 355032 285364 355060
rect 283116 355020 283122 355032
rect 285358 355020 285364 355032
rect 285416 355020 285422 355072
rect 288578 355020 288584 355072
rect 288636 355060 288642 355072
rect 290326 355060 290332 355072
rect 288636 355032 290332 355060
rect 288636 355020 288642 355032
rect 290326 355020 290332 355032
rect 290384 355020 290390 355072
rect 309278 355020 309284 355072
rect 309336 355060 309342 355072
rect 310382 355060 310388 355072
rect 309336 355032 310388 355060
rect 309336 355020 309342 355032
rect 310382 355020 310388 355032
rect 310440 355020 310446 355072
rect 313418 355020 313424 355072
rect 313476 355060 313482 355072
rect 315350 355060 315356 355072
rect 313476 355032 315356 355060
rect 313476 355020 313482 355032
rect 315350 355020 315356 355032
rect 315408 355020 315414 355072
rect 118010 354952 118016 355004
rect 118068 354992 118074 355004
rect 122153 354995 122211 355001
rect 122153 354992 122165 354995
rect 118068 354964 122165 354992
rect 118068 354952 118074 354964
rect 122153 354961 122165 354964
rect 122199 354961 122211 354995
rect 122153 354955 122211 354961
rect 212678 354952 212684 355004
rect 212736 354992 212742 355004
rect 216453 354995 216511 355001
rect 216453 354992 216465 354995
rect 212736 354964 216465 354992
rect 212736 354952 212742 354964
rect 216453 354961 216465 354964
rect 216499 354961 216511 354995
rect 216453 354955 216511 354961
rect 112180 354896 112352 354924
rect 112180 354884 112186 354896
rect 200258 354000 200264 354052
rect 200316 354040 200322 354052
rect 201362 354040 201368 354052
rect 200316 354012 201368 354040
rect 200316 354000 200322 354012
rect 201362 354000 201368 354012
rect 201420 354000 201426 354052
rect 76242 353904 76248 353916
rect 76203 353876 76248 353904
rect 76242 353864 76248 353876
rect 76300 353864 76306 353916
rect 196210 353864 196216 353916
rect 196268 353904 196274 353916
rect 196486 353904 196492 353916
rect 196268 353876 196492 353904
rect 196268 353864 196274 353876
rect 196486 353864 196492 353876
rect 196544 353864 196550 353916
rect 390698 353864 390704 353916
rect 390756 353904 390762 353916
rect 429430 353904 429436 353916
rect 390756 353876 429436 353904
rect 390756 353864 390762 353876
rect 429430 353864 429436 353876
rect 429488 353864 429494 353916
rect 80198 353796 80204 353848
rect 80256 353836 80262 353848
rect 106510 353836 106516 353848
rect 80256 353808 106516 353836
rect 80256 353796 80262 353808
rect 106510 353796 106516 353808
rect 106568 353836 106574 353848
rect 139630 353836 139636 353848
rect 106568 353808 139636 353836
rect 106568 353796 106574 353808
rect 139630 353796 139636 353808
rect 139688 353796 139694 353848
rect 174038 353796 174044 353848
rect 174096 353836 174102 353848
rect 200350 353836 200356 353848
rect 174096 353808 200356 353836
rect 174096 353796 174102 353808
rect 200350 353796 200356 353808
rect 200408 353836 200414 353848
rect 233470 353836 233476 353848
rect 200408 353808 233476 353836
rect 200408 353796 200414 353808
rect 233470 353796 233476 353808
rect 233528 353796 233534 353848
rect 266590 353796 266596 353848
rect 266648 353836 266654 353848
rect 294190 353836 294196 353848
rect 266648 353808 294196 353836
rect 266648 353796 266654 353808
rect 294190 353796 294196 353808
rect 294248 353836 294254 353848
rect 328046 353836 328052 353848
rect 294248 353808 328052 353836
rect 294248 353796 294254 353808
rect 328046 353796 328052 353808
rect 328104 353796 328110 353848
rect 80198 352368 80204 352420
rect 80256 352408 80262 352420
rect 102646 352408 102652 352420
rect 80256 352380 102652 352408
rect 80256 352368 80262 352380
rect 102646 352368 102652 352380
rect 102704 352408 102710 352420
rect 139630 352408 139636 352420
rect 102704 352380 139636 352408
rect 102704 352368 102710 352380
rect 139630 352368 139636 352380
rect 139688 352368 139694 352420
rect 174038 352368 174044 352420
rect 174096 352408 174102 352420
rect 196210 352408 196216 352420
rect 174096 352380 196216 352408
rect 174096 352368 174102 352380
rect 196210 352368 196216 352380
rect 196268 352408 196274 352420
rect 233470 352408 233476 352420
rect 196268 352380 233476 352408
rect 196268 352368 196274 352380
rect 233470 352368 233476 352380
rect 233528 352368 233534 352420
rect 266590 352368 266596 352420
rect 266648 352408 266654 352420
rect 290050 352408 290056 352420
rect 266648 352380 290056 352408
rect 266648 352368 266654 352380
rect 290050 352368 290056 352380
rect 290108 352408 290114 352420
rect 328506 352408 328512 352420
rect 290108 352380 328512 352408
rect 290108 352368 290114 352380
rect 328506 352368 328512 352380
rect 328564 352368 328570 352420
rect 191242 351864 191248 351876
rect 191203 351836 191248 351864
rect 191242 351824 191248 351836
rect 191300 351824 191306 351876
rect 284530 351592 284536 351604
rect 284491 351564 284536 351592
rect 284530 351552 284536 351564
rect 284588 351552 284594 351604
rect 96758 351524 96764 351536
rect 96719 351496 96764 351524
rect 96758 351484 96764 351496
rect 96816 351484 96822 351536
rect 226294 351280 226300 351332
rect 226352 351320 226358 351332
rect 231630 351320 231636 351332
rect 226352 351292 231636 351320
rect 226352 351280 226358 351292
rect 231630 351280 231636 351292
rect 231688 351280 231694 351332
rect 131810 351076 131816 351128
rect 131868 351116 131874 351128
rect 139446 351116 139452 351128
rect 131868 351088 139452 351116
rect 131868 351076 131874 351088
rect 139446 351076 139452 351088
rect 139504 351076 139510 351128
rect 272018 351076 272024 351128
rect 272076 351116 272082 351128
rect 274870 351116 274876 351128
rect 272076 351088 274876 351116
rect 272076 351076 272082 351088
rect 274870 351076 274876 351088
rect 274928 351076 274934 351128
rect 320594 351076 320600 351128
rect 320652 351116 320658 351128
rect 328138 351116 328144 351128
rect 320652 351088 328144 351116
rect 320652 351076 320658 351088
rect 328138 351076 328144 351088
rect 328196 351076 328202 351128
rect 79830 351008 79836 351060
rect 79888 351048 79894 351060
rect 89858 351048 89864 351060
rect 79888 351020 89864 351048
rect 79888 351008 79894 351020
rect 89858 351008 89864 351020
rect 89916 351048 89922 351060
rect 139630 351048 139636 351060
rect 89916 351020 139636 351048
rect 89916 351008 89922 351020
rect 139630 351008 139636 351020
rect 139688 351008 139694 351060
rect 173854 351008 173860 351060
rect 173912 351048 173918 351060
rect 185262 351048 185268 351060
rect 173912 351020 185268 351048
rect 173912 351008 173918 351020
rect 185262 351008 185268 351020
rect 185320 351048 185326 351060
rect 233562 351048 233568 351060
rect 185320 351020 233568 351048
rect 185320 351008 185326 351020
rect 233562 351008 233568 351020
rect 233620 351008 233626 351060
rect 266682 351008 266688 351060
rect 266740 351048 266746 351060
rect 277538 351048 277544 351060
rect 266740 351020 277544 351048
rect 266740 351008 266746 351020
rect 277538 351008 277544 351020
rect 277596 351048 277602 351060
rect 327862 351048 327868 351060
rect 277596 351020 327868 351048
rect 277596 351008 277602 351020
rect 327862 351008 327868 351020
rect 327920 351008 327926 351060
rect 80198 350328 80204 350380
rect 80256 350368 80262 350380
rect 96761 350371 96819 350377
rect 96761 350368 96773 350371
rect 80256 350340 96773 350368
rect 80256 350328 80262 350340
rect 96761 350337 96773 350340
rect 96807 350368 96819 350371
rect 139722 350368 139728 350380
rect 96807 350340 139728 350368
rect 96807 350337 96819 350340
rect 96761 350331 96819 350337
rect 139722 350328 139728 350340
rect 139780 350328 139786 350380
rect 173670 350328 173676 350380
rect 173728 350368 173734 350380
rect 191245 350371 191303 350377
rect 191245 350368 191257 350371
rect 173728 350340 191257 350368
rect 173728 350328 173734 350340
rect 191245 350337 191257 350340
rect 191291 350368 191303 350371
rect 233470 350368 233476 350380
rect 191291 350340 233476 350368
rect 191291 350337 191303 350340
rect 191245 350331 191303 350337
rect 233470 350328 233476 350340
rect 233528 350328 233534 350380
rect 266590 350328 266596 350380
rect 266648 350368 266654 350380
rect 284533 350371 284591 350377
rect 284533 350368 284545 350371
rect 266648 350340 284545 350368
rect 266648 350328 266654 350340
rect 284533 350337 284545 350340
rect 284579 350368 284591 350371
rect 327494 350368 327500 350380
rect 284579 350340 327500 350368
rect 284579 350337 284591 350340
rect 284533 350331 284591 350337
rect 327494 350328 327500 350340
rect 327552 350328 327558 350380
rect 131810 349716 131816 349768
rect 131868 349756 131874 349768
rect 139538 349756 139544 349768
rect 131868 349728 139544 349756
rect 131868 349716 131874 349728
rect 139538 349716 139544 349728
rect 139596 349716 139602 349768
rect 271926 349716 271932 349768
rect 271984 349756 271990 349768
rect 274870 349756 274876 349768
rect 271984 349728 274876 349756
rect 271984 349716 271990 349728
rect 274870 349716 274876 349728
rect 274928 349716 274934 349768
rect 321606 349716 321612 349768
rect 321664 349756 321670 349768
rect 328322 349756 328328 349768
rect 321664 349728 328328 349756
rect 321664 349716 321670 349728
rect 328322 349716 328328 349728
rect 328380 349716 328386 349768
rect 75969 349691 76027 349697
rect 75969 349657 75981 349691
rect 76015 349688 76027 349691
rect 76058 349688 76064 349700
rect 76015 349660 76064 349688
rect 76015 349657 76027 349660
rect 75969 349651 76027 349657
rect 76058 349648 76064 349660
rect 76116 349648 76122 349700
rect 172842 349648 172848 349700
rect 172900 349688 172906 349700
rect 182318 349688 182324 349700
rect 172900 349660 182324 349688
rect 172900 349648 172906 349660
rect 182318 349648 182324 349660
rect 182376 349648 182382 349700
rect 231630 349648 231636 349700
rect 231688 349688 231694 349700
rect 233470 349688 233476 349700
rect 231688 349660 233476 349688
rect 231688 349648 231694 349660
rect 233470 349648 233476 349660
rect 233528 349648 233534 349700
rect 266590 349648 266596 349700
rect 266648 349688 266654 349700
rect 272018 349688 272024 349700
rect 266648 349660 272024 349688
rect 266648 349648 266654 349660
rect 272018 349648 272024 349660
rect 272076 349648 272082 349700
rect 78910 348900 78916 348952
rect 78968 348940 78974 348952
rect 87098 348940 87104 348952
rect 78968 348912 87104 348940
rect 78968 348900 78974 348912
rect 87098 348900 87104 348912
rect 87156 348900 87162 348952
rect 321698 348424 321704 348476
rect 321756 348464 321762 348476
rect 327218 348464 327224 348476
rect 321756 348436 327224 348464
rect 321756 348424 321762 348436
rect 327218 348424 327224 348436
rect 327276 348424 327282 348476
rect 131810 348356 131816 348408
rect 131868 348396 131874 348408
rect 137238 348396 137244 348408
rect 131868 348368 137244 348396
rect 131868 348356 131874 348368
rect 137238 348356 137244 348368
rect 137296 348356 137302 348408
rect 226478 348356 226484 348408
rect 226536 348396 226542 348408
rect 231998 348396 232004 348408
rect 226536 348368 232004 348396
rect 226536 348356 226542 348368
rect 231998 348356 232004 348368
rect 232056 348356 232062 348408
rect 131902 348288 131908 348340
rect 131960 348328 131966 348340
rect 137514 348328 137520 348340
rect 131960 348300 137520 348328
rect 131960 348288 131966 348300
rect 137514 348288 137520 348300
rect 137572 348288 137578 348340
rect 226386 348288 226392 348340
rect 226444 348328 226450 348340
rect 231630 348328 231636 348340
rect 226444 348300 231636 348328
rect 226444 348288 226450 348300
rect 231630 348288 231636 348300
rect 231688 348288 231694 348340
rect 321606 348288 321612 348340
rect 321664 348328 321670 348340
rect 327126 348328 327132 348340
rect 321664 348300 327132 348328
rect 321664 348288 321670 348300
rect 327126 348288 327132 348300
rect 327184 348288 327190 348340
rect 226570 348220 226576 348272
rect 226628 348260 226634 348272
rect 233470 348260 233476 348272
rect 226628 348232 233476 348260
rect 226628 348220 226634 348232
rect 233470 348220 233476 348232
rect 233528 348220 233534 348272
rect 266590 348220 266596 348272
rect 266648 348260 266654 348272
rect 271926 348260 271932 348272
rect 266648 348232 271932 348260
rect 266648 348220 266654 348232
rect 271926 348220 271932 348232
rect 271984 348220 271990 348272
rect 174038 347948 174044 348000
rect 174096 347988 174102 348000
rect 180754 347988 180760 348000
rect 174096 347960 180760 347988
rect 174096 347948 174102 347960
rect 180754 347948 180760 347960
rect 180812 347948 180818 348000
rect 78910 347336 78916 347388
rect 78968 347376 78974 347388
rect 87006 347376 87012 347388
rect 78968 347348 87012 347376
rect 78968 347336 78974 347348
rect 87006 347336 87012 347348
rect 87064 347336 87070 347388
rect 132178 346928 132184 346980
rect 132236 346968 132242 346980
rect 139722 346968 139728 346980
rect 132236 346940 139728 346968
rect 132236 346928 132242 346940
rect 139722 346928 139728 346940
rect 139780 346928 139786 346980
rect 226386 346928 226392 346980
rect 226444 346968 226450 346980
rect 228594 346968 228600 346980
rect 226444 346940 228600 346968
rect 226444 346928 226450 346940
rect 228594 346928 228600 346940
rect 228652 346928 228658 346980
rect 321054 346928 321060 346980
rect 321112 346968 321118 346980
rect 323170 346968 323176 346980
rect 321112 346940 323176 346968
rect 321112 346928 321118 346940
rect 323170 346928 323176 346940
rect 323228 346928 323234 346980
rect 137514 346860 137520 346912
rect 137572 346900 137578 346912
rect 139630 346900 139636 346912
rect 137572 346872 139636 346900
rect 137572 346860 137578 346872
rect 139630 346860 139636 346872
rect 139688 346860 139694 346912
rect 174038 346860 174044 346912
rect 174096 346900 174102 346912
rect 180938 346900 180944 346912
rect 174096 346872 180944 346900
rect 174096 346860 174102 346872
rect 180938 346860 180944 346872
rect 180996 346860 181002 346912
rect 231998 346860 232004 346912
rect 232056 346900 232062 346912
rect 233470 346900 233476 346912
rect 232056 346872 233476 346900
rect 232056 346860 232062 346872
rect 233470 346860 233476 346872
rect 233528 346860 233534 346912
rect 266590 346860 266596 346912
rect 266648 346900 266654 346912
rect 274870 346900 274876 346912
rect 266648 346872 274876 346900
rect 266648 346860 266654 346872
rect 274870 346860 274876 346872
rect 274928 346860 274934 346912
rect 137238 346792 137244 346844
rect 137296 346832 137302 346844
rect 139814 346832 139820 346844
rect 137296 346804 139820 346832
rect 137296 346792 137302 346804
rect 139814 346792 139820 346804
rect 139872 346792 139878 346844
rect 231630 346792 231636 346844
rect 231688 346832 231694 346844
rect 233562 346832 233568 346844
rect 231688 346804 233568 346832
rect 231688 346792 231694 346804
rect 233562 346792 233568 346804
rect 233620 346792 233626 346844
rect 266682 346792 266688 346844
rect 266740 346832 266746 346844
rect 274962 346832 274968 346844
rect 266740 346804 274968 346832
rect 266740 346792 266746 346804
rect 274962 346792 274968 346804
rect 275020 346792 275026 346844
rect 173118 346248 173124 346300
rect 173176 346288 173182 346300
rect 180846 346288 180852 346300
rect 173176 346260 180852 346288
rect 173176 346248 173182 346260
rect 180846 346248 180852 346260
rect 180904 346248 180910 346300
rect 78910 346180 78916 346232
rect 78968 346220 78974 346232
rect 87098 346220 87104 346232
rect 78968 346192 87104 346220
rect 78968 346180 78974 346192
rect 87098 346180 87104 346192
rect 87156 346180 87162 346232
rect 79002 345976 79008 346028
rect 79060 346016 79066 346028
rect 86914 346016 86920 346028
rect 79060 345988 86920 346016
rect 79060 345976 79066 345988
rect 86914 345976 86920 345988
rect 86972 345976 86978 346028
rect 131810 345636 131816 345688
rect 131868 345676 131874 345688
rect 134110 345676 134116 345688
rect 131868 345648 134116 345676
rect 131868 345636 131874 345648
rect 134110 345636 134116 345648
rect 134168 345636 134174 345688
rect 226478 345636 226484 345688
rect 226536 345676 226542 345688
rect 228042 345676 228048 345688
rect 226536 345648 228048 345676
rect 226536 345636 226542 345648
rect 228042 345636 228048 345648
rect 228100 345636 228106 345688
rect 320410 345636 320416 345688
rect 320468 345676 320474 345688
rect 323262 345676 323268 345688
rect 320468 345648 323268 345676
rect 320468 345636 320474 345648
rect 323262 345636 323268 345648
rect 323320 345636 323326 345688
rect 85810 345568 85816 345620
rect 85868 345608 85874 345620
rect 87926 345608 87932 345620
rect 85868 345580 87932 345608
rect 85868 345568 85874 345580
rect 87926 345568 87932 345580
rect 87984 345568 87990 345620
rect 131902 345568 131908 345620
rect 131960 345608 131966 345620
rect 139630 345608 139636 345620
rect 131960 345580 139636 345608
rect 131960 345568 131966 345580
rect 139630 345568 139636 345580
rect 139688 345568 139694 345620
rect 173026 345568 173032 345620
rect 173084 345608 173090 345620
rect 182318 345608 182324 345620
rect 173084 345580 182324 345608
rect 173084 345568 173090 345580
rect 182318 345568 182324 345580
rect 182376 345568 182382 345620
rect 226386 345568 226392 345620
rect 226444 345608 226450 345620
rect 234574 345608 234580 345620
rect 226444 345580 234580 345608
rect 226444 345568 226450 345580
rect 234574 345568 234580 345580
rect 234632 345568 234638 345620
rect 320502 345568 320508 345620
rect 320560 345608 320566 345620
rect 327034 345608 327040 345620
rect 320560 345580 327040 345608
rect 320560 345568 320566 345580
rect 327034 345568 327040 345580
rect 327092 345568 327098 345620
rect 395301 345611 395359 345617
rect 395301 345577 395313 345611
rect 395347 345608 395359 345611
rect 395390 345608 395396 345620
rect 395347 345580 395396 345608
rect 395347 345577 395359 345580
rect 395301 345571 395359 345577
rect 395390 345568 395396 345580
rect 395448 345568 395454 345620
rect 228594 345500 228600 345552
rect 228652 345540 228658 345552
rect 233470 345540 233476 345552
rect 228652 345512 233476 345540
rect 228652 345500 228658 345512
rect 233470 345500 233476 345512
rect 233528 345500 233534 345552
rect 266590 345500 266596 345552
rect 266648 345540 266654 345552
rect 275054 345540 275060 345552
rect 266648 345512 275060 345540
rect 266648 345500 266654 345512
rect 275054 345500 275060 345512
rect 275112 345500 275118 345552
rect 323170 345500 323176 345552
rect 323228 345540 323234 345552
rect 328046 345540 328052 345552
rect 323228 345512 328052 345540
rect 323228 345500 323234 345512
rect 328046 345500 328052 345512
rect 328104 345500 328110 345552
rect 173302 345160 173308 345212
rect 173360 345200 173366 345212
rect 180754 345200 180760 345212
rect 173360 345172 180760 345200
rect 173360 345160 173366 345172
rect 180754 345160 180760 345172
rect 180812 345160 180818 345212
rect 85902 344616 85908 344668
rect 85960 344656 85966 344668
rect 87466 344656 87472 344668
rect 85960 344628 87472 344656
rect 85960 344616 85966 344628
rect 87466 344616 87472 344628
rect 87524 344616 87530 344668
rect 226018 344616 226024 344668
rect 226076 344656 226082 344668
rect 228502 344656 228508 344668
rect 226076 344628 228508 344656
rect 226076 344616 226082 344628
rect 228502 344616 228508 344628
rect 228560 344616 228566 344668
rect 321054 344616 321060 344668
rect 321112 344656 321118 344668
rect 323170 344656 323176 344668
rect 321112 344628 323176 344656
rect 321112 344616 321118 344628
rect 323170 344616 323176 344628
rect 323228 344616 323234 344668
rect 78910 344412 78916 344464
rect 78968 344452 78974 344464
rect 87006 344452 87012 344464
rect 78968 344424 87012 344452
rect 78968 344412 78974 344424
rect 87006 344412 87012 344424
rect 87064 344412 87070 344464
rect 321606 344344 321612 344396
rect 321664 344384 321670 344396
rect 326850 344384 326856 344396
rect 321664 344356 326856 344384
rect 321664 344344 321670 344356
rect 326850 344344 326856 344356
rect 326908 344344 326914 344396
rect 131810 344208 131816 344260
rect 131868 344248 131874 344260
rect 138158 344248 138164 344260
rect 131868 344220 138164 344248
rect 131868 344208 131874 344220
rect 138158 344208 138164 344220
rect 138216 344208 138222 344260
rect 226386 344208 226392 344260
rect 226444 344248 226450 344260
rect 227950 344248 227956 344260
rect 226444 344220 227956 344248
rect 226444 344208 226450 344220
rect 227950 344208 227956 344220
rect 228008 344208 228014 344260
rect 132362 344140 132368 344192
rect 132420 344180 132426 344192
rect 139722 344180 139728 344192
rect 132420 344152 139728 344180
rect 132420 344140 132426 344152
rect 139722 344140 139728 344152
rect 139780 344140 139786 344192
rect 172934 344140 172940 344192
rect 172992 344180 172998 344192
rect 182318 344180 182324 344192
rect 172992 344152 182324 344180
rect 172992 344140 172998 344152
rect 182318 344140 182324 344152
rect 182376 344140 182382 344192
rect 228042 344072 228048 344124
rect 228100 344112 228106 344124
rect 233470 344112 233476 344124
rect 228100 344084 233476 344112
rect 228100 344072 228106 344084
rect 233470 344072 233476 344084
rect 233528 344072 233534 344124
rect 266590 344072 266596 344124
rect 266648 344112 266654 344124
rect 274962 344112 274968 344124
rect 266648 344084 274968 344112
rect 266648 344072 266654 344084
rect 274962 344072 274968 344084
rect 275020 344072 275026 344124
rect 323262 344072 323268 344124
rect 323320 344112 323326 344124
rect 328506 344112 328512 344124
rect 323320 344084 328512 344112
rect 323320 344072 323326 344084
rect 328506 344072 328512 344084
rect 328564 344072 328570 344124
rect 173670 343732 173676 343784
rect 173728 343772 173734 343784
rect 180846 343772 180852 343784
rect 173728 343744 180852 343772
rect 173728 343732 173734 343744
rect 180846 343732 180852 343744
rect 180904 343732 180910 343784
rect 78910 342916 78916 342968
rect 78968 342956 78974 342968
rect 85810 342956 85816 342968
rect 78968 342928 85816 342956
rect 78968 342916 78974 342928
rect 85810 342916 85816 342928
rect 85868 342916 85874 342968
rect 321606 342848 321612 342900
rect 321664 342888 321670 342900
rect 327126 342888 327132 342900
rect 321664 342860 327132 342888
rect 321664 342848 321670 342860
rect 327126 342848 327132 342860
rect 327184 342848 327190 342900
rect 131810 342780 131816 342832
rect 131868 342820 131874 342832
rect 139814 342820 139820 342832
rect 131868 342792 139820 342820
rect 131868 342780 131874 342792
rect 139814 342780 139820 342792
rect 139872 342780 139878 342832
rect 173670 342780 173676 342832
rect 173728 342820 173734 342832
rect 181398 342820 181404 342832
rect 173728 342792 181404 342820
rect 173728 342780 173734 342792
rect 181398 342780 181404 342792
rect 181456 342780 181462 342832
rect 226386 342780 226392 342832
rect 226444 342820 226450 342832
rect 233654 342820 233660 342832
rect 226444 342792 233660 342820
rect 226444 342780 226450 342792
rect 233654 342780 233660 342792
rect 233712 342780 233718 342832
rect 78910 342712 78916 342764
rect 78968 342752 78974 342764
rect 88110 342752 88116 342764
rect 78968 342724 88116 342752
rect 78968 342712 78974 342724
rect 88110 342712 88116 342724
rect 88168 342712 88174 342764
rect 134110 342712 134116 342764
rect 134168 342752 134174 342764
rect 139630 342752 139636 342764
rect 134168 342724 139636 342752
rect 134168 342712 134174 342724
rect 139630 342712 139636 342724
rect 139688 342712 139694 342764
rect 228502 342712 228508 342764
rect 228560 342752 228566 342764
rect 233470 342752 233476 342764
rect 228560 342724 233476 342752
rect 228560 342712 228566 342724
rect 233470 342712 233476 342724
rect 233528 342712 233534 342764
rect 266682 342712 266688 342764
rect 266740 342752 266746 342764
rect 274870 342752 274876 342764
rect 266740 342724 274876 342752
rect 266740 342712 266746 342724
rect 274870 342712 274876 342724
rect 274928 342712 274934 342764
rect 323170 342712 323176 342764
rect 323228 342752 323234 342764
rect 328046 342752 328052 342764
rect 323228 342724 328052 342752
rect 323228 342712 323234 342724
rect 328046 342712 328052 342724
rect 328104 342712 328110 342764
rect 266590 342644 266596 342696
rect 266648 342684 266654 342696
rect 275238 342684 275244 342696
rect 266648 342656 275244 342684
rect 266648 342644 266654 342656
rect 275238 342644 275244 342656
rect 275296 342644 275302 342696
rect 172750 342236 172756 342288
rect 172808 342276 172814 342288
rect 180938 342276 180944 342288
rect 172808 342248 180944 342276
rect 172808 342236 172814 342248
rect 180938 342236 180944 342248
rect 180996 342236 181002 342288
rect 78910 341488 78916 341540
rect 78968 341528 78974 341540
rect 85902 341528 85908 341540
rect 78968 341500 85908 341528
rect 78968 341488 78974 341500
rect 85902 341488 85908 341500
rect 85960 341488 85966 341540
rect 131902 341488 131908 341540
rect 131960 341528 131966 341540
rect 139722 341528 139728 341540
rect 131960 341500 139728 341528
rect 131960 341488 131966 341500
rect 139722 341488 139728 341500
rect 139780 341488 139786 341540
rect 226478 341488 226484 341540
rect 226536 341528 226542 341540
rect 233562 341528 233568 341540
rect 226536 341500 233568 341528
rect 226536 341488 226542 341500
rect 233562 341488 233568 341500
rect 233620 341488 233626 341540
rect 321606 341488 321612 341540
rect 321664 341528 321670 341540
rect 327034 341528 327040 341540
rect 321664 341500 327040 341528
rect 321664 341488 321670 341500
rect 327034 341488 327040 341500
rect 327092 341488 327098 341540
rect 131810 341420 131816 341472
rect 131868 341460 131874 341472
rect 139906 341460 139912 341472
rect 131868 341432 139912 341460
rect 131868 341420 131874 341432
rect 139906 341420 139912 341432
rect 139964 341420 139970 341472
rect 226386 341420 226392 341472
rect 226444 341460 226450 341472
rect 233746 341460 233752 341472
rect 226444 341432 233752 341460
rect 226444 341420 226450 341432
rect 233746 341420 233752 341432
rect 233804 341420 233810 341472
rect 321054 341420 321060 341472
rect 321112 341460 321118 341472
rect 327218 341460 327224 341472
rect 321112 341432 327224 341460
rect 321112 341420 321118 341432
rect 327218 341420 327224 341432
rect 327276 341420 327282 341472
rect 394838 341420 394844 341472
rect 394896 341460 394902 341472
rect 429430 341460 429436 341472
rect 394896 341432 429436 341460
rect 394896 341420 394902 341432
rect 429430 341420 429436 341432
rect 429488 341420 429494 341472
rect 78910 341352 78916 341404
rect 78968 341392 78974 341404
rect 88478 341392 88484 341404
rect 78968 341364 88484 341392
rect 78968 341352 78974 341364
rect 88478 341352 88484 341364
rect 88536 341352 88542 341404
rect 138158 341352 138164 341404
rect 138216 341392 138222 341404
rect 139630 341392 139636 341404
rect 138216 341364 139636 341392
rect 138216 341352 138222 341364
rect 139630 341352 139636 341364
rect 139688 341352 139694 341404
rect 227950 341352 227956 341404
rect 228008 341392 228014 341404
rect 233470 341392 233476 341404
rect 228008 341364 233476 341392
rect 228008 341352 228014 341364
rect 233470 341352 233476 341364
rect 233528 341352 233534 341404
rect 266590 341352 266596 341404
rect 266648 341392 266654 341404
rect 275054 341392 275060 341404
rect 266648 341364 275060 341392
rect 266648 341352 266654 341364
rect 275054 341352 275060 341364
rect 275112 341352 275118 341404
rect 76058 340060 76064 340112
rect 76116 340100 76122 340112
rect 76242 340100 76248 340112
rect 76116 340072 76248 340100
rect 76116 340060 76122 340072
rect 76242 340060 76248 340072
rect 76300 340060 76306 340112
rect 85718 340060 85724 340112
rect 85776 340100 85782 340112
rect 87558 340100 87564 340112
rect 85776 340072 87564 340100
rect 85776 340060 85782 340072
rect 87558 340060 87564 340072
rect 87616 340060 87622 340112
rect 131810 340060 131816 340112
rect 131868 340100 131874 340112
rect 137330 340100 137336 340112
rect 131868 340072 137336 340100
rect 131868 340060 131874 340072
rect 137330 340060 137336 340072
rect 137388 340060 137394 340112
rect 173486 340060 173492 340112
rect 173544 340100 173550 340112
rect 181398 340100 181404 340112
rect 173544 340072 181404 340100
rect 173544 340060 173550 340072
rect 181398 340060 181404 340072
rect 181456 340060 181462 340112
rect 226386 340060 226392 340112
rect 226444 340100 226450 340112
rect 231906 340100 231912 340112
rect 226444 340072 231912 340100
rect 226444 340060 226450 340072
rect 231906 340060 231912 340072
rect 231964 340060 231970 340112
rect 272018 340060 272024 340112
rect 272076 340100 272082 340112
rect 275054 340100 275060 340112
rect 272076 340072 275060 340100
rect 272076 340060 272082 340072
rect 275054 340060 275060 340072
rect 275112 340060 275118 340112
rect 320594 340060 320600 340112
rect 320652 340100 320658 340112
rect 326942 340100 326948 340112
rect 320652 340072 326948 340100
rect 320652 340060 320658 340072
rect 326942 340060 326948 340072
rect 327000 340060 327006 340112
rect 78910 339992 78916 340044
rect 78968 340032 78974 340044
rect 87374 340032 87380 340044
rect 78968 340004 87380 340032
rect 78968 339992 78974 340004
rect 87374 339992 87380 340004
rect 87432 339992 87438 340044
rect 266590 339992 266596 340044
rect 266648 340032 266654 340044
rect 274962 340032 274968 340044
rect 266648 340004 274968 340032
rect 266648 339992 266654 340004
rect 274962 339992 274968 340004
rect 275020 339992 275026 340044
rect 226478 338768 226484 338820
rect 226536 338808 226542 338820
rect 233654 338808 233660 338820
rect 226536 338780 233660 338808
rect 226536 338768 226542 338780
rect 233654 338768 233660 338780
rect 233712 338768 233718 338820
rect 321606 338768 321612 338820
rect 321664 338808 321670 338820
rect 326666 338808 326672 338820
rect 321664 338780 326672 338808
rect 321664 338768 321670 338780
rect 326666 338768 326672 338780
rect 326724 338768 326730 338820
rect 131810 338700 131816 338752
rect 131868 338740 131874 338752
rect 136134 338740 136140 338752
rect 131868 338712 136140 338740
rect 131868 338700 131874 338712
rect 136134 338700 136140 338712
rect 136192 338700 136198 338752
rect 173302 338700 173308 338752
rect 173360 338740 173366 338752
rect 181582 338740 181588 338752
rect 173360 338712 181588 338740
rect 173360 338700 173366 338712
rect 181582 338700 181588 338712
rect 181640 338700 181646 338752
rect 84982 338632 84988 338684
rect 85040 338672 85046 338684
rect 87374 338672 87380 338684
rect 85040 338644 87380 338672
rect 85040 338632 85046 338644
rect 87374 338632 87380 338644
rect 87432 338632 87438 338684
rect 131902 338632 131908 338684
rect 131960 338672 131966 338684
rect 139630 338672 139636 338684
rect 131960 338644 139636 338672
rect 131960 338632 131966 338644
rect 139630 338632 139636 338644
rect 139688 338632 139694 338684
rect 173394 338632 173400 338684
rect 173452 338672 173458 338684
rect 182318 338672 182324 338684
rect 173452 338644 182324 338672
rect 173452 338632 173458 338644
rect 182318 338632 182324 338644
rect 182376 338632 182382 338684
rect 225926 338632 225932 338684
rect 225984 338672 225990 338684
rect 230802 338672 230808 338684
rect 225984 338644 230808 338672
rect 225984 338632 225990 338644
rect 230802 338632 230808 338644
rect 230860 338632 230866 338684
rect 321238 338632 321244 338684
rect 321296 338672 321302 338684
rect 327126 338672 327132 338684
rect 321296 338644 327132 338672
rect 321296 338632 321302 338644
rect 327126 338632 327132 338644
rect 327184 338632 327190 338684
rect 80198 338564 80204 338616
rect 80256 338604 80262 338616
rect 87466 338604 87472 338616
rect 80256 338576 87472 338604
rect 80256 338564 80262 338576
rect 87466 338564 87472 338576
rect 87524 338564 87530 338616
rect 173946 338564 173952 338616
rect 174004 338604 174010 338616
rect 181766 338604 181772 338616
rect 174004 338576 181772 338604
rect 174004 338564 174010 338576
rect 181766 338564 181772 338576
rect 181824 338564 181830 338616
rect 266682 338564 266688 338616
rect 266740 338604 266746 338616
rect 274870 338604 274876 338616
rect 266740 338576 274876 338604
rect 266740 338564 266746 338576
rect 274870 338564 274876 338576
rect 274928 338564 274934 338616
rect 78910 338496 78916 338548
rect 78968 338536 78974 338548
rect 87282 338536 87288 338548
rect 78968 338508 87288 338536
rect 78968 338496 78974 338508
rect 87282 338496 87288 338508
rect 87340 338496 87346 338548
rect 174038 338496 174044 338548
rect 174096 338536 174102 338548
rect 182134 338536 182140 338548
rect 174096 338508 182140 338536
rect 174096 338496 174102 338508
rect 182134 338496 182140 338508
rect 182192 338496 182198 338548
rect 266590 338496 266596 338548
rect 266648 338536 266654 338548
rect 275146 338536 275152 338548
rect 266648 338508 275152 338536
rect 266648 338496 266654 338508
rect 275146 338496 275152 338508
rect 275204 338496 275210 338548
rect 131810 337272 131816 337324
rect 131868 337312 131874 337324
rect 136226 337312 136232 337324
rect 131868 337284 136232 337312
rect 131868 337272 131874 337284
rect 136226 337272 136232 337284
rect 136284 337272 136290 337324
rect 225926 337272 225932 337324
rect 225984 337312 225990 337324
rect 230710 337312 230716 337324
rect 225984 337284 230716 337312
rect 225984 337272 225990 337284
rect 230710 337272 230716 337284
rect 230768 337272 230774 337324
rect 271466 337272 271472 337324
rect 271524 337312 271530 337324
rect 274870 337312 274876 337324
rect 271524 337284 274876 337312
rect 271524 337272 271530 337284
rect 274870 337272 274876 337284
rect 274928 337272 274934 337324
rect 321606 337272 321612 337324
rect 321664 337312 321670 337324
rect 327034 337312 327040 337324
rect 321664 337284 327040 337312
rect 321664 337272 321670 337284
rect 327034 337272 327040 337284
rect 327092 337272 327098 337324
rect 137330 337204 137336 337256
rect 137388 337244 137394 337256
rect 139722 337244 139728 337256
rect 137388 337216 139728 337244
rect 137388 337204 137394 337216
rect 139722 337204 139728 337216
rect 139780 337204 139786 337256
rect 231906 337204 231912 337256
rect 231964 337244 231970 337256
rect 233470 337244 233476 337256
rect 231964 337216 233476 337244
rect 231964 337204 231970 337216
rect 233470 337204 233476 337216
rect 233528 337204 233534 337256
rect 266590 337204 266596 337256
rect 266648 337244 266654 337256
rect 272018 337244 272024 337256
rect 266648 337216 272024 337244
rect 266648 337204 266654 337216
rect 272018 337204 272024 337216
rect 272076 337204 272082 337256
rect 80198 336048 80204 336100
rect 80256 336088 80262 336100
rect 85718 336088 85724 336100
rect 80256 336060 85724 336088
rect 80256 336048 80262 336060
rect 85718 336048 85724 336060
rect 85776 336048 85782 336100
rect 321422 336048 321428 336100
rect 321480 336088 321486 336100
rect 327310 336088 327316 336100
rect 321480 336060 327316 336088
rect 321480 336048 321486 336060
rect 327310 336048 327316 336060
rect 327368 336048 327374 336100
rect 131902 335980 131908 336032
rect 131960 336020 131966 336032
rect 138066 336020 138072 336032
rect 131960 335992 138072 336020
rect 131960 335980 131966 335992
rect 138066 335980 138072 335992
rect 138124 335980 138130 336032
rect 85810 335912 85816 335964
rect 85868 335952 85874 335964
rect 87834 335952 87840 335964
rect 85868 335924 87840 335952
rect 85868 335912 85874 335924
rect 87834 335912 87840 335924
rect 87892 335912 87898 335964
rect 131810 335912 131816 335964
rect 131868 335952 131874 335964
rect 138158 335952 138164 335964
rect 131868 335924 138164 335952
rect 131868 335912 131874 335924
rect 138158 335912 138164 335924
rect 138216 335912 138222 335964
rect 172842 335912 172848 335964
rect 172900 335952 172906 335964
rect 181582 335952 181588 335964
rect 172900 335924 181588 335952
rect 172900 335912 172906 335924
rect 181582 335912 181588 335924
rect 181640 335912 181646 335964
rect 225926 335912 225932 335964
rect 225984 335952 225990 335964
rect 230894 335952 230900 335964
rect 225984 335924 230900 335952
rect 225984 335912 225990 335924
rect 230894 335912 230900 335924
rect 230952 335912 230958 335964
rect 321606 335912 321612 335964
rect 321664 335952 321670 335964
rect 327218 335952 327224 335964
rect 321664 335924 327224 335952
rect 321664 335912 321670 335924
rect 327218 335912 327224 335924
rect 327276 335912 327282 335964
rect 395206 335912 395212 335964
rect 395264 335952 395270 335964
rect 395298 335952 395304 335964
rect 395264 335924 395304 335952
rect 395264 335912 395270 335924
rect 395298 335912 395304 335924
rect 395356 335912 395362 335964
rect 230802 335844 230808 335896
rect 230860 335884 230866 335896
rect 233470 335884 233476 335896
rect 230860 335856 233476 335884
rect 230860 335844 230866 335856
rect 233470 335844 233476 335856
rect 233528 335844 233534 335896
rect 266590 335844 266596 335896
rect 266648 335884 266654 335896
rect 275054 335884 275060 335896
rect 266648 335856 275060 335884
rect 266648 335844 266654 335856
rect 275054 335844 275060 335856
rect 275112 335844 275118 335896
rect 80198 335096 80204 335148
rect 80256 335136 80262 335148
rect 84982 335136 84988 335148
rect 80256 335108 84988 335136
rect 80256 335096 80262 335108
rect 84982 335096 84988 335108
rect 85040 335096 85046 335148
rect 75417 334799 75475 334805
rect 75417 334765 75429 334799
rect 75463 334796 75475 334799
rect 75966 334796 75972 334808
rect 75463 334768 75972 334796
rect 75463 334765 75475 334768
rect 75417 334759 75475 334765
rect 75966 334756 75972 334768
rect 76024 334756 76030 334808
rect 75509 334731 75567 334737
rect 75509 334697 75521 334731
rect 75555 334728 75567 334731
rect 75874 334728 75880 334740
rect 75555 334700 75880 334728
rect 75555 334697 75567 334700
rect 75509 334691 75567 334697
rect 75874 334688 75880 334700
rect 75932 334688 75938 334740
rect 76058 334688 76064 334740
rect 76116 334688 76122 334740
rect 76076 334536 76104 334688
rect 212773 334595 212831 334601
rect 212773 334561 212785 334595
rect 212819 334592 212831 334595
rect 221053 334595 221111 334601
rect 221053 334592 221065 334595
rect 212819 334564 221065 334592
rect 212819 334561 212831 334564
rect 212773 334555 212831 334561
rect 221053 334561 221065 334564
rect 221099 334561 221111 334595
rect 221053 334555 221111 334561
rect 75966 334524 75972 334536
rect 75927 334496 75972 334524
rect 75966 334484 75972 334496
rect 76024 334484 76030 334536
rect 76058 334484 76064 334536
rect 76116 334484 76122 334536
rect 108258 334456 108264 334468
rect 75800 334428 108264 334456
rect 75800 334320 75828 334428
rect 108258 334416 108264 334428
rect 108316 334456 108322 334468
rect 131626 334456 131632 334468
rect 108316 334428 131632 334456
rect 108316 334416 108322 334428
rect 131626 334416 131632 334428
rect 131684 334416 131690 334468
rect 136134 334416 136140 334468
rect 136192 334456 136198 334468
rect 139630 334456 139636 334468
rect 136192 334428 139636 334456
rect 136192 334416 136198 334428
rect 139630 334416 139636 334428
rect 139688 334416 139694 334468
rect 212310 334416 212316 334468
rect 212368 334456 212374 334468
rect 212773 334459 212831 334465
rect 212773 334456 212785 334459
rect 212368 334428 212785 334456
rect 212368 334416 212374 334428
rect 212773 334425 212785 334428
rect 212819 334425 212831 334459
rect 212773 334419 212831 334425
rect 230710 334416 230716 334468
rect 230768 334456 230774 334468
rect 233470 334456 233476 334468
rect 230768 334428 233476 334456
rect 230768 334416 230774 334428
rect 233470 334416 233476 334428
rect 233528 334416 233534 334468
rect 266590 334416 266596 334468
rect 266648 334456 266654 334468
rect 275606 334456 275612 334468
rect 266648 334428 275612 334456
rect 266648 334416 266654 334428
rect 275606 334416 275612 334428
rect 275664 334416 275670 334468
rect 75874 334348 75880 334400
rect 75932 334388 75938 334400
rect 104854 334388 104860 334400
rect 75932 334360 104860 334388
rect 75932 334348 75938 334360
rect 104854 334348 104860 334360
rect 104912 334388 104918 334400
rect 131718 334388 131724 334400
rect 104912 334360 131724 334388
rect 104912 334348 104918 334360
rect 131718 334348 131724 334360
rect 131776 334348 131782 334400
rect 266682 334348 266688 334400
rect 266740 334388 266746 334400
rect 271466 334388 271472 334400
rect 266740 334360 271472 334388
rect 266740 334348 266746 334360
rect 271466 334348 271472 334360
rect 271524 334348 271530 334400
rect 75966 334320 75972 334332
rect 75800 334292 75972 334320
rect 75966 334280 75972 334292
rect 76024 334280 76030 334332
rect 76978 334280 76984 334332
rect 77036 334320 77042 334332
rect 98230 334320 98236 334332
rect 77036 334292 98236 334320
rect 77036 334280 77042 334292
rect 98230 334280 98236 334292
rect 98288 334280 98294 334332
rect 111386 334280 111392 334332
rect 111444 334320 111450 334332
rect 131534 334320 131540 334332
rect 111444 334292 131540 334320
rect 111444 334280 111450 334292
rect 131534 334280 131540 334292
rect 131592 334280 131598 334332
rect 80198 334212 80204 334264
rect 80256 334252 80262 334264
rect 87834 334252 87840 334264
rect 80256 334224 87840 334252
rect 80256 334212 80262 334224
rect 87834 334212 87840 334224
rect 87892 334212 87898 334264
rect 114790 334212 114796 334264
rect 114848 334252 114854 334264
rect 131442 334252 131448 334264
rect 114848 334224 131448 334252
rect 114848 334212 114854 334224
rect 131442 334212 131448 334224
rect 131500 334212 131506 334264
rect 136226 334212 136232 334264
rect 136284 334252 136290 334264
rect 139630 334252 139636 334264
rect 136284 334224 139636 334252
rect 136284 334212 136290 334224
rect 139630 334212 139636 334224
rect 139688 334212 139694 334264
rect 221053 334255 221111 334261
rect 221053 334221 221065 334255
rect 221099 334252 221111 334255
rect 225282 334252 225288 334264
rect 221099 334224 225288 334252
rect 221099 334221 221111 334224
rect 221053 334215 221111 334221
rect 225282 334212 225288 334224
rect 225340 334252 225346 334264
rect 231354 334252 231360 334264
rect 225340 334224 231360 334252
rect 225340 334212 225346 334224
rect 231354 334212 231360 334224
rect 231412 334212 231418 334264
rect 78910 334144 78916 334196
rect 78968 334184 78974 334196
rect 88018 334184 88024 334196
rect 78968 334156 88024 334184
rect 78968 334144 78974 334156
rect 88018 334144 88024 334156
rect 88076 334144 88082 334196
rect 118194 334144 118200 334196
rect 118252 334184 118258 334196
rect 131350 334184 131356 334196
rect 118252 334156 131356 334184
rect 118252 334144 118258 334156
rect 131350 334144 131356 334156
rect 131408 334144 131414 334196
rect 131626 334144 131632 334196
rect 131684 334184 131690 334196
rect 136962 334184 136968 334196
rect 131684 334156 136968 334184
rect 131684 334144 131690 334156
rect 136962 334144 136968 334156
rect 137020 334144 137026 334196
rect 116078 334008 116084 334060
rect 116136 334048 116142 334060
rect 127854 334048 127860 334060
rect 116136 334020 127860 334048
rect 116136 334008 116142 334020
rect 127854 334008 127860 334020
rect 127912 334008 127918 334060
rect 131368 334048 131396 334144
rect 131534 334076 131540 334128
rect 131592 334116 131598 334128
rect 137054 334116 137060 334128
rect 131592 334088 137060 334116
rect 131592 334076 131598 334088
rect 137054 334076 137060 334088
rect 137112 334076 137118 334128
rect 137238 334048 137244 334060
rect 131368 334020 137244 334048
rect 137238 334008 137244 334020
rect 137296 334008 137302 334060
rect 103658 333940 103664 333992
rect 103716 333980 103722 333992
rect 124542 333980 124548 333992
rect 103716 333952 124548 333980
rect 103716 333940 103722 333952
rect 124542 333940 124548 333952
rect 124600 333940 124606 333992
rect 131442 333940 131448 333992
rect 131500 333980 131506 333992
rect 137146 333980 137152 333992
rect 131500 333952 137152 333980
rect 131500 333940 131506 333952
rect 137146 333940 137152 333952
rect 137204 333940 137210 333992
rect 211298 333940 211304 333992
rect 211356 333980 211362 333992
rect 221878 333980 221884 333992
rect 211356 333952 221884 333980
rect 211356 333940 211362 333952
rect 221878 333940 221884 333952
rect 221936 333940 221942 333992
rect 305138 333940 305144 333992
rect 305196 333980 305202 333992
rect 316178 333980 316184 333992
rect 305196 333952 316184 333980
rect 305196 333940 305202 333952
rect 316178 333940 316184 333952
rect 316236 333940 316242 333992
rect 91238 333872 91244 333924
rect 91296 333912 91302 333924
rect 121230 333912 121236 333924
rect 91296 333884 121236 333912
rect 91296 333872 91302 333884
rect 121230 333872 121236 333884
rect 121288 333872 121294 333924
rect 131718 333872 131724 333924
rect 131776 333912 131782 333924
rect 137514 333912 137520 333924
rect 131776 333884 137520 333912
rect 131776 333872 131782 333884
rect 137514 333872 137520 333884
rect 137572 333872 137578 333924
rect 197498 333872 197504 333924
rect 197556 333912 197562 333924
rect 218566 333912 218572 333924
rect 197556 333884 218572 333912
rect 197556 333872 197562 333884
rect 218566 333872 218572 333884
rect 218624 333872 218630 333924
rect 292718 333872 292724 333924
rect 292776 333912 292782 333924
rect 312866 333912 312872 333924
rect 292776 333884 312872 333912
rect 292776 333872 292782 333884
rect 312866 333872 312872 333884
rect 312924 333872 312930 333924
rect 98230 333804 98236 333856
rect 98288 333844 98294 333856
rect 137974 333844 137980 333856
rect 98288 333816 137980 333844
rect 98288 333804 98294 333816
rect 137974 333804 137980 333816
rect 138032 333804 138038 333856
rect 185078 333804 185084 333856
rect 185136 333844 185142 333856
rect 215622 333844 215628 333856
rect 185136 333816 215628 333844
rect 185136 333804 185142 333816
rect 215622 333804 215628 333816
rect 215680 333804 215686 333856
rect 280298 333804 280304 333856
rect 280356 333844 280362 333856
rect 309554 333844 309560 333856
rect 280356 333816 309560 333844
rect 280356 333804 280362 333816
rect 309554 333804 309560 333816
rect 309612 333804 309618 333856
rect 91882 333736 91888 333788
rect 91940 333776 91946 333788
rect 134846 333776 134852 333788
rect 91940 333748 134852 333776
rect 91940 333736 91946 333748
rect 134846 333736 134852 333748
rect 134904 333736 134910 333788
rect 185906 333736 185912 333788
rect 185964 333776 185970 333788
rect 228594 333776 228600 333788
rect 185964 333748 228600 333776
rect 185964 333736 185970 333748
rect 228594 333736 228600 333748
rect 228652 333736 228658 333788
rect 279562 333736 279568 333788
rect 279620 333776 279626 333788
rect 322618 333776 322624 333788
rect 279620 333748 322624 333776
rect 279620 333736 279626 333748
rect 322618 333736 322624 333748
rect 322676 333736 322682 333788
rect 173302 333464 173308 333516
rect 173360 333504 173366 333516
rect 180386 333504 180392 333516
rect 173360 333476 180392 333504
rect 173360 333464 173366 333476
rect 180386 333464 180392 333476
rect 180444 333464 180450 333516
rect 80198 333056 80204 333108
rect 80256 333096 80262 333108
rect 87374 333096 87380 333108
rect 80256 333068 87380 333096
rect 80256 333056 80262 333068
rect 87374 333056 87380 333068
rect 87432 333056 87438 333108
rect 138066 333056 138072 333108
rect 138124 333096 138130 333108
rect 139630 333096 139636 333108
rect 138124 333068 139636 333096
rect 138124 333056 138130 333068
rect 139630 333056 139636 333068
rect 139688 333056 139694 333108
rect 230894 333056 230900 333108
rect 230952 333096 230958 333108
rect 233470 333096 233476 333108
rect 230952 333068 233476 333096
rect 230952 333056 230958 333068
rect 233470 333056 233476 333068
rect 233528 333056 233534 333108
rect 266590 333056 266596 333108
rect 266648 333096 266654 333108
rect 274870 333096 274876 333108
rect 266648 333068 274876 333096
rect 266648 333056 266654 333068
rect 274870 333056 274876 333068
rect 274928 333056 274934 333108
rect 201733 331875 201791 331881
rect 201733 331841 201745 331875
rect 201779 331872 201791 331875
rect 211301 331875 211359 331881
rect 211301 331872 211313 331875
rect 201779 331844 211313 331872
rect 201779 331841 201791 331844
rect 201733 331835 201791 331841
rect 211301 331841 211313 331844
rect 211347 331841 211359 331875
rect 211301 331835 211359 331841
rect 319306 331764 319312 331816
rect 319364 331804 319370 331816
rect 325378 331804 325384 331816
rect 319364 331776 325384 331804
rect 319364 331764 319370 331776
rect 325378 331764 325384 331776
rect 325436 331764 325442 331816
rect 76886 331696 76892 331748
rect 76944 331736 76950 331748
rect 118194 331736 118200 331748
rect 76944 331708 118200 331736
rect 76944 331696 76950 331708
rect 118194 331696 118200 331708
rect 118252 331696 118258 331748
rect 138158 331696 138164 331748
rect 138216 331736 138222 331748
rect 139630 331736 139636 331748
rect 138216 331708 139636 331736
rect 138216 331696 138222 331708
rect 139630 331696 139636 331708
rect 139688 331696 139694 331748
rect 173670 331696 173676 331748
rect 173728 331736 173734 331748
rect 180938 331736 180944 331748
rect 173728 331708 180944 331736
rect 173728 331696 173734 331708
rect 180938 331696 180944 331708
rect 180996 331696 181002 331748
rect 198694 331696 198700 331748
rect 198752 331736 198758 331748
rect 201733 331739 201791 331745
rect 201733 331736 201745 331739
rect 198752 331708 201745 331736
rect 198752 331696 198758 331708
rect 201733 331705 201745 331708
rect 201779 331705 201791 331739
rect 201733 331699 201791 331705
rect 225116 331708 225420 331736
rect 75509 331671 75567 331677
rect 75509 331637 75521 331671
rect 75555 331668 75567 331671
rect 114790 331668 114796 331680
rect 75555 331640 114796 331668
rect 75555 331637 75567 331640
rect 75509 331631 75567 331637
rect 114790 331628 114796 331640
rect 114848 331628 114854 331680
rect 225116 331668 225144 331708
rect 212788 331640 225144 331668
rect 75417 331603 75475 331609
rect 75417 331569 75429 331603
rect 75463 331600 75475 331603
rect 111386 331600 111392 331612
rect 75463 331572 111392 331600
rect 75463 331569 75475 331572
rect 75417 331563 75475 331569
rect 111386 331560 111392 331572
rect 111444 331560 111450 331612
rect 211301 331603 211359 331609
rect 211301 331569 211313 331603
rect 211347 331600 211359 331603
rect 212788 331600 212816 331640
rect 211347 331572 212816 331600
rect 225392 331600 225420 331708
rect 226570 331696 226576 331748
rect 226628 331736 226634 331748
rect 233470 331736 233476 331748
rect 226628 331708 233476 331736
rect 226628 331696 226634 331708
rect 233470 331696 233476 331708
rect 233528 331696 233534 331748
rect 266590 331696 266596 331748
rect 266648 331736 266654 331748
rect 274962 331736 274968 331748
rect 266648 331708 274968 331736
rect 266648 331696 266654 331708
rect 274962 331696 274968 331708
rect 275020 331696 275026 331748
rect 299526 331696 299532 331748
rect 299584 331736 299590 331748
rect 319214 331736 319220 331748
rect 299584 331708 319220 331736
rect 299584 331696 299590 331708
rect 319214 331696 319220 331708
rect 319272 331696 319278 331748
rect 225558 331600 225564 331612
rect 225392 331572 225564 331600
rect 211347 331569 211359 331572
rect 211301 331563 211359 331569
rect 225558 331560 225564 331572
rect 225616 331600 225622 331612
rect 230802 331600 230808 331612
rect 225616 331572 230808 331600
rect 225616 331560 225622 331572
rect 230802 331560 230808 331572
rect 230860 331560 230866 331612
rect 80198 330608 80204 330660
rect 80256 330648 80262 330660
rect 85810 330648 85816 330660
rect 80256 330620 85816 330648
rect 80256 330608 80262 330620
rect 85810 330608 85816 330620
rect 85868 330608 85874 330660
rect 319398 330472 319404 330524
rect 319456 330512 319462 330524
rect 325562 330512 325568 330524
rect 319456 330484 325568 330512
rect 319456 330472 319462 330484
rect 325562 330472 325568 330484
rect 325620 330472 325626 330524
rect 319214 330404 319220 330456
rect 319272 330444 319278 330456
rect 324642 330444 324648 330456
rect 319272 330416 324648 330444
rect 319272 330404 319278 330416
rect 324642 330404 324648 330416
rect 324700 330404 324706 330456
rect 305230 330336 305236 330388
rect 305288 330376 305294 330388
rect 306242 330376 306248 330388
rect 305288 330348 306248 330376
rect 305288 330336 305294 330348
rect 306242 330336 306248 330348
rect 306300 330376 306306 330388
rect 319030 330376 319036 330388
rect 306300 330348 319036 330376
rect 306300 330336 306306 330348
rect 319030 330336 319036 330348
rect 319088 330376 319094 330388
rect 325746 330376 325752 330388
rect 319088 330348 325752 330376
rect 319088 330336 319094 330348
rect 325746 330336 325752 330348
rect 325804 330336 325810 330388
rect 75506 330172 75512 330184
rect 75467 330144 75512 330172
rect 75506 330132 75512 330144
rect 75564 330132 75570 330184
rect 75414 330104 75420 330116
rect 75375 330076 75420 330104
rect 75414 330064 75420 330076
rect 75472 330064 75478 330116
rect 182413 329291 182471 329297
rect 182413 329257 182425 329291
rect 182459 329288 182471 329291
rect 191981 329291 192039 329297
rect 191981 329288 191993 329291
rect 182459 329260 191993 329288
rect 182459 329257 182471 329260
rect 182413 329251 182471 329257
rect 191981 329257 191993 329260
rect 192027 329257 192039 329291
rect 191981 329251 192039 329257
rect 154813 329223 154871 329229
rect 154813 329189 154825 329223
rect 154859 329220 154871 329223
rect 158214 329220 158220 329232
rect 154859 329192 158220 329220
rect 154859 329189 154871 329192
rect 154813 329183 154871 329189
rect 158214 329180 158220 329192
rect 158272 329180 158278 329232
rect 174133 329223 174191 329229
rect 164672 329192 174084 329220
rect 137514 329044 137520 329096
rect 137572 329084 137578 329096
rect 147729 329087 147787 329093
rect 147729 329084 147741 329087
rect 137572 329056 147741 329084
rect 137572 329044 137578 329056
rect 147729 329053 147741 329056
rect 147775 329053 147787 329087
rect 147729 329047 147787 329053
rect 148005 329087 148063 329093
rect 148005 329053 148017 329087
rect 148051 329084 148063 329087
rect 154813 329087 154871 329093
rect 154813 329084 154825 329087
rect 148051 329056 154825 329084
rect 148051 329053 148063 329056
rect 148005 329047 148063 329053
rect 154813 329053 154825 329056
rect 154859 329053 154871 329087
rect 154813 329047 154871 329053
rect 158214 329044 158220 329096
rect 158272 329084 158278 329096
rect 164672 329084 164700 329192
rect 174056 329152 174084 329192
rect 174133 329189 174145 329223
rect 174179 329189 174191 329223
rect 174133 329183 174191 329189
rect 174148 329152 174176 329183
rect 174056 329124 174176 329152
rect 191981 329155 192039 329161
rect 191981 329121 191993 329155
rect 192027 329152 192039 329155
rect 198878 329152 198884 329164
rect 192027 329124 198884 329152
rect 192027 329121 192039 329124
rect 191981 329115 192039 329121
rect 198878 329112 198884 329124
rect 198936 329112 198942 329164
rect 158272 329056 164700 329084
rect 158272 329044 158278 329056
rect 172106 329044 172112 329096
rect 172164 329084 172170 329096
rect 176801 329087 176859 329093
rect 176801 329084 176813 329087
rect 172164 329056 176813 329084
rect 172164 329044 172170 329056
rect 176801 329053 176813 329056
rect 176847 329053 176859 329087
rect 176801 329047 176859 329053
rect 176893 329087 176951 329093
rect 176893 329053 176905 329087
rect 176939 329084 176951 329087
rect 186461 329087 186519 329093
rect 186461 329084 186473 329087
rect 176939 329056 186473 329084
rect 176939 329053 176951 329056
rect 176893 329047 176951 329053
rect 186461 329053 186473 329056
rect 186507 329053 186519 329087
rect 186461 329047 186519 329053
rect 186645 329087 186703 329093
rect 186645 329053 186657 329087
rect 186691 329084 186703 329087
rect 222522 329084 222528 329096
rect 186691 329056 222528 329084
rect 186691 329053 186703 329056
rect 186645 329047 186703 329053
rect 222522 329044 222528 329056
rect 222580 329084 222586 329096
rect 233470 329084 233476 329096
rect 222580 329056 233476 329084
rect 222580 329044 222586 329056
rect 233470 329044 233476 329056
rect 233528 329044 233534 329096
rect 266590 329044 266596 329096
rect 266648 329084 266654 329096
rect 316546 329084 316552 329096
rect 266648 329056 316552 329084
rect 266648 329044 266654 329056
rect 316546 329044 316552 329056
rect 316604 329084 316610 329096
rect 328414 329084 328420 329096
rect 316604 329056 328420 329084
rect 316604 329044 316610 329056
rect 328414 329044 328420 329056
rect 328472 329044 328478 329096
rect 78910 328976 78916 329028
rect 78968 329016 78974 329028
rect 128498 329016 128504 329028
rect 78968 328988 128504 329016
rect 78968 328976 78974 328988
rect 128498 328976 128504 328988
rect 128556 329016 128562 329028
rect 140366 329016 140372 329028
rect 128556 328988 140372 329016
rect 128556 328976 128562 328988
rect 140366 328976 140372 328988
rect 140424 328976 140430 329028
rect 231354 328976 231360 329028
rect 231412 329016 231418 329028
rect 255550 329016 255556 329028
rect 231412 328988 255556 329016
rect 231412 328976 231418 328988
rect 255550 328976 255556 328988
rect 255608 329016 255614 329028
rect 305230 329016 305236 329028
rect 255608 328988 305236 329016
rect 255608 328976 255614 328988
rect 305230 328976 305236 328988
rect 305288 328976 305294 329028
rect 325194 328976 325200 329028
rect 325252 329016 325258 329028
rect 429430 329016 429436 329028
rect 325252 328988 429436 329016
rect 325252 328976 325258 328988
rect 429430 328976 429436 328988
rect 429488 328976 429494 329028
rect 208722 328908 208728 328960
rect 208780 328948 208786 328960
rect 225190 328948 225196 328960
rect 208780 328920 225196 328948
rect 208780 328908 208786 328920
rect 225190 328908 225196 328920
rect 225248 328948 225254 328960
rect 231078 328948 231084 328960
rect 225248 328920 231084 328948
rect 225248 328908 225254 328920
rect 231078 328908 231084 328920
rect 231136 328908 231142 328960
rect 302470 328908 302476 328960
rect 302528 328948 302534 328960
rect 303114 328948 303120 328960
rect 302528 328920 303120 328948
rect 302528 328908 302534 328920
rect 303114 328908 303120 328920
rect 303172 328948 303178 328960
rect 319122 328948 319128 328960
rect 303172 328920 319128 328948
rect 303172 328908 303178 328920
rect 319122 328908 319128 328920
rect 319180 328948 319186 328960
rect 325654 328948 325660 328960
rect 319180 328920 325660 328948
rect 319180 328908 319186 328920
rect 325654 328908 325660 328920
rect 325712 328908 325718 328960
rect 174133 328883 174191 328889
rect 174133 328849 174145 328883
rect 174179 328880 174191 328883
rect 182413 328883 182471 328889
rect 182413 328880 182425 328883
rect 174179 328852 182425 328880
rect 174179 328849 174191 328852
rect 174133 328843 174191 328849
rect 182413 328849 182425 328852
rect 182459 328849 182471 328883
rect 182413 328843 182471 328849
rect 342490 327616 342496 327668
rect 342548 327656 342554 327668
rect 346446 327656 346452 327668
rect 342548 327628 346452 327656
rect 342548 327616 342554 327628
rect 346446 327616 346452 327628
rect 346504 327616 346510 327668
rect 395114 327616 395120 327668
rect 395172 327656 395178 327668
rect 395206 327656 395212 327668
rect 395172 327628 395212 327656
rect 395172 327616 395178 327628
rect 395206 327616 395212 327628
rect 395264 327616 395270 327668
rect 76058 327548 76064 327600
rect 76116 327588 76122 327600
rect 100990 327588 100996 327600
rect 76116 327560 100996 327588
rect 76116 327548 76122 327560
rect 100990 327548 100996 327560
rect 101048 327548 101054 327600
rect 156282 327548 156288 327600
rect 156340 327588 156346 327600
rect 156834 327588 156840 327600
rect 156340 327560 156840 327588
rect 156340 327548 156346 327560
rect 156834 327548 156840 327560
rect 156892 327588 156898 327600
rect 194830 327588 194836 327600
rect 156892 327560 194836 327588
rect 156892 327548 156898 327560
rect 194830 327548 194836 327560
rect 194888 327548 194894 327600
rect 241474 327548 241480 327600
rect 241532 327588 241538 327600
rect 252882 327588 252888 327600
rect 241532 327560 252888 327588
rect 241532 327548 241538 327560
rect 252882 327548 252888 327560
rect 252940 327548 252946 327600
rect 254814 327548 254820 327600
rect 254872 327588 254878 327600
rect 302470 327588 302476 327600
rect 254872 327560 302476 327588
rect 254872 327548 254878 327560
rect 302470 327548 302476 327560
rect 302528 327548 302534 327600
rect 339914 327548 339920 327600
rect 339972 327588 339978 327600
rect 356014 327588 356020 327600
rect 339972 327560 356020 327588
rect 339972 327548 339978 327560
rect 356014 327548 356020 327560
rect 356072 327548 356078 327600
rect 65478 327480 65484 327532
rect 65536 327520 65542 327532
rect 69434 327520 69440 327532
rect 65536 327492 69440 327520
rect 65536 327480 65542 327492
rect 69434 327480 69440 327492
rect 69492 327480 69498 327532
rect 137698 327480 137704 327532
rect 137756 327520 137762 327532
rect 137974 327520 137980 327532
rect 137756 327492 137980 327520
rect 137756 327480 137762 327492
rect 137974 327480 137980 327492
rect 138032 327520 138038 327532
rect 155914 327520 155920 327532
rect 138032 327492 155920 327520
rect 138032 327480 138038 327492
rect 155914 327480 155920 327492
rect 155972 327520 155978 327532
rect 163369 327523 163427 327529
rect 163369 327520 163381 327523
rect 155972 327492 163381 327520
rect 155972 327480 155978 327492
rect 163369 327489 163381 327492
rect 163415 327489 163427 327523
rect 163369 327483 163427 327489
rect 168337 327523 168395 327529
rect 168337 327489 168349 327523
rect 168383 327520 168395 327523
rect 181033 327523 181091 327529
rect 181033 327520 181045 327523
rect 168383 327492 181045 327520
rect 168383 327489 168395 327492
rect 168337 327483 168395 327489
rect 181033 327489 181045 327492
rect 181079 327489 181091 327523
rect 181033 327483 181091 327489
rect 238622 327480 238628 327532
rect 238680 327520 238686 327532
rect 249938 327520 249944 327532
rect 238680 327492 249944 327520
rect 238680 327480 238686 327492
rect 249938 327480 249944 327492
rect 249996 327480 250002 327532
rect 250030 327480 250036 327532
rect 250088 327520 250094 327532
rect 250766 327520 250772 327532
rect 250088 327492 250772 327520
rect 250088 327480 250094 327492
rect 250766 327480 250772 327492
rect 250824 327520 250830 327532
rect 288670 327520 288676 327532
rect 250824 327492 288676 327520
rect 250824 327480 250830 327492
rect 288670 327480 288676 327492
rect 288728 327520 288734 327532
rect 289958 327520 289964 327532
rect 288728 327492 289964 327520
rect 288728 327480 288734 327492
rect 289958 327480 289964 327492
rect 290016 327480 290022 327532
rect 337154 327480 337160 327532
rect 337212 327520 337218 327532
rect 352794 327520 352800 327532
rect 337212 327492 352800 327520
rect 337212 327480 337218 327492
rect 352794 327480 352800 327492
rect 352852 327480 352858 327532
rect 66858 327412 66864 327464
rect 66916 327452 66922 327464
rect 70630 327452 70636 327464
rect 66916 327424 70636 327452
rect 66916 327412 66922 327424
rect 70630 327412 70636 327424
rect 70688 327412 70694 327464
rect 154810 327412 154816 327464
rect 154868 327452 154874 327464
rect 168245 327455 168303 327461
rect 168245 327452 168257 327455
rect 154868 327424 168257 327452
rect 154868 327412 154874 327424
rect 168245 327421 168257 327424
rect 168291 327421 168303 327455
rect 168245 327415 168303 327421
rect 174041 327455 174099 327461
rect 174041 327421 174053 327455
rect 174087 327452 174099 327455
rect 183793 327455 183851 327461
rect 183793 327452 183805 327455
rect 174087 327424 183805 327452
rect 174087 327421 174099 327424
rect 174041 327415 174099 327421
rect 183793 327421 183805 327424
rect 183839 327421 183851 327455
rect 192070 327452 192076 327464
rect 183793 327415 183851 327421
rect 191996 327424 192076 327452
rect 59222 327344 59228 327396
rect 59280 327384 59286 327396
rect 63638 327384 63644 327396
rect 59280 327356 63644 327384
rect 59280 327344 59286 327356
rect 63638 327344 63644 327356
rect 63696 327344 63702 327396
rect 66306 327344 66312 327396
rect 66364 327384 66370 327396
rect 67502 327384 67508 327396
rect 66364 327356 67508 327384
rect 66364 327344 66370 327356
rect 67502 327344 67508 327356
rect 67560 327344 67566 327396
rect 69066 327344 69072 327396
rect 69124 327384 69130 327396
rect 72654 327384 72660 327396
rect 69124 327356 72660 327384
rect 69124 327344 69130 327356
rect 72654 327344 72660 327356
rect 72712 327344 72718 327396
rect 151958 327344 151964 327396
rect 152016 327384 152022 327396
rect 165206 327384 165212 327396
rect 152016 327356 165212 327384
rect 152016 327344 152022 327356
rect 165206 327344 165212 327356
rect 165264 327344 165270 327396
rect 181033 327387 181091 327393
rect 181033 327353 181045 327387
rect 181079 327384 181091 327387
rect 191996 327384 192024 327424
rect 192070 327412 192076 327424
rect 192128 327452 192134 327464
rect 196213 327455 196271 327461
rect 196213 327452 196225 327455
rect 192128 327424 196225 327452
rect 192128 327412 192134 327424
rect 196213 327421 196225 327424
rect 196259 327421 196271 327455
rect 196213 327415 196271 327421
rect 231998 327412 232004 327464
rect 232056 327452 232062 327464
rect 248650 327452 248656 327464
rect 232056 327424 248656 327452
rect 232056 327412 232062 327424
rect 248650 327412 248656 327424
rect 248708 327412 248714 327464
rect 248742 327412 248748 327464
rect 248800 327452 248806 327464
rect 249846 327452 249852 327464
rect 248800 327424 249852 327452
rect 248800 327412 248806 327424
rect 249846 327412 249852 327424
rect 249904 327452 249910 327464
rect 285910 327452 285916 327464
rect 249904 327424 285916 327452
rect 249904 327412 249910 327424
rect 285910 327412 285916 327424
rect 285968 327412 285974 327464
rect 338626 327412 338632 327464
rect 338684 327452 338690 327464
rect 353622 327452 353628 327464
rect 338684 327424 353628 327452
rect 338684 327412 338690 327424
rect 353622 327412 353628 327424
rect 353680 327412 353686 327464
rect 181079 327356 192024 327384
rect 181079 327353 181091 327356
rect 181033 327347 181091 327353
rect 238990 327344 238996 327396
rect 239048 327384 239054 327396
rect 239910 327384 239916 327396
rect 239048 327356 239916 327384
rect 239048 327344 239054 327356
rect 239910 327344 239916 327356
rect 239968 327344 239974 327396
rect 244418 327344 244424 327396
rect 244476 327384 244482 327396
rect 246902 327384 246908 327396
rect 244476 327356 246908 327384
rect 244476 327344 244482 327356
rect 246902 327344 246908 327356
rect 246960 327344 246966 327396
rect 258221 327387 258279 327393
rect 258221 327353 258233 327387
rect 258267 327384 258279 327387
rect 281770 327384 281776 327396
rect 258267 327356 281776 327384
rect 258267 327353 258279 327356
rect 258221 327347 258279 327353
rect 281770 327344 281776 327356
rect 281828 327384 281834 327396
rect 282230 327384 282236 327396
rect 281828 327356 282236 327384
rect 281828 327344 281834 327356
rect 282230 327344 282236 327356
rect 282288 327344 282294 327396
rect 332922 327344 332928 327396
rect 332980 327384 332986 327396
rect 333658 327384 333664 327396
rect 332980 327356 333664 327384
rect 332980 327344 332986 327356
rect 333658 327344 333664 327356
rect 333716 327344 333722 327396
rect 334210 327344 334216 327396
rect 334268 327384 334274 327396
rect 335222 327384 335228 327396
rect 334268 327356 335228 327384
rect 334268 327344 334274 327356
rect 335222 327344 335228 327356
rect 335280 327344 335286 327396
rect 341478 327344 341484 327396
rect 341536 327384 341542 327396
rect 357578 327384 357584 327396
rect 341536 327356 357584 327384
rect 341536 327344 341542 327356
rect 357578 327344 357584 327356
rect 357636 327344 357642 327396
rect 60234 327276 60240 327328
rect 60292 327316 60298 327328
rect 65018 327316 65024 327328
rect 60292 327288 65024 327316
rect 60292 327276 60298 327288
rect 65018 327276 65024 327288
rect 65076 327276 65082 327328
rect 66490 327276 66496 327328
rect 66548 327316 66554 327328
rect 68514 327316 68520 327328
rect 66548 327288 68520 327316
rect 66548 327276 66554 327288
rect 68514 327276 68520 327288
rect 68572 327276 68578 327328
rect 151314 327276 151320 327328
rect 151372 327316 151378 327328
rect 163182 327316 163188 327328
rect 151372 327288 163188 327316
rect 151372 327276 151378 327288
rect 163182 327276 163188 327288
rect 163240 327276 163246 327328
rect 163369 327319 163427 327325
rect 163369 327285 163381 327319
rect 163415 327316 163427 327319
rect 168337 327319 168395 327325
rect 168337 327316 168349 327319
rect 163415 327288 168349 327316
rect 163415 327285 163427 327288
rect 163369 327279 163427 327285
rect 168337 327285 168349 327288
rect 168383 327285 168395 327319
rect 168337 327279 168395 327285
rect 245338 327276 245344 327328
rect 245396 327316 245402 327328
rect 247914 327316 247920 327328
rect 245396 327288 247920 327316
rect 245396 327276 245402 327288
rect 247914 327276 247920 327288
rect 247972 327276 247978 327328
rect 261162 327316 261168 327328
rect 248024 327288 261168 327316
rect 68422 327208 68428 327260
rect 68480 327248 68486 327260
rect 71642 327248 71648 327260
rect 68480 327220 71648 327248
rect 68480 327208 68486 327220
rect 71642 327208 71648 327220
rect 71700 327208 71706 327260
rect 149382 327208 149388 327260
rect 149440 327248 149446 327260
rect 163274 327248 163280 327260
rect 149440 327220 163280 327248
rect 149440 327208 149446 327220
rect 163274 327208 163280 327220
rect 163332 327208 163338 327260
rect 168245 327251 168303 327257
rect 168245 327217 168257 327251
rect 168291 327248 168303 327251
rect 174041 327251 174099 327257
rect 174041 327248 174053 327251
rect 168291 327220 174053 327248
rect 168291 327217 168303 327220
rect 168245 327211 168303 327217
rect 174041 327217 174053 327220
rect 174087 327217 174099 327251
rect 174041 327211 174099 327217
rect 247362 327208 247368 327260
rect 247420 327248 247426 327260
rect 248024 327248 248052 327288
rect 261162 327276 261168 327288
rect 261220 327276 261226 327328
rect 339546 327276 339552 327328
rect 339604 327316 339610 327328
rect 345897 327319 345955 327325
rect 345897 327316 345909 327319
rect 339604 327288 345909 327316
rect 339604 327276 339610 327288
rect 345897 327285 345909 327288
rect 345943 327285 345955 327319
rect 345897 327279 345955 327285
rect 348013 327319 348071 327325
rect 348013 327285 348025 327319
rect 348059 327316 348071 327319
rect 351966 327316 351972 327328
rect 348059 327288 351972 327316
rect 348059 327285 348071 327288
rect 348013 327279 348071 327285
rect 351966 327276 351972 327288
rect 352024 327276 352030 327328
rect 247420 327220 248052 327248
rect 248101 327251 248159 327257
rect 247420 327208 247426 327220
rect 248101 327217 248113 327251
rect 248147 327248 248159 327251
rect 258402 327248 258408 327260
rect 248147 327220 258408 327248
rect 248147 327217 248159 327220
rect 248101 327211 248159 327217
rect 258402 327208 258408 327220
rect 258460 327208 258466 327260
rect 344790 327208 344796 327260
rect 344848 327248 344854 327260
rect 358314 327248 358320 327260
rect 344848 327220 358320 327248
rect 344848 327208 344854 327220
rect 358314 327208 358320 327220
rect 358372 327208 358378 327260
rect 62350 327140 62356 327192
rect 62408 327180 62414 327192
rect 66582 327180 66588 327192
rect 62408 327152 66588 327180
rect 62408 327140 62414 327152
rect 66582 327140 66588 327152
rect 66640 327140 66646 327192
rect 154166 327140 154172 327192
rect 154224 327180 154230 327192
rect 168058 327180 168064 327192
rect 154224 327152 168064 327180
rect 154224 327140 154230 327152
rect 168058 327140 168064 327152
rect 168116 327140 168122 327192
rect 247178 327140 247184 327192
rect 247236 327180 247242 327192
rect 258954 327180 258960 327192
rect 247236 327152 258960 327180
rect 247236 327140 247242 327152
rect 258954 327140 258960 327152
rect 259012 327140 259018 327192
rect 342398 327140 342404 327192
rect 342456 327180 342462 327192
rect 355554 327180 355560 327192
rect 342456 327152 355560 327180
rect 342456 327140 342462 327152
rect 355554 327140 355560 327152
rect 355612 327140 355618 327192
rect 150762 327072 150768 327124
rect 150820 327112 150826 327124
rect 164562 327112 164568 327124
rect 150820 327084 164568 327112
rect 150820 327072 150826 327084
rect 164562 327072 164568 327084
rect 164620 327072 164626 327124
rect 194830 327072 194836 327124
rect 194888 327112 194894 327124
rect 232090 327112 232096 327124
rect 194888 327084 232096 327112
rect 194888 327072 194894 327084
rect 232090 327072 232096 327084
rect 232148 327112 232154 327124
rect 250030 327112 250036 327124
rect 232148 327084 250036 327112
rect 232148 327072 232154 327084
rect 250030 327072 250036 327084
rect 250088 327072 250094 327124
rect 250122 327072 250128 327124
rect 250180 327112 250186 327124
rect 264014 327112 264020 327124
rect 250180 327084 264020 327112
rect 250180 327072 250186 327084
rect 264014 327072 264020 327084
rect 264072 327072 264078 327124
rect 289958 327072 289964 327124
rect 290016 327112 290022 327124
rect 325286 327112 325292 327124
rect 290016 327084 325292 327112
rect 290016 327072 290022 327084
rect 325286 327072 325292 327084
rect 325344 327072 325350 327124
rect 341202 327072 341208 327124
rect 341260 327112 341266 327124
rect 358406 327112 358412 327124
rect 341260 327084 358412 327112
rect 341260 327072 341266 327084
rect 358406 327072 358412 327084
rect 358464 327072 358470 327124
rect 64374 327004 64380 327056
rect 64432 327044 64438 327056
rect 69158 327044 69164 327056
rect 64432 327016 69164 327044
rect 64432 327004 64438 327016
rect 69158 327004 69164 327016
rect 69216 327004 69222 327056
rect 153246 327004 153252 327056
rect 153304 327044 153310 327056
rect 165114 327044 165120 327056
rect 153304 327016 165120 327044
rect 153304 327004 153310 327016
rect 165114 327004 165120 327016
rect 165172 327004 165178 327056
rect 196213 327047 196271 327053
rect 196213 327013 196225 327047
rect 196259 327044 196271 327047
rect 233470 327044 233476 327056
rect 196259 327016 233476 327044
rect 196259 327013 196271 327016
rect 196213 327007 196271 327013
rect 233470 327004 233476 327016
rect 233528 327044 233534 327056
rect 248650 327044 248656 327056
rect 233528 327016 248656 327044
rect 233528 327004 233534 327016
rect 248650 327004 248656 327016
rect 248708 327004 248714 327056
rect 248742 327004 248748 327056
rect 248800 327044 248806 327056
rect 263094 327044 263100 327056
rect 248800 327016 263100 327044
rect 248800 327004 248806 327016
rect 263094 327004 263100 327016
rect 263152 327004 263158 327056
rect 285910 327004 285916 327056
rect 285968 327044 285974 327056
rect 324550 327044 324556 327056
rect 285968 327016 324556 327044
rect 285968 327004 285974 327016
rect 324550 327004 324556 327016
rect 324608 327004 324614 327056
rect 339914 327004 339920 327056
rect 339972 327044 339978 327056
rect 356750 327044 356756 327056
rect 339972 327016 356756 327044
rect 339972 327004 339978 327016
rect 356750 327004 356756 327016
rect 356808 327004 356814 327056
rect 137606 326936 137612 326988
rect 137664 326976 137670 326988
rect 154810 326976 154816 326988
rect 137664 326948 154816 326976
rect 137664 326936 137670 326948
rect 154810 326936 154816 326948
rect 154868 326936 154874 326988
rect 154902 326936 154908 326988
rect 154960 326976 154966 326988
rect 162357 326979 162415 326985
rect 162357 326976 162369 326979
rect 154960 326948 162369 326976
rect 154960 326936 154966 326948
rect 162357 326945 162369 326948
rect 162403 326945 162415 326979
rect 162357 326939 162415 326945
rect 183793 326979 183851 326985
rect 183793 326945 183805 326979
rect 183839 326976 183851 326979
rect 187930 326976 187936 326988
rect 183839 326948 187936 326976
rect 183839 326945 183851 326948
rect 183793 326939 183851 326945
rect 187930 326936 187936 326948
rect 187988 326976 187994 326988
rect 230710 326976 230716 326988
rect 187988 326948 230716 326976
rect 187988 326936 187994 326948
rect 230710 326936 230716 326948
rect 230768 326976 230774 326988
rect 231998 326976 232004 326988
rect 230768 326948 232004 326976
rect 230768 326936 230774 326948
rect 231998 326936 232004 326948
rect 232056 326936 232062 326988
rect 244602 326936 244608 326988
rect 244660 326976 244666 326988
rect 248101 326979 248159 326985
rect 248101 326976 248113 326979
rect 244660 326948 248113 326976
rect 244660 326936 244666 326948
rect 248101 326945 248113 326948
rect 248147 326945 248159 326979
rect 248101 326939 248159 326945
rect 248282 326936 248288 326988
rect 248340 326976 248346 326988
rect 268614 326976 268620 326988
rect 248340 326948 268620 326976
rect 248340 326936 248346 326948
rect 268614 326936 268620 326948
rect 268672 326936 268678 326988
rect 282230 326936 282236 326988
rect 282288 326976 282294 326988
rect 325470 326976 325476 326988
rect 282288 326948 325476 326976
rect 282288 326936 282294 326948
rect 325470 326936 325476 326948
rect 325528 326936 325534 326988
rect 338534 326936 338540 326988
rect 338592 326976 338598 326988
rect 355186 326976 355192 326988
rect 338592 326948 355192 326976
rect 338592 326936 338598 326948
rect 355186 326936 355192 326948
rect 355244 326936 355250 326988
rect 100990 326868 100996 326920
rect 101048 326908 101054 326920
rect 136870 326908 136876 326920
rect 101048 326880 136876 326908
rect 101048 326868 101054 326880
rect 136870 326868 136876 326880
rect 136928 326868 136934 326920
rect 154258 326868 154264 326920
rect 154316 326908 154322 326920
rect 326574 326908 326580 326920
rect 154316 326880 326580 326908
rect 154316 326868 154322 326880
rect 326574 326868 326580 326880
rect 326632 326868 326638 326920
rect 335682 326868 335688 326920
rect 335740 326908 335746 326920
rect 336786 326908 336792 326920
rect 335740 326880 336792 326908
rect 335740 326868 335746 326880
rect 336786 326868 336792 326880
rect 336844 326868 336850 326920
rect 345897 326911 345955 326917
rect 345897 326877 345909 326911
rect 345943 326908 345955 326911
rect 354358 326908 354364 326920
rect 345943 326880 354364 326908
rect 345943 326877 345955 326880
rect 345897 326871 345955 326877
rect 354358 326868 354364 326880
rect 354416 326868 354422 326920
rect 354453 326911 354511 326917
rect 354453 326877 354465 326911
rect 354499 326908 354511 326911
rect 363834 326908 363840 326920
rect 354499 326880 363840 326908
rect 354499 326877 354511 326880
rect 354453 326871 354511 326877
rect 363834 326868 363840 326880
rect 363892 326868 363898 326920
rect 153522 326800 153528 326852
rect 153580 326840 153586 326852
rect 167322 326840 167328 326852
rect 153580 326812 167328 326840
rect 153580 326800 153586 326812
rect 167322 326800 167328 326812
rect 167380 326800 167386 326852
rect 243130 326800 243136 326852
rect 243188 326840 243194 326852
rect 243188 326812 253112 326840
rect 243188 326800 243194 326812
rect 57198 326732 57204 326784
rect 57256 326772 57262 326784
rect 62258 326772 62264 326784
rect 57256 326744 62264 326772
rect 57256 326732 57262 326744
rect 62258 326732 62264 326744
rect 62316 326732 62322 326784
rect 152050 326732 152056 326784
rect 152108 326772 152114 326784
rect 166126 326772 166132 326784
rect 152108 326744 166132 326772
rect 152108 326732 152114 326744
rect 166126 326732 166132 326744
rect 166184 326732 166190 326784
rect 239542 326732 239548 326784
rect 239600 326772 239606 326784
rect 239600 326744 243912 326772
rect 239600 326732 239606 326744
rect 73853 326707 73911 326713
rect 73853 326673 73865 326707
rect 73899 326704 73911 326707
rect 74310 326704 74316 326716
rect 73899 326676 74316 326704
rect 73899 326673 73911 326676
rect 73853 326667 73911 326673
rect 74310 326664 74316 326676
rect 74368 326704 74374 326716
rect 76886 326704 76892 326716
rect 74368 326676 76892 326704
rect 74368 326664 74374 326676
rect 76886 326664 76892 326676
rect 76944 326664 76950 326716
rect 144598 326664 144604 326716
rect 144656 326704 144662 326716
rect 155546 326704 155552 326716
rect 144656 326676 155552 326704
rect 144656 326664 144662 326676
rect 155546 326664 155552 326676
rect 155604 326664 155610 326716
rect 156190 326664 156196 326716
rect 156248 326704 156254 326716
rect 169990 326704 169996 326716
rect 156248 326676 169996 326704
rect 156248 326664 156254 326676
rect 169990 326664 169996 326676
rect 170048 326664 170054 326716
rect 241934 326664 241940 326716
rect 241992 326704 241998 326716
rect 242762 326704 242768 326716
rect 241992 326676 242768 326704
rect 241992 326664 241998 326676
rect 242762 326664 242768 326676
rect 242820 326664 242826 326716
rect 243884 326704 243912 326744
rect 245890 326732 245896 326784
rect 245948 326772 245954 326784
rect 252977 326775 253035 326781
rect 252977 326772 252989 326775
rect 245948 326744 252989 326772
rect 245948 326732 245954 326744
rect 252977 326741 252989 326744
rect 253023 326741 253035 326775
rect 252977 326735 253035 326741
rect 250030 326704 250036 326716
rect 243884 326676 250036 326704
rect 250030 326664 250036 326676
rect 250088 326664 250094 326716
rect 253084 326704 253112 326812
rect 255458 326800 255464 326852
rect 255516 326840 255522 326852
rect 256286 326840 256292 326852
rect 255516 326812 256292 326840
rect 255516 326800 255522 326812
rect 256286 326800 256292 326812
rect 256344 326800 256350 326852
rect 256930 326800 256936 326852
rect 256988 326840 256994 326852
rect 262082 326840 262088 326852
rect 256988 326812 262088 326840
rect 256988 326800 256994 326812
rect 262082 326800 262088 326812
rect 262140 326800 262146 326852
rect 340834 326800 340840 326852
rect 340892 326840 340898 326852
rect 352797 326843 352855 326849
rect 352797 326840 352809 326843
rect 340892 326812 352809 326840
rect 340892 326800 340898 326812
rect 352797 326809 352809 326812
rect 352843 326809 352855 326843
rect 352797 326803 352855 326809
rect 253161 326775 253219 326781
rect 253161 326741 253173 326775
rect 253207 326772 253219 326775
rect 260150 326772 260156 326784
rect 253207 326744 260156 326772
rect 253207 326741 253219 326744
rect 253161 326735 253219 326741
rect 260150 326732 260156 326744
rect 260208 326732 260214 326784
rect 341570 326732 341576 326784
rect 341628 326772 341634 326784
rect 354174 326772 354180 326784
rect 341628 326744 354180 326772
rect 341628 326732 341634 326744
rect 354174 326732 354180 326744
rect 354232 326732 354238 326784
rect 257298 326704 257304 326716
rect 253084 326676 257304 326704
rect 257298 326664 257304 326676
rect 257356 326664 257362 326716
rect 343962 326664 343968 326716
rect 344020 326704 344026 326716
rect 356934 326704 356940 326716
rect 344020 326676 356940 326704
rect 344020 326664 344026 326676
rect 356934 326664 356940 326676
rect 356992 326664 356998 326716
rect 63362 326596 63368 326648
rect 63420 326636 63426 326648
rect 66766 326636 66772 326648
rect 63420 326608 66772 326636
rect 63420 326596 63426 326608
rect 66766 326596 66772 326608
rect 66824 326596 66830 326648
rect 145518 326596 145524 326648
rect 145576 326636 145582 326648
rect 157570 326636 157576 326648
rect 145576 326608 157576 326636
rect 145576 326596 145582 326608
rect 157570 326596 157576 326608
rect 157628 326596 157634 326648
rect 162357 326639 162415 326645
rect 162357 326605 162369 326639
rect 162403 326636 162415 326639
rect 169070 326636 169076 326648
rect 162403 326608 169076 326636
rect 162403 326605 162415 326608
rect 162357 326599 162415 326605
rect 169070 326596 169076 326608
rect 169128 326596 169134 326648
rect 246350 326596 246356 326648
rect 246408 326636 246414 326648
rect 258218 326636 258224 326648
rect 246408 326608 258224 326636
rect 246408 326596 246414 326608
rect 258218 326596 258224 326608
rect 258276 326596 258282 326648
rect 343226 326596 343232 326648
rect 343284 326636 343290 326648
rect 355646 326636 355652 326648
rect 343284 326608 355652 326636
rect 343284 326596 343290 326608
rect 355646 326596 355652 326608
rect 355704 326596 355710 326648
rect 58210 326528 58216 326580
rect 58268 326568 58274 326580
rect 62442 326568 62448 326580
rect 58268 326540 62448 326568
rect 58268 326528 58274 326540
rect 62442 326528 62448 326540
rect 62500 326528 62506 326580
rect 150394 326528 150400 326580
rect 150452 326568 150458 326580
rect 161618 326568 161624 326580
rect 150452 326540 161624 326568
rect 150452 326528 150458 326540
rect 161618 326528 161624 326540
rect 161676 326528 161682 326580
rect 337062 326528 337068 326580
rect 337120 326568 337126 326580
rect 338353 326571 338411 326577
rect 338353 326568 338365 326571
rect 337120 326540 338365 326568
rect 337120 326528 337126 326540
rect 338353 326537 338365 326540
rect 338399 326537 338411 326571
rect 338353 326531 338411 326537
rect 347921 326571 347979 326577
rect 347921 326537 347933 326571
rect 347967 326568 347979 326571
rect 348013 326571 348071 326577
rect 348013 326568 348025 326571
rect 347967 326540 348025 326568
rect 347967 326537 347979 326540
rect 347921 326531 347979 326537
rect 348013 326537 348025 326540
rect 348059 326537 348071 326571
rect 348013 326531 348071 326537
rect 29141 326503 29199 326509
rect 29141 326469 29153 326503
rect 29187 326500 29199 326503
rect 31993 326503 32051 326509
rect 31993 326500 32005 326503
rect 29187 326472 32005 326500
rect 29187 326469 29199 326472
rect 29141 326463 29199 326469
rect 31993 326469 32005 326472
rect 32039 326469 32051 326503
rect 31993 326463 32051 326469
rect 32085 326503 32143 326509
rect 32085 326469 32097 326503
rect 32131 326500 32143 326503
rect 32131 326472 38844 326500
rect 32131 326469 32143 326472
rect 32085 326463 32143 326469
rect 14694 326392 14700 326444
rect 14752 326432 14758 326444
rect 19573 326435 19631 326441
rect 19573 326432 19585 326435
rect 14752 326404 19585 326432
rect 14752 326392 14758 326404
rect 19573 326401 19585 326404
rect 19619 326401 19631 326435
rect 38816 326432 38844 326472
rect 148462 326460 148468 326512
rect 148520 326500 148526 326512
rect 160238 326500 160244 326512
rect 148520 326472 160244 326500
rect 148520 326460 148526 326472
rect 160238 326460 160244 326472
rect 160296 326460 160302 326512
rect 248834 326460 248840 326512
rect 248892 326500 248898 326512
rect 258221 326503 258279 326509
rect 258221 326500 258233 326503
rect 248892 326472 258233 326500
rect 248892 326460 248898 326472
rect 258221 326469 258233 326472
rect 258267 326469 258279 326503
rect 258221 326463 258279 326469
rect 345618 326460 345624 326512
rect 345676 326500 345682 326512
rect 345676 326472 350724 326500
rect 345676 326460 345682 326472
rect 58213 326435 58271 326441
rect 58213 326432 58225 326435
rect 38816 326404 58225 326432
rect 19573 326395 19631 326401
rect 58213 326401 58225 326404
rect 58259 326401 58271 326435
rect 58213 326395 58271 326401
rect 61338 326392 61344 326444
rect 61396 326432 61402 326444
rect 66398 326432 66404 326444
rect 61396 326404 66404 326432
rect 61396 326392 61402 326404
rect 66398 326392 66404 326404
rect 66456 326392 66462 326444
rect 147910 326392 147916 326444
rect 147968 326432 147974 326444
rect 148738 326432 148744 326444
rect 147968 326404 148744 326432
rect 147968 326392 147974 326404
rect 148738 326392 148744 326404
rect 148796 326392 148802 326444
rect 152326 326392 152332 326444
rect 152384 326432 152390 326444
rect 163090 326432 163096 326444
rect 152384 326404 163096 326432
rect 152384 326392 152390 326404
rect 163090 326392 163096 326404
rect 163148 326392 163154 326444
rect 338353 326435 338411 326441
rect 338353 326401 338365 326435
rect 338399 326432 338411 326435
rect 347921 326435 347979 326441
rect 347921 326432 347933 326435
rect 338399 326404 347933 326432
rect 338399 326401 338411 326404
rect 338353 326395 338411 326401
rect 347921 326401 347933 326404
rect 347967 326401 347979 326435
rect 347921 326395 347979 326401
rect 74034 326324 74040 326376
rect 74092 326364 74098 326376
rect 76058 326364 76064 326376
rect 74092 326336 76064 326364
rect 74092 326324 74098 326336
rect 76058 326324 76064 326336
rect 76116 326324 76122 326376
rect 145150 326324 145156 326376
rect 145208 326364 145214 326376
rect 145886 326364 145892 326376
rect 145208 326336 145892 326364
rect 145208 326324 145214 326336
rect 145886 326324 145892 326336
rect 145944 326324 145950 326376
rect 147450 326324 147456 326376
rect 147508 326364 147514 326376
rect 156926 326364 156932 326376
rect 147508 326336 156932 326364
rect 147508 326324 147514 326336
rect 156926 326324 156932 326336
rect 156984 326324 156990 326376
rect 242486 326324 242492 326376
rect 242544 326364 242550 326376
rect 250214 326364 250220 326376
rect 242544 326336 250220 326364
rect 242544 326324 242550 326336
rect 250214 326324 250220 326336
rect 250272 326324 250278 326376
rect 350696 326364 350724 326472
rect 354453 326367 354511 326373
rect 354453 326364 354465 326367
rect 350696 326336 354465 326364
rect 354453 326333 354465 326336
rect 354499 326333 354511 326367
rect 354453 326327 354511 326333
rect 19573 326299 19631 326305
rect 19573 326265 19585 326299
rect 19619 326296 19631 326299
rect 29141 326299 29199 326305
rect 29141 326296 29153 326299
rect 19619 326268 29153 326296
rect 19619 326265 19631 326268
rect 19573 326259 19631 326265
rect 29141 326265 29153 326268
rect 29187 326265 29199 326299
rect 29141 326259 29199 326265
rect 67781 326299 67839 326305
rect 67781 326265 67793 326299
rect 67827 326296 67839 326299
rect 73853 326299 73911 326305
rect 73853 326296 73865 326299
rect 67827 326268 73865 326296
rect 67827 326265 67839 326268
rect 67781 326259 67839 326265
rect 73853 326265 73865 326268
rect 73899 326265 73911 326299
rect 73853 326259 73911 326265
rect 75782 326256 75788 326308
rect 75840 326296 75846 326308
rect 76978 326296 76984 326308
rect 75840 326268 76984 326296
rect 75840 326256 75846 326268
rect 76978 326256 76984 326268
rect 77036 326256 77042 326308
rect 136870 326256 136876 326308
rect 136928 326296 136934 326308
rect 156282 326296 156288 326308
rect 136928 326268 156288 326296
rect 136928 326256 136934 326268
rect 156282 326256 156288 326268
rect 156340 326256 156346 326308
rect 161526 326256 161532 326308
rect 161584 326296 161590 326308
rect 162262 326296 162268 326308
rect 161584 326268 162268 326296
rect 161584 326256 161590 326268
rect 162262 326256 162268 326268
rect 162320 326256 162326 326308
rect 254906 326256 254912 326308
rect 254964 326296 254970 326308
rect 259230 326296 259236 326308
rect 254964 326268 259236 326296
rect 254964 326256 254970 326268
rect 259230 326256 259236 326268
rect 259288 326256 259294 326308
rect 137698 326228 137704 326240
rect 137659 326200 137704 326228
rect 137698 326188 137704 326200
rect 137756 326188 137762 326240
rect 58213 326163 58271 326169
rect 58213 326129 58225 326163
rect 58259 326160 58271 326163
rect 67781 326163 67839 326169
rect 67781 326160 67793 326163
rect 58259 326132 67793 326160
rect 58259 326129 58271 326132
rect 58213 326123 58271 326129
rect 67781 326129 67793 326132
rect 67827 326129 67839 326163
rect 67781 326123 67839 326129
rect 352797 325211 352855 325217
rect 352797 325177 352809 325211
rect 352843 325208 352855 325211
rect 352886 325208 352892 325220
rect 352843 325180 352892 325208
rect 352843 325177 352855 325180
rect 352797 325171 352855 325177
rect 352886 325168 352892 325180
rect 352944 325168 352950 325220
rect 325286 324828 325292 324880
rect 325344 324868 325350 324880
rect 343870 324868 343876 324880
rect 325344 324840 343876 324868
rect 325344 324828 325350 324840
rect 343870 324828 343876 324840
rect 343928 324868 343934 324880
rect 347182 324868 347188 324880
rect 343928 324840 347188 324868
rect 343928 324828 343934 324840
rect 347182 324828 347188 324840
rect 347240 324828 347246 324880
rect 210010 323468 210016 323520
rect 210068 323508 210074 323520
rect 211298 323508 211304 323520
rect 210068 323480 211304 323508
rect 210068 323468 210074 323480
rect 211298 323468 211304 323480
rect 211356 323468 211362 323520
rect 279102 323468 279108 323520
rect 279160 323508 279166 323520
rect 280298 323508 280304 323520
rect 279160 323480 280304 323508
rect 279160 323468 279166 323480
rect 280298 323468 280304 323480
rect 280356 323468 280362 323520
rect 291522 323468 291528 323520
rect 291580 323508 291586 323520
rect 292718 323508 292724 323520
rect 291580 323480 292724 323508
rect 291580 323468 291586 323480
rect 292718 323468 292724 323480
rect 292776 323468 292782 323520
rect 304034 323468 304040 323520
rect 304092 323508 304098 323520
rect 305138 323508 305144 323520
rect 304092 323480 305144 323508
rect 304092 323468 304098 323480
rect 305138 323468 305144 323480
rect 305196 323468 305202 323520
rect 324734 323468 324740 323520
rect 324792 323508 324798 323520
rect 325746 323508 325752 323520
rect 324792 323480 325752 323508
rect 324792 323468 324798 323480
rect 325746 323468 325752 323480
rect 325804 323508 325810 323520
rect 346998 323508 347004 323520
rect 325804 323480 347004 323508
rect 325804 323468 325810 323480
rect 346998 323468 347004 323480
rect 347056 323508 347062 323520
rect 351230 323508 351236 323520
rect 347056 323480 351236 323508
rect 347056 323468 347062 323480
rect 351230 323468 351236 323480
rect 351288 323468 351294 323520
rect 344330 323400 344336 323452
rect 344388 323440 344394 323452
rect 348010 323440 348016 323452
rect 344388 323412 348016 323440
rect 344388 323400 344394 323412
rect 348010 323400 348016 323412
rect 348068 323400 348074 323452
rect 325562 322108 325568 322160
rect 325620 322148 325626 322160
rect 344330 322148 344336 322160
rect 325620 322120 344336 322148
rect 325620 322108 325626 322120
rect 344330 322108 344336 322120
rect 344388 322108 344394 322160
rect 346446 322040 346452 322092
rect 346504 322080 346510 322092
rect 350402 322080 350408 322092
rect 346504 322052 350408 322080
rect 346504 322040 346510 322052
rect 350402 322040 350408 322052
rect 350460 322040 350466 322092
rect 395114 320748 395120 320800
rect 395172 320788 395178 320800
rect 395206 320788 395212 320800
rect 395172 320760 395212 320788
rect 395172 320748 395178 320760
rect 395206 320748 395212 320760
rect 395264 320748 395270 320800
rect 324826 320680 324832 320732
rect 324884 320720 324890 320732
rect 325654 320720 325660 320732
rect 324884 320692 325660 320720
rect 324884 320680 324890 320692
rect 325654 320680 325660 320692
rect 325712 320720 325718 320732
rect 346446 320720 346452 320732
rect 325712 320692 346452 320720
rect 325712 320680 325718 320692
rect 346446 320680 346452 320692
rect 346504 320680 346510 320732
rect 62258 320612 62264 320664
rect 62316 320652 62322 320664
rect 63270 320652 63276 320664
rect 62316 320624 63276 320652
rect 62316 320612 62322 320624
rect 63270 320612 63276 320624
rect 63328 320612 63334 320664
rect 248926 320612 248932 320664
rect 248984 320652 248990 320664
rect 256930 320652 256936 320664
rect 248984 320624 256936 320652
rect 248984 320612 248990 320624
rect 256930 320612 256936 320624
rect 256988 320612 256994 320664
rect 337154 320612 337160 320664
rect 337212 320652 337218 320664
rect 337522 320652 337528 320664
rect 337212 320624 337528 320652
rect 337212 320612 337218 320624
rect 337522 320612 337528 320624
rect 337580 320612 337586 320664
rect 339270 320612 339276 320664
rect 339328 320652 339334 320664
rect 339546 320652 339552 320664
rect 339328 320624 339552 320652
rect 339328 320612 339334 320624
rect 339546 320612 339552 320624
rect 339604 320612 339610 320664
rect 339914 320612 339920 320664
rect 339972 320652 339978 320664
rect 340558 320652 340564 320664
rect 339972 320624 340564 320652
rect 339972 320612 339978 320624
rect 340558 320612 340564 320624
rect 340616 320612 340622 320664
rect 66858 320584 66864 320596
rect 63472 320556 66864 320584
rect 58762 320476 58768 320528
rect 58820 320516 58826 320528
rect 63472 320516 63500 320556
rect 66858 320544 66864 320556
rect 66916 320544 66922 320596
rect 248742 320544 248748 320596
rect 248800 320584 248806 320596
rect 249202 320584 249208 320596
rect 248800 320556 249208 320584
rect 248800 320544 248806 320556
rect 249202 320544 249208 320556
rect 249260 320544 249266 320596
rect 346078 320544 346084 320596
rect 346136 320584 346142 320596
rect 349390 320584 349396 320596
rect 346136 320556 349396 320584
rect 346136 320544 346142 320556
rect 349390 320544 349396 320556
rect 349448 320544 349454 320596
rect 58820 320488 63500 320516
rect 58820 320476 58826 320488
rect 63638 320476 63644 320528
rect 63696 320516 63702 320528
rect 65018 320516 65024 320528
rect 63696 320488 65024 320516
rect 63696 320476 63702 320488
rect 65018 320476 65024 320488
rect 65076 320476 65082 320528
rect 336970 320476 336976 320528
rect 337028 320516 337034 320528
rect 351598 320516 351604 320528
rect 337028 320488 351604 320516
rect 337028 320476 337034 320488
rect 351598 320476 351604 320488
rect 351656 320476 351662 320528
rect 60602 320408 60608 320460
rect 60660 320448 60666 320460
rect 69066 320448 69072 320460
rect 60660 320420 69072 320448
rect 60660 320408 60666 320420
rect 69066 320408 69072 320420
rect 69124 320408 69130 320460
rect 338350 320408 338356 320460
rect 338408 320448 338414 320460
rect 352242 320448 352248 320460
rect 338408 320420 352248 320448
rect 338408 320408 338414 320420
rect 352242 320408 352248 320420
rect 352300 320408 352306 320460
rect 59682 320340 59688 320392
rect 59740 320380 59746 320392
rect 68422 320380 68428 320392
rect 59740 320352 68428 320380
rect 59740 320340 59746 320352
rect 68422 320340 68428 320352
rect 68480 320340 68486 320392
rect 247914 320340 247920 320392
rect 247972 320380 247978 320392
rect 257114 320380 257120 320392
rect 247972 320352 257120 320380
rect 247972 320340 247978 320352
rect 257114 320340 257120 320352
rect 257172 320340 257178 320392
rect 335590 320340 335596 320392
rect 335648 320380 335654 320392
rect 350678 320380 350684 320392
rect 335648 320352 350684 320380
rect 335648 320340 335654 320352
rect 350678 320340 350684 320352
rect 350736 320340 350742 320392
rect 57014 320272 57020 320324
rect 57072 320312 57078 320324
rect 66490 320312 66496 320324
rect 57072 320284 66496 320312
rect 57072 320272 57078 320284
rect 66490 320272 66496 320284
rect 66548 320272 66554 320324
rect 243130 320272 243136 320324
rect 243188 320312 243194 320324
rect 243774 320312 243780 320324
rect 243188 320284 243780 320312
rect 243188 320272 243194 320284
rect 243774 320272 243780 320284
rect 243832 320272 243838 320324
rect 245890 320272 245896 320324
rect 245948 320312 245954 320324
rect 246442 320312 246448 320324
rect 245948 320284 246448 320312
rect 245948 320272 245954 320284
rect 246442 320272 246448 320284
rect 246500 320272 246506 320324
rect 334210 320272 334216 320324
rect 334268 320312 334274 320324
rect 349758 320312 349764 320324
rect 334268 320284 349764 320312
rect 334268 320272 334274 320284
rect 349758 320272 349764 320284
rect 349816 320272 349822 320324
rect 56094 320204 56100 320256
rect 56152 320244 56158 320256
rect 66306 320244 66312 320256
rect 56152 320216 66312 320244
rect 56152 320204 56158 320216
rect 66306 320204 66312 320216
rect 66364 320204 66370 320256
rect 156926 320204 156932 320256
rect 156984 320244 156990 320256
rect 159962 320244 159968 320256
rect 156984 320216 159968 320244
rect 156984 320204 156990 320216
rect 159962 320204 159968 320216
rect 160020 320204 160026 320256
rect 246902 320204 246908 320256
rect 246960 320244 246966 320256
rect 256286 320244 256292 320256
rect 246960 320216 256292 320244
rect 246960 320204 246966 320216
rect 256286 320204 256292 320216
rect 256344 320204 256350 320256
rect 332830 320204 332836 320256
rect 332888 320244 332894 320256
rect 348010 320244 348016 320256
rect 332888 320216 348016 320244
rect 332888 320204 332894 320216
rect 348010 320204 348016 320216
rect 348068 320204 348074 320256
rect 62350 320136 62356 320188
rect 62408 320176 62414 320188
rect 74770 320176 74776 320188
rect 62408 320148 74776 320176
rect 62408 320136 62414 320148
rect 74770 320136 74776 320148
rect 74828 320136 74834 320188
rect 246258 320136 246264 320188
rect 246316 320176 246322 320188
rect 254906 320176 254912 320188
rect 246316 320148 254912 320176
rect 246316 320136 246322 320148
rect 254906 320136 254912 320148
rect 254964 320136 254970 320188
rect 331450 320136 331456 320188
rect 331508 320176 331514 320188
rect 347274 320176 347280 320188
rect 331508 320148 347280 320176
rect 331508 320136 331514 320148
rect 347274 320136 347280 320148
rect 347332 320136 347338 320188
rect 61430 320068 61436 320120
rect 61488 320108 61494 320120
rect 73390 320108 73396 320120
rect 61488 320080 73396 320108
rect 61488 320068 61494 320080
rect 73390 320068 73396 320080
rect 73448 320068 73454 320120
rect 149290 320068 149296 320120
rect 149348 320108 149354 320120
rect 161526 320108 161532 320120
rect 149348 320080 161532 320108
rect 149348 320068 149354 320080
rect 161526 320068 161532 320080
rect 161584 320068 161590 320120
rect 243590 320068 243596 320120
rect 243648 320108 243654 320120
rect 255458 320108 255464 320120
rect 243648 320080 255464 320108
rect 243648 320068 243654 320080
rect 255458 320068 255464 320080
rect 255516 320068 255522 320120
rect 335682 320068 335688 320120
rect 335740 320108 335746 320120
rect 350954 320108 350960 320120
rect 335740 320080 350960 320108
rect 335740 320068 335746 320080
rect 350954 320068 350960 320080
rect 351012 320068 351018 320120
rect 55266 320000 55272 320052
rect 55324 320040 55330 320052
rect 66674 320040 66680 320052
rect 55324 320012 66680 320040
rect 55324 320000 55330 320012
rect 66674 320000 66680 320012
rect 66732 320000 66738 320052
rect 147910 320000 147916 320052
rect 147968 320040 147974 320052
rect 147968 320012 152832 320040
rect 147968 320000 147974 320012
rect 57934 319932 57940 319984
rect 57992 319972 57998 319984
rect 69342 319972 69348 319984
rect 57992 319944 69348 319972
rect 57992 319932 57998 319944
rect 69342 319932 69348 319944
rect 69400 319932 69406 319984
rect 62442 319864 62448 319916
rect 62500 319904 62506 319916
rect 64098 319904 64104 319916
rect 62500 319876 64104 319904
rect 62500 319864 62506 319876
rect 64098 319864 64104 319876
rect 64156 319864 64162 319916
rect 145150 319864 145156 319916
rect 145208 319904 145214 319916
rect 152804 319904 152832 320012
rect 238990 320000 238996 320052
rect 239048 320040 239054 320052
rect 252790 320040 252796 320052
rect 239048 320012 252796 320040
rect 239048 320000 239054 320012
rect 252790 320000 252796 320012
rect 252848 320000 252854 320052
rect 334302 320000 334308 320052
rect 334360 320040 334366 320052
rect 349390 320040 349396 320052
rect 334360 320012 349396 320040
rect 334360 320000 334366 320012
rect 349390 320000 349396 320012
rect 349448 320000 349454 320052
rect 241934 319932 241940 319984
rect 241992 319972 241998 319984
rect 255550 319972 255556 319984
rect 241992 319944 255556 319972
rect 241992 319932 241998 319944
rect 255550 319932 255556 319944
rect 255608 319932 255614 319984
rect 332922 319932 332928 319984
rect 332980 319972 332986 319984
rect 348562 319972 348568 319984
rect 332980 319944 348568 319972
rect 332980 319932 332986 319944
rect 348562 319932 348568 319944
rect 348620 319932 348626 319984
rect 161710 319904 161716 319916
rect 145208 319876 152648 319904
rect 152804 319876 161716 319904
rect 145208 319864 145214 319876
rect 66766 319796 66772 319848
rect 66824 319836 66830 319848
rect 68606 319836 68612 319848
rect 66824 319808 68612 319836
rect 66824 319796 66830 319808
rect 68606 319796 68612 319808
rect 68664 319796 68670 319848
rect 152620 319768 152648 319876
rect 161710 319864 161716 319876
rect 161768 319864 161774 319916
rect 250214 319864 250220 319916
rect 250272 319904 250278 319916
rect 254446 319904 254452 319916
rect 250272 319876 254452 319904
rect 250272 319864 250278 319876
rect 254446 319864 254452 319876
rect 254504 319864 254510 319916
rect 159042 319768 159048 319780
rect 152620 319740 159048 319768
rect 159042 319728 159048 319740
rect 159100 319728 159106 319780
rect 250030 319728 250036 319780
rect 250088 319768 250094 319780
rect 251778 319768 251784 319780
rect 250088 319740 251784 319768
rect 250088 319728 250094 319740
rect 251778 319728 251784 319740
rect 251836 319728 251842 319780
rect 338534 319592 338540 319644
rect 338592 319632 338598 319644
rect 339546 319632 339552 319644
rect 338592 319604 339552 319632
rect 338592 319592 338598 319604
rect 339546 319592 339552 319604
rect 339604 319592 339610 319644
rect 249938 319456 249944 319508
rect 249996 319496 250002 319508
rect 250950 319496 250956 319508
rect 249996 319468 250956 319496
rect 249996 319456 250002 319468
rect 250950 319456 250956 319468
rect 251008 319456 251014 319508
rect 341128 319400 341892 319428
rect 65110 319320 65116 319372
rect 65168 319360 65174 319372
rect 65938 319360 65944 319372
rect 65168 319332 65944 319360
rect 65168 319320 65174 319332
rect 65938 319320 65944 319332
rect 65996 319320 66002 319372
rect 152050 319320 152056 319372
rect 152108 319360 152114 319372
rect 152786 319360 152792 319372
rect 152108 319332 152792 319360
rect 152108 319320 152114 319332
rect 152786 319320 152792 319332
rect 152844 319320 152850 319372
rect 155546 319320 155552 319372
rect 155604 319360 155610 319372
rect 157294 319360 157300 319372
rect 155604 319332 157300 319360
rect 155604 319320 155610 319332
rect 157294 319320 157300 319332
rect 157352 319320 157358 319372
rect 161618 319320 161624 319372
rect 161676 319360 161682 319372
rect 162630 319360 162636 319372
rect 161676 319332 162636 319360
rect 161676 319320 161682 319332
rect 162630 319320 162636 319332
rect 162688 319320 162694 319372
rect 325378 319320 325384 319372
rect 325436 319360 325442 319372
rect 341128 319360 341156 319400
rect 325436 319332 341156 319360
rect 325436 319320 325442 319332
rect 341202 319320 341208 319372
rect 341260 319360 341266 319372
rect 341754 319360 341760 319372
rect 341260 319332 341760 319360
rect 341260 319320 341266 319332
rect 341754 319320 341760 319332
rect 341812 319320 341818 319372
rect 341864 319360 341892 319400
rect 345158 319360 345164 319372
rect 341864 319332 345164 319360
rect 345158 319320 345164 319332
rect 345216 319360 345222 319372
rect 348102 319360 348108 319372
rect 345216 319332 348108 319360
rect 345216 319320 345222 319332
rect 348102 319320 348108 319332
rect 348160 319320 348166 319372
rect 163090 318504 163096 318556
rect 163148 318544 163154 318556
rect 164102 318544 164108 318556
rect 163148 318516 164108 318544
rect 163148 318504 163154 318516
rect 164102 318504 164108 318516
rect 164160 318504 164166 318556
rect 231078 317892 231084 317944
rect 231136 317932 231142 317944
rect 231354 317932 231360 317944
rect 231136 317904 231360 317932
rect 231136 317892 231142 317904
rect 231354 317892 231360 317904
rect 231412 317932 231418 317944
rect 246166 317932 246172 317944
rect 231412 317904 246172 317932
rect 231412 317892 231418 317904
rect 246166 317892 246172 317904
rect 246224 317932 246230 317944
rect 254814 317932 254820 317944
rect 246224 317904 254820 317932
rect 246224 317892 246230 317904
rect 254814 317892 254820 317904
rect 254872 317892 254878 317944
rect 137701 316643 137759 316649
rect 137701 316609 137713 316643
rect 137747 316640 137759 316643
rect 137790 316640 137796 316652
rect 137747 316612 137796 316640
rect 137747 316609 137759 316612
rect 137701 316603 137759 316609
rect 137790 316600 137796 316612
rect 137848 316600 137854 316652
rect 325470 316600 325476 316652
rect 325528 316640 325534 316652
rect 343042 316640 343048 316652
rect 325528 316612 343048 316640
rect 325528 316600 325534 316612
rect 343042 316600 343048 316612
rect 343100 316640 343106 316652
rect 429430 316640 429436 316652
rect 343100 316612 429436 316640
rect 343100 316600 343106 316612
rect 429430 316600 429436 316612
rect 429488 316600 429494 316652
rect 38798 315852 38804 315904
rect 38856 315892 38862 315904
rect 55082 315892 55088 315904
rect 38856 315864 55088 315892
rect 38856 315852 38862 315864
rect 55082 315852 55088 315864
rect 55140 315852 55146 315904
rect 357670 315852 357676 315904
rect 357728 315892 357734 315904
rect 358314 315892 358320 315904
rect 357728 315864 358320 315892
rect 357728 315852 357734 315864
rect 358314 315852 358320 315864
rect 358372 315892 358378 315904
rect 405970 315892 405976 315904
rect 358372 315864 405976 315892
rect 358372 315852 358378 315864
rect 405970 315852 405976 315864
rect 406028 315852 406034 315904
rect 352886 315172 352892 315224
rect 352944 315212 352950 315224
rect 353070 315212 353076 315224
rect 352944 315184 353076 315212
rect 352944 315172 352950 315184
rect 353070 315172 353076 315184
rect 353128 315172 353134 315224
rect 38430 313744 38436 313796
rect 38488 313784 38494 313796
rect 51586 313784 51592 313796
rect 38488 313756 51592 313784
rect 38488 313744 38494 313756
rect 51586 313744 51592 313756
rect 51644 313744 51650 313796
rect 356198 313744 356204 313796
rect 356256 313784 356262 313796
rect 405970 313784 405976 313796
rect 356256 313756 405976 313784
rect 356256 313744 356262 313756
rect 405970 313744 405976 313756
rect 406028 313744 406034 313796
rect 76978 313540 76984 313592
rect 77036 313580 77042 313592
rect 81670 313580 81676 313592
rect 77036 313552 81676 313580
rect 77036 313540 77042 313552
rect 81670 313540 81676 313552
rect 81728 313540 81734 313592
rect 165114 313064 165120 313116
rect 165172 313104 165178 313116
rect 175510 313104 175516 313116
rect 165172 313076 175516 313104
rect 165172 313064 165178 313076
rect 175510 313064 175516 313076
rect 175568 313064 175574 313116
rect 258954 313064 258960 313116
rect 259012 313104 259018 313116
rect 270270 313104 270276 313116
rect 259012 313076 270276 313104
rect 259012 313064 259018 313076
rect 270270 313064 270276 313076
rect 270328 313064 270334 313116
rect 76150 312452 76156 312504
rect 76208 312492 76214 312504
rect 76978 312492 76984 312504
rect 76208 312464 76984 312492
rect 76208 312452 76214 312464
rect 76978 312452 76984 312464
rect 77036 312452 77042 312504
rect 137790 311092 137796 311144
rect 137848 311092 137854 311144
rect 136962 310820 136968 310872
rect 137020 310860 137026 310872
rect 137808 310860 137836 311092
rect 395022 311024 395028 311076
rect 395080 311064 395086 311076
rect 395206 311064 395212 311076
rect 395080 311036 395212 311064
rect 395080 311024 395086 311036
rect 395206 311024 395212 311036
rect 395264 311024 395270 311076
rect 137020 310832 137836 310860
rect 137020 310820 137026 310832
rect 38798 310276 38804 310328
rect 38856 310316 38862 310328
rect 54070 310316 54076 310328
rect 38856 310288 54076 310316
rect 38856 310276 38862 310288
rect 54070 310276 54076 310288
rect 54128 310276 54134 310328
rect 356934 310276 356940 310328
rect 356992 310316 356998 310328
rect 405970 310316 405976 310328
rect 356992 310288 405976 310316
rect 356992 310276 356998 310288
rect 405970 310276 405976 310288
rect 406028 310276 406034 310328
rect 137698 309664 137704 309716
rect 137756 309704 137762 309716
rect 145518 309704 145524 309716
rect 137756 309676 145524 309704
rect 137756 309664 137762 309676
rect 145518 309664 145524 309676
rect 145576 309664 145582 309716
rect 231446 309664 231452 309716
rect 231504 309704 231510 309716
rect 240646 309704 240652 309716
rect 231504 309676 240652 309704
rect 231504 309664 231510 309676
rect 240646 309664 240652 309676
rect 240704 309664 240710 309716
rect 325378 309664 325384 309716
rect 325436 309704 325442 309716
rect 334210 309704 334216 309716
rect 325436 309676 334216 309704
rect 325436 309664 325442 309676
rect 334210 309664 334216 309676
rect 334268 309664 334274 309716
rect 356290 309664 356296 309716
rect 356348 309704 356354 309716
rect 356934 309704 356940 309716
rect 356348 309676 356940 309704
rect 356348 309664 356354 309676
rect 356934 309664 356940 309676
rect 356992 309664 356998 309716
rect 38798 308236 38804 308288
rect 38856 308276 38862 308288
rect 51218 308276 51224 308288
rect 38856 308248 51224 308276
rect 38856 308236 38862 308248
rect 51218 308236 51224 308248
rect 51276 308236 51282 308288
rect 136410 308236 136416 308288
rect 136468 308276 136474 308288
rect 136962 308276 136968 308288
rect 136468 308248 136968 308276
rect 136468 308236 136474 308248
rect 136962 308236 136968 308248
rect 137020 308236 137026 308288
rect 356198 308236 356204 308288
rect 356256 308276 356262 308288
rect 405970 308276 405976 308288
rect 356256 308248 405976 308276
rect 356256 308236 356262 308248
rect 405970 308236 405976 308248
rect 406028 308236 406034 308288
rect 352702 306876 352708 306928
rect 352760 306916 352766 306928
rect 352886 306916 352892 306928
rect 352760 306888 352892 306916
rect 352760 306876 352766 306888
rect 352886 306876 352892 306888
rect 352944 306876 352950 306928
rect 38798 306196 38804 306248
rect 38856 306236 38862 306248
rect 54070 306236 54076 306248
rect 38856 306208 54076 306236
rect 38856 306196 38862 306208
rect 54070 306196 54076 306208
rect 54128 306196 54134 306248
rect 354910 306196 354916 306248
rect 354968 306236 354974 306248
rect 355646 306236 355652 306248
rect 354968 306208 355652 306236
rect 354968 306196 354974 306208
rect 355646 306196 355652 306208
rect 355704 306236 355710 306248
rect 406062 306236 406068 306248
rect 355704 306208 406068 306236
rect 355704 306196 355710 306208
rect 406062 306196 406068 306208
rect 406120 306196 406126 306248
rect 73390 305380 73396 305432
rect 73448 305420 73454 305432
rect 75506 305420 75512 305432
rect 73448 305392 75512 305420
rect 73448 305380 73454 305392
rect 75506 305380 75512 305392
rect 75564 305380 75570 305432
rect 51862 304196 51868 304208
rect 49764 304168 51868 304196
rect 38614 304088 38620 304140
rect 38672 304128 38678 304140
rect 49764 304128 49792 304168
rect 51862 304156 51868 304168
rect 51920 304156 51926 304208
rect 232090 304156 232096 304208
rect 232148 304196 232154 304208
rect 232734 304196 232740 304208
rect 232148 304168 232740 304196
rect 232148 304156 232154 304168
rect 232734 304156 232740 304168
rect 232792 304156 232798 304208
rect 38672 304100 49792 304128
rect 38672 304088 38678 304100
rect 356198 304088 356204 304140
rect 356256 304128 356262 304140
rect 405970 304128 405976 304140
rect 356256 304100 405976 304128
rect 356256 304088 356262 304100
rect 405970 304088 405976 304100
rect 406028 304088 406034 304140
rect 231998 301368 232004 301420
rect 232056 301408 232062 301420
rect 233470 301408 233476 301420
rect 232056 301380 233476 301408
rect 232056 301368 232062 301380
rect 233470 301368 233476 301380
rect 233528 301408 233534 301420
rect 234114 301408 234120 301420
rect 233528 301380 234120 301408
rect 233528 301368 233534 301380
rect 234114 301368 234120 301380
rect 234172 301368 234178 301420
rect 38798 300620 38804 300672
rect 38856 300660 38862 300672
rect 50298 300660 50304 300672
rect 38856 300632 50304 300660
rect 38856 300620 38862 300632
rect 50298 300620 50304 300632
rect 50356 300620 50362 300672
rect 355554 300620 355560 300672
rect 355612 300660 355618 300672
rect 405970 300660 405976 300672
rect 355612 300632 405976 300660
rect 355612 300620 355618 300632
rect 405970 300620 405976 300632
rect 406028 300620 406034 300672
rect 355002 300008 355008 300060
rect 355060 300048 355066 300060
rect 355554 300048 355560 300060
rect 355060 300020 355560 300048
rect 355060 300008 355066 300020
rect 355554 300008 355560 300020
rect 355612 300008 355618 300060
rect 136410 298648 136416 298700
rect 136468 298688 136474 298700
rect 136870 298688 136876 298700
rect 136468 298660 136876 298688
rect 136468 298648 136474 298660
rect 136870 298648 136876 298660
rect 136928 298648 136934 298700
rect 38246 298580 38252 298632
rect 38304 298620 38310 298632
rect 51678 298620 51684 298632
rect 38304 298592 51684 298620
rect 38304 298580 38310 298592
rect 51678 298580 51684 298592
rect 51736 298580 51742 298632
rect 356198 298580 356204 298632
rect 356256 298620 356262 298632
rect 405970 298620 405976 298632
rect 356256 298592 405976 298620
rect 356256 298580 356262 298592
rect 405970 298580 405976 298592
rect 406028 298580 406034 298632
rect 74218 297152 74224 297204
rect 74276 297192 74282 297204
rect 81670 297192 81676 297204
rect 74276 297164 81676 297192
rect 74276 297152 74282 297164
rect 81670 297152 81676 297164
rect 81728 297152 81734 297204
rect 167874 297152 167880 297204
rect 167932 297192 167938 297204
rect 175510 297192 175516 297204
rect 167932 297164 175516 297192
rect 167932 297152 167938 297164
rect 175510 297152 175516 297164
rect 175568 297152 175574 297204
rect 261714 297152 261720 297204
rect 261772 297192 261778 297204
rect 269350 297192 269356 297204
rect 261772 297164 269356 297192
rect 261772 297152 261778 297164
rect 269350 297152 269356 297164
rect 269408 297152 269414 297204
rect 137790 295860 137796 295912
rect 137848 295900 137854 295912
rect 145426 295900 145432 295912
rect 137848 295872 145432 295900
rect 137848 295860 137854 295872
rect 145426 295860 145432 295872
rect 145484 295860 145490 295912
rect 231538 295860 231544 295912
rect 231596 295900 231602 295912
rect 240922 295900 240928 295912
rect 231596 295872 240928 295900
rect 231596 295860 231602 295872
rect 240922 295860 240928 295872
rect 240980 295860 240986 295912
rect 325470 295860 325476 295912
rect 325528 295900 325534 295912
rect 334210 295900 334216 295912
rect 325528 295872 334216 295900
rect 325528 295860 325534 295872
rect 334210 295860 334216 295872
rect 334268 295860 334274 295912
rect 353530 295792 353536 295844
rect 353588 295832 353594 295844
rect 354174 295832 354180 295844
rect 353588 295804 354180 295832
rect 353588 295792 353594 295804
rect 354174 295792 354180 295804
rect 354232 295792 354238 295844
rect 38798 295112 38804 295164
rect 38856 295152 38862 295164
rect 51310 295152 51316 295164
rect 38856 295124 51316 295152
rect 38856 295112 38862 295124
rect 51310 295112 51316 295124
rect 51368 295112 51374 295164
rect 353530 295112 353536 295164
rect 353588 295152 353594 295164
rect 405970 295152 405976 295164
rect 353588 295124 405976 295152
rect 353588 295112 353594 295124
rect 405970 295112 405976 295124
rect 406028 295112 406034 295164
rect 38430 293752 38436 293804
rect 38488 293792 38494 293804
rect 52598 293792 52604 293804
rect 38488 293764 52604 293792
rect 38488 293752 38494 293764
rect 52598 293752 52604 293764
rect 52656 293752 52662 293804
rect 356198 293752 356204 293804
rect 356256 293792 356262 293804
rect 405970 293792 405976 293804
rect 356256 293764 405976 293792
rect 356256 293752 356262 293764
rect 405970 293752 405976 293764
rect 406028 293752 406034 293804
rect 427866 293208 427872 293260
rect 427924 293248 427930 293260
rect 428786 293248 428792 293260
rect 427924 293220 428792 293248
rect 427924 293208 427930 293220
rect 428786 293208 428792 293220
rect 428844 293208 428850 293260
rect 427682 293140 427688 293192
rect 427740 293180 427746 293192
rect 429890 293180 429896 293192
rect 427740 293152 429896 293180
rect 427740 293140 427746 293152
rect 429890 293140 429896 293152
rect 429948 293140 429954 293192
rect 352702 291752 352708 291764
rect 352663 291724 352708 291752
rect 352702 291712 352708 291724
rect 352760 291712 352766 291764
rect 395022 291712 395028 291764
rect 395080 291752 395086 291764
rect 395206 291752 395212 291764
rect 395080 291724 395212 291752
rect 395080 291712 395086 291724
rect 395206 291712 395212 291724
rect 395264 291712 395270 291764
rect 38522 291644 38528 291696
rect 38580 291684 38586 291696
rect 50022 291684 50028 291696
rect 38580 291656 50028 291684
rect 38580 291644 38586 291656
rect 50022 291644 50028 291656
rect 50080 291644 50086 291696
rect 50022 291236 50028 291288
rect 50080 291276 50086 291288
rect 51494 291276 51500 291288
rect 50080 291248 51500 291276
rect 50080 291236 50086 291248
rect 51494 291236 51500 291248
rect 51552 291236 51558 291288
rect 386653 291279 386711 291285
rect 386653 291245 386665 291279
rect 386699 291276 386711 291279
rect 396221 291279 396279 291285
rect 396221 291276 396233 291279
rect 386699 291248 396233 291276
rect 386699 291245 386711 291248
rect 386653 291239 386711 291245
rect 396221 291245 396233 291248
rect 396267 291245 396279 291279
rect 396221 291239 396279 291245
rect 367333 291211 367391 291217
rect 367333 291177 367345 291211
rect 367379 291208 367391 291211
rect 376901 291211 376959 291217
rect 376901 291208 376913 291211
rect 367379 291180 376913 291208
rect 367379 291177 367391 291180
rect 367333 291171 367391 291177
rect 376901 291177 376913 291180
rect 376947 291177 376959 291211
rect 376901 291171 376959 291177
rect 379845 291143 379903 291149
rect 379845 291109 379857 291143
rect 379891 291140 379903 291143
rect 386653 291143 386711 291149
rect 386653 291140 386665 291143
rect 379891 291112 386665 291140
rect 379891 291109 379903 291112
rect 379845 291103 379903 291109
rect 386653 291109 386665 291112
rect 386699 291109 386711 291143
rect 386653 291103 386711 291109
rect 362457 291075 362515 291081
rect 362457 291041 362469 291075
rect 362503 291072 362515 291075
rect 367333 291075 367391 291081
rect 367333 291072 367345 291075
rect 362503 291044 367345 291072
rect 362503 291041 362515 291044
rect 362457 291035 362515 291041
rect 367333 291041 367345 291044
rect 367379 291041 367391 291075
rect 367333 291035 367391 291041
rect 396221 291075 396279 291081
rect 396221 291041 396233 291075
rect 396267 291072 396279 291075
rect 398981 291075 399039 291081
rect 398981 291072 398993 291075
rect 396267 291044 398993 291072
rect 396267 291041 396279 291044
rect 396221 291035 396279 291041
rect 398981 291041 398993 291044
rect 399027 291041 399039 291075
rect 398981 291035 399039 291041
rect 399073 291075 399131 291081
rect 399073 291041 399085 291075
rect 399119 291072 399131 291075
rect 399119 291044 400312 291072
rect 399119 291041 399131 291044
rect 399073 291035 399131 291041
rect 352705 291007 352763 291013
rect 352705 290973 352717 291007
rect 352751 291004 352763 291007
rect 352981 291007 353039 291013
rect 352981 291004 352993 291007
rect 352751 290976 352993 291004
rect 352751 290973 352763 290976
rect 352705 290967 352763 290973
rect 352981 290973 352993 290976
rect 353027 291004 353039 291007
rect 357673 291007 357731 291013
rect 357673 291004 357685 291007
rect 353027 290976 357685 291004
rect 353027 290973 353039 290976
rect 352981 290967 353039 290973
rect 357673 290973 357685 290976
rect 357719 290973 357731 291007
rect 357673 290967 357731 290973
rect 376901 291007 376959 291013
rect 376901 290973 376913 291007
rect 376947 291004 376959 291007
rect 379661 291007 379719 291013
rect 379661 291004 379673 291007
rect 376947 290976 379673 291004
rect 376947 290973 376959 290976
rect 376901 290967 376959 290973
rect 379661 290973 379673 290976
rect 379707 290973 379719 291007
rect 400284 291004 400312 291044
rect 405970 291004 405976 291016
rect 400284 290976 405976 291004
rect 379661 290967 379719 290973
rect 405970 290964 405976 290976
rect 406028 290964 406034 291016
rect 357673 290871 357731 290877
rect 357673 290837 357685 290871
rect 357719 290868 357731 290871
rect 362457 290871 362515 290877
rect 362457 290868 362469 290871
rect 357719 290840 362469 290868
rect 357719 290837 357731 290840
rect 357673 290831 357731 290837
rect 362457 290837 362469 290840
rect 362503 290837 362515 290871
rect 362457 290831 362515 290837
rect 230710 289060 230716 289112
rect 230768 289100 230774 289112
rect 236046 289100 236052 289112
rect 230768 289072 236052 289100
rect 230768 289060 230774 289072
rect 236046 289060 236052 289072
rect 236104 289060 236110 289112
rect 54530 289032 54536 289044
rect 48568 289004 54536 289032
rect 38522 288924 38528 288976
rect 38580 288964 38586 288976
rect 48568 288964 48596 289004
rect 54530 288992 54536 289004
rect 54588 288992 54594 289044
rect 38580 288936 48596 288964
rect 38580 288924 38586 288936
rect 356198 288924 356204 288976
rect 356256 288964 356262 288976
rect 405970 288964 405976 288976
rect 356256 288936 405976 288964
rect 356256 288924 356262 288936
rect 405970 288924 405976 288936
rect 406028 288924 406034 288976
rect 395114 288896 395120 288908
rect 395075 288868 395120 288896
rect 395114 288856 395120 288868
rect 395172 288856 395178 288908
rect 261714 286544 261720 286596
rect 261772 286584 261778 286596
rect 266590 286584 266596 286596
rect 261772 286556 266596 286584
rect 261772 286544 261778 286556
rect 266590 286544 266596 286556
rect 266648 286544 266654 286596
rect 168058 286204 168064 286256
rect 168116 286244 168122 286256
rect 172750 286244 172756 286256
rect 168116 286216 172756 286244
rect 168116 286204 168122 286216
rect 172750 286204 172756 286216
rect 172808 286204 172814 286256
rect 38522 285456 38528 285508
rect 38580 285496 38586 285508
rect 49930 285496 49936 285508
rect 38580 285468 49936 285496
rect 38580 285456 38586 285468
rect 49930 285456 49936 285468
rect 49988 285456 49994 285508
rect 353714 285456 353720 285508
rect 353772 285496 353778 285508
rect 405970 285496 405976 285508
rect 353772 285468 405976 285496
rect 353772 285456 353778 285468
rect 405970 285456 405976 285468
rect 406028 285456 406034 285508
rect 427958 283552 427964 283604
rect 428016 283592 428022 283604
rect 429430 283592 429436 283604
rect 428016 283564 429436 283592
rect 428016 283552 428022 283564
rect 429430 283552 429436 283564
rect 429488 283552 429494 283604
rect 141654 283484 141660 283536
rect 141712 283524 141718 283536
rect 145610 283524 145616 283536
rect 141712 283496 145616 283524
rect 141712 283484 141718 283496
rect 145610 283484 145616 283496
rect 145668 283484 145674 283536
rect 231814 283484 231820 283536
rect 231872 283524 231878 283536
rect 240922 283524 240928 283536
rect 231872 283496 240928 283524
rect 231872 283484 231878 283496
rect 240922 283484 240928 283496
rect 240980 283484 240986 283536
rect 325194 283484 325200 283536
rect 325252 283524 325258 283536
rect 334210 283524 334216 283536
rect 325252 283496 334216 283524
rect 325252 283484 325258 283496
rect 334210 283484 334216 283496
rect 334268 283484 334274 283536
rect 38522 283416 38528 283468
rect 38580 283456 38586 283468
rect 52046 283456 52052 283468
rect 38580 283428 52052 283456
rect 38580 283416 38586 283428
rect 52046 283416 52052 283428
rect 52104 283416 52110 283468
rect 356198 283416 356204 283468
rect 356256 283456 356262 283468
rect 405970 283456 405976 283468
rect 356256 283428 405976 283456
rect 356256 283416 356262 283428
rect 405970 283416 405976 283428
rect 406028 283416 406034 283468
rect 231630 282804 231636 282856
rect 231688 282844 231694 282856
rect 236230 282844 236236 282856
rect 231688 282816 236236 282844
rect 231688 282804 231694 282816
rect 236230 282804 236236 282816
rect 236288 282804 236294 282856
rect 324550 282736 324556 282788
rect 324608 282776 324614 282788
rect 330070 282776 330076 282788
rect 324608 282748 330076 282776
rect 324608 282736 324614 282748
rect 330070 282736 330076 282748
rect 330128 282736 330134 282788
rect 136870 282328 136876 282380
rect 136928 282368 136934 282380
rect 142390 282368 142396 282380
rect 136928 282340 142396 282368
rect 136928 282328 136934 282340
rect 142390 282328 142396 282340
rect 142448 282368 142454 282380
rect 143034 282368 143040 282380
rect 142448 282340 143040 282368
rect 142448 282328 142454 282340
rect 143034 282328 143040 282340
rect 143092 282328 143098 282380
rect 236230 282056 236236 282108
rect 236288 282096 236294 282108
rect 236874 282096 236880 282108
rect 236288 282068 236880 282096
rect 236288 282056 236294 282068
rect 236874 282056 236880 282068
rect 236932 282056 236938 282108
rect 395117 282099 395175 282105
rect 395117 282065 395129 282099
rect 395163 282096 395175 282099
rect 395298 282096 395304 282108
rect 395163 282068 395304 282096
rect 395163 282065 395175 282068
rect 395117 282059 395175 282065
rect 395298 282056 395304 282068
rect 395356 282056 395362 282108
rect 74126 280628 74132 280680
rect 74184 280668 74190 280680
rect 81670 280668 81676 280680
rect 74184 280640 81676 280668
rect 74184 280628 74190 280640
rect 81670 280628 81676 280640
rect 81728 280628 81734 280680
rect 172750 280628 172756 280680
rect 172808 280668 172814 280680
rect 175786 280668 175792 280680
rect 172808 280640 175792 280668
rect 172808 280628 172814 280640
rect 175786 280628 175792 280640
rect 175844 280628 175850 280680
rect 266590 280628 266596 280680
rect 266648 280668 266654 280680
rect 270270 280668 270276 280680
rect 266648 280640 270276 280668
rect 266648 280628 266654 280640
rect 270270 280628 270276 280640
rect 270328 280628 270334 280680
rect 38062 279948 38068 280000
rect 38120 279988 38126 280000
rect 48550 279988 48556 280000
rect 38120 279960 48556 279988
rect 38120 279948 38126 279960
rect 48550 279948 48556 279960
rect 48608 279948 48614 280000
rect 13590 279336 13596 279388
rect 13648 279376 13654 279388
rect 18098 279376 18104 279388
rect 13648 279348 18104 279376
rect 13648 279336 13654 279348
rect 18098 279336 18104 279348
rect 18156 279336 18162 279388
rect 352978 279376 352984 279388
rect 352939 279348 352984 279376
rect 352978 279336 352984 279348
rect 353036 279336 353042 279388
rect 38614 279268 38620 279320
rect 38672 279308 38678 279320
rect 52598 279308 52604 279320
rect 38672 279280 52604 279308
rect 38672 279268 38678 279280
rect 52598 279268 52604 279280
rect 52656 279268 52662 279320
rect 356198 279268 356204 279320
rect 356256 279308 356262 279320
rect 405970 279308 405976 279320
rect 356256 279280 405976 279308
rect 356256 279268 356262 279280
rect 405970 279268 405976 279280
rect 406028 279268 406034 279320
rect 395114 279200 395120 279252
rect 395172 279240 395178 279252
rect 395298 279240 395304 279252
rect 395172 279212 395304 279240
rect 395172 279200 395178 279212
rect 395298 279200 395304 279212
rect 395356 279200 395362 279252
rect 51494 277908 51500 277960
rect 51552 277948 51558 277960
rect 51678 277948 51684 277960
rect 51552 277920 51684 277948
rect 51552 277908 51558 277920
rect 51678 277908 51684 277920
rect 51736 277908 51742 277960
rect 137514 275120 137520 275172
rect 137572 275160 137578 275172
rect 155914 275160 155920 275172
rect 137572 275132 155920 275160
rect 137572 275120 137578 275132
rect 155914 275120 155920 275132
rect 155972 275120 155978 275172
rect 234114 275120 234120 275172
rect 234172 275160 234178 275172
rect 249110 275160 249116 275172
rect 234172 275132 249116 275160
rect 234172 275120 234178 275132
rect 249110 275120 249116 275132
rect 249168 275120 249174 275172
rect 138618 275052 138624 275104
rect 138676 275092 138682 275104
rect 155270 275092 155276 275104
rect 138676 275064 155276 275092
rect 138676 275052 138682 275064
rect 155270 275052 155276 275064
rect 155328 275052 155334 275104
rect 339638 274984 339644 275036
rect 339696 275024 339702 275036
rect 351230 275024 351236 275036
rect 339696 274996 351236 275024
rect 339696 274984 339702 274996
rect 351230 274984 351236 274996
rect 351288 274984 351294 275036
rect 149750 274916 149756 274968
rect 149808 274956 149814 274968
rect 160514 274956 160520 274968
rect 149808 274928 160520 274956
rect 149808 274916 149814 274928
rect 160514 274916 160520 274928
rect 160572 274916 160578 274968
rect 337614 274916 337620 274968
rect 337672 274956 337678 274968
rect 339086 274956 339092 274968
rect 337672 274928 339092 274956
rect 337672 274916 337678 274928
rect 339086 274916 339092 274928
rect 339144 274916 339150 274968
rect 341018 274916 341024 274968
rect 341076 274956 341082 274968
rect 352150 274956 352156 274968
rect 341076 274928 352156 274956
rect 341076 274916 341082 274928
rect 352150 274916 352156 274928
rect 352208 274916 352214 274968
rect 151958 274848 151964 274900
rect 152016 274888 152022 274900
rect 154813 274891 154871 274897
rect 152016 274860 154672 274888
rect 152016 274848 152022 274860
rect 153430 274780 153436 274832
rect 153488 274820 153494 274832
rect 154534 274820 154540 274832
rect 153488 274792 154540 274820
rect 153488 274780 153494 274792
rect 154534 274780 154540 274792
rect 154592 274780 154598 274832
rect 154644 274820 154672 274860
rect 154813 274857 154825 274891
rect 154859 274888 154871 274891
rect 162722 274888 162728 274900
rect 154859 274860 162728 274888
rect 154859 274857 154871 274860
rect 154813 274851 154871 274857
rect 162722 274848 162728 274860
rect 162780 274848 162786 274900
rect 247914 274848 247920 274900
rect 247972 274888 247978 274900
rect 249570 274888 249576 274900
rect 247972 274860 249576 274888
rect 247972 274848 247978 274860
rect 249570 274848 249576 274860
rect 249628 274848 249634 274900
rect 338258 274848 338264 274900
rect 338316 274888 338322 274900
rect 349574 274888 349580 274900
rect 338316 274860 349580 274888
rect 338316 274848 338322 274860
rect 349574 274848 349580 274860
rect 349632 274848 349638 274900
rect 163274 274820 163280 274832
rect 154644 274792 163280 274820
rect 163274 274780 163280 274792
rect 163332 274780 163338 274832
rect 244050 274780 244056 274832
rect 244108 274820 244114 274832
rect 254446 274820 254452 274832
rect 244108 274792 254452 274820
rect 244108 274780 244114 274792
rect 254446 274780 254452 274792
rect 254504 274780 254510 274832
rect 334118 274780 334124 274832
rect 334176 274820 334182 274832
rect 346170 274820 346176 274832
rect 334176 274792 346176 274820
rect 334176 274780 334182 274792
rect 346170 274780 346176 274792
rect 346228 274780 346234 274832
rect 63086 274712 63092 274764
rect 63144 274752 63150 274764
rect 65018 274752 65024 274764
rect 63144 274724 65024 274752
rect 63144 274712 63150 274724
rect 65018 274712 65024 274724
rect 65076 274712 65082 274764
rect 151038 274712 151044 274764
rect 151096 274752 151102 274764
rect 151774 274752 151780 274764
rect 151096 274724 151780 274752
rect 151096 274712 151102 274724
rect 151774 274712 151780 274724
rect 151832 274712 151838 274764
rect 152234 274712 152240 274764
rect 152292 274752 152298 274764
rect 153338 274752 153344 274764
rect 152292 274724 153344 274752
rect 152292 274712 152298 274724
rect 153338 274712 153344 274724
rect 153396 274712 153402 274764
rect 154074 274712 154080 274764
rect 154132 274752 154138 274764
rect 154626 274752 154632 274764
rect 154132 274724 154632 274752
rect 154132 274712 154138 274724
rect 154626 274712 154632 274724
rect 154684 274712 154690 274764
rect 154721 274755 154779 274761
rect 154721 274721 154733 274755
rect 154767 274752 154779 274755
rect 162078 274752 162084 274764
rect 154767 274724 162084 274752
rect 154767 274721 154779 274724
rect 154721 274715 154779 274721
rect 162078 274712 162084 274724
rect 162136 274712 162142 274764
rect 243038 274712 243044 274764
rect 243096 274752 243102 274764
rect 255734 274752 255740 274764
rect 243096 274724 255740 274752
rect 243096 274712 243102 274724
rect 255734 274712 255740 274724
rect 255792 274712 255798 274764
rect 336878 274712 336884 274764
rect 336936 274752 336942 274764
rect 348746 274752 348752 274764
rect 336936 274724 348752 274752
rect 336936 274712 336942 274724
rect 348746 274712 348752 274724
rect 348804 274712 348810 274764
rect 34566 274644 34572 274696
rect 34624 274684 34630 274696
rect 47078 274684 47084 274696
rect 34624 274656 47084 274684
rect 34624 274644 34630 274656
rect 47078 274644 47084 274656
rect 47136 274644 47142 274696
rect 59682 274644 59688 274696
rect 59740 274684 59746 274696
rect 60878 274684 60884 274696
rect 59740 274656 60884 274684
rect 59740 274644 59746 274656
rect 60878 274644 60884 274656
rect 60936 274644 60942 274696
rect 147818 274644 147824 274696
rect 147876 274684 147882 274696
rect 161434 274684 161440 274696
rect 147876 274656 161440 274684
rect 147876 274644 147882 274656
rect 161434 274644 161440 274656
rect 161492 274644 161498 274696
rect 240278 274644 240284 274696
rect 240336 274684 240342 274696
rect 254538 274684 254544 274696
rect 240336 274656 254544 274684
rect 240336 274644 240342 274656
rect 254538 274644 254544 274656
rect 254596 274644 254602 274696
rect 335406 274644 335412 274696
rect 335464 274684 335470 274696
rect 346998 274684 347004 274696
rect 335464 274656 347004 274684
rect 335464 274644 335470 274656
rect 346998 274644 347004 274656
rect 347056 274644 347062 274696
rect 29230 274576 29236 274628
rect 29288 274616 29294 274628
rect 46618 274616 46624 274628
rect 29288 274588 46624 274616
rect 29288 274576 29294 274588
rect 46618 274576 46624 274588
rect 46676 274576 46682 274628
rect 62350 274576 62356 274628
rect 62408 274616 62414 274628
rect 63546 274616 63552 274628
rect 62408 274588 63552 274616
rect 62408 274576 62414 274588
rect 63546 274576 63552 274588
rect 63604 274576 63610 274628
rect 65018 274576 65024 274628
rect 65076 274616 65082 274628
rect 68606 274616 68612 274628
rect 65076 274588 68612 274616
rect 65076 274576 65082 274588
rect 68606 274576 68612 274588
rect 68664 274576 68670 274628
rect 145058 274576 145064 274628
rect 145116 274616 145122 274628
rect 160238 274616 160244 274628
rect 145116 274588 160244 274616
rect 145116 274576 145122 274588
rect 160238 274576 160244 274588
rect 160296 274576 160302 274628
rect 241658 274576 241664 274628
rect 241716 274616 241722 274628
rect 255090 274616 255096 274628
rect 241716 274588 255096 274616
rect 241716 274576 241722 274588
rect 255090 274576 255096 274588
rect 255148 274576 255154 274628
rect 256194 274576 256200 274628
rect 256252 274616 256258 274628
rect 256930 274616 256936 274628
rect 256252 274588 256936 274616
rect 256252 274576 256258 274588
rect 256930 274576 256936 274588
rect 256988 274576 256994 274628
rect 335498 274576 335504 274628
rect 335556 274616 335562 274628
rect 348102 274616 348108 274628
rect 335556 274588 348108 274616
rect 335556 274576 335562 274588
rect 348102 274576 348108 274588
rect 348160 274576 348166 274628
rect 26562 274508 26568 274560
rect 26620 274548 26626 274560
rect 46526 274548 46532 274560
rect 26620 274520 46532 274548
rect 26620 274508 26626 274520
rect 46526 274508 46532 274520
rect 46584 274508 46590 274560
rect 146438 274508 146444 274560
rect 146496 274548 146502 274560
rect 160882 274548 160888 274560
rect 146496 274520 160888 274548
rect 146496 274508 146502 274520
rect 160882 274508 160888 274520
rect 160940 274508 160946 274560
rect 238898 274508 238904 274560
rect 238956 274548 238962 274560
rect 254262 274548 254268 274560
rect 238956 274520 254268 274548
rect 238956 274508 238962 274520
rect 254262 274508 254268 274520
rect 254320 274508 254326 274560
rect 332738 274508 332744 274560
rect 332796 274548 332802 274560
rect 345342 274548 345348 274560
rect 332796 274520 345348 274548
rect 332796 274508 332802 274520
rect 345342 274508 345348 274520
rect 345400 274508 345406 274560
rect 23894 274440 23900 274492
rect 23952 274480 23958 274492
rect 46434 274480 46440 274492
rect 23952 274452 46440 274480
rect 23952 274440 23958 274452
rect 46434 274440 46440 274452
rect 46492 274440 46498 274492
rect 57014 274440 57020 274492
rect 57072 274480 57078 274492
rect 67134 274480 67140 274492
rect 57072 274452 67140 274480
rect 57072 274440 57078 274452
rect 67134 274440 67140 274452
rect 67192 274440 67198 274492
rect 143678 274440 143684 274492
rect 143736 274480 143742 274492
rect 159318 274480 159324 274492
rect 143736 274452 159324 274480
rect 143736 274440 143742 274452
rect 159318 274440 159324 274452
rect 159376 274440 159382 274492
rect 159594 274440 159600 274492
rect 159652 274480 159658 274492
rect 164562 274480 164568 274492
rect 159652 274452 164568 274480
rect 159652 274440 159658 274452
rect 164562 274440 164568 274452
rect 164620 274440 164626 274492
rect 237518 274440 237524 274492
rect 237576 274480 237582 274492
rect 237576 274452 247684 274480
rect 237576 274440 237582 274452
rect 149198 274372 149204 274424
rect 149256 274412 149262 274424
rect 154721 274415 154779 274421
rect 154721 274412 154733 274415
rect 149256 274384 154733 274412
rect 149256 274372 149262 274384
rect 154721 274381 154733 274384
rect 154767 274381 154779 274415
rect 154721 274375 154779 274381
rect 149106 274304 149112 274356
rect 149164 274344 149170 274356
rect 156834 274344 156840 274356
rect 149164 274316 156840 274344
rect 149164 274304 149170 274316
rect 156834 274304 156840 274316
rect 156892 274304 156898 274356
rect 245338 274304 245344 274356
rect 245396 274344 245402 274356
rect 245798 274344 245804 274356
rect 245396 274316 245804 274344
rect 245396 274304 245402 274316
rect 245798 274304 245804 274316
rect 245856 274304 245862 274356
rect 247656 274344 247684 274452
rect 247730 274440 247736 274492
rect 247788 274480 247794 274492
rect 248558 274480 248564 274492
rect 247788 274452 248564 274480
rect 247788 274440 247794 274452
rect 248558 274440 248564 274452
rect 248616 274440 248622 274492
rect 345158 274440 345164 274492
rect 345216 274480 345222 274492
rect 365306 274480 365312 274492
rect 345216 274452 365312 274480
rect 345216 274440 345222 274452
rect 365306 274440 365312 274452
rect 365364 274440 365370 274492
rect 369906 274440 369912 274492
rect 369964 274480 369970 274492
rect 410202 274480 410208 274492
rect 369964 274452 410208 274480
rect 369964 274440 369970 274452
rect 410202 274440 410208 274452
rect 410260 274440 410266 274492
rect 253434 274344 253440 274356
rect 247656 274316 253440 274344
rect 253434 274304 253440 274316
rect 253492 274304 253498 274356
rect 150486 274236 150492 274288
rect 150544 274276 150550 274288
rect 154813 274279 154871 274285
rect 154813 274276 154825 274279
rect 150544 274248 154825 274276
rect 150544 274236 150550 274248
rect 154813 274245 154825 274248
rect 154859 274245 154871 274279
rect 154813 274239 154871 274245
rect 341754 274236 341760 274288
rect 341812 274276 341818 274288
rect 344606 274276 344612 274288
rect 341812 274248 344612 274276
rect 341812 274236 341818 274248
rect 344606 274236 344612 274248
rect 344664 274236 344670 274288
rect 254814 274168 254820 274220
rect 254872 274208 254878 274220
rect 258310 274208 258316 274220
rect 254872 274180 258316 274208
rect 254872 274168 254878 274180
rect 258310 274168 258316 274180
rect 258368 274168 258374 274220
rect 249018 274032 249024 274084
rect 249076 274072 249082 274084
rect 249938 274072 249944 274084
rect 249076 274044 249944 274072
rect 249076 274032 249082 274044
rect 249938 274032 249944 274044
rect 249996 274032 250002 274084
rect 60234 273964 60240 274016
rect 60292 274004 60298 274016
rect 63270 274004 63276 274016
rect 60292 273976 63276 274004
rect 60292 273964 60298 273976
rect 63270 273964 63276 273976
rect 63328 273964 63334 274016
rect 250674 273964 250680 274016
rect 250732 274004 250738 274016
rect 256378 274004 256384 274016
rect 250732 273976 256384 274004
rect 250732 273964 250738 273976
rect 256378 273964 256384 273976
rect 256436 273964 256442 274016
rect 344330 273964 344336 274016
rect 344388 274004 344394 274016
rect 347366 274004 347372 274016
rect 344388 273976 347372 274004
rect 344388 273964 344394 273976
rect 347366 273964 347372 273976
rect 347424 273964 347430 274016
rect 62994 273896 63000 273948
rect 63052 273936 63058 273948
rect 65938 273936 65944 273948
rect 63052 273908 65944 273936
rect 63052 273896 63058 273908
rect 65938 273896 65944 273908
rect 65996 273896 66002 273948
rect 246534 273896 246540 273948
rect 246592 273936 246598 273948
rect 247178 273936 247184 273948
rect 246592 273908 247184 273936
rect 246592 273896 246598 273908
rect 247178 273896 247184 273908
rect 247236 273896 247242 273948
rect 253434 273896 253440 273948
rect 253492 273936 253498 273948
rect 257574 273936 257580 273948
rect 253492 273908 257580 273936
rect 253492 273896 253498 273908
rect 257574 273896 257580 273908
rect 257632 273896 257638 273948
rect 343502 273896 343508 273948
rect 343560 273936 343566 273948
rect 347274 273936 347280 273948
rect 343560 273908 347280 273936
rect 343560 273896 343566 273908
rect 347274 273896 347280 273908
rect 347332 273896 347338 273948
rect 61614 273828 61620 273880
rect 61672 273868 61678 273880
rect 64098 273868 64104 273880
rect 61672 273840 64104 273868
rect 61672 273828 61678 273840
rect 64098 273828 64104 273840
rect 64156 273828 64162 273880
rect 66398 273828 66404 273880
rect 66456 273868 66462 273880
rect 70354 273868 70360 273880
rect 66456 273840 70360 273868
rect 66456 273828 66462 273840
rect 70354 273828 70360 273840
rect 70412 273828 70418 273880
rect 234114 273828 234120 273880
rect 234172 273868 234178 273880
rect 234758 273868 234764 273880
rect 234172 273840 234764 273868
rect 234172 273828 234178 273840
rect 234758 273828 234764 273840
rect 234816 273828 234822 273880
rect 243498 273828 243504 273880
rect 243556 273868 243562 273880
rect 250766 273868 250772 273880
rect 243556 273840 250772 273868
rect 243556 273828 243562 273840
rect 250766 273828 250772 273840
rect 250824 273828 250830 273880
rect 339270 273828 339276 273880
rect 339328 273868 339334 273880
rect 341846 273868 341852 273880
rect 339328 273840 341852 273868
rect 339328 273828 339334 273840
rect 341846 273828 341852 273840
rect 341904 273828 341910 273880
rect 342398 273828 342404 273880
rect 342456 273868 342462 273880
rect 344514 273868 344520 273880
rect 342456 273840 344520 273868
rect 342456 273828 342462 273840
rect 344514 273828 344520 273840
rect 344572 273828 344578 273880
rect 21226 273760 21232 273812
rect 21284 273800 21290 273812
rect 22238 273800 22244 273812
rect 21284 273772 22244 273800
rect 21284 273760 21290 273772
rect 22238 273760 22244 273772
rect 22296 273760 22302 273812
rect 61430 273760 61436 273812
rect 61488 273800 61494 273812
rect 62258 273800 62264 273812
rect 61488 273772 62264 273800
rect 61488 273760 61494 273772
rect 62258 273760 62264 273772
rect 62316 273760 62322 273812
rect 63638 273760 63644 273812
rect 63696 273800 63702 273812
rect 67686 273800 67692 273812
rect 63696 273772 67692 273800
rect 63696 273760 63702 273772
rect 67686 273760 67692 273772
rect 67744 273760 67750 273812
rect 162354 273760 162360 273812
rect 162412 273800 162418 273812
rect 163918 273800 163924 273812
rect 162412 273772 163924 273800
rect 162412 273760 162418 273772
rect 163918 273760 163924 273772
rect 163976 273760 163982 273812
rect 338166 273760 338172 273812
rect 338224 273800 338230 273812
rect 338994 273800 339000 273812
rect 338224 273772 339000 273800
rect 338224 273760 338230 273772
rect 338994 273760 339000 273772
rect 339052 273760 339058 273812
rect 340098 273760 340104 273812
rect 340156 273800 340162 273812
rect 340926 273800 340932 273812
rect 340156 273772 340932 273800
rect 340156 273760 340162 273772
rect 340926 273760 340932 273772
rect 340984 273760 340990 273812
rect 348654 273760 348660 273812
rect 348712 273800 348718 273812
rect 350402 273800 350408 273812
rect 348712 273772 350408 273800
rect 348712 273760 348718 273772
rect 350402 273760 350408 273772
rect 350460 273760 350466 273812
rect 13038 273692 13044 273744
rect 13096 273732 13102 273744
rect 31898 273732 31904 273744
rect 13096 273704 31904 273732
rect 13096 273692 13102 273704
rect 31898 273692 31904 273704
rect 31956 273692 31962 273744
rect 138066 273692 138072 273744
rect 138124 273732 138130 273744
rect 141654 273732 141660 273744
rect 138124 273704 141660 273732
rect 138124 273692 138130 273704
rect 141654 273692 141660 273704
rect 141712 273692 141718 273744
rect 247270 273692 247276 273744
rect 247328 273732 247334 273744
rect 252146 273732 252152 273744
rect 247328 273704 252152 273732
rect 247328 273692 247334 273704
rect 252146 273692 252152 273704
rect 252204 273692 252210 273744
rect 31898 273012 31904 273064
rect 31956 273052 31962 273064
rect 46710 273052 46716 273064
rect 31956 273024 46716 273052
rect 31956 273012 31962 273024
rect 46710 273012 46716 273024
rect 46768 273012 46774 273064
rect 51405 272511 51463 272517
rect 51405 272477 51417 272511
rect 51451 272508 51463 272511
rect 51494 272508 51500 272520
rect 51451 272480 51500 272508
rect 51451 272477 51463 272480
rect 51405 272471 51463 272477
rect 51494 272468 51500 272480
rect 51552 272468 51558 272520
rect 352794 272400 352800 272452
rect 352852 272440 352858 272452
rect 352978 272440 352984 272452
rect 352852 272412 352984 272440
rect 352852 272400 352858 272412
rect 352978 272400 352984 272412
rect 353036 272400 353042 272452
rect 51402 269720 51408 269732
rect 51363 269692 51408 269720
rect 51402 269680 51408 269692
rect 51460 269680 51466 269732
rect 88386 269612 88392 269664
rect 88444 269652 88450 269664
rect 182410 269652 182416 269664
rect 88444 269624 182416 269652
rect 88444 269612 88450 269624
rect 182410 269612 182416 269624
rect 182468 269652 182474 269664
rect 276434 269652 276440 269664
rect 182468 269624 276440 269652
rect 182468 269612 182474 269624
rect 276434 269612 276440 269624
rect 276492 269612 276498 269664
rect 290694 269612 290700 269664
rect 290752 269652 290758 269664
rect 395390 269652 395396 269664
rect 290752 269624 395396 269652
rect 290752 269612 290758 269624
rect 395390 269612 395396 269624
rect 395448 269612 395454 269664
rect 427590 269612 427596 269664
rect 427648 269652 427654 269664
rect 429430 269652 429436 269664
rect 427648 269624 429436 269652
rect 427648 269612 427654 269624
rect 429430 269612 429436 269624
rect 429488 269612 429494 269664
rect 102646 269544 102652 269596
rect 102704 269584 102710 269596
rect 196670 269584 196676 269596
rect 102704 269556 196676 269584
rect 102704 269544 102710 269556
rect 196670 269544 196676 269556
rect 196728 269584 196734 269596
rect 197498 269584 197504 269596
rect 196728 269556 197504 269584
rect 196728 269544 196734 269556
rect 197498 269544 197504 269556
rect 197556 269544 197562 269596
rect 189494 269476 189500 269528
rect 189552 269516 189558 269528
rect 283518 269516 283524 269528
rect 189552 269488 283524 269516
rect 189552 269476 189558 269488
rect 283518 269476 283524 269488
rect 283576 269476 283582 269528
rect 127762 269340 127768 269392
rect 127820 269380 127826 269392
rect 131166 269380 131172 269392
rect 127820 269352 131172 269380
rect 127820 269340 127826 269352
rect 131166 269340 131172 269352
rect 131224 269340 131230 269392
rect 95562 269000 95568 269052
rect 95620 269040 95626 269052
rect 109730 269040 109736 269052
rect 95620 269012 109736 269040
rect 95620 269000 95626 269012
rect 109730 269000 109736 269012
rect 109788 269000 109794 269052
rect 189310 269000 189316 269052
rect 189368 269040 189374 269052
rect 203754 269040 203760 269052
rect 189368 269012 203760 269040
rect 189368 269000 189374 269012
rect 203754 269000 203760 269012
rect 203812 269000 203818 269052
rect 284530 269000 284536 269052
rect 284588 269040 284594 269052
rect 297778 269040 297784 269052
rect 284588 269012 297784 269040
rect 284588 269000 284594 269012
rect 297778 269000 297784 269012
rect 297836 269000 297842 269052
rect 95470 268932 95476 268984
rect 95528 268972 95534 268984
rect 174866 268972 174872 268984
rect 95528 268944 174872 268972
rect 95528 268932 95534 268944
rect 174866 268932 174872 268944
rect 174924 268972 174930 268984
rect 189494 268972 189500 268984
rect 174924 268944 189500 268972
rect 174924 268932 174930 268944
rect 189494 268932 189500 268944
rect 189552 268932 189558 268984
rect 197498 268932 197504 268984
rect 197556 268972 197562 268984
rect 264474 268972 264480 268984
rect 197556 268944 264480 268972
rect 197556 268932 197562 268944
rect 264474 268932 264480 268944
rect 264532 268972 264538 268984
rect 290694 268972 290700 268984
rect 264532 268944 290700 268972
rect 264532 268932 264538 268944
rect 290694 268932 290700 268944
rect 290752 268932 290758 268984
rect 114790 268524 114796 268576
rect 114848 268564 114854 268576
rect 116906 268564 116912 268576
rect 114848 268536 116912 268564
rect 114848 268524 114854 268536
rect 116906 268524 116912 268536
rect 116964 268524 116970 268576
rect 209918 268252 209924 268304
rect 209976 268292 209982 268304
rect 210930 268292 210936 268304
rect 209976 268264 210936 268292
rect 209976 268252 209982 268264
rect 210930 268252 210936 268264
rect 210988 268252 210994 268304
rect 303758 268252 303764 268304
rect 303816 268292 303822 268304
rect 304954 268292 304960 268304
rect 303816 268264 304960 268292
rect 303816 268252 303822 268264
rect 304954 268252 304960 268264
rect 305012 268252 305018 268304
rect 51310 267844 51316 267896
rect 51368 267884 51374 267896
rect 52046 267884 52052 267896
rect 51368 267856 52052 267884
rect 51368 267844 51374 267856
rect 52046 267844 52052 267856
rect 52104 267844 52110 267896
rect 354910 267844 354916 267896
rect 354968 267884 354974 267896
rect 355830 267884 355836 267896
rect 354968 267856 355836 267884
rect 354968 267844 354974 267856
rect 355830 267844 355836 267856
rect 355888 267844 355894 267896
rect 333382 266824 333388 266876
rect 333440 266864 333446 266876
rect 334118 266864 334124 266876
rect 333440 266836 334124 266864
rect 333440 266824 333446 266836
rect 334118 266824 334124 266836
rect 334176 266824 334182 266876
rect 334394 266824 334400 266876
rect 334452 266864 334458 266876
rect 335406 266864 335412 266876
rect 334452 266836 335412 266864
rect 334452 266824 334458 266836
rect 335406 266824 335412 266836
rect 335464 266824 335470 266876
rect 337522 266824 337528 266876
rect 337580 266864 337586 266876
rect 338258 266864 338264 266876
rect 337580 266836 338264 266864
rect 337580 266824 337586 266836
rect 338258 266824 338264 266836
rect 338316 266824 338322 266876
rect 347274 266824 347280 266876
rect 347332 266864 347338 266876
rect 348930 266864 348936 266876
rect 347332 266836 348936 266864
rect 347332 266824 347338 266836
rect 348930 266824 348936 266836
rect 348988 266824 348994 266876
rect 64834 266756 64840 266808
rect 64892 266796 64898 266808
rect 69342 266796 69348 266808
rect 64892 266768 69348 266796
rect 64892 266756 64898 266768
rect 69342 266756 69348 266768
rect 69400 266756 69406 266808
rect 245706 266756 245712 266808
rect 245764 266796 245770 266808
rect 253621 266799 253679 266805
rect 253621 266796 253633 266799
rect 245764 266768 253633 266796
rect 245764 266756 245770 266768
rect 253621 266765 253633 266768
rect 253667 266765 253679 266799
rect 253621 266759 253679 266765
rect 344514 266756 344520 266808
rect 344572 266796 344578 266808
rect 347918 266796 347924 266808
rect 344572 266768 347924 266796
rect 344572 266756 344578 266768
rect 347918 266756 347924 266768
rect 347976 266756 347982 266808
rect 59498 266688 59504 266740
rect 59556 266728 59562 266740
rect 71090 266728 71096 266740
rect 59556 266700 71096 266728
rect 59556 266688 59562 266700
rect 71090 266688 71096 266700
rect 71148 266688 71154 266740
rect 153246 266688 153252 266740
rect 153304 266728 153310 266740
rect 162354 266728 162360 266740
rect 153304 266700 162360 266728
rect 153304 266688 153310 266700
rect 162354 266688 162360 266700
rect 162412 266688 162418 266740
rect 246258 266688 246264 266740
rect 246316 266728 246322 266740
rect 256194 266728 256200 266740
rect 246316 266700 256200 266728
rect 246316 266688 246322 266700
rect 256194 266688 256200 266700
rect 256252 266688 256258 266740
rect 60878 266620 60884 266672
rect 60936 266660 60942 266672
rect 72102 266660 72108 266672
rect 60936 266632 72108 266660
rect 60936 266620 60942 266632
rect 72102 266620 72108 266632
rect 72160 266620 72166 266672
rect 150578 266620 150584 266672
rect 150636 266660 150642 266672
rect 161710 266660 161716 266672
rect 150636 266632 161716 266660
rect 150636 266620 150642 266632
rect 161710 266620 161716 266632
rect 161768 266620 161774 266672
rect 245798 266620 245804 266672
rect 245856 266660 245862 266672
rect 256930 266660 256936 266672
rect 245856 266632 256936 266660
rect 245856 266620 245862 266632
rect 256930 266620 256936 266632
rect 256988 266620 256994 266672
rect 62258 266552 62264 266604
rect 62316 266592 62322 266604
rect 74218 266592 74224 266604
rect 62316 266564 74224 266592
rect 62316 266552 62322 266564
rect 74218 266552 74224 266564
rect 74276 266552 74282 266604
rect 244418 266552 244424 266604
rect 244476 266592 244482 266604
rect 255550 266592 255556 266604
rect 244476 266564 255556 266592
rect 244476 266552 244482 266564
rect 255550 266552 255556 266564
rect 255608 266552 255614 266604
rect 57658 266484 57664 266536
rect 57716 266524 57722 266536
rect 60234 266524 60240 266536
rect 57716 266496 60240 266524
rect 57716 266484 57722 266496
rect 60234 266484 60240 266496
rect 60292 266484 60298 266536
rect 143034 266484 143040 266536
rect 143092 266524 143098 266536
rect 155730 266524 155736 266536
rect 143092 266496 155736 266524
rect 143092 266484 143098 266496
rect 155730 266484 155736 266496
rect 155788 266484 155794 266536
rect 247638 266484 247644 266536
rect 247696 266524 247702 266536
rect 253434 266524 253440 266536
rect 247696 266496 253440 266524
rect 247696 266484 247702 266496
rect 253434 266484 253440 266496
rect 253492 266484 253498 266536
rect 259690 266524 259696 266536
rect 253544 266496 259696 266524
rect 56738 266416 56744 266468
rect 56796 266456 56802 266468
rect 67962 266456 67968 266468
rect 56796 266428 67968 266456
rect 56796 266416 56802 266428
rect 67962 266416 67968 266428
rect 68020 266416 68026 266468
rect 153338 266416 153344 266468
rect 153396 266456 153402 266468
rect 165942 266456 165948 266468
rect 153396 266428 165948 266456
rect 153396 266416 153402 266428
rect 165942 266416 165948 266428
rect 166000 266416 166006 266468
rect 247178 266416 247184 266468
rect 247236 266456 247242 266468
rect 253544 266456 253572 266496
rect 259690 266484 259696 266496
rect 259748 266484 259754 266536
rect 344606 266484 344612 266536
rect 344664 266524 344670 266536
rect 346814 266524 346820 266536
rect 344664 266496 346820 266524
rect 344664 266484 344670 266496
rect 346814 266484 346820 266496
rect 346872 266484 346878 266536
rect 247236 266428 253572 266456
rect 253621 266459 253679 266465
rect 247236 266416 247242 266428
rect 253621 266425 253633 266459
rect 253667 266456 253679 266459
rect 258310 266456 258316 266468
rect 253667 266428 258316 266456
rect 253667 266425 253679 266428
rect 253621 266419 253679 266425
rect 258310 266416 258316 266428
rect 258368 266416 258374 266468
rect 341846 266416 341852 266468
rect 341904 266456 341910 266468
rect 343778 266456 343784 266468
rect 341904 266428 343784 266456
rect 341904 266416 341910 266428
rect 343778 266416 343784 266428
rect 343836 266416 343842 266468
rect 55358 266348 55364 266400
rect 55416 266388 55422 266400
rect 66950 266388 66956 266400
rect 55416 266360 66956 266388
rect 55416 266348 55422 266360
rect 66950 266348 66956 266360
rect 67008 266348 67014 266400
rect 151866 266348 151872 266400
rect 151924 266388 151930 266400
rect 164562 266388 164568 266400
rect 151924 266360 164568 266388
rect 151924 266348 151930 266360
rect 164562 266348 164568 266360
rect 164620 266348 164626 266400
rect 236874 266348 236880 266400
rect 236932 266388 236938 266400
rect 250030 266388 250036 266400
rect 236932 266360 250036 266388
rect 236932 266348 236938 266360
rect 250030 266348 250036 266360
rect 250088 266348 250094 266400
rect 252977 266391 253035 266397
rect 252977 266388 252989 266391
rect 250140 266360 252989 266388
rect 58118 266280 58124 266332
rect 58176 266320 58182 266332
rect 70078 266320 70084 266332
rect 58176 266292 70084 266320
rect 58176 266280 58182 266292
rect 70078 266280 70084 266292
rect 70136 266280 70142 266332
rect 153154 266280 153160 266332
rect 153212 266320 153218 266332
rect 167322 266320 167328 266332
rect 153212 266292 167328 266320
rect 153212 266280 153218 266292
rect 167322 266280 167328 266292
rect 167380 266280 167386 266332
rect 247086 266280 247092 266332
rect 247144 266320 247150 266332
rect 250140 266320 250168 266360
rect 252977 266357 252989 266360
rect 253023 266357 253035 266391
rect 252977 266351 253035 266357
rect 247144 266292 250168 266320
rect 247144 266280 247150 266292
rect 250766 266280 250772 266332
rect 250824 266320 250830 266332
rect 252790 266320 252796 266332
rect 250824 266292 252796 266320
rect 250824 266280 250830 266292
rect 252790 266280 252796 266292
rect 252848 266280 252854 266332
rect 262450 266320 262456 266332
rect 252900 266292 262456 266320
rect 60786 266212 60792 266264
rect 60844 266252 60850 266264
rect 73114 266252 73120 266264
rect 60844 266224 73120 266252
rect 60844 266212 60850 266224
rect 73114 266212 73120 266224
rect 73172 266212 73178 266264
rect 154534 266212 154540 266264
rect 154592 266252 154598 266264
rect 168702 266252 168708 266264
rect 154592 266224 168708 266252
rect 154592 266212 154598 266224
rect 168702 266212 168708 266224
rect 168760 266212 168766 266264
rect 248558 266212 248564 266264
rect 248616 266252 248622 266264
rect 252900 266252 252928 266292
rect 262450 266280 262456 266292
rect 262508 266280 262514 266332
rect 347366 266280 347372 266332
rect 347424 266320 347430 266332
rect 349942 266320 349948 266332
rect 347424 266292 349948 266320
rect 347424 266280 347430 266292
rect 349942 266280 349948 266292
rect 350000 266280 350006 266332
rect 248616 266224 252928 266252
rect 252977 266255 253035 266261
rect 248616 266212 248622 266224
rect 252977 266221 252989 266255
rect 253023 266252 253035 266255
rect 261070 266252 261076 266264
rect 253023 266224 261076 266252
rect 253023 266221 253035 266224
rect 252977 266215 253035 266221
rect 261070 266212 261076 266224
rect 261128 266212 261134 266264
rect 340834 266212 340840 266264
rect 340892 266252 340898 266264
rect 345802 266252 345808 266264
rect 340892 266224 345808 266252
rect 340892 266212 340898 266224
rect 345802 266212 345808 266224
rect 345860 266212 345866 266264
rect 63546 266144 63552 266196
rect 63604 266184 63610 266196
rect 75230 266184 75236 266196
rect 63604 266156 75236 266184
rect 63604 266144 63610 266156
rect 75230 266144 75236 266156
rect 75288 266144 75294 266196
rect 154626 266144 154632 266196
rect 154684 266184 154690 266196
rect 170082 266184 170088 266196
rect 154684 266156 170088 266184
rect 154684 266144 154690 266156
rect 170082 266144 170088 266156
rect 170140 266144 170146 266196
rect 244878 266144 244884 266196
rect 244936 266184 244942 266196
rect 250674 266184 250680 266196
rect 244936 266156 250680 266184
rect 244936 266144 244942 266156
rect 250674 266144 250680 266156
rect 250732 266144 250738 266196
rect 263830 266184 263836 266196
rect 250784 266156 263836 266184
rect 151774 266076 151780 266128
rect 151832 266116 151838 266128
rect 163090 266116 163096 266128
rect 151832 266088 163096 266116
rect 151832 266076 151838 266088
rect 163090 266076 163096 266088
rect 163148 266076 163154 266128
rect 248466 266076 248472 266128
rect 248524 266116 248530 266128
rect 250784 266116 250812 266156
rect 263830 266144 263836 266156
rect 263888 266144 263894 266196
rect 338534 266144 338540 266196
rect 338592 266184 338598 266196
rect 348654 266184 348660 266196
rect 338592 266156 348660 266184
rect 338592 266144 338598 266156
rect 348654 266144 348660 266156
rect 348712 266144 348718 266196
rect 248524 266088 250812 266116
rect 248524 266076 248530 266088
rect 61798 265872 61804 265924
rect 61856 265912 61862 265924
rect 66582 265912 66588 265924
rect 61856 265884 66588 265912
rect 61856 265872 61862 265884
rect 66582 265872 66588 265884
rect 66640 265872 66646 265924
rect 59682 265736 59688 265788
rect 59740 265776 59746 265788
rect 63086 265776 63092 265788
rect 59740 265748 63092 265776
rect 59740 265736 59746 265748
rect 63086 265736 63092 265748
rect 63144 265736 63150 265788
rect 251870 265736 251876 265788
rect 251928 265776 251934 265788
rect 258954 265776 258960 265788
rect 251928 265748 258960 265776
rect 251928 265736 251934 265748
rect 258954 265736 258960 265748
rect 259012 265736 259018 265788
rect 58670 265668 58676 265720
rect 58728 265708 58734 265720
rect 61614 265708 61620 265720
rect 58728 265680 61620 265708
rect 58728 265668 58734 265680
rect 61614 265668 61620 265680
rect 61672 265668 61678 265720
rect 157846 265668 157852 265720
rect 157904 265708 157910 265720
rect 165114 265708 165120 265720
rect 157904 265680 165120 265708
rect 157904 265668 157910 265680
rect 165114 265668 165120 265680
rect 165172 265668 165178 265720
rect 338994 265668 339000 265720
rect 339052 265708 339058 265720
rect 342674 265708 342680 265720
rect 339052 265680 342680 265708
rect 339052 265668 339058 265680
rect 342674 265668 342680 265680
rect 342732 265668 342738 265720
rect 60694 265600 60700 265652
rect 60752 265640 60758 265652
rect 62994 265640 63000 265652
rect 60752 265612 63000 265640
rect 60752 265600 60758 265612
rect 62994 265600 63000 265612
rect 63052 265600 63058 265652
rect 154718 265600 154724 265652
rect 154776 265640 154782 265652
rect 159594 265640 159600 265652
rect 154776 265612 159600 265640
rect 154776 265600 154782 265612
rect 159594 265600 159600 265612
rect 159652 265600 159658 265652
rect 249018 265600 249024 265652
rect 249076 265640 249082 265652
rect 254814 265640 254820 265652
rect 249076 265612 254820 265640
rect 249076 265600 249082 265612
rect 254814 265600 254820 265612
rect 254872 265600 254878 265652
rect 340926 265600 340932 265652
rect 340984 265640 340990 265652
rect 344790 265640 344796 265652
rect 340984 265612 344796 265640
rect 340984 265600 340990 265612
rect 344790 265600 344796 265612
rect 344848 265600 344854 265652
rect 62810 265532 62816 265584
rect 62868 265572 62874 265584
rect 63638 265572 63644 265584
rect 62868 265544 63644 265572
rect 62868 265532 62874 265544
rect 63638 265532 63644 265544
rect 63696 265532 63702 265584
rect 63822 265532 63828 265584
rect 63880 265572 63886 265584
rect 65018 265572 65024 265584
rect 63880 265544 65024 265572
rect 63880 265532 63886 265544
rect 65018 265532 65024 265544
rect 65076 265532 65082 265584
rect 67134 265532 67140 265584
rect 67192 265572 67198 265584
rect 68974 265572 68980 265584
rect 67192 265544 68980 265572
rect 67192 265532 67198 265544
rect 68974 265532 68980 265544
rect 69032 265532 69038 265584
rect 156834 265532 156840 265584
rect 156892 265572 156898 265584
rect 158950 265572 158956 265584
rect 156892 265544 158956 265572
rect 156892 265532 156898 265544
rect 158950 265532 158956 265544
rect 159008 265532 159014 265584
rect 339086 265532 339092 265584
rect 339144 265572 339150 265584
rect 341662 265572 341668 265584
rect 339144 265544 341668 265572
rect 339144 265532 339150 265544
rect 341662 265532 341668 265544
rect 341720 265532 341726 265584
rect 77254 264036 77260 264088
rect 77312 264076 77318 264088
rect 123254 264076 123260 264088
rect 77312 264048 123260 264076
rect 77312 264036 77318 264048
rect 123254 264036 123260 264048
rect 123312 264076 123318 264088
rect 124358 264076 124364 264088
rect 123312 264048 124364 264076
rect 123312 264036 123318 264048
rect 124358 264036 124364 264048
rect 124416 264036 124422 264088
rect 310750 264036 310756 264088
rect 310808 264076 310814 264088
rect 312038 264076 312044 264088
rect 310808 264048 312044 264076
rect 310808 264036 310814 264048
rect 312038 264036 312044 264048
rect 312096 264076 312102 264088
rect 327310 264076 327316 264088
rect 312096 264048 327316 264076
rect 312096 264036 312102 264048
rect 327310 264036 327316 264048
rect 327368 264036 327374 264088
rect 203113 263807 203171 263813
rect 203113 263773 203125 263807
rect 203159 263804 203171 263807
rect 212681 263807 212739 263813
rect 212681 263804 212693 263807
rect 203159 263776 212693 263804
rect 203159 263773 203171 263776
rect 203113 263767 203171 263773
rect 212681 263773 212693 263776
rect 212727 263773 212739 263807
rect 212681 263767 212739 263773
rect 154813 263739 154871 263745
rect 154813 263705 154825 263739
rect 154859 263736 154871 263739
rect 164381 263739 164439 263745
rect 164381 263736 164393 263739
rect 154859 263708 164393 263736
rect 154859 263705 154871 263708
rect 154813 263699 154871 263705
rect 164381 263705 164393 263708
rect 164427 263705 164439 263739
rect 164381 263699 164439 263705
rect 174133 263671 174191 263677
rect 174133 263637 174145 263671
rect 174179 263668 174191 263671
rect 183701 263671 183759 263677
rect 183701 263668 183713 263671
rect 174179 263640 183713 263668
rect 174179 263637 174191 263640
rect 174133 263631 174191 263637
rect 183701 263637 183713 263640
rect 183747 263637 183759 263671
rect 203113 263671 203171 263677
rect 203113 263668 203125 263671
rect 183701 263631 183759 263637
rect 196136 263640 203125 263668
rect 154442 263560 154448 263612
rect 154500 263600 154506 263612
rect 154813 263603 154871 263609
rect 154813 263600 154825 263603
rect 154500 263572 154825 263600
rect 154500 263560 154506 263572
rect 154813 263569 154825 263572
rect 154859 263569 154871 263603
rect 196136 263600 196164 263640
rect 203113 263637 203125 263640
rect 203159 263637 203171 263671
rect 241661 263671 241719 263677
rect 241661 263668 241673 263671
rect 203113 263631 203171 263637
rect 225024 263640 225236 263668
rect 154813 263563 154871 263569
rect 187764 263572 196164 263600
rect 212681 263603 212739 263609
rect 164381 263535 164439 263541
rect 164381 263501 164393 263535
rect 164427 263532 164439 263535
rect 167233 263535 167291 263541
rect 164427 263504 164562 263532
rect 164427 263501 164439 263504
rect 164381 263495 164439 263501
rect 73850 263464 73856 263476
rect 73811 263436 73856 263464
rect 73850 263424 73856 263436
rect 73908 263424 73914 263476
rect 74034 263424 74040 263476
rect 74092 263424 74098 263476
rect 124358 263424 124364 263476
rect 124416 263464 124422 263476
rect 140274 263464 140280 263476
rect 124416 263436 140280 263464
rect 124416 263424 124422 263436
rect 140274 263424 140280 263436
rect 140332 263424 140338 263476
rect 164534 263464 164562 263504
rect 167233 263501 167245 263535
rect 167279 263532 167291 263535
rect 174133 263535 174191 263541
rect 167279 263504 174084 263532
rect 167279 263501 167291 263504
rect 167233 263495 167291 263501
rect 167141 263467 167199 263473
rect 167141 263464 167153 263467
rect 164534 263436 167153 263464
rect 167141 263433 167153 263436
rect 167187 263433 167199 263467
rect 174056 263464 174084 263504
rect 174133 263501 174145 263535
rect 174179 263501 174191 263535
rect 174133 263495 174191 263501
rect 183701 263535 183759 263541
rect 183701 263501 183713 263535
rect 183747 263532 183759 263535
rect 186461 263535 186519 263541
rect 186461 263532 186473 263535
rect 183747 263504 186473 263532
rect 183747 263501 183759 263504
rect 183701 263495 183759 263501
rect 186461 263501 186473 263504
rect 186507 263501 186519 263535
rect 186461 263495 186519 263501
rect 186553 263535 186611 263541
rect 186553 263501 186565 263535
rect 186599 263532 186611 263535
rect 187764 263532 187792 263572
rect 212681 263569 212693 263603
rect 212727 263600 212739 263603
rect 215533 263603 215591 263609
rect 212727 263572 215484 263600
rect 212727 263569 212739 263572
rect 212681 263563 212739 263569
rect 186599 263504 187792 263532
rect 186599 263501 186611 263504
rect 186553 263495 186611 263501
rect 174148 263464 174176 263495
rect 174056 263436 174176 263464
rect 215456 263464 215484 263572
rect 215533 263569 215545 263603
rect 215579 263600 215591 263603
rect 225024 263600 225052 263640
rect 215579 263572 225052 263600
rect 215579 263569 215591 263572
rect 215533 263563 215591 263569
rect 225208 263532 225236 263640
rect 234684 263640 241673 263668
rect 234684 263532 234712 263640
rect 241661 263637 241673 263640
rect 241707 263637 241719 263671
rect 241661 263631 241719 263637
rect 312133 263671 312191 263677
rect 312133 263637 312145 263671
rect 312179 263668 312191 263671
rect 321701 263671 321759 263677
rect 321701 263668 321713 263671
rect 312179 263640 321713 263668
rect 312179 263637 312191 263640
rect 312133 263631 312191 263637
rect 321701 263637 321713 263640
rect 321747 263637 321759 263671
rect 321701 263631 321759 263637
rect 321793 263671 321851 263677
rect 321793 263637 321805 263671
rect 321839 263668 321851 263671
rect 331361 263671 331419 263677
rect 331361 263668 331373 263671
rect 321839 263640 331373 263668
rect 321839 263637 321851 263640
rect 321793 263631 321851 263637
rect 331361 263637 331373 263640
rect 331407 263637 331419 263671
rect 331361 263631 331419 263637
rect 336896 263640 337016 263668
rect 241753 263603 241811 263609
rect 241753 263569 241765 263603
rect 241799 263600 241811 263603
rect 250585 263603 250643 263609
rect 250585 263600 250597 263603
rect 241799 263572 250597 263600
rect 241799 263569 241811 263572
rect 241753 263563 241811 263569
rect 250585 263569 250597 263572
rect 250631 263569 250643 263603
rect 250585 263563 250643 263569
rect 267234 263560 267240 263612
rect 267292 263600 267298 263612
rect 310750 263600 310756 263612
rect 267292 263572 310756 263600
rect 267292 263560 267298 263572
rect 310750 263560 310756 263572
rect 310808 263560 310814 263612
rect 336896 263609 336924 263640
rect 336988 263609 337016 263640
rect 336881 263603 336939 263609
rect 336881 263569 336893 263603
rect 336927 263569 336939 263603
rect 336881 263563 336939 263569
rect 336973 263603 337031 263609
rect 336973 263569 336985 263603
rect 337019 263569 337031 263603
rect 336973 263563 337031 263569
rect 358406 263560 358412 263612
rect 358464 263560 358470 263612
rect 225208 263504 234712 263532
rect 241661 263535 241719 263541
rect 241661 263501 241673 263535
rect 241707 263532 241719 263535
rect 241707 263504 241796 263532
rect 241707 263501 241719 263504
rect 241661 263495 241719 263501
rect 241768 263473 241796 263504
rect 249938 263492 249944 263544
rect 249996 263532 250002 263544
rect 341113 263535 341171 263541
rect 341113 263532 341125 263535
rect 249996 263504 341125 263532
rect 249996 263492 250002 263504
rect 341113 263501 341125 263504
rect 341159 263501 341171 263535
rect 341113 263495 341171 263501
rect 341297 263535 341355 263541
rect 341297 263501 341309 263535
rect 341343 263532 341355 263535
rect 358424 263532 358452 263560
rect 341343 263504 358452 263532
rect 341343 263501 341355 263504
rect 341297 263495 341355 263501
rect 215533 263467 215591 263473
rect 215533 263464 215545 263467
rect 215456 263436 215545 263464
rect 167141 263427 167199 263433
rect 215533 263433 215545 263436
rect 215579 263433 215591 263467
rect 215533 263427 215591 263433
rect 241753 263467 241811 263473
rect 241753 263433 241765 263467
rect 241799 263433 241811 263467
rect 241753 263427 241811 263433
rect 272757 263467 272815 263473
rect 272757 263433 272769 263467
rect 272803 263464 272815 263467
rect 277633 263467 277691 263473
rect 277633 263464 277645 263467
rect 272803 263436 277645 263464
rect 272803 263433 272815 263436
rect 272757 263427 272815 263433
rect 277633 263433 277645 263436
rect 277679 263433 277691 263467
rect 277633 263427 277691 263433
rect 287201 263467 287259 263473
rect 287201 263433 287213 263467
rect 287247 263464 287259 263467
rect 296953 263467 297011 263473
rect 296953 263464 296965 263467
rect 287247 263436 296965 263464
rect 287247 263433 287259 263436
rect 287201 263427 287259 263433
rect 296953 263433 296965 263436
rect 296999 263433 297011 263467
rect 296953 263427 297011 263433
rect 302657 263467 302715 263473
rect 302657 263433 302669 263467
rect 302703 263464 302715 263467
rect 312133 263467 312191 263473
rect 312133 263464 312145 263467
rect 302703 263436 312145 263464
rect 302703 263433 302715 263436
rect 302657 263427 302715 263433
rect 312133 263433 312145 263436
rect 312179 263433 312191 263467
rect 312133 263427 312191 263433
rect 331361 263467 331419 263473
rect 331361 263433 331373 263467
rect 331407 263464 331419 263467
rect 336881 263467 336939 263473
rect 336881 263464 336893 263467
rect 331407 263436 336893 263464
rect 331407 263433 331419 263436
rect 331361 263427 331419 263433
rect 336881 263433 336893 263436
rect 336927 263433 336939 263467
rect 336881 263427 336939 263433
rect 336973 263467 337031 263473
rect 336973 263433 336985 263467
rect 337019 263464 337031 263467
rect 358406 263464 358412 263476
rect 337019 263436 358412 263464
rect 337019 263433 337031 263436
rect 336973 263427 337031 263433
rect 358406 263424 358412 263436
rect 358464 263424 358470 263476
rect 74052 263396 74080 263424
rect 369538 263396 369544 263408
rect 74052 263368 369544 263396
rect 369538 263356 369544 263368
rect 369596 263356 369602 263408
rect 250585 263331 250643 263337
rect 250585 263297 250597 263331
rect 250631 263328 250643 263331
rect 272757 263331 272815 263337
rect 272757 263328 272769 263331
rect 250631 263300 272769 263328
rect 250631 263297 250643 263300
rect 250585 263291 250643 263297
rect 272757 263297 272769 263300
rect 272803 263297 272815 263331
rect 272757 263291 272815 263297
rect 277633 263263 277691 263269
rect 277633 263229 277645 263263
rect 277679 263260 277691 263263
rect 287201 263263 287259 263269
rect 287201 263260 287213 263263
rect 277679 263232 287213 263260
rect 277679 263229 277691 263232
rect 277633 263223 277691 263229
rect 287201 263229 287213 263232
rect 287247 263229 287259 263263
rect 287201 263223 287259 263229
rect 296953 263263 297011 263269
rect 296953 263229 296965 263263
rect 296999 263260 297011 263263
rect 302657 263263 302715 263269
rect 302657 263260 302669 263263
rect 296999 263232 302669 263260
rect 296999 263229 297011 263232
rect 296953 263223 297011 263229
rect 302657 263229 302669 263232
rect 302703 263229 302715 263263
rect 302657 263223 302715 263229
rect 225926 262880 225932 262932
rect 225984 262920 225990 262932
rect 233470 262920 233476 262932
rect 225984 262892 233476 262920
rect 225984 262880 225990 262892
rect 233470 262880 233476 262892
rect 233528 262880 233534 262932
rect 132086 262744 132092 262796
rect 132144 262784 132150 262796
rect 139814 262784 139820 262796
rect 132144 262756 139820 262784
rect 132144 262744 132150 262756
rect 139814 262744 139820 262756
rect 139872 262744 139878 262796
rect 237797 262787 237855 262793
rect 237797 262753 237809 262787
rect 237843 262784 237855 262787
rect 263833 262787 263891 262793
rect 263833 262784 263845 262787
rect 237843 262756 263845 262784
rect 237843 262753 237855 262756
rect 237797 262747 237855 262753
rect 263833 262753 263845 262756
rect 263879 262753 263891 262787
rect 263833 262747 263891 262753
rect 13314 262676 13320 262728
rect 13372 262716 13378 262728
rect 372850 262716 372856 262728
rect 13372 262688 372856 262716
rect 13372 262676 13378 262688
rect 372850 262676 372856 262688
rect 372908 262676 372914 262728
rect 13406 262608 13412 262660
rect 13464 262648 13470 262660
rect 381130 262648 381136 262660
rect 13464 262620 381136 262648
rect 13464 262608 13470 262620
rect 381130 262608 381136 262620
rect 381188 262608 381194 262660
rect 13498 262540 13504 262592
rect 13556 262580 13562 262592
rect 385270 262580 385276 262592
rect 13556 262552 385276 262580
rect 13556 262540 13562 262552
rect 385270 262540 385276 262552
rect 385328 262540 385334 262592
rect 47078 262472 47084 262524
rect 47136 262512 47142 262524
rect 49194 262512 49200 262524
rect 47136 262484 49200 262512
rect 47136 262472 47142 262484
rect 49194 262472 49200 262484
rect 49252 262512 49258 262524
rect 73853 262515 73911 262521
rect 73853 262512 73865 262515
rect 49252 262484 73865 262512
rect 49252 262472 49258 262484
rect 73853 262481 73865 262484
rect 73899 262481 73911 262515
rect 73853 262475 73911 262481
rect 228594 262268 228600 262320
rect 228652 262308 228658 262320
rect 237797 262311 237855 262317
rect 237797 262308 237809 262311
rect 228652 262280 237809 262308
rect 228652 262268 228658 262280
rect 237797 262277 237809 262280
rect 237843 262277 237855 262311
rect 237797 262271 237855 262277
rect 263833 262311 263891 262317
rect 263833 262277 263845 262311
rect 263879 262308 263891 262311
rect 369722 262308 369728 262320
rect 263879 262280 369728 262308
rect 263879 262277 263891 262280
rect 263833 262271 263891 262277
rect 369722 262268 369728 262280
rect 369780 262268 369786 262320
rect 360430 261996 360436 262048
rect 360488 262036 360494 262048
rect 360798 262036 360804 262048
rect 360488 262008 360804 262036
rect 360488 261996 360494 262008
rect 360798 261996 360804 262008
rect 360856 262036 360862 262048
rect 422530 262036 422536 262048
rect 360856 262008 422536 262036
rect 360856 261996 360862 262008
rect 422530 261996 422536 262008
rect 422588 261996 422594 262048
rect 79738 261384 79744 261436
rect 79796 261424 79802 261436
rect 87190 261424 87196 261436
rect 79796 261396 87196 261424
rect 79796 261384 79802 261396
rect 87190 261384 87196 261396
rect 87248 261384 87254 261436
rect 131994 261384 132000 261436
rect 132052 261424 132058 261436
rect 140366 261424 140372 261436
rect 132052 261396 140372 261424
rect 132052 261384 132058 261396
rect 140366 261384 140372 261396
rect 140424 261384 140430 261436
rect 225834 261384 225840 261436
rect 225892 261424 225898 261436
rect 233470 261424 233476 261436
rect 225892 261396 233476 261424
rect 225892 261384 225898 261396
rect 233470 261384 233476 261396
rect 233528 261384 233534 261436
rect 95562 261316 95568 261368
rect 95620 261356 95626 261368
rect 96206 261356 96212 261368
rect 95620 261328 96212 261356
rect 95620 261316 95626 261328
rect 96206 261316 96212 261328
rect 96264 261316 96270 261368
rect 203846 261248 203852 261300
rect 203904 261288 203910 261300
rect 209918 261288 209924 261300
rect 203904 261260 209924 261288
rect 203904 261248 203910 261260
rect 209918 261248 209924 261260
rect 209976 261248 209982 261300
rect 297870 261248 297876 261300
rect 297928 261288 297934 261300
rect 303758 261288 303764 261300
rect 297928 261260 303764 261288
rect 297928 261248 297934 261260
rect 303758 261248 303764 261260
rect 303816 261248 303822 261300
rect 189310 260840 189316 260892
rect 189368 260880 189374 260892
rect 190506 260880 190512 260892
rect 189368 260852 190512 260880
rect 189368 260840 189374 260852
rect 190506 260840 190512 260852
rect 190564 260840 190570 260892
rect 217186 260636 217192 260688
rect 217244 260676 217250 260688
rect 225190 260676 225196 260688
rect 217244 260648 225196 260676
rect 217244 260636 217250 260648
rect 225190 260636 225196 260648
rect 225248 260636 225254 260688
rect 311210 260636 311216 260688
rect 311268 260676 311274 260688
rect 319214 260676 319220 260688
rect 311268 260648 319220 260676
rect 311268 260636 311274 260648
rect 319214 260636 319220 260648
rect 319272 260636 319278 260688
rect 123530 260568 123536 260620
rect 123588 260608 123594 260620
rect 127762 260608 127768 260620
rect 123588 260580 127768 260608
rect 123588 260568 123594 260580
rect 127762 260568 127768 260580
rect 127820 260568 127826 260620
rect 110190 260432 110196 260484
rect 110248 260472 110254 260484
rect 114790 260472 114796 260484
rect 110248 260444 114796 260472
rect 110248 260432 110254 260444
rect 114790 260432 114796 260444
rect 114848 260432 114854 260484
rect 79738 260024 79744 260076
rect 79796 260064 79802 260076
rect 85074 260064 85080 260076
rect 79796 260036 85080 260064
rect 79796 260024 79802 260036
rect 85074 260024 85080 260036
rect 85132 260024 85138 260076
rect 132362 260024 132368 260076
rect 132420 260064 132426 260076
rect 140366 260064 140372 260076
rect 132420 260036 140372 260064
rect 132420 260024 132426 260036
rect 140366 260024 140372 260036
rect 140424 260024 140430 260076
rect 226294 260024 226300 260076
rect 226352 260064 226358 260076
rect 233470 260064 233476 260076
rect 226352 260036 233476 260064
rect 226352 260024 226358 260036
rect 233470 260024 233476 260036
rect 233528 260024 233534 260076
rect 360522 259276 360528 259328
rect 360580 259316 360586 259328
rect 419770 259316 419776 259328
rect 360580 259288 419776 259316
rect 360580 259276 360586 259288
rect 419770 259276 419776 259288
rect 419828 259276 419834 259328
rect 79738 258664 79744 258716
rect 79796 258704 79802 258716
rect 84430 258704 84436 258716
rect 79796 258676 84436 258704
rect 79796 258664 79802 258676
rect 84430 258664 84436 258676
rect 84488 258664 84494 258716
rect 132638 258596 132644 258648
rect 132696 258636 132702 258648
rect 140550 258636 140556 258648
rect 132696 258608 140556 258636
rect 132696 258596 132702 258608
rect 140550 258596 140556 258608
rect 140608 258596 140614 258648
rect 226202 258596 226208 258648
rect 226260 258636 226266 258648
rect 233470 258636 233476 258648
rect 226260 258608 233476 258636
rect 226260 258596 226266 258608
rect 233470 258596 233476 258608
rect 233528 258596 233534 258648
rect 324550 258596 324556 258648
rect 324608 258636 324614 258648
rect 328414 258636 328420 258648
rect 324608 258608 328420 258636
rect 324608 258596 324614 258608
rect 328414 258596 328420 258608
rect 328472 258596 328478 258648
rect 321238 258392 321244 258444
rect 321296 258432 321302 258444
rect 327218 258432 327224 258444
rect 321296 258404 327224 258432
rect 321296 258392 321302 258404
rect 327218 258392 327224 258404
rect 327276 258392 327282 258444
rect 131350 257304 131356 257356
rect 131408 257344 131414 257356
rect 135122 257344 135128 257356
rect 131408 257316 135128 257344
rect 131408 257304 131414 257316
rect 135122 257304 135128 257316
rect 135180 257304 135186 257356
rect 132270 257236 132276 257288
rect 132328 257276 132334 257288
rect 140550 257276 140556 257288
rect 132328 257248 140556 257276
rect 132328 257236 132334 257248
rect 140550 257236 140556 257248
rect 140608 257236 140614 257288
rect 179190 257236 179196 257288
rect 179248 257276 179254 257288
rect 182318 257276 182324 257288
rect 179248 257248 182324 257276
rect 179248 257236 179254 257248
rect 182318 257236 182324 257248
rect 182376 257236 182382 257288
rect 226110 257236 226116 257288
rect 226168 257276 226174 257288
rect 233470 257276 233476 257288
rect 226168 257248 233476 257276
rect 226168 257236 226174 257248
rect 233470 257236 233476 257248
rect 233528 257236 233534 257288
rect 267142 257236 267148 257288
rect 267200 257276 267206 257288
rect 274870 257276 274876 257288
rect 267200 257248 274876 257276
rect 267200 257236 267206 257248
rect 274870 257236 274876 257248
rect 274928 257236 274934 257288
rect 321054 257168 321060 257220
rect 321112 257208 321118 257220
rect 326758 257208 326764 257220
rect 321112 257180 326764 257208
rect 321112 257168 321118 257180
rect 326758 257168 326764 257180
rect 326816 257168 326822 257220
rect 360614 257168 360620 257220
rect 360672 257208 360678 257220
rect 417010 257208 417016 257220
rect 360672 257180 417016 257208
rect 360672 257168 360678 257180
rect 417010 257168 417016 257180
rect 417068 257168 417074 257220
rect 85074 256828 85080 256880
rect 85132 256868 85138 256880
rect 87190 256868 87196 256880
rect 85132 256840 87196 256868
rect 85132 256828 85138 256840
rect 87190 256828 87196 256840
rect 87248 256828 87254 256880
rect 131718 256488 131724 256540
rect 131776 256528 131782 256540
rect 132362 256528 132368 256540
rect 131776 256500 132368 256528
rect 131776 256488 131782 256500
rect 132362 256488 132368 256500
rect 132420 256488 132426 256540
rect 225650 256488 225656 256540
rect 225708 256528 225714 256540
rect 226294 256528 226300 256540
rect 225708 256500 226300 256528
rect 225708 256488 225714 256500
rect 226294 256488 226300 256500
rect 226352 256488 226358 256540
rect 181030 256080 181036 256132
rect 181088 256120 181094 256132
rect 181674 256120 181680 256132
rect 181088 256092 181680 256120
rect 181088 256080 181094 256092
rect 181674 256080 181680 256092
rect 181732 256080 181738 256132
rect 136226 255944 136232 255996
rect 136284 255984 136290 255996
rect 140550 255984 140556 255996
rect 136284 255956 140556 255984
rect 136284 255944 136290 255956
rect 140550 255944 140556 255956
rect 140608 255944 140614 255996
rect 174038 255944 174044 255996
rect 174096 255984 174102 255996
rect 181030 255984 181036 255996
rect 174096 255956 181036 255984
rect 174096 255944 174102 255956
rect 181030 255944 181036 255956
rect 181088 255944 181094 255996
rect 229974 255944 229980 255996
rect 230032 255984 230038 255996
rect 233470 255984 233476 255996
rect 230032 255956 233476 255984
rect 230032 255944 230038 255956
rect 233470 255944 233476 255956
rect 233528 255944 233534 255996
rect 79738 255876 79744 255928
rect 79796 255916 79802 255928
rect 87374 255916 87380 255928
rect 79796 255888 87380 255916
rect 79796 255876 79802 255888
rect 87374 255876 87380 255888
rect 87432 255876 87438 255928
rect 132362 255876 132368 255928
rect 132420 255916 132426 255928
rect 139538 255916 139544 255928
rect 132420 255888 139544 255916
rect 132420 255876 132426 255888
rect 139538 255876 139544 255888
rect 139596 255876 139602 255928
rect 178270 255876 178276 255928
rect 178328 255916 178334 255928
rect 182318 255916 182324 255928
rect 178328 255888 182324 255916
rect 178328 255876 178334 255888
rect 182318 255876 182324 255888
rect 182376 255876 182382 255928
rect 226294 255876 226300 255928
rect 226352 255916 226358 255928
rect 233562 255916 233568 255928
rect 226352 255888 233568 255916
rect 226352 255876 226358 255888
rect 233562 255876 233568 255888
rect 233620 255876 233626 255928
rect 266590 255876 266596 255928
rect 266648 255916 266654 255928
rect 275698 255916 275704 255928
rect 266648 255888 275704 255916
rect 266648 255876 266654 255888
rect 275698 255876 275704 255888
rect 275756 255876 275762 255928
rect 80290 255808 80296 255860
rect 80348 255848 80354 255860
rect 87190 255848 87196 255860
rect 80348 255820 87196 255848
rect 80348 255808 80354 255820
rect 87190 255808 87196 255820
rect 87248 255808 87254 255860
rect 320686 255808 320692 255860
rect 320744 255848 320750 255860
rect 327218 255848 327224 255860
rect 320744 255820 327224 255848
rect 320744 255808 320750 255820
rect 327218 255808 327224 255820
rect 327276 255808 327282 255860
rect 84430 255740 84436 255792
rect 84488 255780 84494 255792
rect 87282 255780 87288 255792
rect 84488 255752 87288 255780
rect 84488 255740 84494 255752
rect 87282 255740 87288 255752
rect 87340 255740 87346 255792
rect 320870 255604 320876 255656
rect 320928 255644 320934 255656
rect 324550 255644 324556 255656
rect 320928 255616 324556 255644
rect 320928 255604 320934 255616
rect 324550 255604 324556 255616
rect 324608 255604 324614 255656
rect 173118 255536 173124 255588
rect 173176 255576 173182 255588
rect 222706 255576 222712 255588
rect 173176 255548 222712 255576
rect 173176 255536 173182 255548
rect 222706 255536 222712 255548
rect 222764 255536 222770 255588
rect 226294 254584 226300 254636
rect 226352 254624 226358 254636
rect 234114 254624 234120 254636
rect 226352 254596 234120 254624
rect 226352 254584 226358 254596
rect 234114 254584 234120 254596
rect 234172 254584 234178 254636
rect 131442 254516 131448 254568
rect 131500 254556 131506 254568
rect 135030 254556 135036 254568
rect 131500 254528 135036 254556
rect 131500 254516 131506 254528
rect 135030 254516 135036 254528
rect 135088 254516 135094 254568
rect 173302 254516 173308 254568
rect 173360 254556 173366 254568
rect 182318 254556 182324 254568
rect 173360 254528 182324 254556
rect 173360 254516 173366 254528
rect 182318 254516 182324 254528
rect 182376 254516 182382 254568
rect 225558 254516 225564 254568
rect 225616 254556 225622 254568
rect 234298 254556 234304 254568
rect 225616 254528 234304 254556
rect 225616 254516 225622 254528
rect 234298 254516 234304 254528
rect 234356 254516 234362 254568
rect 131350 254448 131356 254500
rect 131408 254488 131414 254500
rect 134938 254488 134944 254500
rect 131408 254460 134944 254488
rect 131408 254448 131414 254460
rect 134938 254448 134944 254460
rect 134996 254448 135002 254500
rect 137514 254448 137520 254500
rect 137572 254488 137578 254500
rect 140550 254488 140556 254500
rect 137572 254460 140556 254488
rect 137572 254448 137578 254460
rect 140550 254448 140556 254460
rect 140608 254448 140614 254500
rect 173762 254448 173768 254500
rect 173820 254488 173826 254500
rect 176154 254488 176160 254500
rect 173820 254460 176160 254488
rect 173820 254448 173826 254460
rect 176154 254448 176160 254460
rect 176212 254448 176218 254500
rect 176246 254448 176252 254500
rect 176304 254488 176310 254500
rect 181582 254488 181588 254500
rect 176304 254460 181588 254488
rect 176304 254448 176310 254460
rect 181582 254448 181588 254460
rect 181640 254448 181646 254500
rect 266590 254448 266596 254500
rect 266648 254488 266654 254500
rect 272754 254488 272760 254500
rect 266648 254460 272760 254488
rect 266648 254448 266654 254460
rect 272754 254448 272760 254460
rect 272812 254448 272818 254500
rect 321606 253632 321612 253684
rect 321664 253672 321670 253684
rect 328046 253672 328052 253684
rect 321664 253644 328052 253672
rect 321664 253632 321670 253644
rect 328046 253632 328052 253644
rect 328104 253632 328110 253684
rect 172934 253224 172940 253276
rect 172992 253264 172998 253276
rect 174774 253264 174780 253276
rect 172992 253236 174780 253264
rect 172992 253224 172998 253236
rect 174774 253224 174780 253236
rect 174832 253224 174838 253276
rect 266590 253156 266596 253208
rect 266648 253196 266654 253208
rect 274226 253196 274232 253208
rect 266648 253168 274232 253196
rect 266648 253156 266654 253168
rect 274226 253156 274232 253168
rect 274284 253156 274290 253208
rect 79738 253088 79744 253140
rect 79796 253128 79802 253140
rect 79796 253100 84476 253128
rect 79796 253088 79802 253100
rect 84448 252992 84476 253100
rect 131350 253088 131356 253140
rect 131408 253128 131414 253140
rect 138894 253128 138900 253140
rect 131408 253100 138900 253128
rect 131408 253088 131414 253100
rect 138894 253088 138900 253100
rect 138952 253088 138958 253140
rect 178914 253088 178920 253140
rect 178972 253128 178978 253140
rect 181766 253128 181772 253140
rect 178972 253100 181772 253128
rect 178972 253088 178978 253100
rect 181766 253088 181772 253100
rect 181824 253088 181830 253140
rect 225374 253088 225380 253140
rect 225432 253128 225438 253140
rect 230066 253128 230072 253140
rect 225432 253100 230072 253128
rect 225432 253088 225438 253100
rect 230066 253088 230072 253100
rect 230124 253088 230130 253140
rect 231446 253088 231452 253140
rect 231504 253128 231510 253140
rect 234206 253128 234212 253140
rect 231504 253100 234212 253128
rect 231504 253088 231510 253100
rect 234206 253088 234212 253100
rect 234264 253088 234270 253140
rect 267878 253088 267884 253140
rect 267936 253128 267942 253140
rect 274870 253128 274876 253140
rect 267936 253100 274876 253128
rect 267936 253088 267942 253100
rect 274870 253088 274876 253100
rect 274928 253088 274934 253140
rect 267418 253020 267424 253072
rect 267476 253060 267482 253072
rect 267694 253060 267700 253072
rect 267476 253032 267700 253060
rect 267476 253020 267482 253032
rect 267694 253020 267700 253032
rect 267752 253020 267758 253072
rect 321606 253020 321612 253072
rect 321664 253060 321670 253072
rect 328414 253060 328420 253072
rect 321664 253032 328420 253060
rect 321664 253020 321670 253032
rect 328414 253020 328420 253032
rect 328472 253020 328478 253072
rect 361166 253020 361172 253072
rect 361224 253060 361230 253072
rect 414250 253060 414256 253072
rect 361224 253032 414256 253060
rect 361224 253020 361230 253032
rect 414250 253020 414256 253032
rect 414308 253020 414314 253072
rect 87282 252992 87288 253004
rect 84448 252964 87288 252992
rect 87282 252952 87288 252964
rect 87340 252952 87346 253004
rect 79830 252884 79836 252936
rect 79888 252924 79894 252936
rect 87190 252924 87196 252936
rect 79888 252896 87196 252924
rect 79888 252884 79894 252896
rect 87190 252884 87196 252896
rect 87248 252884 87254 252936
rect 321606 252000 321612 252052
rect 321664 252040 321670 252052
rect 327218 252040 327224 252052
rect 321664 252012 327224 252040
rect 321664 252000 321670 252012
rect 327218 252000 327224 252012
rect 327276 252000 327282 252052
rect 173670 251864 173676 251916
rect 173728 251904 173734 251916
rect 180294 251904 180300 251916
rect 173728 251876 180300 251904
rect 173728 251864 173734 251876
rect 180294 251864 180300 251876
rect 180352 251864 180358 251916
rect 131350 251796 131356 251848
rect 131408 251836 131414 251848
rect 136318 251836 136324 251848
rect 131408 251808 136324 251836
rect 131408 251796 131414 251808
rect 136318 251796 136324 251808
rect 136376 251796 136382 251848
rect 179006 251796 179012 251848
rect 179064 251836 179070 251848
rect 181582 251836 181588 251848
rect 179064 251808 181588 251836
rect 179064 251796 179070 251808
rect 181582 251796 181588 251808
rect 181640 251796 181646 251848
rect 79738 251728 79744 251780
rect 79796 251768 79802 251780
rect 79796 251740 85764 251768
rect 79796 251728 79802 251740
rect 85736 251700 85764 251740
rect 173578 251728 173584 251780
rect 173636 251768 173642 251780
rect 181766 251768 181772 251780
rect 173636 251740 181772 251768
rect 173636 251728 173642 251740
rect 181766 251728 181772 251740
rect 181824 251728 181830 251780
rect 225742 251728 225748 251780
rect 225800 251768 225806 251780
rect 234114 251768 234120 251780
rect 225800 251740 234120 251768
rect 225800 251728 225806 251740
rect 234114 251728 234120 251740
rect 234172 251728 234178 251780
rect 266590 251728 266596 251780
rect 266648 251768 266654 251780
rect 272846 251768 272852 251780
rect 266648 251740 272852 251768
rect 266648 251728 266654 251740
rect 272846 251728 272852 251740
rect 272904 251728 272910 251780
rect 87190 251700 87196 251712
rect 85736 251672 87196 251700
rect 87190 251660 87196 251672
rect 87248 251660 87254 251712
rect 13130 251456 13136 251508
rect 13188 251496 13194 251508
rect 17546 251496 17552 251508
rect 13188 251468 17552 251496
rect 13188 251456 13194 251468
rect 17546 251456 17552 251468
rect 17604 251456 17610 251508
rect 222798 250980 222804 251032
rect 222856 251020 222862 251032
rect 233470 251020 233476 251032
rect 222856 250992 233476 251020
rect 222856 250980 222862 250992
rect 233470 250980 233476 250992
rect 233528 250980 233534 251032
rect 320594 250572 320600 250624
rect 320652 250612 320658 250624
rect 327126 250612 327132 250624
rect 320652 250584 327132 250612
rect 320652 250572 320658 250584
rect 327126 250572 327132 250584
rect 327184 250572 327190 250624
rect 79738 250368 79744 250420
rect 79796 250408 79802 250420
rect 79796 250380 85764 250408
rect 79796 250368 79802 250380
rect 85736 250272 85764 250380
rect 173670 250300 173676 250352
rect 173728 250340 173734 250352
rect 182318 250340 182324 250352
rect 173728 250312 182324 250340
rect 173728 250300 173734 250312
rect 182318 250300 182324 250312
rect 182376 250300 182382 250352
rect 87190 250272 87196 250284
rect 85736 250244 87196 250272
rect 87190 250232 87196 250244
rect 87248 250232 87254 250284
rect 135122 250232 135128 250284
rect 135180 250272 135186 250284
rect 140550 250272 140556 250284
rect 135180 250244 140556 250272
rect 135180 250232 135186 250244
rect 140550 250232 140556 250244
rect 140608 250232 140614 250284
rect 173394 250232 173400 250284
rect 173452 250272 173458 250284
rect 181490 250272 181496 250284
rect 173452 250244 181496 250272
rect 173452 250232 173458 250244
rect 181490 250232 181496 250244
rect 181548 250232 181554 250284
rect 226386 250232 226392 250284
rect 226444 250272 226450 250284
rect 233470 250272 233476 250284
rect 226444 250244 233476 250272
rect 226444 250232 226450 250244
rect 233470 250232 233476 250244
rect 233528 250232 233534 250284
rect 267510 250232 267516 250284
rect 267568 250272 267574 250284
rect 274870 250272 274876 250284
rect 267568 250244 274876 250272
rect 267568 250232 267574 250244
rect 274870 250232 274876 250244
rect 274928 250232 274934 250284
rect 361442 250232 361448 250284
rect 361500 250272 361506 250284
rect 412870 250272 412876 250284
rect 361500 250244 412876 250272
rect 361500 250232 361506 250244
rect 412870 250232 412876 250244
rect 412928 250232 412934 250284
rect 77254 249552 77260 249604
rect 77312 249592 77318 249604
rect 87190 249592 87196 249604
rect 77312 249564 87196 249592
rect 77312 249552 77318 249564
rect 87190 249552 87196 249564
rect 87248 249552 87254 249604
rect 321054 249484 321060 249536
rect 321112 249524 321118 249536
rect 327218 249524 327224 249536
rect 321112 249496 327224 249524
rect 321112 249484 321118 249496
rect 327218 249484 327224 249496
rect 327276 249484 327282 249536
rect 173302 249416 173308 249468
rect 173360 249456 173366 249468
rect 179190 249456 179196 249468
rect 173360 249428 179196 249456
rect 173360 249416 173366 249428
rect 179190 249416 179196 249428
rect 179248 249416 179254 249468
rect 321606 249076 321612 249128
rect 321664 249116 321670 249128
rect 328414 249116 328420 249128
rect 321664 249088 328420 249116
rect 321664 249076 321670 249088
rect 328414 249076 328420 249088
rect 328472 249076 328478 249128
rect 131994 248940 132000 248992
rect 132052 248980 132058 248992
rect 136134 248980 136140 248992
rect 132052 248952 136140 248980
rect 132052 248940 132058 248952
rect 136134 248940 136140 248952
rect 136192 248940 136198 248992
rect 174038 248940 174044 248992
rect 174096 248980 174102 248992
rect 182226 248980 182232 248992
rect 174096 248952 182232 248980
rect 174096 248940 174102 248952
rect 182226 248940 182232 248952
rect 182284 248940 182290 248992
rect 225374 248940 225380 248992
rect 225432 248980 225438 248992
rect 227306 248980 227312 248992
rect 225432 248952 227312 248980
rect 225432 248940 225438 248952
rect 227306 248940 227312 248952
rect 227364 248940 227370 248992
rect 173486 248872 173492 248924
rect 173544 248912 173550 248924
rect 181950 248912 181956 248924
rect 173544 248884 181956 248912
rect 173544 248872 173550 248884
rect 181950 248872 181956 248884
rect 182008 248872 182014 248924
rect 267602 248872 267608 248924
rect 267660 248912 267666 248924
rect 274962 248912 274968 248924
rect 267660 248884 274968 248912
rect 267660 248872 267666 248884
rect 274962 248872 274968 248884
rect 275020 248872 275026 248924
rect 173762 248804 173768 248856
rect 173820 248844 173826 248856
rect 181858 248844 181864 248856
rect 173820 248816 181864 248844
rect 173820 248804 173826 248816
rect 181858 248804 181864 248816
rect 181916 248804 181922 248856
rect 267694 248804 267700 248856
rect 267752 248844 267758 248856
rect 274870 248844 274876 248856
rect 267752 248816 274876 248844
rect 267752 248804 267758 248816
rect 274870 248804 274876 248816
rect 274928 248804 274934 248856
rect 266590 248736 266596 248788
rect 266648 248776 266654 248788
rect 275054 248776 275060 248788
rect 266648 248748 275060 248776
rect 266648 248736 266654 248748
rect 275054 248736 275060 248748
rect 275112 248736 275118 248788
rect 77254 248192 77260 248244
rect 77312 248232 77318 248244
rect 87190 248232 87196 248244
rect 77312 248204 87196 248232
rect 77312 248192 77318 248204
rect 87190 248192 87196 248204
rect 87248 248192 87254 248244
rect 173302 247852 173308 247904
rect 173360 247892 173366 247904
rect 178270 247892 178276 247904
rect 173360 247864 178276 247892
rect 173360 247852 173366 247864
rect 178270 247852 178276 247864
rect 178328 247852 178334 247904
rect 321606 247648 321612 247700
rect 321664 247688 321670 247700
rect 328414 247688 328420 247700
rect 321664 247660 328420 247688
rect 321664 247648 321670 247660
rect 328414 247648 328420 247660
rect 328472 247648 328478 247700
rect 77254 247512 77260 247564
rect 77312 247552 77318 247564
rect 88478 247552 88484 247564
rect 77312 247524 88484 247552
rect 77312 247512 77318 247524
rect 88478 247512 88484 247524
rect 88536 247512 88542 247564
rect 173854 247512 173860 247564
rect 173912 247552 173918 247564
rect 182318 247552 182324 247564
rect 173912 247524 182324 247552
rect 173912 247512 173918 247524
rect 182318 247512 182324 247524
rect 182376 247512 182382 247564
rect 266590 247512 266596 247564
rect 266648 247552 266654 247564
rect 275882 247552 275888 247564
rect 266648 247524 275888 247552
rect 266648 247512 266654 247524
rect 275882 247512 275888 247524
rect 275940 247512 275946 247564
rect 321790 247512 321796 247564
rect 321848 247552 321854 247564
rect 328414 247552 328420 247564
rect 321848 247524 328420 247552
rect 321848 247512 321854 247524
rect 328414 247512 328420 247524
rect 328472 247512 328478 247564
rect 267694 247444 267700 247496
rect 267752 247484 267758 247496
rect 274870 247484 274876 247496
rect 267752 247456 274876 247484
rect 267752 247444 267758 247456
rect 274870 247444 274876 247456
rect 274928 247444 274934 247496
rect 135030 247308 135036 247360
rect 135088 247348 135094 247360
rect 140642 247348 140648 247360
rect 135088 247320 140648 247348
rect 135088 247308 135094 247320
rect 140642 247308 140648 247320
rect 140700 247308 140706 247360
rect 173670 246900 173676 246952
rect 173728 246940 173734 246952
rect 176246 246940 176252 246952
rect 173728 246912 176252 246940
rect 173728 246900 173734 246912
rect 176246 246900 176252 246912
rect 176304 246900 176310 246952
rect 321238 246220 321244 246272
rect 321296 246260 321302 246272
rect 321296 246232 321836 246260
rect 321296 246220 321302 246232
rect 78910 246152 78916 246204
rect 78968 246192 78974 246204
rect 87190 246192 87196 246204
rect 78968 246164 87196 246192
rect 78968 246152 78974 246164
rect 87190 246152 87196 246164
rect 87248 246152 87254 246204
rect 134938 246152 134944 246204
rect 134996 246192 135002 246204
rect 140550 246192 140556 246204
rect 134996 246164 140556 246192
rect 134996 246152 135002 246164
rect 140550 246152 140556 246164
rect 140608 246152 140614 246204
rect 173946 246152 173952 246204
rect 174004 246192 174010 246204
rect 181674 246192 181680 246204
rect 174004 246164 181680 246192
rect 174004 246152 174010 246164
rect 181674 246152 181680 246164
rect 181732 246152 181738 246204
rect 267786 246152 267792 246204
rect 267844 246192 267850 246204
rect 274870 246192 274876 246204
rect 267844 246164 274876 246192
rect 267844 246152 267850 246164
rect 274870 246152 274876 246164
rect 274928 246152 274934 246204
rect 321808 246192 321836 246232
rect 327862 246192 327868 246204
rect 321808 246164 327868 246192
rect 327862 246152 327868 246164
rect 327920 246152 327926 246204
rect 427498 246152 427504 246204
rect 427556 246192 427562 246204
rect 429430 246192 429436 246204
rect 427556 246164 429436 246192
rect 427556 246152 427562 246164
rect 429430 246152 429436 246164
rect 429488 246152 429494 246204
rect 131350 246084 131356 246136
rect 131408 246124 131414 246136
rect 136226 246124 136232 246136
rect 131408 246096 136232 246124
rect 131408 246084 131414 246096
rect 136226 246084 136232 246096
rect 136284 246084 136290 246136
rect 266590 246084 266596 246136
rect 266648 246124 266654 246136
rect 274410 246124 274416 246136
rect 266648 246096 274416 246124
rect 266648 246084 266654 246096
rect 274410 246084 274416 246096
rect 274468 246084 274474 246136
rect 225374 245472 225380 245524
rect 225432 245512 225438 245524
rect 229974 245512 229980 245524
rect 225432 245484 229980 245512
rect 225432 245472 225438 245484
rect 229974 245472 229980 245484
rect 230032 245472 230038 245524
rect 321698 244860 321704 244912
rect 321756 244900 321762 244912
rect 323170 244900 323176 244912
rect 321756 244872 323176 244900
rect 321756 244860 321762 244872
rect 323170 244860 323176 244872
rect 323228 244860 323234 244912
rect 80198 244792 80204 244844
rect 80256 244832 80262 244844
rect 87190 244832 87196 244844
rect 80256 244804 87196 244832
rect 80256 244792 80262 244804
rect 87190 244792 87196 244804
rect 87248 244792 87254 244844
rect 321606 244792 321612 244844
rect 321664 244832 321670 244844
rect 321664 244804 321836 244832
rect 321664 244792 321670 244804
rect 78910 244724 78916 244776
rect 78968 244764 78974 244776
rect 87282 244764 87288 244776
rect 78968 244736 87288 244764
rect 78968 244724 78974 244736
rect 87282 244724 87288 244736
rect 87340 244724 87346 244776
rect 131350 244724 131356 244776
rect 131408 244764 131414 244776
rect 137514 244764 137520 244776
rect 131408 244736 137520 244764
rect 131408 244724 131414 244736
rect 137514 244724 137520 244736
rect 137572 244724 137578 244776
rect 225558 244724 225564 244776
rect 225616 244764 225622 244776
rect 232734 244764 232740 244776
rect 225616 244736 232740 244764
rect 225616 244724 225622 244736
rect 232734 244724 232740 244736
rect 232792 244724 232798 244776
rect 272754 244724 272760 244776
rect 272812 244764 272818 244776
rect 274870 244764 274876 244776
rect 272812 244736 274876 244764
rect 272812 244724 272818 244736
rect 274870 244724 274876 244736
rect 274928 244724 274934 244776
rect 321808 244764 321836 244804
rect 327862 244764 327868 244776
rect 321808 244736 327868 244764
rect 327862 244724 327868 244736
rect 327920 244724 327926 244776
rect 176154 244656 176160 244708
rect 176212 244696 176218 244708
rect 182042 244696 182048 244708
rect 176212 244668 182048 244696
rect 176212 244656 176218 244668
rect 182042 244656 182048 244668
rect 182100 244656 182106 244708
rect 230066 244656 230072 244708
rect 230124 244696 230130 244708
rect 233562 244696 233568 244708
rect 230124 244668 233568 244696
rect 230124 244656 230130 244668
rect 233562 244656 233568 244668
rect 233620 244656 233626 244708
rect 173302 244384 173308 244436
rect 173360 244424 173366 244436
rect 178914 244424 178920 244436
rect 173360 244396 178920 244424
rect 173360 244384 173366 244396
rect 178914 244384 178920 244396
rect 178972 244384 178978 244436
rect 321606 243432 321612 243484
rect 321664 243472 321670 243484
rect 327034 243472 327040 243484
rect 321664 243444 327040 243472
rect 321664 243432 321670 243444
rect 327034 243432 327040 243444
rect 327092 243432 327098 243484
rect 136318 243364 136324 243416
rect 136376 243404 136382 243416
rect 140642 243404 140648 243416
rect 136376 243376 140648 243404
rect 136376 243364 136382 243376
rect 140642 243364 140648 243376
rect 140700 243364 140706 243416
rect 174774 243364 174780 243416
rect 174832 243404 174838 243416
rect 181030 243404 181036 243416
rect 174832 243376 181036 243404
rect 174832 243364 174838 243376
rect 181030 243364 181036 243376
rect 181088 243364 181094 243416
rect 226386 243364 226392 243416
rect 226444 243404 226450 243416
rect 232826 243404 232832 243416
rect 226444 243376 232832 243404
rect 226444 243364 226450 243376
rect 232826 243364 232832 243376
rect 232884 243364 232890 243416
rect 272846 243364 272852 243416
rect 272904 243404 272910 243416
rect 275790 243404 275796 243416
rect 272904 243376 275796 243404
rect 272904 243364 272910 243376
rect 275790 243364 275796 243376
rect 275848 243364 275854 243416
rect 323170 243364 323176 243416
rect 323228 243404 323234 243416
rect 327862 243404 327868 243416
rect 323228 243376 327868 243404
rect 323228 243364 323234 243376
rect 327862 243364 327868 243376
rect 327920 243364 327926 243416
rect 132638 243296 132644 243348
rect 132696 243336 132702 243348
rect 140458 243336 140464 243348
rect 132696 243308 140464 243336
rect 132696 243296 132702 243308
rect 140458 243296 140464 243308
rect 140516 243296 140522 243348
rect 267878 243228 267884 243280
rect 267936 243268 267942 243280
rect 274318 243268 274324 243280
rect 267936 243240 274324 243268
rect 267936 243228 267942 243240
rect 274318 243228 274324 243240
rect 274376 243228 274382 243280
rect 131902 243160 131908 243212
rect 131960 243200 131966 243212
rect 140550 243200 140556 243212
rect 131960 243172 140556 243200
rect 131960 243160 131966 243172
rect 140550 243160 140556 243172
rect 140608 243160 140614 243212
rect 226294 243092 226300 243144
rect 226352 243132 226358 243144
rect 231446 243132 231452 243144
rect 226352 243104 231452 243132
rect 226352 243092 226358 243104
rect 231446 243092 231452 243104
rect 231504 243092 231510 243144
rect 172934 242752 172940 242804
rect 172992 242792 172998 242804
rect 179006 242792 179012 242804
rect 172992 242764 179012 242792
rect 172992 242752 172998 242764
rect 179006 242752 179012 242764
rect 179064 242752 179070 242804
rect 321606 242208 321612 242260
rect 321664 242248 321670 242260
rect 327218 242248 327224 242260
rect 321664 242220 327224 242248
rect 321664 242208 321670 242220
rect 327218 242208 327224 242220
rect 327276 242208 327282 242260
rect 79002 242140 79008 242192
rect 79060 242180 79066 242192
rect 87282 242180 87288 242192
rect 79060 242152 87288 242180
rect 79060 242140 79066 242152
rect 87282 242140 87288 242152
rect 87340 242140 87346 242192
rect 79094 242072 79100 242124
rect 79152 242112 79158 242124
rect 87190 242112 87196 242124
rect 79152 242084 87196 242112
rect 79152 242072 79158 242084
rect 87190 242072 87196 242084
rect 87248 242072 87254 242124
rect 320502 242072 320508 242124
rect 320560 242112 320566 242124
rect 327126 242112 327132 242124
rect 320560 242084 327132 242112
rect 320560 242072 320566 242084
rect 327126 242072 327132 242084
rect 327184 242072 327190 242124
rect 123070 241596 123076 241648
rect 123128 241636 123134 241648
rect 124312 241636 124318 241648
rect 123128 241608 124318 241636
rect 123128 241596 123134 241608
rect 124312 241596 124318 241608
rect 124370 241596 124376 241648
rect 78910 240576 78916 240628
rect 78968 240616 78974 240628
rect 87374 240616 87380 240628
rect 78968 240588 87380 240616
rect 78968 240576 78974 240588
rect 87374 240576 87380 240588
rect 87432 240576 87438 240628
rect 133374 240576 133380 240628
rect 133432 240616 133438 240628
rect 140550 240616 140556 240628
rect 133432 240588 140556 240616
rect 133432 240576 133438 240588
rect 140550 240576 140556 240588
rect 140608 240576 140614 240628
rect 227214 240576 227220 240628
rect 227272 240616 227278 240628
rect 233470 240616 233476 240628
rect 227272 240588 233476 240616
rect 227272 240576 227278 240588
rect 233470 240576 233476 240588
rect 233528 240576 233534 240628
rect 267878 240576 267884 240628
rect 267936 240616 267942 240628
rect 275606 240616 275612 240628
rect 267936 240588 275612 240616
rect 267936 240576 267942 240588
rect 275606 240576 275612 240588
rect 275664 240576 275670 240628
rect 389870 240576 389876 240628
rect 389928 240616 389934 240628
rect 390698 240616 390704 240628
rect 389928 240588 390704 240616
rect 389928 240576 389934 240588
rect 390698 240576 390704 240588
rect 390756 240576 390762 240628
rect 393826 240576 393832 240628
rect 393884 240616 393890 240628
rect 394838 240616 394844 240628
rect 393884 240588 394844 240616
rect 393884 240576 393890 240588
rect 394838 240576 394844 240588
rect 394896 240576 394902 240628
rect 13314 240508 13320 240560
rect 13372 240548 13378 240560
rect 17454 240548 17460 240560
rect 13372 240520 17460 240548
rect 13372 240508 13378 240520
rect 17454 240508 17460 240520
rect 17512 240508 17518 240560
rect 368618 239896 368624 239948
rect 368676 239936 368682 239948
rect 377818 239936 377824 239948
rect 368676 239908 377824 239936
rect 368676 239896 368682 239908
rect 377818 239896 377824 239908
rect 377876 239896 377882 239948
rect 314890 239828 314896 239880
rect 314948 239868 314954 239880
rect 316086 239868 316092 239880
rect 314948 239840 316092 239868
rect 314948 239828 314954 239840
rect 316086 239828 316092 239840
rect 316144 239828 316150 239880
rect 185630 239284 185636 239336
rect 185688 239324 185694 239336
rect 186458 239324 186464 239336
rect 185688 239296 186464 239324
rect 185688 239284 185694 239296
rect 186458 239284 186464 239296
rect 186516 239284 186522 239336
rect 279654 239284 279660 239336
rect 279712 239324 279718 239336
rect 280298 239324 280304 239336
rect 279712 239296 280304 239324
rect 279712 239284 279718 239296
rect 280298 239284 280304 239296
rect 280356 239284 280362 239336
rect 132178 239216 132184 239268
rect 132236 239256 132242 239268
rect 140550 239256 140556 239268
rect 132236 239228 140556 239256
rect 132236 239216 132242 239228
rect 140550 239216 140556 239228
rect 140608 239216 140614 239268
rect 226018 239216 226024 239268
rect 226076 239256 226082 239268
rect 233470 239256 233476 239268
rect 226076 239228 233476 239256
rect 226076 239216 226082 239228
rect 233470 239216 233476 239228
rect 233528 239216 233534 239268
rect 267878 239216 267884 239268
rect 267936 239256 267942 239268
rect 275514 239256 275520 239268
rect 267936 239228 275520 239256
rect 267936 239216 267942 239228
rect 275514 239216 275520 239228
rect 275572 239216 275578 239268
rect 136134 239148 136140 239200
rect 136192 239188 136198 239200
rect 140182 239188 140188 239200
rect 136192 239160 140188 239188
rect 136192 239148 136198 239160
rect 140182 239148 140188 239160
rect 140240 239148 140246 239200
rect 227306 239148 227312 239200
rect 227364 239188 227370 239200
rect 233562 239188 233568 239200
rect 227364 239160 233568 239188
rect 227364 239148 227370 239160
rect 233562 239148 233568 239160
rect 233620 239148 233626 239200
rect 267510 239148 267516 239200
rect 267568 239188 267574 239200
rect 274134 239188 274140 239200
rect 267568 239160 274140 239188
rect 267568 239148 267574 239160
rect 274134 239148 274140 239160
rect 274192 239148 274198 239200
rect 136962 238604 136968 238656
rect 137020 238644 137026 238656
rect 142390 238644 142396 238656
rect 137020 238616 142396 238644
rect 137020 238604 137026 238616
rect 142390 238604 142396 238616
rect 142448 238644 142454 238656
rect 142758 238644 142764 238656
rect 142448 238616 142764 238644
rect 142448 238604 142454 238616
rect 142758 238604 142764 238616
rect 142816 238604 142822 238656
rect 294190 238604 294196 238656
rect 294248 238644 294254 238656
rect 325194 238644 325200 238656
rect 294248 238616 325200 238644
rect 294248 238604 294254 238616
rect 325194 238604 325200 238616
rect 325252 238604 325258 238656
rect 200166 238536 200172 238588
rect 200224 238576 200230 238588
rect 230894 238576 230900 238588
rect 200224 238548 230900 238576
rect 200224 238536 200230 238548
rect 230894 238536 230900 238548
rect 230952 238536 230958 238588
rect 286922 238536 286928 238588
rect 286980 238576 286986 238588
rect 325562 238576 325568 238588
rect 286980 238548 325568 238576
rect 286980 238536 286986 238548
rect 325562 238536 325568 238548
rect 325620 238536 325626 238588
rect 127854 237176 127860 237228
rect 127912 237216 127918 237228
rect 140366 237216 140372 237228
rect 127912 237188 140372 237216
rect 127912 237176 127918 237188
rect 140366 237176 140372 237188
rect 140424 237176 140430 237228
rect 172934 237176 172940 237228
rect 172992 237216 172998 237228
rect 219762 237216 219768 237228
rect 172992 237188 219768 237216
rect 172992 237176 172998 237188
rect 219762 237176 219768 237188
rect 219820 237216 219826 237228
rect 233470 237216 233476 237228
rect 219820 237188 233476 237216
rect 219820 237176 219826 237188
rect 233470 237176 233476 237188
rect 233528 237176 233534 237228
rect 267326 237176 267332 237228
rect 267384 237216 267390 237228
rect 316270 237216 316276 237228
rect 267384 237188 316276 237216
rect 267384 237176 267390 237188
rect 316270 237176 316276 237188
rect 316328 237176 316334 237228
rect 78910 236564 78916 236616
rect 78968 236604 78974 236616
rect 127854 236604 127860 236616
rect 78968 236576 127860 236604
rect 78968 236564 78974 236576
rect 127854 236564 127860 236576
rect 127912 236604 127918 236616
rect 128130 236604 128136 236616
rect 127912 236576 128136 236604
rect 127912 236564 127918 236576
rect 128130 236564 128136 236576
rect 128188 236564 128194 236616
rect 316270 236564 316276 236616
rect 316328 236604 316334 236616
rect 328414 236604 328420 236616
rect 316328 236576 328420 236604
rect 316328 236564 316334 236576
rect 328414 236564 328420 236576
rect 328472 236564 328478 236616
rect 297686 236332 297692 236344
rect 262560 236304 297692 236332
rect 262560 236208 262588 236304
rect 297686 236292 297692 236304
rect 297744 236292 297750 236344
rect 262542 236156 262548 236208
rect 262600 236156 262606 236208
rect 203754 235816 203760 235868
rect 203812 235856 203818 235868
rect 230802 235856 230808 235868
rect 203812 235828 230808 235856
rect 203812 235816 203818 235828
rect 230802 235816 230808 235828
rect 230860 235856 230866 235868
rect 231998 235856 232004 235868
rect 230860 235828 232004 235856
rect 230860 235816 230866 235828
rect 231998 235816 232004 235828
rect 232056 235816 232062 235868
rect 297686 235816 297692 235868
rect 297744 235856 297750 235868
rect 325378 235856 325384 235868
rect 297744 235828 325384 235856
rect 297744 235816 297750 235828
rect 325378 235816 325384 235828
rect 325436 235816 325442 235868
rect 136962 235204 136968 235256
rect 137020 235244 137026 235256
rect 137146 235244 137152 235256
rect 137020 235216 137152 235244
rect 137020 235204 137026 235216
rect 137146 235204 137152 235216
rect 137204 235244 137210 235256
rect 148646 235244 148652 235256
rect 137204 235216 148652 235244
rect 137204 235204 137210 235216
rect 148646 235204 148652 235216
rect 148704 235244 148710 235256
rect 150670 235244 150676 235256
rect 148704 235216 150676 235244
rect 148704 235204 148710 235216
rect 150670 235204 150676 235216
rect 150728 235204 150734 235256
rect 149198 235136 149204 235188
rect 149256 235176 149262 235188
rect 196486 235176 196492 235188
rect 149256 235148 196492 235176
rect 149256 235136 149262 235148
rect 196486 235136 196492 235148
rect 196544 235136 196550 235188
rect 231998 235136 232004 235188
rect 232056 235176 232062 235188
rect 244970 235176 244976 235188
rect 232056 235148 244976 235176
rect 232056 235136 232062 235148
rect 244970 235136 244976 235148
rect 245028 235176 245034 235188
rect 262542 235176 262548 235188
rect 245028 235148 262548 235176
rect 245028 235136 245034 235148
rect 262542 235136 262548 235148
rect 262600 235136 262606 235188
rect 363834 235068 363840 235120
rect 363892 235108 363898 235120
rect 368710 235108 368716 235120
rect 363892 235080 368716 235108
rect 363892 235068 363898 235080
rect 368710 235068 368716 235080
rect 368768 235068 368774 235120
rect 113502 234496 113508 234508
rect 73592 234468 113508 234496
rect 46894 234388 46900 234440
rect 46952 234428 46958 234440
rect 73482 234428 73488 234440
rect 46952 234400 73488 234428
rect 46952 234388 46958 234400
rect 73482 234388 73488 234400
rect 73540 234428 73546 234440
rect 73592 234428 73620 234468
rect 113502 234456 113508 234468
rect 113560 234496 113566 234508
rect 137330 234496 137336 234508
rect 113560 234468 137336 234496
rect 113560 234456 113566 234468
rect 137330 234456 137336 234468
rect 137388 234496 137394 234508
rect 139262 234496 139268 234508
rect 137388 234468 139268 234496
rect 137388 234456 137394 234468
rect 139262 234456 139268 234468
rect 139320 234456 139326 234508
rect 73540 234400 73620 234428
rect 73540 234388 73546 234400
rect 74402 234388 74408 234440
rect 74460 234428 74466 234440
rect 117090 234428 117096 234440
rect 74460 234400 117096 234428
rect 74460 234388 74466 234400
rect 117090 234388 117096 234400
rect 117148 234428 117154 234440
rect 137698 234428 137704 234440
rect 117148 234400 137704 234428
rect 117148 234388 117154 234400
rect 137698 234388 137704 234400
rect 137756 234388 137762 234440
rect 207250 234388 207256 234440
rect 207308 234428 207314 234440
rect 231170 234428 231176 234440
rect 207308 234400 231176 234428
rect 207308 234388 207314 234400
rect 231170 234388 231176 234400
rect 231228 234428 231234 234440
rect 231814 234428 231820 234440
rect 231228 234400 231820 234428
rect 231228 234388 231234 234400
rect 231814 234388 231820 234400
rect 231872 234388 231878 234440
rect 302010 234388 302016 234440
rect 302068 234428 302074 234440
rect 324550 234428 324556 234440
rect 302068 234400 324556 234428
rect 302068 234388 302074 234400
rect 324550 234388 324556 234400
rect 324608 234388 324614 234440
rect 346538 234388 346544 234440
rect 346596 234428 346602 234440
rect 360522 234428 360528 234440
rect 346596 234400 360528 234428
rect 346596 234388 346602 234400
rect 360522 234388 360528 234400
rect 360580 234388 360586 234440
rect 221050 233776 221056 233828
rect 221108 233816 221114 233828
rect 222154 233816 222160 233828
rect 221108 233788 222160 233816
rect 221108 233776 221114 233788
rect 222154 233776 222160 233788
rect 222212 233776 222218 233828
rect 324550 233776 324556 233828
rect 324608 233816 324614 233828
rect 324734 233816 324740 233828
rect 324608 233788 324740 233816
rect 324608 233776 324614 233788
rect 324734 233776 324740 233788
rect 324792 233816 324798 233828
rect 345434 233816 345440 233828
rect 324792 233788 345440 233816
rect 324792 233776 324798 233788
rect 345434 233776 345440 233788
rect 345492 233816 345498 233828
rect 346538 233816 346544 233828
rect 345492 233788 346544 233816
rect 345492 233776 345498 233788
rect 346538 233776 346544 233788
rect 346596 233776 346602 233828
rect 138158 233708 138164 233760
rect 138216 233748 138222 233760
rect 146806 233748 146812 233760
rect 138216 233720 146812 233748
rect 138216 233708 138222 233720
rect 146806 233708 146812 233720
rect 146864 233708 146870 233760
rect 150578 233708 150584 233760
rect 150636 233748 150642 233760
rect 162262 233748 162268 233760
rect 150636 233720 162268 233748
rect 150636 233708 150642 233720
rect 162262 233708 162268 233720
rect 162320 233708 162326 233760
rect 234758 233708 234764 233760
rect 234816 233748 234822 233760
rect 241474 233748 241480 233760
rect 234816 233720 241480 233748
rect 234816 233708 234822 233720
rect 241474 233708 241480 233720
rect 241532 233708 241538 233760
rect 248926 233708 248932 233760
rect 248984 233748 248990 233760
rect 262082 233748 262088 233760
rect 248984 233720 262088 233748
rect 248984 233708 248990 233720
rect 262082 233708 262088 233720
rect 262140 233708 262146 233760
rect 268614 233708 268620 233760
rect 268672 233748 268678 233760
rect 368894 233748 368900 233760
rect 268672 233720 368900 233748
rect 268672 233708 268678 233720
rect 368894 233708 368900 233720
rect 368952 233708 368958 233760
rect 427406 233708 427412 233760
rect 427464 233748 427470 233760
rect 429798 233748 429804 233760
rect 427464 233720 429804 233748
rect 427464 233708 427470 233720
rect 429798 233708 429804 233720
rect 429856 233708 429862 233760
rect 62258 233640 62264 233692
rect 62316 233680 62322 233692
rect 74218 233680 74224 233692
rect 62316 233652 74224 233680
rect 62316 233640 62322 233652
rect 74218 233640 74224 233652
rect 74276 233640 74282 233692
rect 157478 233640 157484 233692
rect 157536 233680 157542 233692
rect 169990 233680 169996 233692
rect 157536 233652 169996 233680
rect 157536 233640 157542 233652
rect 169990 233640 169996 233652
rect 170048 233640 170054 233692
rect 246258 233640 246264 233692
rect 246316 233680 246322 233692
rect 259230 233680 259236 233692
rect 246316 233652 259236 233680
rect 246316 233640 246322 233652
rect 259230 233640 259236 233652
rect 259288 233640 259294 233692
rect 322618 233640 322624 233692
rect 322676 233680 322682 233692
rect 368710 233680 368716 233692
rect 322676 233652 368716 233680
rect 322676 233640 322682 233652
rect 368710 233640 368716 233652
rect 368768 233640 368774 233692
rect 66950 233612 66956 233624
rect 56664 233584 66956 233612
rect 55358 233164 55364 233216
rect 55416 233204 55422 233216
rect 56664 233204 56692 233584
rect 66950 233572 66956 233584
rect 67008 233572 67014 233624
rect 160974 233572 160980 233624
rect 161032 233612 161038 233624
rect 163182 233612 163188 233624
rect 161032 233584 163188 233612
rect 161032 233572 161038 233584
rect 163182 233572 163188 233584
rect 163240 233572 163246 233624
rect 244418 233572 244424 233624
rect 244476 233612 244482 233624
rect 256286 233612 256292 233624
rect 244476 233584 256292 233612
rect 244476 233572 244482 233584
rect 256286 233572 256292 233584
rect 256344 233572 256350 233624
rect 323814 233572 323820 233624
rect 323872 233612 323878 233624
rect 368802 233612 368808 233624
rect 323872 233584 368808 233612
rect 323872 233572 323878 233584
rect 368802 233572 368808 233584
rect 368860 233572 368866 233624
rect 62810 233504 62816 233556
rect 62868 233544 62874 233556
rect 65846 233544 65852 233556
rect 62868 233516 65852 233544
rect 62868 233504 62874 233516
rect 65846 233504 65852 233516
rect 65904 233504 65910 233556
rect 153338 233504 153344 233556
rect 153396 233544 153402 233556
rect 166126 233544 166132 233556
rect 153396 233516 166132 233544
rect 153396 233504 153402 233516
rect 166126 233504 166132 233516
rect 166184 233504 166190 233556
rect 248006 233504 248012 233556
rect 248064 233544 248070 233556
rect 261162 233544 261168 233556
rect 248064 233516 261168 233544
rect 248064 233504 248070 233516
rect 261162 233504 261168 233516
rect 261220 233504 261226 233556
rect 64834 233436 64840 233488
rect 64892 233476 64898 233488
rect 67226 233476 67232 233488
rect 64892 233448 67232 233476
rect 64892 233436 64898 233448
rect 67226 233436 67232 233448
rect 67284 233436 67290 233488
rect 151958 233436 151964 233488
rect 152016 233476 152022 233488
rect 165206 233476 165212 233488
rect 152016 233448 165212 233476
rect 152016 233436 152022 233448
rect 165206 233436 165212 233448
rect 165264 233436 165270 233488
rect 250674 233436 250680 233488
rect 250732 233476 250738 233488
rect 264014 233476 264020 233488
rect 250732 233448 264020 233476
rect 250732 233436 250738 233448
rect 264014 233436 264020 233448
rect 264072 233436 264078 233488
rect 63822 233368 63828 233420
rect 63880 233408 63886 233420
rect 67134 233408 67140 233420
rect 63880 233380 67140 233408
rect 63880 233368 63886 233380
rect 67134 233368 67140 233380
rect 67192 233368 67198 233420
rect 154718 233368 154724 233420
rect 154776 233408 154782 233420
rect 167230 233408 167236 233420
rect 154776 233380 167236 233408
rect 154776 233368 154782 233380
rect 167230 233368 167236 233380
rect 167288 233368 167294 233420
rect 61798 233300 61804 233352
rect 61856 233340 61862 233352
rect 65754 233340 65760 233352
rect 61856 233312 65760 233340
rect 61856 233300 61862 233312
rect 65754 233300 65760 233312
rect 65812 233300 65818 233352
rect 75230 233340 75236 233352
rect 69912 233312 75236 233340
rect 56738 233232 56744 233284
rect 56796 233272 56802 233284
rect 67962 233272 67968 233284
rect 56796 233244 67968 233272
rect 56796 233232 56802 233244
rect 67962 233232 67968 233244
rect 68020 233232 68026 233284
rect 55416 233176 56692 233204
rect 55416 233164 55422 233176
rect 63638 233164 63644 233216
rect 63696 233204 63702 233216
rect 69912 233204 69940 233312
rect 75230 233300 75236 233312
rect 75288 233300 75294 233352
rect 150486 233300 150492 233352
rect 150544 233340 150550 233352
rect 156837 233343 156895 233349
rect 156837 233340 156849 233343
rect 150544 233312 156849 233340
rect 150544 233300 150550 233312
rect 156837 233309 156849 233312
rect 156883 233309 156895 233343
rect 156837 233303 156895 233309
rect 231446 233300 231452 233352
rect 231504 233340 231510 233352
rect 234758 233340 234764 233352
rect 231504 233312 234764 233340
rect 231504 233300 231510 233312
rect 234758 233300 234764 233312
rect 234816 233300 234822 233352
rect 249846 233300 249852 233352
rect 249904 233340 249910 233352
rect 263094 233340 263100 233352
rect 249904 233312 263100 233340
rect 249904 233300 249910 233312
rect 263094 233300 263100 233312
rect 263152 233300 263158 233352
rect 341018 233300 341024 233352
rect 341076 233340 341082 233352
rect 346814 233340 346820 233352
rect 341076 233312 346820 233340
rect 341076 233300 341082 233312
rect 346814 233300 346820 233312
rect 346872 233300 346878 233352
rect 151866 233232 151872 233284
rect 151924 233272 151930 233284
rect 164562 233272 164568 233284
rect 151924 233244 164568 233272
rect 151924 233232 151930 233244
rect 164562 233232 164568 233244
rect 164620 233232 164626 233284
rect 231722 233232 231728 233284
rect 231780 233272 231786 233284
rect 243038 233272 243044 233284
rect 231780 233244 243044 233272
rect 231780 233232 231786 233244
rect 243038 233232 243044 233244
rect 243096 233232 243102 233284
rect 245338 233232 245344 233284
rect 245396 233272 245402 233284
rect 258402 233272 258408 233284
rect 245396 233244 258408 233272
rect 245396 233232 245402 233244
rect 258402 233232 258408 233244
rect 258460 233232 258466 233284
rect 63696 233176 69940 233204
rect 63696 233164 63702 233176
rect 154626 233164 154632 233216
rect 154684 233204 154690 233216
rect 168058 233204 168064 233216
rect 154684 233176 168064 233204
rect 154684 233164 154690 233176
rect 168058 233164 168064 233176
rect 168116 233164 168122 233216
rect 231630 233164 231636 233216
rect 231688 233204 231694 233216
rect 242118 233204 242124 233216
rect 231688 233176 242124 233204
rect 231688 233164 231694 233176
rect 242118 233164 242124 233176
rect 242176 233164 242182 233216
rect 244326 233164 244332 233216
rect 244384 233204 244390 233216
rect 257298 233204 257304 233216
rect 244384 233176 257304 233204
rect 244384 233164 244390 233176
rect 257298 233164 257304 233176
rect 257356 233164 257362 233216
rect 58118 233096 58124 233148
rect 58176 233136 58182 233148
rect 70078 233136 70084 233148
rect 58176 233108 70084 233136
rect 58176 233096 58182 233108
rect 70078 233096 70084 233108
rect 70136 233096 70142 233148
rect 144598 233096 144604 233148
rect 144656 233136 144662 233148
rect 165114 233136 165120 233148
rect 144656 233108 165120 233136
rect 144656 233096 144662 233108
rect 165114 233096 165120 233108
rect 165172 233096 165178 233148
rect 238622 233096 238628 233148
rect 238680 233136 238686 233148
rect 258954 233136 258960 233148
rect 238680 233108 258960 233136
rect 238680 233096 238686 233108
rect 258954 233096 258960 233108
rect 259012 233096 259018 233148
rect 60786 233028 60792 233080
rect 60844 233068 60850 233080
rect 72102 233068 72108 233080
rect 60844 233040 72108 233068
rect 60844 233028 60850 233040
rect 72102 233028 72108 233040
rect 72160 233028 72166 233080
rect 74126 233028 74132 233080
rect 74184 233068 74190 233080
rect 75138 233068 75144 233080
rect 74184 233040 75144 233068
rect 74184 233028 74190 233040
rect 75138 233028 75144 233040
rect 75196 233068 75202 233080
rect 105130 233068 105136 233080
rect 75196 233040 105136 233068
rect 75196 233028 75202 233040
rect 105130 233028 105136 233040
rect 105188 233068 105194 233080
rect 137146 233068 137152 233080
rect 105188 233040 137152 233068
rect 105188 233028 105194 233040
rect 137146 233028 137152 233040
rect 137204 233028 137210 233080
rect 145242 233028 145248 233080
rect 145300 233068 145306 233080
rect 352886 233068 352892 233080
rect 145300 233040 352892 233068
rect 145300 233028 145306 233040
rect 352886 233028 352892 233040
rect 352944 233028 352950 233080
rect 340926 232960 340932 233012
rect 340984 233000 340990 233012
rect 347918 233000 347924 233012
rect 340984 232972 347924 233000
rect 340984 232960 340990 232972
rect 347918 232960 347924 232972
rect 347976 232960 347982 233012
rect 60878 232892 60884 232944
rect 60936 232932 60942 232944
rect 73114 232932 73120 232944
rect 60936 232904 73120 232932
rect 60936 232892 60942 232904
rect 73114 232892 73120 232904
rect 73172 232892 73178 232944
rect 156837 232935 156895 232941
rect 156837 232901 156849 232935
rect 156883 232932 156895 232935
rect 163274 232932 163280 232944
rect 156883 232904 163280 232932
rect 156883 232901 156895 232904
rect 156837 232895 156895 232901
rect 163274 232892 163280 232904
rect 163332 232892 163338 232944
rect 247086 232892 247092 232944
rect 247144 232932 247150 232944
rect 260150 232932 260156 232944
rect 247144 232904 260156 232932
rect 247144 232892 247150 232904
rect 260150 232892 260156 232904
rect 260208 232892 260214 232944
rect 59498 232824 59504 232876
rect 59556 232864 59562 232876
rect 71090 232864 71096 232876
rect 59556 232836 71096 232864
rect 59556 232824 59562 232836
rect 71090 232824 71096 232836
rect 71148 232824 71154 232876
rect 156006 232824 156012 232876
rect 156064 232864 156070 232876
rect 169070 232864 169076 232876
rect 156064 232836 169076 232864
rect 156064 232824 156070 232836
rect 169070 232824 169076 232836
rect 169128 232824 169134 232876
rect 160054 232756 160060 232808
rect 160112 232796 160118 232808
rect 161802 232796 161808 232808
rect 160112 232768 161808 232796
rect 160112 232756 160118 232768
rect 161802 232756 161808 232768
rect 161860 232756 161866 232808
rect 58670 232620 58676 232672
rect 58728 232660 58734 232672
rect 63178 232660 63184 232672
rect 58728 232632 63184 232660
rect 58728 232620 58734 232632
rect 63178 232620 63184 232632
rect 63236 232620 63242 232672
rect 156098 232620 156104 232672
rect 156156 232660 156162 232672
rect 158214 232660 158220 232672
rect 156156 232632 158220 232660
rect 156156 232620 156162 232632
rect 158214 232620 158220 232632
rect 158272 232620 158278 232672
rect 57658 232552 57664 232604
rect 57716 232592 57722 232604
rect 61614 232592 61620 232604
rect 57716 232564 61620 232592
rect 57716 232552 57722 232564
rect 61614 232552 61620 232564
rect 61672 232552 61678 232604
rect 157110 232552 157116 232604
rect 157168 232592 157174 232604
rect 159042 232592 159048 232604
rect 157168 232564 159048 232592
rect 157168 232552 157174 232564
rect 159042 232552 159048 232564
rect 159100 232552 159106 232604
rect 59682 232484 59688 232536
rect 59740 232524 59746 232536
rect 62994 232524 63000 232536
rect 59740 232496 63000 232524
rect 59740 232484 59746 232496
rect 62994 232484 63000 232496
rect 63052 232484 63058 232536
rect 65938 232484 65944 232536
rect 65996 232524 66002 232536
rect 68514 232524 68520 232536
rect 65996 232496 68520 232524
rect 65996 232484 66002 232496
rect 68514 232484 68520 232496
rect 68572 232484 68578 232536
rect 155178 232484 155184 232536
rect 155236 232524 155242 232536
rect 157570 232524 157576 232536
rect 155236 232496 157576 232524
rect 155236 232484 155242 232496
rect 157570 232484 157576 232496
rect 157628 232484 157634 232536
rect 158122 232484 158128 232536
rect 158180 232524 158186 232536
rect 160330 232524 160336 232536
rect 158180 232496 160336 232524
rect 158180 232484 158186 232496
rect 160330 232484 160336 232496
rect 160388 232484 160394 232536
rect 248282 232484 248288 232536
rect 248340 232524 248346 232536
rect 250122 232524 250128 232536
rect 248340 232496 250128 232524
rect 248340 232484 248346 232496
rect 250122 232484 250128 232496
rect 250180 232484 250186 232536
rect 338994 232484 339000 232536
rect 339052 232524 339058 232536
rect 341662 232524 341668 232536
rect 339052 232496 341668 232524
rect 339052 232484 339058 232496
rect 341662 232484 341668 232496
rect 341720 232484 341726 232536
rect 342858 232484 342864 232536
rect 342916 232524 342922 232536
rect 345802 232524 345808 232536
rect 342916 232496 345808 232524
rect 342916 232484 342922 232496
rect 345802 232484 345808 232496
rect 345860 232484 345866 232536
rect 346722 232484 346728 232536
rect 346780 232524 346786 232536
rect 349942 232524 349948 232536
rect 346780 232496 349948 232524
rect 346780 232484 346786 232496
rect 349942 232484 349948 232496
rect 350000 232484 350006 232536
rect 60694 232416 60700 232468
rect 60752 232456 60758 232468
rect 63086 232456 63092 232468
rect 60752 232428 63092 232456
rect 60752 232416 60758 232428
rect 63086 232416 63092 232428
rect 63144 232416 63150 232468
rect 67318 232416 67324 232468
rect 67376 232456 67382 232468
rect 68974 232456 68980 232468
rect 67376 232428 68980 232456
rect 67376 232416 67382 232428
rect 68974 232416 68980 232428
rect 69032 232416 69038 232468
rect 154258 232416 154264 232468
rect 154316 232456 154322 232468
rect 156374 232456 156380 232468
rect 154316 232428 156380 232456
rect 154316 232416 154322 232428
rect 156374 232416 156380 232428
rect 156432 232416 156438 232468
rect 158858 232416 158864 232468
rect 158916 232456 158922 232468
rect 160974 232456 160980 232468
rect 158916 232428 160980 232456
rect 158916 232416 158922 232428
rect 160974 232416 160980 232428
rect 161032 232416 161038 232468
rect 161986 232416 161992 232468
rect 162044 232456 162050 232468
rect 162998 232456 163004 232468
rect 162044 232428 163004 232456
rect 162044 232416 162050 232428
rect 162998 232416 163004 232428
rect 163056 232416 163062 232468
rect 239542 232416 239548 232468
rect 239600 232456 239606 232468
rect 240278 232456 240284 232468
rect 239600 232428 240284 232456
rect 239600 232416 239606 232428
rect 240278 232416 240284 232428
rect 240336 232416 240342 232468
rect 249938 232416 249944 232468
rect 249996 232456 250002 232468
rect 252882 232456 252888 232468
rect 249996 232428 252888 232456
rect 249996 232416 250002 232428
rect 252882 232416 252888 232428
rect 252940 232416 252946 232468
rect 333382 232416 333388 232468
rect 333440 232456 333446 232468
rect 334118 232456 334124 232468
rect 333440 232428 334124 232456
rect 333440 232416 333446 232428
rect 334118 232416 334124 232428
rect 334176 232416 334182 232468
rect 334394 232416 334400 232468
rect 334452 232456 334458 232468
rect 335406 232456 335412 232468
rect 334452 232428 335412 232456
rect 334452 232416 334458 232428
rect 335406 232416 335412 232428
rect 335464 232416 335470 232468
rect 338534 232416 338540 232468
rect 338592 232456 338598 232468
rect 339638 232456 339644 232468
rect 338592 232428 339644 232456
rect 338592 232416 338598 232428
rect 339638 232416 339644 232428
rect 339696 232416 339702 232468
rect 342950 232416 342956 232468
rect 343008 232456 343014 232468
rect 344790 232456 344796 232468
rect 343008 232428 344796 232456
rect 343008 232416 343014 232428
rect 344790 232416 344796 232428
rect 344848 232416 344854 232468
rect 346630 232416 346636 232468
rect 346688 232456 346694 232468
rect 348930 232456 348936 232468
rect 346688 232428 348936 232456
rect 346688 232416 346694 232428
rect 348930 232416 348936 232428
rect 348988 232416 348994 232468
rect 134846 232348 134852 232400
rect 134904 232388 134910 232400
rect 368894 232388 368900 232400
rect 134904 232360 368900 232388
rect 134904 232348 134910 232360
rect 368894 232348 368900 232360
rect 368952 232348 368958 232400
rect 265854 232280 265860 232332
rect 265912 232320 265918 232332
rect 368710 232320 368716 232332
rect 265912 232292 368716 232320
rect 265912 232280 265918 232292
rect 368710 232280 368716 232292
rect 368768 232280 368774 232332
rect 326574 232212 326580 232264
rect 326632 232252 326638 232264
rect 368802 232252 368808 232264
rect 326632 232224 368808 232252
rect 326632 232212 326638 232224
rect 368802 232212 368808 232224
rect 368860 232212 368866 232264
rect 354910 232008 354916 232060
rect 354968 232048 354974 232060
rect 355830 232048 355836 232060
rect 354968 232020 355836 232048
rect 354968 232008 354974 232020
rect 355830 232008 355836 232020
rect 355888 232008 355894 232060
rect 239634 231668 239640 231720
rect 239692 231708 239698 231720
rect 324642 231708 324648 231720
rect 239692 231680 324648 231708
rect 239692 231668 239698 231680
rect 324642 231668 324648 231680
rect 324700 231668 324706 231720
rect 345158 231668 345164 231720
rect 345216 231708 345222 231720
rect 360706 231708 360712 231720
rect 345216 231680 360712 231708
rect 345216 231668 345222 231680
rect 360706 231668 360712 231680
rect 360764 231668 360770 231720
rect 369998 231464 370004 231516
rect 370056 231464 370062 231516
rect 369906 231260 369912 231312
rect 369964 231300 369970 231312
rect 370016 231300 370044 231464
rect 369964 231272 370044 231300
rect 369964 231260 369970 231272
rect 222614 230988 222620 231040
rect 222672 231028 222678 231040
rect 222798 231028 222804 231040
rect 222672 231000 222804 231028
rect 222672 230988 222678 231000
rect 222798 230988 222804 231000
rect 222856 230988 222862 231040
rect 325562 230988 325568 231040
rect 325620 231028 325626 231040
rect 343962 231028 343968 231040
rect 325620 231000 343968 231028
rect 325620 230988 325626 231000
rect 343962 230988 343968 231000
rect 344020 231028 344026 231040
rect 345158 231028 345164 231040
rect 344020 231000 345164 231028
rect 344020 230988 344026 231000
rect 345158 230988 345164 231000
rect 345216 230988 345222 231040
rect 12854 230920 12860 230972
rect 12912 230960 12918 230972
rect 16166 230960 16172 230972
rect 12912 230932 16172 230960
rect 12912 230920 12918 230932
rect 16166 230920 16172 230932
rect 16224 230920 16230 230972
rect 47078 230920 47084 230972
rect 47136 230960 47142 230972
rect 368894 230960 368900 230972
rect 47136 230932 368900 230960
rect 47136 230920 47142 230932
rect 368894 230920 368900 230932
rect 368952 230920 368958 230972
rect 76794 230852 76800 230904
rect 76852 230892 76858 230904
rect 368710 230892 368716 230904
rect 76852 230864 368716 230892
rect 76852 230852 76858 230864
rect 368710 230852 368716 230864
rect 368768 230852 368774 230904
rect 134754 230784 134760 230836
rect 134812 230824 134818 230836
rect 368802 230824 368808 230836
rect 134812 230796 368808 230824
rect 134812 230784 134818 230796
rect 368802 230784 368808 230796
rect 368860 230784 368866 230836
rect 115986 230376 115992 230428
rect 116044 230416 116050 230428
rect 127210 230416 127216 230428
rect 116044 230388 127216 230416
rect 116044 230376 116050 230388
rect 127210 230376 127216 230388
rect 127268 230376 127274 230428
rect 210010 230376 210016 230428
rect 210068 230416 210074 230428
rect 221050 230416 221056 230428
rect 210068 230388 221056 230416
rect 210068 230376 210074 230388
rect 221050 230376 221056 230388
rect 221108 230376 221114 230428
rect 304034 230376 304040 230428
rect 304092 230416 304098 230428
rect 314890 230416 314896 230428
rect 304092 230388 314896 230416
rect 304092 230376 304098 230388
rect 314890 230376 314896 230388
rect 314948 230376 314954 230428
rect 103474 230308 103480 230360
rect 103532 230348 103538 230360
rect 123070 230348 123076 230360
rect 103532 230320 123076 230348
rect 103532 230308 103538 230320
rect 123070 230308 123076 230320
rect 123128 230308 123134 230360
rect 197498 230308 197504 230360
rect 197556 230348 197562 230360
rect 218290 230348 218296 230360
rect 197556 230320 218296 230348
rect 197556 230308 197562 230320
rect 218290 230308 218296 230320
rect 218348 230308 218354 230360
rect 291522 230308 291528 230360
rect 291580 230348 291586 230360
rect 312130 230348 312136 230360
rect 291580 230320 312136 230348
rect 291580 230308 291586 230320
rect 312130 230308 312136 230320
rect 312188 230308 312194 230360
rect 339638 230308 339644 230360
rect 339696 230348 339702 230360
rect 343137 230351 343195 230357
rect 343137 230348 343149 230351
rect 339696 230320 343149 230348
rect 339696 230308 339702 230320
rect 343137 230317 343149 230320
rect 343183 230317 343195 230351
rect 343137 230311 343195 230317
rect 91054 230240 91060 230292
rect 91112 230280 91118 230292
rect 120310 230280 120316 230292
rect 91112 230252 120316 230280
rect 91112 230240 91118 230252
rect 120310 230240 120316 230252
rect 120368 230240 120374 230292
rect 185078 230240 185084 230292
rect 185136 230280 185142 230292
rect 214150 230280 214156 230292
rect 185136 230252 214156 230280
rect 185136 230240 185142 230252
rect 214150 230240 214156 230252
rect 214208 230240 214214 230292
rect 279102 230240 279108 230292
rect 279160 230280 279166 230292
rect 307990 230280 307996 230292
rect 279160 230252 307996 230280
rect 279160 230240 279166 230252
rect 307990 230240 307996 230252
rect 308048 230240 308054 230292
rect 343778 230240 343784 230292
rect 343836 230280 343842 230292
rect 360798 230280 360804 230292
rect 343836 230252 360804 230280
rect 343836 230240 343842 230252
rect 360798 230240 360804 230252
rect 360856 230240 360862 230292
rect 324642 229628 324648 229680
rect 324700 229668 324706 229680
rect 325470 229668 325476 229680
rect 324700 229640 325476 229668
rect 324700 229628 324706 229640
rect 325470 229628 325476 229640
rect 325528 229668 325534 229680
rect 343042 229668 343048 229680
rect 325528 229640 343048 229668
rect 325528 229628 325534 229640
rect 343042 229628 343048 229640
rect 343100 229668 343106 229680
rect 343778 229668 343784 229680
rect 343100 229640 343784 229668
rect 343100 229628 343106 229640
rect 343778 229628 343784 229640
rect 343836 229628 343842 229680
rect 22238 229560 22244 229612
rect 22296 229600 22302 229612
rect 368710 229600 368716 229612
rect 22296 229572 368716 229600
rect 22296 229560 22302 229572
rect 368710 229560 368716 229572
rect 368768 229560 368774 229612
rect 74034 228404 74040 228456
rect 74092 228444 74098 228456
rect 368710 228444 368716 228456
rect 74092 228416 368716 228444
rect 74092 228404 74098 228416
rect 368710 228404 368716 228416
rect 368768 228404 368774 228456
rect 47078 228336 47084 228388
rect 47136 228376 47142 228388
rect 368802 228376 368808 228388
rect 47136 228348 368808 228376
rect 47136 228336 47142 228348
rect 368802 228336 368808 228348
rect 368860 228336 368866 228388
rect 34014 228268 34020 228320
rect 34072 228308 34078 228320
rect 368710 228308 368716 228320
rect 34072 228280 368716 228308
rect 34072 228268 34078 228280
rect 368710 228268 368716 228280
rect 368768 228268 368774 228320
rect 305138 227656 305144 227708
rect 305196 227696 305202 227708
rect 322986 227696 322992 227708
rect 305196 227668 322992 227696
rect 305196 227656 305202 227668
rect 322986 227656 322992 227668
rect 323044 227656 323050 227708
rect 346998 227656 347004 227708
rect 347056 227696 347062 227708
rect 360430 227696 360436 227708
rect 347056 227668 360436 227696
rect 347056 227656 347062 227668
rect 360430 227656 360436 227668
rect 360488 227656 360494 227708
rect 222430 227588 222436 227640
rect 222488 227628 222494 227640
rect 222614 227628 222620 227640
rect 222488 227600 222620 227628
rect 222488 227588 222494 227600
rect 222614 227588 222620 227600
rect 222672 227588 222678 227640
rect 280298 227588 280304 227640
rect 280356 227628 280362 227640
rect 353070 227628 353076 227640
rect 280356 227600 353076 227628
rect 280356 227588 280362 227600
rect 353070 227588 353076 227600
rect 353128 227588 353134 227640
rect 186458 227520 186464 227572
rect 186516 227560 186522 227572
rect 369078 227560 369084 227572
rect 186516 227532 369084 227560
rect 186516 227520 186522 227532
rect 369078 227520 369084 227532
rect 369136 227520 369142 227572
rect 322986 226976 322992 227028
rect 323044 227016 323050 227028
rect 346998 227016 347004 227028
rect 323044 226988 347004 227016
rect 323044 226976 323050 226988
rect 346998 226976 347004 226988
rect 347056 226976 347062 227028
rect 76794 226908 76800 226960
rect 76852 226948 76858 226960
rect 368802 226948 368808 226960
rect 76852 226920 368808 226948
rect 76852 226908 76858 226920
rect 368802 226908 368808 226920
rect 368860 226908 368866 226960
rect 34566 226840 34572 226892
rect 34624 226880 34630 226892
rect 368710 226880 368716 226892
rect 34624 226852 368716 226880
rect 34624 226840 34630 226852
rect 368710 226840 368716 226852
rect 368768 226840 368774 226892
rect 240278 226228 240284 226280
rect 240336 226268 240342 226280
rect 353254 226268 353260 226280
rect 240336 226240 353260 226268
rect 240336 226228 240342 226240
rect 353254 226228 353260 226240
rect 353312 226228 353318 226280
rect 231354 226160 231360 226212
rect 231412 226200 231418 226212
rect 353162 226200 353168 226212
rect 231412 226172 353168 226200
rect 231412 226160 231418 226172
rect 353162 226160 353168 226172
rect 353220 226160 353226 226212
rect 137606 226092 137612 226144
rect 137664 226132 137670 226144
rect 353346 226132 353352 226144
rect 137664 226104 353352 226132
rect 137664 226092 137670 226104
rect 353346 226092 353352 226104
rect 353404 226092 353410 226144
rect 324550 225684 324556 225736
rect 324608 225724 324614 225736
rect 325378 225724 325384 225736
rect 324608 225696 325384 225724
rect 324608 225684 324614 225696
rect 325378 225684 325384 225696
rect 325436 225724 325442 225736
rect 345710 225724 345716 225736
rect 325436 225696 345716 225724
rect 325436 225684 325442 225696
rect 345710 225684 345716 225696
rect 345768 225684 345774 225736
rect 172014 225616 172020 225668
rect 172072 225656 172078 225668
rect 368802 225656 368808 225668
rect 172072 225628 368808 225656
rect 172072 225616 172078 225628
rect 368802 225616 368808 225628
rect 368860 225616 368866 225668
rect 137514 225548 137520 225600
rect 137572 225588 137578 225600
rect 368710 225588 368716 225600
rect 137572 225560 368716 225588
rect 137572 225548 137578 225560
rect 368710 225548 368716 225560
rect 368768 225548 368774 225600
rect 134754 225480 134760 225532
rect 134812 225520 134818 225532
rect 368894 225520 368900 225532
rect 134812 225492 368900 225520
rect 134812 225480 134818 225492
rect 368894 225480 368900 225492
rect 368952 225480 368958 225532
rect 251226 225412 251232 225464
rect 251284 225452 251290 225464
rect 253986 225452 253992 225464
rect 251284 225424 253992 225452
rect 251284 225412 251290 225424
rect 253986 225412 253992 225424
rect 254044 225412 254050 225464
rect 254998 225412 255004 225464
rect 255056 225452 255062 225464
rect 257482 225452 257488 225464
rect 255056 225424 257488 225452
rect 255056 225412 255062 225424
rect 257482 225412 257488 225424
rect 257540 225412 257546 225464
rect 338350 225412 338356 225464
rect 338408 225452 338414 225464
rect 338408 225424 341340 225452
rect 338408 225412 338414 225424
rect 62350 225344 62356 225396
rect 62408 225384 62414 225396
rect 63638 225384 63644 225396
rect 62408 225356 63644 225384
rect 62408 225344 62414 225356
rect 63638 225344 63644 225356
rect 63696 225344 63702 225396
rect 249202 225344 249208 225396
rect 249260 225384 249266 225396
rect 252146 225384 252152 225396
rect 249260 225356 252152 225384
rect 249260 225344 249266 225356
rect 252146 225344 252152 225356
rect 252204 225344 252210 225396
rect 252238 225344 252244 225396
rect 252296 225384 252302 225396
rect 254814 225384 254820 225396
rect 252296 225356 254820 225384
rect 252296 225344 252302 225356
rect 254814 225344 254820 225356
rect 254872 225344 254878 225396
rect 256010 225344 256016 225396
rect 256068 225384 256074 225396
rect 258402 225384 258408 225396
rect 256068 225356 258408 225384
rect 256068 225344 256074 225356
rect 258402 225344 258408 225356
rect 258460 225344 258466 225396
rect 337154 225344 337160 225396
rect 337212 225384 337218 225396
rect 338994 225384 339000 225396
rect 337212 225356 339000 225384
rect 337212 225344 337218 225356
rect 338994 225344 339000 225356
rect 339052 225344 339058 225396
rect 340190 225344 340196 225396
rect 340248 225384 340254 225396
rect 341018 225384 341024 225396
rect 340248 225356 341024 225384
rect 340248 225344 340254 225356
rect 341018 225344 341024 225356
rect 341076 225344 341082 225396
rect 341312 225384 341340 225424
rect 341386 225412 341392 225464
rect 341444 225452 341450 225464
rect 346630 225452 346636 225464
rect 341444 225424 346636 225452
rect 341444 225412 341450 225424
rect 346630 225412 346636 225424
rect 346688 225412 346694 225464
rect 341312 225356 341432 225384
rect 56094 225276 56100 225328
rect 56152 225316 56158 225328
rect 56738 225316 56744 225328
rect 56152 225288 56744 225316
rect 56152 225276 56158 225288
rect 56738 225276 56744 225288
rect 56796 225276 56802 225328
rect 59682 225276 59688 225328
rect 59740 225316 59746 225328
rect 60786 225316 60792 225328
rect 59740 225288 60792 225316
rect 59740 225276 59746 225288
rect 60786 225276 60792 225288
rect 60844 225276 60850 225328
rect 61430 225276 61436 225328
rect 61488 225316 61494 225328
rect 62258 225316 62264 225328
rect 61488 225288 62264 225316
rect 61488 225276 61494 225288
rect 62258 225276 62264 225288
rect 62316 225276 62322 225328
rect 63178 225276 63184 225328
rect 63236 225316 63242 225328
rect 64098 225316 64104 225328
rect 63236 225288 64104 225316
rect 63236 225276 63242 225288
rect 64098 225276 64104 225288
rect 64156 225276 64162 225328
rect 65754 225276 65760 225328
rect 65812 225316 65818 225328
rect 66766 225316 66772 225328
rect 65812 225288 66772 225316
rect 65812 225276 65818 225288
rect 66766 225276 66772 225288
rect 66824 225276 66830 225328
rect 68514 225276 68520 225328
rect 68572 225316 68578 225328
rect 70354 225316 70360 225328
rect 68572 225288 70360 225316
rect 68572 225276 68578 225288
rect 70354 225276 70360 225288
rect 70412 225276 70418 225328
rect 153706 225276 153712 225328
rect 153764 225316 153770 225328
rect 154718 225316 154724 225328
rect 153764 225288 154724 225316
rect 153764 225276 153770 225288
rect 154718 225276 154724 225288
rect 154776 225276 154782 225328
rect 155454 225276 155460 225328
rect 155512 225316 155518 225328
rect 156098 225316 156104 225328
rect 155512 225288 156104 225316
rect 155512 225276 155518 225288
rect 156098 225276 156104 225288
rect 156156 225276 156162 225328
rect 156374 225276 156380 225328
rect 156432 225316 156438 225328
rect 157478 225316 157484 225328
rect 156432 225288 157484 225316
rect 156432 225276 156438 225288
rect 157478 225276 157484 225288
rect 157536 225276 157542 225328
rect 228594 225276 228600 225328
rect 228652 225316 228658 225328
rect 341297 225319 341355 225325
rect 341297 225316 341309 225319
rect 228652 225288 341309 225316
rect 228652 225276 228658 225288
rect 341297 225285 341309 225288
rect 341343 225285 341355 225319
rect 341297 225279 341355 225285
rect 61614 225208 61620 225260
rect 61672 225248 61678 225260
rect 63270 225248 63276 225260
rect 61672 225220 63276 225248
rect 61672 225208 61678 225220
rect 63270 225208 63276 225220
rect 63328 225208 63334 225260
rect 65846 225208 65852 225260
rect 65904 225248 65910 225260
rect 67686 225248 67692 225260
rect 65904 225220 67692 225248
rect 65904 225208 65910 225220
rect 67686 225208 67692 225220
rect 67744 225208 67750 225260
rect 254078 225208 254084 225260
rect 254136 225248 254142 225260
rect 256654 225248 256660 225260
rect 254136 225220 256660 225248
rect 254136 225208 254142 225220
rect 256654 225208 256660 225220
rect 256712 225208 256718 225260
rect 339546 225208 339552 225260
rect 339604 225248 339610 225260
rect 341205 225251 341263 225257
rect 341205 225248 341217 225251
rect 339604 225220 341217 225248
rect 339604 225208 339610 225220
rect 341205 225217 341217 225220
rect 341251 225217 341263 225251
rect 341404 225248 341432 225356
rect 342030 225344 342036 225396
rect 342088 225384 342094 225396
rect 346722 225384 346728 225396
rect 342088 225356 346728 225384
rect 342088 225344 342094 225356
rect 346722 225344 346728 225356
rect 346780 225344 346786 225396
rect 341481 225319 341539 225325
rect 341481 225285 341493 225319
rect 341527 225316 341539 225319
rect 368710 225316 368716 225328
rect 341527 225288 368716 225316
rect 341527 225285 341539 225288
rect 341481 225279 341539 225285
rect 368710 225276 368716 225288
rect 368768 225276 368774 225328
rect 343502 225248 343508 225260
rect 341404 225220 343508 225248
rect 341205 225211 341263 225217
rect 343502 225208 343508 225220
rect 343560 225208 343566 225260
rect 345897 225251 345955 225257
rect 345897 225217 345909 225251
rect 345943 225248 345955 225251
rect 351598 225248 351604 225260
rect 345943 225220 351604 225248
rect 345943 225217 345955 225220
rect 345897 225211 345955 225217
rect 351598 225208 351604 225220
rect 351656 225208 351662 225260
rect 151038 225140 151044 225192
rect 151096 225180 151102 225192
rect 151866 225180 151872 225192
rect 151096 225152 151872 225180
rect 151096 225140 151102 225152
rect 151866 225140 151872 225152
rect 151924 225140 151930 225192
rect 162998 225140 163004 225192
rect 163056 225180 163062 225192
rect 164378 225180 164384 225192
rect 163056 225152 164384 225180
rect 163056 225140 163062 225152
rect 164378 225140 164384 225152
rect 164436 225140 164442 225192
rect 252606 225140 252612 225192
rect 252664 225180 252670 225192
rect 255734 225180 255740 225192
rect 252664 225152 255740 225180
rect 252664 225140 252670 225152
rect 255734 225140 255740 225152
rect 255792 225140 255798 225192
rect 338994 225140 339000 225192
rect 339052 225180 339058 225192
rect 342950 225180 342956 225192
rect 339052 225152 342956 225180
rect 339052 225140 339058 225152
rect 342950 225140 342956 225152
rect 343008 225140 343014 225192
rect 352242 225180 352248 225192
rect 348672 225152 352248 225180
rect 63086 225072 63092 225124
rect 63144 225112 63150 225124
rect 65938 225112 65944 225124
rect 63144 225084 65944 225112
rect 63144 225072 63150 225084
rect 65938 225072 65944 225084
rect 65996 225072 66002 225124
rect 335406 225072 335412 225124
rect 335464 225112 335470 225124
rect 348562 225112 348568 225124
rect 335464 225084 348568 225112
rect 335464 225072 335470 225084
rect 348562 225072 348568 225084
rect 348620 225072 348626 225124
rect 58762 225004 58768 225056
rect 58820 225044 58826 225056
rect 59498 225044 59504 225056
rect 58820 225016 59504 225044
rect 58820 225004 58826 225016
rect 59498 225004 59504 225016
rect 59556 225004 59562 225056
rect 337706 225004 337712 225056
rect 337764 225044 337770 225056
rect 342582 225044 342588 225056
rect 337764 225016 342588 225044
rect 337764 225004 337770 225016
rect 342582 225004 342588 225016
rect 342640 225004 342646 225056
rect 342674 225004 342680 225056
rect 342732 225044 342738 225056
rect 348672 225044 348700 225152
rect 352242 225140 352248 225152
rect 352300 225140 352306 225192
rect 342732 225016 348700 225044
rect 342732 225004 342738 225016
rect 62994 224936 63000 224988
rect 63052 224976 63058 224988
rect 65018 224976 65024 224988
rect 63052 224948 65024 224976
rect 63052 224936 63058 224948
rect 65018 224936 65024 224948
rect 65076 224936 65082 224988
rect 334118 224936 334124 224988
rect 334176 224976 334182 224988
rect 348010 224976 348016 224988
rect 334176 224948 348016 224976
rect 334176 224936 334182 224948
rect 348010 224936 348016 224948
rect 348068 224936 348074 224988
rect 335498 224868 335504 224920
rect 335556 224908 335562 224920
rect 349390 224908 349396 224920
rect 335556 224880 349396 224908
rect 335556 224868 335562 224880
rect 349390 224868 349396 224880
rect 349448 224868 349454 224920
rect 149290 224800 149296 224852
rect 149348 224840 149354 224852
rect 150578 224840 150584 224852
rect 149348 224812 150584 224840
rect 149348 224800 149354 224812
rect 150578 224800 150584 224812
rect 150636 224800 150642 224852
rect 332738 224800 332744 224852
rect 332796 224840 332802 224852
rect 335593 224843 335651 224849
rect 335593 224840 335605 224843
rect 332796 224812 335605 224840
rect 332796 224800 332802 224812
rect 335593 224809 335605 224812
rect 335639 224809 335651 224843
rect 335593 224803 335651 224809
rect 340834 224800 340840 224852
rect 340892 224840 340898 224852
rect 341294 224840 341300 224852
rect 340892 224812 341300 224840
rect 340892 224800 340898 224812
rect 341294 224800 341300 224812
rect 341352 224800 341358 224852
rect 57014 224732 57020 224784
rect 57072 224772 57078 224784
rect 67318 224772 67324 224784
rect 57072 224744 67324 224772
rect 57072 224732 57078 224744
rect 67318 224732 67324 224744
rect 67376 224732 67382 224784
rect 341205 224775 341263 224781
rect 341205 224741 341217 224775
rect 341251 224772 341263 224775
rect 342858 224772 342864 224784
rect 341251 224744 342864 224772
rect 341251 224741 341263 224744
rect 341205 224735 341263 224741
rect 342858 224732 342864 224744
rect 342916 224732 342922 224784
rect 343042 224732 343048 224784
rect 343100 224772 343106 224784
rect 360614 224772 360620 224784
rect 343100 224744 360620 224772
rect 343100 224732 343106 224744
rect 360614 224732 360620 224744
rect 360672 224732 360678 224784
rect 338258 224596 338264 224648
rect 338316 224636 338322 224648
rect 350678 224636 350684 224648
rect 338316 224608 350684 224636
rect 338316 224596 338322 224608
rect 350678 224596 350684 224608
rect 350736 224596 350742 224648
rect 67226 224528 67232 224580
rect 67284 224568 67290 224580
rect 69434 224568 69440 224580
rect 67284 224540 69440 224568
rect 67284 224528 67290 224540
rect 69434 224528 69440 224540
rect 69492 224528 69498 224580
rect 339638 224528 339644 224580
rect 339696 224568 339702 224580
rect 345897 224571 345955 224577
rect 345897 224568 345909 224571
rect 339696 224540 345909 224568
rect 339696 224528 339702 224540
rect 345897 224537 345909 224540
rect 345943 224537 345955 224571
rect 345897 224531 345955 224537
rect 336878 224460 336884 224512
rect 336936 224500 336942 224512
rect 349758 224500 349764 224512
rect 336936 224472 349764 224500
rect 336936 224460 336942 224472
rect 349758 224460 349764 224472
rect 349816 224460 349822 224512
rect 335593 224435 335651 224441
rect 335593 224401 335605 224435
rect 335639 224432 335651 224435
rect 347274 224432 347280 224444
rect 335639 224404 347280 224432
rect 335639 224401 335651 224404
rect 335593 224395 335651 224401
rect 347274 224392 347280 224404
rect 347332 224392 347338 224444
rect 160974 224324 160980 224376
rect 161032 224364 161038 224376
rect 161710 224364 161716 224376
rect 161032 224336 161716 224364
rect 161032 224324 161038 224336
rect 161710 224324 161716 224336
rect 161768 224324 161774 224376
rect 325654 224324 325660 224376
rect 325712 224364 325718 224376
rect 343042 224364 343048 224376
rect 325712 224336 343048 224364
rect 325712 224324 325718 224336
rect 343042 224324 343048 224336
rect 343100 224324 343106 224376
rect 343137 224367 343195 224373
rect 343137 224333 343149 224367
rect 343183 224364 343195 224367
rect 348013 224367 348071 224373
rect 348013 224364 348025 224367
rect 343183 224336 348025 224364
rect 343183 224333 343195 224336
rect 343137 224327 343195 224333
rect 348013 224333 348025 224336
rect 348059 224333 348071 224367
rect 348013 224327 348071 224333
rect 67134 224256 67140 224308
rect 67192 224296 67198 224308
rect 68606 224296 68612 224308
rect 67192 224268 68612 224296
rect 67192 224256 67198 224268
rect 68606 224256 68612 224268
rect 68664 224256 68670 224308
rect 325378 224256 325384 224308
rect 325436 224296 325442 224308
rect 325746 224296 325752 224308
rect 325436 224268 325752 224296
rect 325436 224256 325442 224268
rect 325746 224256 325752 224268
rect 325804 224296 325810 224308
rect 344238 224296 344244 224308
rect 325804 224268 344244 224296
rect 325804 224256 325810 224268
rect 344238 224256 344244 224268
rect 344296 224256 344302 224308
rect 158214 224188 158220 224240
rect 158272 224228 158278 224240
rect 159042 224228 159048 224240
rect 158272 224200 159048 224228
rect 158272 224188 158278 224200
rect 159042 224188 159048 224200
rect 159100 224188 159106 224240
rect 325194 224188 325200 224240
rect 325252 224228 325258 224240
rect 325838 224228 325844 224240
rect 325252 224200 325844 224228
rect 325252 224188 325258 224200
rect 325838 224188 325844 224200
rect 325896 224228 325902 224240
rect 345158 224228 345164 224240
rect 325896 224200 345164 224228
rect 325896 224188 325902 224200
rect 345158 224188 345164 224200
rect 345216 224188 345222 224240
rect 243590 224120 243596 224172
rect 243648 224160 243654 224172
rect 244418 224160 244424 224172
rect 243648 224132 244424 224160
rect 243648 224120 243654 224132
rect 244418 224120 244424 224132
rect 244476 224120 244482 224172
rect 322618 224120 322624 224172
rect 322676 224160 322682 224172
rect 368802 224160 368808 224172
rect 322676 224132 368808 224160
rect 322676 224120 322682 224132
rect 368802 224120 368808 224132
rect 368860 224120 368866 224172
rect 369078 223712 369084 223764
rect 369136 223752 369142 223764
rect 369354 223752 369360 223764
rect 369136 223724 369360 223752
rect 369136 223712 369142 223724
rect 369354 223712 369360 223724
rect 369412 223712 369418 223764
rect 348013 223075 348071 223081
rect 348013 223041 348025 223075
rect 348059 223072 348071 223075
rect 351276 223072 351282 223084
rect 348059 223044 351282 223072
rect 348059 223041 348071 223044
rect 348013 223035 348071 223041
rect 351276 223032 351282 223044
rect 351334 223032 351340 223084
rect 363834 222896 363840 222948
rect 363892 222936 363898 222948
rect 368894 222936 368900 222948
rect 363892 222908 368900 222936
rect 363892 222896 363898 222908
rect 368894 222896 368900 222908
rect 368952 222896 368958 222948
rect 323814 222828 323820 222880
rect 323872 222868 323878 222880
rect 368710 222868 368716 222880
rect 323872 222840 368716 222868
rect 323872 222828 323878 222840
rect 368710 222828 368716 222840
rect 368768 222828 368774 222880
rect 322710 222760 322716 222812
rect 322768 222800 322774 222812
rect 368802 222800 368808 222812
rect 322768 222772 368808 222800
rect 322768 222760 322774 222772
rect 368802 222760 368808 222772
rect 368860 222760 368866 222812
rect 250122 222692 250128 222744
rect 250180 222732 250186 222744
rect 250950 222732 250956 222744
rect 250180 222704 250956 222732
rect 250180 222692 250186 222704
rect 250950 222692 250956 222704
rect 251008 222692 251014 222744
rect 34566 221740 34572 221792
rect 34624 221780 34630 221792
rect 34934 221780 34940 221792
rect 34624 221752 34940 221780
rect 34624 221740 34630 221752
rect 34934 221740 34940 221752
rect 34992 221740 34998 221792
rect 34014 221672 34020 221724
rect 34072 221712 34078 221724
rect 34750 221712 34756 221724
rect 34072 221684 34756 221712
rect 34072 221672 34078 221684
rect 34750 221672 34756 221684
rect 34808 221672 34814 221724
rect 361074 221468 361080 221520
rect 361132 221508 361138 221520
rect 368894 221508 368900 221520
rect 361132 221480 368900 221508
rect 361132 221468 361138 221480
rect 368894 221468 368900 221480
rect 368952 221468 368958 221520
rect 325194 221400 325200 221452
rect 325252 221440 325258 221452
rect 368802 221440 368808 221452
rect 325252 221412 368808 221440
rect 325252 221400 325258 221412
rect 368802 221400 368808 221412
rect 368860 221400 368866 221452
rect 322894 221332 322900 221384
rect 322952 221372 322958 221384
rect 368710 221372 368716 221384
rect 322952 221344 368716 221372
rect 322952 221332 322958 221344
rect 368710 221332 368716 221344
rect 368768 221332 368774 221384
rect 325286 220584 325292 220636
rect 325344 220624 325350 220636
rect 353438 220624 353444 220636
rect 325344 220596 353444 220624
rect 325344 220584 325350 220596
rect 353438 220584 353444 220596
rect 353496 220584 353502 220636
rect 34658 220516 34664 220568
rect 34716 220556 34722 220568
rect 34934 220556 34940 220568
rect 34716 220528 34940 220556
rect 34716 220516 34722 220528
rect 34934 220516 34940 220528
rect 34992 220516 34998 220568
rect 325378 220516 325384 220568
rect 325436 220556 325442 220568
rect 368802 220556 368808 220568
rect 325436 220528 368808 220556
rect 325436 220516 325442 220528
rect 368802 220516 368808 220528
rect 368860 220516 368866 220568
rect 34750 220448 34756 220500
rect 34808 220488 34814 220500
rect 34845 220491 34903 220497
rect 34845 220488 34857 220491
rect 34808 220460 34857 220488
rect 34808 220448 34814 220460
rect 34845 220457 34857 220460
rect 34891 220457 34903 220491
rect 34845 220451 34903 220457
rect 322802 220448 322808 220500
rect 322860 220488 322866 220500
rect 368710 220488 368716 220500
rect 322860 220460 368716 220488
rect 322860 220448 322866 220460
rect 368710 220448 368716 220460
rect 368768 220448 368774 220500
rect 51862 220012 51868 220024
rect 47832 219984 51868 220012
rect 38062 219904 38068 219956
rect 38120 219944 38126 219956
rect 47832 219944 47860 219984
rect 51862 219972 51868 219984
rect 51920 219972 51926 220024
rect 359694 219972 359700 220024
rect 359752 220012 359758 220024
rect 368894 220012 368900 220024
rect 359752 219984 368900 220012
rect 359752 219972 359758 219984
rect 368894 219972 368900 219984
rect 368952 219972 368958 220024
rect 38120 219916 47860 219944
rect 38120 219904 38126 219916
rect 76150 219496 76156 219548
rect 76208 219536 76214 219548
rect 81670 219536 81676 219548
rect 76208 219508 81676 219536
rect 76208 219496 76214 219508
rect 81670 219496 81676 219508
rect 81728 219496 81734 219548
rect 369078 219468 369084 219480
rect 369039 219440 369084 219468
rect 369078 219428 369084 219440
rect 369136 219428 369142 219480
rect 13038 219360 13044 219412
rect 13096 219400 13102 219412
rect 16350 219400 16356 219412
rect 13096 219372 16356 219400
rect 13096 219360 13102 219372
rect 16350 219360 16356 219372
rect 16408 219360 16414 219412
rect 368894 219360 368900 219412
rect 368952 219400 368958 219412
rect 369262 219400 369268 219412
rect 368952 219372 369268 219400
rect 368952 219360 368958 219372
rect 369262 219360 369268 219372
rect 369320 219360 369326 219412
rect 369354 219360 369360 219412
rect 369412 219400 369418 219412
rect 369412 219372 369457 219400
rect 369412 219360 369418 219372
rect 165114 219224 165120 219276
rect 165172 219264 165178 219276
rect 179282 219264 179288 219276
rect 165172 219236 179288 219264
rect 165172 219224 165178 219236
rect 179282 219224 179288 219236
rect 179340 219224 179346 219276
rect 258954 219224 258960 219276
rect 259012 219264 259018 219276
rect 272938 219264 272944 219276
rect 259012 219236 272944 219264
rect 259012 219224 259018 219236
rect 272938 219224 272944 219236
rect 272996 219224 273002 219276
rect 368986 218952 368992 219004
rect 369044 218992 369050 219004
rect 369170 218992 369176 219004
rect 369044 218964 369176 218992
rect 369044 218952 369050 218964
rect 369170 218952 369176 218964
rect 369228 218952 369234 219004
rect 365214 218680 365220 218732
rect 365272 218720 365278 218732
rect 368802 218720 368808 218732
rect 365272 218692 368808 218720
rect 365272 218680 365278 218692
rect 368802 218680 368808 218692
rect 368860 218680 368866 218732
rect 352794 218612 352800 218664
rect 352852 218652 352858 218664
rect 368710 218652 368716 218664
rect 352852 218624 368716 218652
rect 352852 218612 352858 218624
rect 368710 218612 368716 218624
rect 368768 218612 368774 218664
rect 394838 218612 394844 218664
rect 394896 218652 394902 218664
rect 405970 218652 405976 218664
rect 394896 218624 405976 218652
rect 394896 218612 394902 218624
rect 405970 218612 405976 218624
rect 406028 218612 406034 218664
rect 352886 218476 352892 218528
rect 352944 218516 352950 218528
rect 368802 218516 368808 218528
rect 352944 218488 368808 218516
rect 352944 218476 352950 218488
rect 368802 218476 368808 218488
rect 368860 218476 368866 218528
rect 352978 217184 352984 217236
rect 353036 217224 353042 217236
rect 368710 217224 368716 217236
rect 353036 217196 368716 217224
rect 353036 217184 353042 217196
rect 368710 217184 368716 217196
rect 368768 217184 368774 217236
rect 38522 217116 38528 217168
rect 38580 217156 38586 217168
rect 53242 217156 53248 217168
rect 38580 217128 53248 217156
rect 38580 217116 38586 217128
rect 53242 217116 53248 217128
rect 53300 217116 53306 217168
rect 353346 217116 353352 217168
rect 353404 217156 353410 217168
rect 368802 217156 368808 217168
rect 353404 217128 368808 217156
rect 353404 217116 353410 217128
rect 368802 217116 368808 217128
rect 368860 217116 368866 217168
rect 358406 217048 358412 217100
rect 358464 217088 358470 217100
rect 368710 217088 368716 217100
rect 358464 217060 368716 217088
rect 358464 217048 358470 217060
rect 368710 217048 368716 217060
rect 368768 217048 368774 217100
rect 369078 216884 369084 216896
rect 369039 216856 369084 216884
rect 369078 216844 369084 216856
rect 369136 216844 369142 216896
rect 369078 216708 369084 216760
rect 369136 216748 369142 216760
rect 369357 216751 369415 216757
rect 369357 216748 369369 216751
rect 369136 216720 369369 216748
rect 369136 216708 369142 216720
rect 369357 216717 369369 216720
rect 369403 216717 369415 216751
rect 369357 216711 369415 216717
rect 137606 215824 137612 215876
rect 137664 215864 137670 215876
rect 145150 215864 145156 215876
rect 137664 215836 145156 215864
rect 137664 215824 137670 215836
rect 145150 215824 145156 215836
rect 145208 215824 145214 215876
rect 231354 215824 231360 215876
rect 231412 215864 231418 215876
rect 240922 215864 240928 215876
rect 231412 215836 240928 215864
rect 231412 215824 231418 215836
rect 240922 215824 240928 215836
rect 240980 215824 240986 215876
rect 325286 215824 325292 215876
rect 325344 215864 325350 215876
rect 334210 215864 334216 215876
rect 325344 215836 334216 215864
rect 325344 215824 325350 215836
rect 334210 215824 334216 215836
rect 334268 215824 334274 215876
rect 353162 215756 353168 215808
rect 353220 215796 353226 215808
rect 368986 215796 368992 215808
rect 353220 215768 368992 215796
rect 353220 215756 353226 215768
rect 368986 215756 368992 215768
rect 369044 215756 369050 215808
rect 353254 215688 353260 215740
rect 353312 215728 353318 215740
rect 368710 215728 368716 215740
rect 353312 215700 368716 215728
rect 353312 215688 353318 215700
rect 368710 215688 368716 215700
rect 368768 215688 368774 215740
rect 358314 215620 358320 215672
rect 358372 215660 358378 215672
rect 368802 215660 368808 215672
rect 358372 215632 368808 215660
rect 358372 215620 358378 215632
rect 368802 215620 368808 215632
rect 368860 215620 368866 215672
rect 368989 214575 369047 214581
rect 368989 214541 369001 214575
rect 369035 214572 369047 214575
rect 369814 214572 369820 214584
rect 369035 214544 369820 214572
rect 369035 214541 369047 214544
rect 368989 214535 369047 214541
rect 369814 214532 369820 214544
rect 369872 214532 369878 214584
rect 51678 214504 51684 214516
rect 48476 214476 51684 214504
rect 38522 214396 38528 214448
rect 38580 214436 38586 214448
rect 48476 214436 48504 214476
rect 51678 214464 51684 214476
rect 51736 214464 51742 214516
rect 74218 214464 74224 214516
rect 74276 214504 74282 214516
rect 74402 214504 74408 214516
rect 74276 214476 74408 214504
rect 74276 214464 74282 214476
rect 74402 214464 74408 214476
rect 74460 214464 74466 214516
rect 38580 214408 48504 214436
rect 38580 214396 38586 214408
rect 353070 214396 353076 214448
rect 353128 214436 353134 214448
rect 368710 214436 368716 214448
rect 353128 214408 368716 214436
rect 353128 214396 353134 214408
rect 368710 214396 368716 214408
rect 368768 214396 368774 214448
rect 368986 214436 368992 214448
rect 368947 214408 368992 214436
rect 368986 214396 368992 214408
rect 369044 214396 369050 214448
rect 361166 214260 361172 214312
rect 361224 214300 361230 214312
rect 368894 214300 368900 214312
rect 361224 214272 368900 214300
rect 361224 214260 361230 214272
rect 368894 214260 368900 214272
rect 368952 214260 368958 214312
rect 356198 214056 356204 214108
rect 356256 214096 356262 214108
rect 405970 214096 405976 214108
rect 356256 214068 405976 214096
rect 356256 214056 356262 214068
rect 405970 214056 405976 214068
rect 406028 214056 406034 214108
rect 355094 213988 355100 214040
rect 355152 214028 355158 214040
rect 394838 214028 394844 214040
rect 355152 214000 394844 214028
rect 355152 213988 355158 214000
rect 394838 213988 394844 214000
rect 394896 213988 394902 214040
rect 365306 213920 365312 213972
rect 365364 213960 365370 213972
rect 368894 213960 368900 213972
rect 365364 213932 368900 213960
rect 365364 213920 365370 213932
rect 368894 213920 368900 213932
rect 368952 213920 368958 213972
rect 34842 213892 34848 213904
rect 34803 213864 34848 213892
rect 34842 213852 34848 213864
rect 34900 213852 34906 213904
rect 353438 213036 353444 213088
rect 353496 213076 353502 213088
rect 368710 213076 368716 213088
rect 353496 213048 368716 213076
rect 353496 213036 353502 213048
rect 368710 213036 368716 213048
rect 368768 213036 368774 213088
rect 262358 211744 262364 211796
rect 262416 211784 262422 211796
rect 268614 211784 268620 211796
rect 262416 211756 268620 211784
rect 262416 211744 262422 211756
rect 268614 211744 268620 211756
rect 268672 211744 268678 211796
rect 167966 211676 167972 211728
rect 168024 211716 168030 211728
rect 174774 211716 174780 211728
rect 168024 211688 174780 211716
rect 168024 211676 168030 211688
rect 174774 211676 174780 211688
rect 174832 211676 174838 211728
rect 369906 211608 369912 211660
rect 369964 211648 369970 211660
rect 370734 211648 370740 211660
rect 369964 211620 370740 211648
rect 369964 211608 369970 211620
rect 370734 211608 370740 211620
rect 370792 211608 370798 211660
rect 38706 210928 38712 210980
rect 38764 210968 38770 210980
rect 54070 210968 54076 210980
rect 38764 210940 54076 210968
rect 38764 210928 38770 210940
rect 54070 210928 54076 210940
rect 54128 210928 54134 210980
rect 354910 210928 354916 210980
rect 354968 210968 354974 210980
rect 405970 210968 405976 210980
rect 354968 210940 405976 210968
rect 354968 210928 354974 210940
rect 405970 210928 405976 210940
rect 406028 210928 406034 210980
rect 378278 210316 378284 210368
rect 378336 210356 378342 210368
rect 383890 210356 383896 210368
rect 378336 210328 383896 210356
rect 378336 210316 378342 210328
rect 383890 210316 383896 210328
rect 383948 210316 383954 210368
rect 369170 209840 369176 209892
rect 369228 209880 369234 209892
rect 369814 209880 369820 209892
rect 369228 209852 369820 209880
rect 369228 209840 369234 209852
rect 369814 209840 369820 209852
rect 369872 209840 369878 209892
rect 174774 209636 174780 209688
rect 174832 209676 174838 209688
rect 178914 209676 178920 209688
rect 174832 209648 178920 209676
rect 174832 209636 174838 209648
rect 178914 209636 178920 209648
rect 178972 209636 178978 209688
rect 38522 209568 38528 209620
rect 38580 209608 38586 209620
rect 51402 209608 51408 209620
rect 38580 209580 51408 209608
rect 38580 209568 38586 209580
rect 51402 209568 51408 209580
rect 51460 209568 51466 209620
rect 356014 209568 356020 209620
rect 356072 209608 356078 209620
rect 405970 209608 405976 209620
rect 356072 209580 405976 209608
rect 356072 209568 356078 209580
rect 405970 209568 405976 209580
rect 406028 209568 406034 209620
rect 368986 209500 368992 209552
rect 369044 209540 369050 209552
rect 369262 209540 369268 209552
rect 369044 209512 369268 209540
rect 369044 209500 369050 209512
rect 369262 209500 369268 209512
rect 369320 209500 369326 209552
rect 427314 208820 427320 208872
rect 427372 208860 427378 208872
rect 429614 208860 429620 208872
rect 427372 208832 429620 208860
rect 427372 208820 427378 208832
rect 429614 208820 429620 208832
rect 429672 208820 429678 208872
rect 13038 208140 13044 208192
rect 13096 208180 13102 208192
rect 16442 208180 16448 208192
rect 13096 208152 16448 208180
rect 13096 208140 13102 208152
rect 16442 208140 16448 208152
rect 16500 208140 16506 208192
rect 268614 207460 268620 207512
rect 268672 207500 268678 207512
rect 272938 207500 272944 207512
rect 268672 207472 272944 207500
rect 268672 207460 268678 207472
rect 272938 207460 272944 207472
rect 272996 207460 273002 207512
rect 34842 206888 34848 206900
rect 34803 206860 34848 206888
rect 34842 206848 34848 206860
rect 34900 206848 34906 206900
rect 38522 206780 38528 206832
rect 38580 206820 38586 206832
rect 51402 206820 51408 206832
rect 38580 206792 51408 206820
rect 38580 206780 38586 206792
rect 51402 206780 51408 206792
rect 51460 206780 51466 206832
rect 355002 206780 355008 206832
rect 355060 206820 355066 206832
rect 405970 206820 405976 206832
rect 355060 206792 405976 206820
rect 355060 206780 355066 206792
rect 405970 206780 405976 206792
rect 406028 206780 406034 206832
rect 38522 204740 38528 204792
rect 38580 204780 38586 204792
rect 51402 204780 51408 204792
rect 38580 204752 51408 204780
rect 38580 204740 38586 204752
rect 51402 204740 51408 204752
rect 51460 204740 51466 204792
rect 136870 204740 136876 204792
rect 136928 204780 136934 204792
rect 145334 204780 145340 204792
rect 136928 204752 145340 204780
rect 136928 204740 136934 204752
rect 145334 204740 145340 204752
rect 145392 204740 145398 204792
rect 231998 204740 232004 204792
rect 232056 204780 232062 204792
rect 239634 204780 239640 204792
rect 232056 204752 239640 204780
rect 232056 204740 232062 204752
rect 239634 204740 239640 204752
rect 239692 204740 239698 204792
rect 356198 204740 356204 204792
rect 356256 204780 356262 204792
rect 406062 204780 406068 204792
rect 356256 204752 406068 204780
rect 356256 204740 356262 204752
rect 406062 204740 406068 204752
rect 406120 204740 406126 204792
rect 34842 204712 34848 204724
rect 34803 204684 34848 204712
rect 34842 204672 34848 204684
rect 34900 204672 34906 204724
rect 368986 204672 368992 204724
rect 369044 204712 369050 204724
rect 369170 204712 369176 204724
rect 369044 204684 369176 204712
rect 369044 204672 369050 204684
rect 369170 204672 369176 204684
rect 369228 204672 369234 204724
rect 74310 203312 74316 203364
rect 74368 203352 74374 203364
rect 81670 203352 81676 203364
rect 74368 203324 81676 203352
rect 74368 203312 74374 203324
rect 81670 203312 81676 203324
rect 81728 203312 81734 203364
rect 137790 202020 137796 202072
rect 137848 202060 137854 202072
rect 145426 202060 145432 202072
rect 137848 202032 145432 202060
rect 137848 202020 137854 202032
rect 145426 202020 145432 202032
rect 145484 202020 145490 202072
rect 231446 202020 231452 202072
rect 231504 202060 231510 202072
rect 240646 202060 240652 202072
rect 231504 202032 240652 202060
rect 231504 202020 231510 202032
rect 240646 202020 240652 202032
rect 240704 202020 240710 202072
rect 325470 202020 325476 202072
rect 325528 202060 325534 202072
rect 334210 202060 334216 202072
rect 325528 202032 334216 202060
rect 325528 202020 325534 202032
rect 334210 202020 334216 202032
rect 334268 202020 334274 202072
rect 38522 201272 38528 201324
rect 38580 201312 38586 201324
rect 51494 201312 51500 201324
rect 38580 201284 51500 201312
rect 38580 201272 38586 201284
rect 51494 201272 51500 201284
rect 51552 201272 51558 201324
rect 353530 201272 353536 201324
rect 353588 201312 353594 201324
rect 405970 201312 405976 201324
rect 353588 201284 405976 201312
rect 353588 201272 353594 201284
rect 405970 201272 405976 201284
rect 406028 201272 406034 201324
rect 368894 199912 368900 199964
rect 368952 199952 368958 199964
rect 369170 199952 369176 199964
rect 368952 199924 369176 199952
rect 368952 199912 368958 199924
rect 369170 199912 369176 199924
rect 369228 199912 369234 199964
rect 427130 199708 427136 199760
rect 427188 199748 427194 199760
rect 428786 199748 428792 199760
rect 427188 199720 428792 199748
rect 427188 199708 427194 199720
rect 428786 199708 428792 199720
rect 428844 199708 428850 199760
rect 369814 199476 369820 199488
rect 369775 199448 369820 199476
rect 369814 199436 369820 199448
rect 369872 199436 369878 199488
rect 13314 199300 13320 199352
rect 13372 199340 13378 199352
rect 17638 199340 17644 199352
rect 13372 199312 17644 199340
rect 13372 199300 13378 199312
rect 17638 199300 17644 199312
rect 17696 199300 17702 199352
rect 38522 199232 38528 199284
rect 38580 199272 38586 199284
rect 51770 199272 51776 199284
rect 38580 199244 51776 199272
rect 38580 199232 38586 199244
rect 51770 199232 51776 199244
rect 51828 199232 51834 199284
rect 355922 199232 355928 199284
rect 355980 199272 355986 199284
rect 405970 199272 405976 199284
rect 355980 199244 405976 199272
rect 355980 199232 355986 199244
rect 405970 199232 405976 199244
rect 406028 199232 406034 199284
rect 13038 197736 13044 197788
rect 13096 197776 13102 197788
rect 16258 197776 16264 197788
rect 13096 197748 16264 197776
rect 13096 197736 13102 197748
rect 16258 197736 16264 197748
rect 16316 197736 16322 197788
rect 427682 196512 427688 196564
rect 427740 196552 427746 196564
rect 429522 196552 429528 196564
rect 427740 196524 429528 196552
rect 427740 196512 427746 196524
rect 429522 196512 429528 196524
rect 429580 196512 429586 196564
rect 38522 195764 38528 195816
rect 38580 195804 38586 195816
rect 51310 195804 51316 195816
rect 38580 195776 51316 195804
rect 38580 195764 38586 195776
rect 51310 195764 51316 195776
rect 51368 195764 51374 195816
rect 352702 195764 352708 195816
rect 352760 195804 352766 195816
rect 405970 195804 405976 195816
rect 352760 195776 405976 195804
rect 352760 195764 352766 195776
rect 405970 195764 405976 195776
rect 406028 195764 406034 195816
rect 369906 195260 369912 195272
rect 369740 195232 369912 195260
rect 369740 195204 369768 195232
rect 369906 195220 369912 195232
rect 369964 195220 369970 195272
rect 368986 195152 368992 195204
rect 369044 195192 369050 195204
rect 369354 195192 369360 195204
rect 369044 195164 369360 195192
rect 369044 195152 369050 195164
rect 369354 195152 369360 195164
rect 369412 195152 369418 195204
rect 369722 195152 369728 195204
rect 369780 195152 369786 195204
rect 38798 195084 38804 195136
rect 38856 195124 38862 195136
rect 51310 195124 51316 195136
rect 38856 195096 51316 195124
rect 38856 195084 38862 195096
rect 51310 195084 51316 195096
rect 51368 195084 51374 195136
rect 356198 195084 356204 195136
rect 356256 195124 356262 195136
rect 406062 195124 406068 195136
rect 356256 195096 406068 195124
rect 356256 195084 356262 195096
rect 406062 195084 406068 195096
rect 406120 195084 406126 195136
rect 230802 194472 230808 194524
rect 230860 194512 230866 194524
rect 235310 194512 235316 194524
rect 230860 194484 235316 194512
rect 230860 194472 230866 194484
rect 235310 194472 235316 194484
rect 235368 194472 235374 194524
rect 369817 192407 369875 192413
rect 369817 192373 369829 192407
rect 369863 192404 369875 192407
rect 369906 192404 369912 192416
rect 369863 192376 369912 192404
rect 369863 192373 369875 192376
rect 369817 192367 369875 192373
rect 369906 192364 369912 192376
rect 369964 192364 369970 192416
rect 369817 192271 369875 192277
rect 369817 192237 369829 192271
rect 369863 192268 369875 192271
rect 369906 192268 369912 192280
rect 369863 192240 369912 192268
rect 369863 192237 369875 192240
rect 369817 192231 369875 192237
rect 369906 192228 369912 192240
rect 369964 192228 369970 192280
rect 38798 191616 38804 191668
rect 38856 191656 38862 191668
rect 49930 191656 49936 191668
rect 38856 191628 49936 191656
rect 38856 191616 38862 191628
rect 49930 191616 49936 191628
rect 49988 191616 49994 191668
rect 352886 191616 352892 191668
rect 352944 191656 352950 191668
rect 405970 191656 405976 191668
rect 352944 191628 405976 191656
rect 352944 191616 352950 191628
rect 405970 191616 405976 191628
rect 406028 191616 406034 191668
rect 426854 189848 426860 189900
rect 426912 189888 426918 189900
rect 429338 189888 429344 189900
rect 426912 189860 429344 189888
rect 426912 189848 426918 189860
rect 429338 189848 429344 189860
rect 429396 189848 429402 189900
rect 13406 189644 13412 189696
rect 13464 189684 13470 189696
rect 17086 189684 17092 189696
rect 13464 189656 17092 189684
rect 13464 189644 13470 189656
rect 17086 189644 17092 189656
rect 17144 189644 17150 189696
rect 38062 189576 38068 189628
rect 38120 189616 38126 189628
rect 51770 189616 51776 189628
rect 38120 189588 51776 189616
rect 38120 189576 38126 189588
rect 51770 189576 51776 189588
rect 51828 189576 51834 189628
rect 355186 189576 355192 189628
rect 355244 189616 355250 189628
rect 405970 189616 405976 189628
rect 355244 189588 405976 189616
rect 355244 189576 355250 189588
rect 405970 189576 405976 189588
rect 406028 189576 406034 189628
rect 324550 188896 324556 188948
rect 324608 188936 324614 188948
rect 330070 188936 330076 188948
rect 324608 188908 330076 188936
rect 324608 188896 324614 188908
rect 330070 188896 330076 188908
rect 330128 188896 330134 188948
rect 231998 188760 232004 188812
rect 232056 188800 232062 188812
rect 236230 188800 236236 188812
rect 232056 188772 236236 188800
rect 232056 188760 232062 188772
rect 236230 188760 236236 188772
rect 236288 188760 236294 188812
rect 137790 188284 137796 188336
rect 137848 188324 137854 188336
rect 142390 188324 142396 188336
rect 137848 188296 142396 188324
rect 137848 188284 137854 188296
rect 142390 188284 142396 188296
rect 142448 188324 142454 188336
rect 143034 188324 143040 188336
rect 142448 188296 143040 188324
rect 142448 188284 142454 188296
rect 143034 188284 143040 188296
rect 143092 188284 143098 188336
rect 236230 188284 236236 188336
rect 236288 188324 236294 188336
rect 236874 188324 236880 188336
rect 236288 188296 236880 188324
rect 236288 188284 236294 188296
rect 236874 188284 236880 188296
rect 236932 188284 236938 188336
rect 138894 188216 138900 188268
rect 138952 188256 138958 188268
rect 145610 188256 145616 188268
rect 138952 188228 145616 188256
rect 138952 188216 138958 188228
rect 145610 188216 145616 188228
rect 145668 188216 145674 188268
rect 232734 188216 232740 188268
rect 232792 188256 232798 188268
rect 240922 188256 240928 188268
rect 232792 188228 240928 188256
rect 232792 188216 232798 188228
rect 240922 188216 240928 188228
rect 240980 188216 240986 188268
rect 326574 188216 326580 188268
rect 326632 188256 326638 188268
rect 334210 188256 334216 188268
rect 326632 188228 334216 188256
rect 326632 188216 326638 188228
rect 334210 188216 334216 188228
rect 334268 188216 334274 188268
rect 75414 186788 75420 186840
rect 75472 186828 75478 186840
rect 81670 186828 81676 186840
rect 75472 186800 81676 186828
rect 75472 186788 75478 186800
rect 81670 186788 81676 186800
rect 81728 186788 81734 186840
rect 169254 186788 169260 186840
rect 169312 186828 169318 186840
rect 178914 186828 178920 186840
rect 169312 186800 178920 186828
rect 169312 186788 169318 186800
rect 178914 186788 178920 186800
rect 178972 186788 178978 186840
rect 263094 186788 263100 186840
rect 263152 186828 263158 186840
rect 272938 186828 272944 186840
rect 263152 186800 272944 186828
rect 263152 186788 263158 186800
rect 272938 186788 272944 186800
rect 272996 186788 273002 186840
rect 13038 186652 13044 186704
rect 13096 186692 13102 186704
rect 16074 186692 16080 186704
rect 13096 186664 16080 186692
rect 13096 186652 13102 186664
rect 16074 186652 16080 186664
rect 16132 186652 16138 186704
rect 38062 186108 38068 186160
rect 38120 186148 38126 186160
rect 48550 186148 48556 186160
rect 38120 186120 48556 186148
rect 38120 186108 38126 186120
rect 48550 186108 48556 186120
rect 48608 186108 48614 186160
rect 352794 186108 352800 186160
rect 352852 186148 352858 186160
rect 405970 186148 405976 186160
rect 352852 186120 405976 186148
rect 352852 186108 352858 186120
rect 405970 186108 405976 186120
rect 406028 186108 406034 186160
rect 369078 185428 369084 185480
rect 369136 185468 369142 185480
rect 369722 185468 369728 185480
rect 369136 185440 369728 185468
rect 369136 185428 369142 185440
rect 369722 185428 369728 185440
rect 369780 185428 369786 185480
rect 38798 184000 38804 184052
rect 38856 184040 38862 184052
rect 51402 184040 51408 184052
rect 38856 184012 51408 184040
rect 38856 184000 38862 184012
rect 51402 184000 51408 184012
rect 51460 184000 51466 184052
rect 356198 184000 356204 184052
rect 356256 184040 356262 184052
rect 405970 184040 405976 184052
rect 356256 184012 405976 184040
rect 356256 184000 356262 184012
rect 405970 184000 405976 184012
rect 406028 184000 406034 184052
rect 34382 183184 34388 183236
rect 34440 183224 34446 183236
rect 34934 183224 34940 183236
rect 34440 183196 34940 183224
rect 34440 183184 34446 183196
rect 34934 183184 34940 183196
rect 34992 183184 34998 183236
rect 369814 182748 369820 182760
rect 369775 182720 369820 182748
rect 369814 182708 369820 182720
rect 369872 182708 369878 182760
rect 34566 182640 34572 182692
rect 34624 182680 34630 182692
rect 34750 182680 34756 182692
rect 34624 182652 34756 182680
rect 34624 182640 34630 182652
rect 34750 182640 34756 182652
rect 34808 182640 34814 182692
rect 261070 182028 261076 182080
rect 261128 182068 261134 182080
rect 267510 182068 267516 182080
rect 261128 182040 267516 182068
rect 261128 182028 261134 182040
rect 267510 182028 267516 182040
rect 267568 182028 267574 182080
rect 21594 181280 21600 181332
rect 21652 181320 21658 181332
rect 34382 181320 34388 181332
rect 21652 181292 34388 181320
rect 21652 181280 21658 181292
rect 34382 181280 34388 181292
rect 34440 181280 34446 181332
rect 59682 181280 59688 181332
rect 59740 181320 59746 181332
rect 60878 181320 60884 181332
rect 59740 181292 60884 181320
rect 59740 181280 59746 181292
rect 60878 181280 60884 181292
rect 60936 181280 60942 181332
rect 61430 181280 61436 181332
rect 61488 181320 61494 181332
rect 62166 181320 62172 181332
rect 61488 181292 62172 181320
rect 61488 181280 61494 181292
rect 62166 181280 62172 181292
rect 62224 181280 62230 181332
rect 245338 181280 245344 181332
rect 245396 181320 245402 181332
rect 245798 181320 245804 181332
rect 245396 181292 245804 181320
rect 245396 181280 245402 181292
rect 245798 181280 245804 181292
rect 245856 181280 245862 181332
rect 247730 181280 247736 181332
rect 247788 181320 247794 181332
rect 248374 181320 248380 181332
rect 247788 181292 248380 181320
rect 247788 181280 247794 181292
rect 248374 181280 248380 181292
rect 248432 181280 248438 181332
rect 337614 181280 337620 181332
rect 337672 181320 337678 181332
rect 341110 181320 341116 181332
rect 337672 181292 341116 181320
rect 337672 181280 337678 181292
rect 341110 181280 341116 181292
rect 341168 181280 341174 181332
rect 344974 181280 344980 181332
rect 345032 181320 345038 181332
rect 359694 181320 359700 181332
rect 345032 181292 359700 181320
rect 345032 181280 345038 181292
rect 359694 181280 359700 181292
rect 359752 181280 359758 181332
rect 370734 181280 370740 181332
rect 370792 181320 370798 181332
rect 410202 181320 410208 181332
rect 370792 181292 410208 181320
rect 370792 181280 370798 181292
rect 410202 181280 410208 181292
rect 410260 181280 410266 181332
rect 60786 181212 60792 181264
rect 60844 181252 60850 181264
rect 65018 181252 65024 181264
rect 60844 181224 65024 181252
rect 60844 181212 60850 181224
rect 65018 181212 65024 181224
rect 65076 181212 65082 181264
rect 338258 181212 338264 181264
rect 338316 181252 338322 181264
rect 341754 181252 341760 181264
rect 338316 181224 341760 181252
rect 338316 181212 338322 181224
rect 341754 181212 341760 181224
rect 341812 181212 341818 181264
rect 343502 181212 343508 181264
rect 343560 181252 343566 181264
rect 343560 181224 346676 181252
rect 343560 181212 343566 181224
rect 59406 181144 59412 181196
rect 59464 181184 59470 181196
rect 64098 181184 64104 181196
rect 59464 181156 64104 181184
rect 59464 181144 59470 181156
rect 64098 181144 64104 181156
rect 64156 181144 64162 181196
rect 149750 181144 149756 181196
rect 149808 181184 149814 181196
rect 159594 181184 159600 181196
rect 149808 181156 159600 181184
rect 149808 181144 149814 181156
rect 159594 181144 159600 181156
rect 159652 181144 159658 181196
rect 344330 181144 344336 181196
rect 344388 181184 344394 181196
rect 345345 181187 345403 181193
rect 345345 181184 345357 181187
rect 344388 181156 345357 181184
rect 344388 181144 344394 181156
rect 345345 181153 345357 181156
rect 345391 181153 345403 181187
rect 346648 181184 346676 181224
rect 347274 181212 347280 181264
rect 347332 181252 347338 181264
rect 350402 181252 350408 181264
rect 347332 181224 350408 181252
rect 347332 181212 347338 181224
rect 350402 181212 350408 181224
rect 350460 181212 350466 181264
rect 348102 181184 348108 181196
rect 346648 181156 348108 181184
rect 345345 181147 345403 181153
rect 348102 181144 348108 181156
rect 348160 181144 348166 181196
rect 149198 181076 149204 181128
rect 149256 181116 149262 181128
rect 158950 181116 158956 181128
rect 149256 181088 158956 181116
rect 149256 181076 149262 181088
rect 158950 181076 158956 181088
rect 159008 181076 159014 181128
rect 248466 181076 248472 181128
rect 248524 181116 248530 181128
rect 257574 181116 257580 181128
rect 248524 181088 257580 181116
rect 248524 181076 248530 181088
rect 257574 181076 257580 181088
rect 257632 181076 257638 181128
rect 339638 181076 339644 181128
rect 339696 181116 339702 181128
rect 351230 181116 351236 181128
rect 339696 181088 351236 181116
rect 339696 181076 339702 181088
rect 351230 181076 351236 181088
rect 351288 181076 351294 181128
rect 151958 181008 151964 181060
rect 152016 181048 152022 181060
rect 163274 181048 163280 181060
rect 152016 181020 163280 181048
rect 152016 181008 152022 181020
rect 163274 181008 163280 181020
rect 163332 181008 163338 181060
rect 243498 181008 243504 181060
rect 243556 181048 243562 181060
rect 252790 181048 252796 181060
rect 243556 181020 252796 181048
rect 243556 181008 243562 181020
rect 252790 181008 252796 181020
rect 252848 181008 252854 181060
rect 334118 181008 334124 181060
rect 334176 181048 334182 181060
rect 346170 181048 346176 181060
rect 334176 181020 346176 181048
rect 334176 181008 334182 181020
rect 346170 181008 346176 181020
rect 346228 181008 346234 181060
rect 66398 180940 66404 180992
rect 66456 180980 66462 180992
rect 70354 180980 70360 180992
rect 66456 180952 70360 180980
rect 66456 180940 66462 180952
rect 70354 180940 70360 180952
rect 70412 180940 70418 180992
rect 150302 180940 150308 180992
rect 150360 180980 150366 180992
rect 162722 180980 162728 180992
rect 150360 180952 162728 180980
rect 150360 180940 150366 180952
rect 162722 180940 162728 180952
rect 162780 180940 162786 180992
rect 244050 180940 244056 180992
rect 244108 180980 244114 180992
rect 253434 180980 253440 180992
rect 244108 180952 253440 180980
rect 244108 180940 244114 180952
rect 253434 180940 253440 180952
rect 253492 180940 253498 180992
rect 335498 180940 335504 180992
rect 335556 180980 335562 180992
rect 346998 180980 347004 180992
rect 335556 180952 347004 180980
rect 335556 180940 335562 180952
rect 346998 180940 347004 180952
rect 347056 180940 347062 180992
rect 34658 180872 34664 180924
rect 34716 180912 34722 180924
rect 46986 180912 46992 180924
rect 34716 180884 46992 180912
rect 34716 180872 34722 180884
rect 46986 180872 46992 180884
rect 47044 180872 47050 180924
rect 62350 180872 62356 180924
rect 62408 180912 62414 180924
rect 63546 180912 63552 180924
rect 62408 180884 63552 180912
rect 62408 180872 62414 180884
rect 63546 180872 63552 180884
rect 63604 180872 63610 180924
rect 147818 180872 147824 180924
rect 147876 180912 147882 180924
rect 161434 180912 161440 180924
rect 147876 180884 161440 180912
rect 147876 180872 147882 180884
rect 161434 180872 161440 180884
rect 161492 180872 161498 180924
rect 241658 180872 241664 180924
rect 241716 180912 241722 180924
rect 255090 180912 255096 180924
rect 241716 180884 255096 180912
rect 241716 180872 241722 180884
rect 255090 180872 255096 180884
rect 255148 180872 255154 180924
rect 336878 180872 336884 180924
rect 336936 180912 336942 180924
rect 348746 180912 348752 180924
rect 336936 180884 348752 180912
rect 336936 180872 336942 180884
rect 348746 180872 348752 180884
rect 348804 180872 348810 180924
rect 31806 180804 31812 180856
rect 31864 180844 31870 180856
rect 46710 180844 46716 180856
rect 31864 180816 46716 180844
rect 31864 180804 31870 180816
rect 46710 180804 46716 180816
rect 46768 180804 46774 180856
rect 64926 180804 64932 180856
rect 64984 180844 64990 180856
rect 68606 180844 68612 180856
rect 64984 180816 68612 180844
rect 64984 180804 64990 180816
rect 68606 180804 68612 180816
rect 68664 180804 68670 180856
rect 149198 180804 149204 180856
rect 149256 180844 149262 180856
rect 162078 180844 162084 180856
rect 149256 180816 162084 180844
rect 149256 180804 149262 180816
rect 162078 180804 162084 180816
rect 162136 180804 162142 180856
rect 243038 180804 243044 180856
rect 243096 180844 243102 180856
rect 255734 180844 255740 180856
rect 243096 180816 255740 180844
rect 243096 180804 243102 180816
rect 255734 180804 255740 180816
rect 255792 180804 255798 180856
rect 338258 180804 338264 180856
rect 338316 180844 338322 180856
rect 349574 180844 349580 180856
rect 338316 180816 349580 180844
rect 338316 180804 338322 180816
rect 349574 180804 349580 180816
rect 349632 180804 349638 180856
rect 29506 180736 29512 180788
rect 29564 180776 29570 180788
rect 46618 180776 46624 180788
rect 29564 180748 46624 180776
rect 29564 180736 29570 180748
rect 46618 180736 46624 180748
rect 46676 180736 46682 180788
rect 65018 180736 65024 180788
rect 65076 180776 65082 180788
rect 69434 180776 69440 180788
rect 65076 180748 69440 180776
rect 65076 180736 65082 180748
rect 69434 180736 69440 180748
rect 69492 180736 69498 180788
rect 145058 180736 145064 180788
rect 145116 180776 145122 180788
rect 160238 180776 160244 180788
rect 145116 180748 160244 180776
rect 145116 180736 145122 180748
rect 160238 180736 160244 180748
rect 160296 180736 160302 180788
rect 240278 180736 240284 180788
rect 240336 180776 240342 180788
rect 254538 180776 254544 180788
rect 240336 180748 254544 180776
rect 240336 180736 240342 180748
rect 254538 180736 254544 180748
rect 254596 180736 254602 180788
rect 340926 180736 340932 180788
rect 340984 180776 340990 180788
rect 345253 180779 345311 180785
rect 345253 180776 345265 180779
rect 340984 180748 345265 180776
rect 340984 180736 340990 180748
rect 345253 180745 345265 180748
rect 345299 180745 345311 180779
rect 345253 180739 345311 180745
rect 345345 180779 345403 180785
rect 345345 180745 345357 180779
rect 345391 180776 345403 180779
rect 349390 180776 349396 180788
rect 345391 180748 349396 180776
rect 345391 180745 345403 180748
rect 345345 180739 345403 180745
rect 349390 180736 349396 180748
rect 349448 180736 349454 180788
rect 26930 180668 26936 180720
rect 26988 180708 26994 180720
rect 46526 180708 46532 180720
rect 26988 180680 46532 180708
rect 26988 180668 26994 180680
rect 46526 180668 46532 180680
rect 46584 180668 46590 180720
rect 146438 180668 146444 180720
rect 146496 180708 146502 180720
rect 160882 180708 160888 180720
rect 146496 180680 160888 180708
rect 146496 180668 146502 180680
rect 160882 180668 160888 180680
rect 160940 180668 160946 180720
rect 237518 180668 237524 180720
rect 237576 180708 237582 180720
rect 253526 180708 253532 180720
rect 237576 180680 253532 180708
rect 237576 180668 237582 180680
rect 253526 180668 253532 180680
rect 253584 180668 253590 180720
rect 332738 180668 332744 180720
rect 332796 180708 332802 180720
rect 345434 180708 345440 180720
rect 332796 180680 345440 180708
rect 332796 180668 332802 180680
rect 345434 180668 345440 180680
rect 345492 180668 345498 180720
rect 24170 180600 24176 180652
rect 24228 180640 24234 180652
rect 46434 180640 46440 180652
rect 24228 180612 46440 180640
rect 24228 180600 24234 180612
rect 46434 180600 46440 180612
rect 46492 180600 46498 180652
rect 57014 180600 57020 180652
rect 57072 180640 57078 180652
rect 67134 180640 67140 180652
rect 57072 180612 67140 180640
rect 57072 180600 57078 180612
rect 67134 180600 67140 180612
rect 67192 180600 67198 180652
rect 143678 180600 143684 180652
rect 143736 180640 143742 180652
rect 159318 180640 159324 180652
rect 143736 180612 159324 180640
rect 143736 180600 143742 180612
rect 159318 180600 159324 180612
rect 159376 180600 159382 180652
rect 238898 180600 238904 180652
rect 238956 180640 238962 180652
rect 254170 180640 254176 180652
rect 238956 180612 254176 180640
rect 238956 180600 238962 180612
rect 254170 180600 254176 180612
rect 254228 180600 254234 180652
rect 335406 180600 335412 180652
rect 335464 180640 335470 180652
rect 348010 180640 348016 180652
rect 335464 180612 348016 180640
rect 335464 180600 335470 180612
rect 348010 180600 348016 180612
rect 348068 180600 348074 180652
rect 254814 180532 254820 180584
rect 254872 180572 254878 180584
rect 256930 180572 256936 180584
rect 254872 180544 256936 180572
rect 254872 180532 254878 180544
rect 256930 180532 256936 180544
rect 256988 180532 256994 180584
rect 345253 180575 345311 180581
rect 345253 180541 345265 180575
rect 345299 180572 345311 180575
rect 352150 180572 352156 180584
rect 345299 180544 352156 180572
rect 345299 180541 345311 180544
rect 345253 180535 345311 180541
rect 352150 180532 352156 180544
rect 352208 180532 352214 180584
rect 340098 180328 340104 180380
rect 340156 180368 340162 180380
rect 341018 180368 341024 180380
rect 340156 180340 341024 180368
rect 340156 180328 340162 180340
rect 341018 180328 341024 180340
rect 341076 180328 341082 180380
rect 341662 180192 341668 180244
rect 341720 180232 341726 180244
rect 345986 180232 345992 180244
rect 341720 180204 345992 180232
rect 341720 180192 341726 180204
rect 345986 180192 345992 180204
rect 346044 180192 346050 180244
rect 60602 180124 60608 180176
rect 60660 180164 60666 180176
rect 65938 180164 65944 180176
rect 60660 180136 65944 180164
rect 60660 180124 60666 180136
rect 65938 180124 65944 180136
rect 65996 180124 66002 180176
rect 63270 180096 63276 180108
rect 57860 180068 63276 180096
rect 57860 180040 57888 180068
rect 63270 180056 63276 180068
rect 63328 180056 63334 180108
rect 57842 179988 57848 180040
rect 57900 179988 57906 180040
rect 62258 179988 62264 180040
rect 62316 180028 62322 180040
rect 66766 180028 66772 180040
rect 62316 180000 66772 180028
rect 62316 179988 62322 180000
rect 66766 179988 66772 180000
rect 66824 179988 66830 180040
rect 340834 179988 340840 180040
rect 340892 180028 340898 180040
rect 345250 180028 345256 180040
rect 340892 180000 345256 180028
rect 340892 179988 340898 180000
rect 345250 179988 345256 180000
rect 345308 179988 345314 180040
rect 63638 179920 63644 179972
rect 63696 179960 63702 179972
rect 67686 179960 67692 179972
rect 63696 179932 67692 179960
rect 63696 179920 63702 179932
rect 67686 179920 67692 179932
rect 67744 179920 67750 179972
rect 152234 179920 152240 179972
rect 152292 179960 152298 179972
rect 153246 179960 153252 179972
rect 152292 179932 153252 179960
rect 152292 179920 152298 179932
rect 153246 179920 153252 179932
rect 153304 179920 153310 179972
rect 153430 179920 153436 179972
rect 153488 179960 153494 179972
rect 154626 179960 154632 179972
rect 153488 179932 154632 179960
rect 153488 179920 153494 179932
rect 154626 179920 154632 179932
rect 154684 179920 154690 179972
rect 342398 179920 342404 179972
rect 342456 179960 342462 179972
rect 345894 179960 345900 179972
rect 342456 179932 345900 179960
rect 342456 179920 342462 179932
rect 345894 179920 345900 179932
rect 345952 179920 345958 179972
rect 230986 179716 230992 179768
rect 231044 179756 231050 179768
rect 232734 179756 232740 179768
rect 231044 179728 232740 179756
rect 231044 179716 231050 179728
rect 232734 179716 232740 179728
rect 232792 179716 232798 179768
rect 324550 179444 324556 179496
rect 324608 179484 324614 179496
rect 326574 179484 326580 179496
rect 324608 179456 326580 179484
rect 324608 179444 324614 179456
rect 326574 179444 326580 179456
rect 326632 179444 326638 179496
rect 273858 178492 273864 178544
rect 273916 178532 273922 178544
rect 276250 178532 276256 178544
rect 273916 178504 276256 178532
rect 273916 178492 273922 178504
rect 276250 178492 276256 178504
rect 276308 178492 276314 178544
rect 369078 175840 369084 175892
rect 369136 175880 369142 175892
rect 369906 175880 369912 175892
rect 369136 175852 369912 175880
rect 369136 175840 369142 175852
rect 369906 175840 369912 175852
rect 369964 175840 369970 175892
rect 13038 175772 13044 175824
rect 13096 175812 13102 175824
rect 16074 175812 16080 175824
rect 13096 175784 16080 175812
rect 13096 175772 13102 175784
rect 16074 175772 16080 175784
rect 16132 175772 16138 175824
rect 88386 175772 88392 175824
rect 88444 175812 88450 175824
rect 182410 175812 182416 175824
rect 88444 175784 182416 175812
rect 88444 175772 88450 175784
rect 182410 175772 182416 175784
rect 182468 175812 182474 175824
rect 182962 175812 182968 175824
rect 182468 175784 182968 175812
rect 182468 175772 182474 175784
rect 182962 175772 182968 175784
rect 183020 175812 183026 175824
rect 276434 175812 276440 175824
rect 183020 175784 276440 175812
rect 183020 175772 183026 175784
rect 276434 175772 276440 175784
rect 276492 175772 276498 175824
rect 95470 175704 95476 175756
rect 95528 175744 95534 175756
rect 174866 175744 174872 175756
rect 95528 175716 174872 175744
rect 95528 175704 95534 175716
rect 174866 175704 174872 175716
rect 174924 175704 174930 175756
rect 189310 175704 189316 175756
rect 189368 175744 189374 175756
rect 189494 175744 189500 175756
rect 189368 175716 189500 175744
rect 189368 175704 189374 175716
rect 189494 175704 189500 175716
rect 189552 175744 189558 175756
rect 283518 175744 283524 175756
rect 189552 175716 283524 175744
rect 189552 175704 189558 175716
rect 283518 175704 283524 175716
rect 283576 175704 283582 175756
rect 196670 175636 196676 175688
rect 196728 175676 196734 175688
rect 264474 175676 264480 175688
rect 196728 175648 264480 175676
rect 196728 175636 196734 175648
rect 264474 175636 264480 175648
rect 264532 175676 264538 175688
rect 290694 175676 290700 175688
rect 264532 175648 290700 175676
rect 264532 175636 264538 175648
rect 290694 175636 290700 175648
rect 290752 175636 290758 175688
rect 96758 175160 96764 175212
rect 96816 175200 96822 175212
rect 109730 175200 109736 175212
rect 96816 175172 109736 175200
rect 96816 175160 96822 175172
rect 109730 175160 109736 175172
rect 109788 175160 109794 175212
rect 112674 175160 112680 175212
rect 112732 175200 112738 175212
rect 116906 175200 116912 175212
rect 112732 175172 116912 175200
rect 112732 175160 112738 175172
rect 116906 175160 116912 175172
rect 116964 175160 116970 175212
rect 174866 175160 174872 175212
rect 174924 175200 174930 175212
rect 176154 175200 176160 175212
rect 174924 175172 176160 175200
rect 174924 175160 174930 175172
rect 176154 175160 176160 175172
rect 176212 175200 176218 175212
rect 189310 175200 189316 175212
rect 176212 175172 189316 175200
rect 176212 175160 176218 175172
rect 189310 175160 189316 175172
rect 189368 175160 189374 175212
rect 190598 175160 190604 175212
rect 190656 175200 190662 175212
rect 203754 175200 203760 175212
rect 190656 175172 203760 175200
rect 190656 175160 190662 175172
rect 203754 175160 203760 175172
rect 203812 175160 203818 175212
rect 102646 175092 102652 175144
rect 102704 175132 102710 175144
rect 174774 175132 174780 175144
rect 102704 175104 174780 175132
rect 102704 175092 102710 175104
rect 174774 175092 174780 175104
rect 174832 175132 174838 175144
rect 196670 175132 196676 175144
rect 174832 175104 196676 175132
rect 174832 175092 174838 175104
rect 196670 175092 196676 175104
rect 196728 175092 196734 175144
rect 285818 175092 285824 175144
rect 285876 175132 285882 175144
rect 297778 175132 297784 175144
rect 285876 175104 297784 175132
rect 285876 175092 285882 175104
rect 297778 175092 297784 175104
rect 297836 175092 297842 175144
rect 354910 175092 354916 175144
rect 354968 175132 354974 175144
rect 355830 175132 355836 175144
rect 354968 175104 355836 175132
rect 354968 175092 354974 175104
rect 355830 175092 355836 175104
rect 355888 175092 355894 175144
rect 206514 174752 206520 174804
rect 206572 174792 206578 174804
rect 210930 174792 210936 174804
rect 206572 174764 210936 174792
rect 206572 174752 206578 174764
rect 210930 174752 210936 174764
rect 210988 174752 210994 174804
rect 129234 174412 129240 174464
rect 129292 174452 129298 174464
rect 131166 174452 131172 174464
rect 129292 174424 131172 174452
rect 129292 174412 129298 174424
rect 131166 174412 131172 174424
rect 131224 174412 131230 174464
rect 300354 174412 300360 174464
rect 300412 174452 300418 174464
rect 304954 174452 304960 174464
rect 300412 174424 304960 174452
rect 300412 174412 300418 174424
rect 304954 174412 304960 174424
rect 305012 174412 305018 174464
rect 57842 172984 57848 173036
rect 57900 173024 57906 173036
rect 58118 173024 58124 173036
rect 57900 172996 58124 173024
rect 57900 172984 57906 172996
rect 58118 172984 58124 172996
rect 58176 172984 58182 173036
rect 58670 172984 58676 173036
rect 58728 173024 58734 173036
rect 59406 173024 59412 173036
rect 58728 172996 59412 173024
rect 58728 172984 58734 172996
rect 59406 172984 59412 172996
rect 59464 172984 59470 173036
rect 59682 172984 59688 173036
rect 59740 173024 59746 173036
rect 60786 173024 60792 173036
rect 59740 172996 60792 173024
rect 59740 172984 59746 172996
rect 60786 172984 60792 172996
rect 60844 172984 60850 173036
rect 62810 172984 62816 173036
rect 62868 173024 62874 173036
rect 63638 173024 63644 173036
rect 62868 172996 63644 173024
rect 62868 172984 62874 172996
rect 63638 172984 63644 172996
rect 63696 172984 63702 173036
rect 63822 172984 63828 173036
rect 63880 173024 63886 173036
rect 64926 173024 64932 173036
rect 63880 172996 64932 173024
rect 63880 172984 63886 172996
rect 64926 172984 64932 172996
rect 64984 172984 64990 173036
rect 67134 172984 67140 173036
rect 67192 173024 67198 173036
rect 68974 173024 68980 173036
rect 67192 172996 68980 173024
rect 67192 172984 67198 172996
rect 68974 172984 68980 172996
rect 69032 172984 69038 173036
rect 153154 172984 153160 173036
rect 153212 173024 153218 173036
rect 153338 173024 153344 173036
rect 153212 172996 153344 173024
rect 153212 172984 153218 172996
rect 153338 172984 153344 172996
rect 153396 172984 153402 173036
rect 159594 172984 159600 173036
rect 159652 173024 159658 173036
rect 160330 173024 160336 173036
rect 159652 172996 160336 173024
rect 159652 172984 159658 172996
rect 160330 172984 160336 172996
rect 160388 172984 160394 173036
rect 253434 172984 253440 173036
rect 253492 173024 253498 173036
rect 254170 173024 254176 173036
rect 253492 172996 254176 173024
rect 253492 172984 253498 172996
rect 254170 172984 254176 172996
rect 254228 172984 254234 173036
rect 333382 172984 333388 173036
rect 333440 173024 333446 173036
rect 334118 173024 334124 173036
rect 333440 172996 334124 173024
rect 333440 172984 333446 172996
rect 334118 172984 334124 172996
rect 334176 172984 334182 173036
rect 341754 172984 341760 173036
rect 341812 173024 341818 173036
rect 342674 173024 342680 173036
rect 341812 172996 342680 173024
rect 341812 172984 341818 172996
rect 342674 172984 342680 172996
rect 342732 172984 342738 173036
rect 345986 172984 345992 173036
rect 346044 173024 346050 173036
rect 346814 173024 346820 173036
rect 346044 172996 346820 173024
rect 346044 172984 346050 172996
rect 346814 172984 346820 172996
rect 346872 172984 346878 173036
rect 427590 172984 427596 173036
rect 427648 173024 427654 173036
rect 429890 173024 429896 173036
rect 427648 172996 429896 173024
rect 427648 172984 427654 172996
rect 429890 172984 429896 172996
rect 429948 172984 429954 173036
rect 154718 172916 154724 172968
rect 154776 172956 154782 172968
rect 164654 172956 164660 172968
rect 154776 172928 164660 172956
rect 154776 172916 154782 172928
rect 164654 172916 164660 172928
rect 164712 172916 164718 172968
rect 246258 172916 246264 172968
rect 246316 172956 246322 172968
rect 254814 172956 254820 172968
rect 246316 172928 254820 172956
rect 246316 172916 246322 172928
rect 254814 172916 254820 172928
rect 254872 172916 254878 172968
rect 254909 172959 254967 172965
rect 254909 172925 254921 172959
rect 254955 172956 254967 172959
rect 258678 172956 258684 172968
rect 254955 172928 258684 172956
rect 254955 172925 254967 172928
rect 254909 172919 254967 172925
rect 258678 172916 258684 172928
rect 258736 172916 258742 172968
rect 341018 172916 341024 172968
rect 341076 172956 341082 172968
rect 344790 172956 344796 172968
rect 341076 172928 344796 172956
rect 341076 172916 341082 172928
rect 344790 172916 344796 172928
rect 344848 172916 344854 172968
rect 345894 172916 345900 172968
rect 345952 172956 345958 172968
rect 347918 172956 347924 172968
rect 345952 172928 347924 172956
rect 345952 172916 345958 172928
rect 347918 172916 347924 172928
rect 347976 172916 347982 172968
rect 153338 172848 153344 172900
rect 153396 172888 153402 172900
rect 163918 172888 163924 172900
rect 153396 172860 163924 172888
rect 153396 172848 153402 172860
rect 163918 172848 163924 172860
rect 163976 172848 163982 172900
rect 244878 172848 244884 172900
rect 244936 172888 244942 172900
rect 256746 172888 256752 172900
rect 244936 172860 256752 172888
rect 244936 172848 244942 172860
rect 256746 172848 256752 172860
rect 256804 172848 256810 172900
rect 334394 172848 334400 172900
rect 334452 172888 334458 172900
rect 335498 172888 335504 172900
rect 334452 172860 335504 172888
rect 334452 172848 334458 172860
rect 335498 172848 335504 172860
rect 335556 172848 335562 172900
rect 339546 172848 339552 172900
rect 339604 172888 339610 172900
rect 343778 172888 343784 172900
rect 339604 172860 343784 172888
rect 339604 172848 339610 172860
rect 343778 172848 343784 172860
rect 343836 172848 343842 172900
rect 59498 172780 59504 172832
rect 59556 172820 59562 172832
rect 71090 172820 71096 172832
rect 59556 172792 71096 172820
rect 59556 172780 59562 172792
rect 71090 172780 71096 172792
rect 71148 172780 71154 172832
rect 150394 172780 150400 172832
rect 150452 172820 150458 172832
rect 161710 172820 161716 172832
rect 150452 172792 161716 172820
rect 150452 172780 150458 172792
rect 161710 172780 161716 172792
rect 161768 172780 161774 172832
rect 60878 172712 60884 172764
rect 60936 172752 60942 172764
rect 72102 172752 72108 172764
rect 60936 172724 72108 172752
rect 60936 172712 60942 172724
rect 72102 172712 72108 172724
rect 72160 172712 72166 172764
rect 151314 172712 151320 172764
rect 151372 172752 151378 172764
rect 163090 172752 163096 172764
rect 151372 172724 163096 172752
rect 151372 172712 151378 172724
rect 163090 172712 163096 172724
rect 163148 172712 163154 172764
rect 244418 172712 244424 172764
rect 244476 172752 244482 172764
rect 255550 172752 255556 172764
rect 244476 172724 255556 172752
rect 244476 172712 244482 172724
rect 255550 172712 255556 172724
rect 255608 172712 255614 172764
rect 57934 172644 57940 172696
rect 57992 172684 57998 172696
rect 70078 172684 70084 172696
rect 57992 172656 70084 172684
rect 57992 172644 57998 172656
rect 70078 172644 70084 172656
rect 70136 172644 70142 172696
rect 143034 172644 143040 172696
rect 143092 172684 143098 172696
rect 155730 172684 155736 172696
rect 143092 172656 155736 172684
rect 143092 172644 143098 172656
rect 155730 172644 155736 172656
rect 155788 172644 155794 172696
rect 157846 172644 157852 172696
rect 157904 172684 157910 172696
rect 165114 172684 165120 172696
rect 157904 172656 165120 172684
rect 157904 172644 157910 172656
rect 165114 172644 165120 172656
rect 165172 172644 165178 172696
rect 245522 172644 245528 172696
rect 245580 172684 245586 172696
rect 258310 172684 258316 172696
rect 245580 172656 258316 172684
rect 245580 172644 245586 172656
rect 258310 172644 258316 172656
rect 258368 172644 258374 172696
rect 55358 172576 55364 172628
rect 55416 172616 55422 172628
rect 66950 172616 66956 172628
rect 55416 172588 66956 172616
rect 55416 172576 55422 172588
rect 66950 172576 66956 172588
rect 67008 172576 67014 172628
rect 153246 172576 153252 172628
rect 153304 172616 153310 172628
rect 165850 172616 165856 172628
rect 153304 172588 165856 172616
rect 153304 172576 153310 172588
rect 165850 172576 165856 172588
rect 165908 172576 165914 172628
rect 246810 172576 246816 172628
rect 246868 172616 246874 172628
rect 259690 172616 259696 172628
rect 246868 172588 259696 172616
rect 246868 172576 246874 172588
rect 259690 172576 259696 172588
rect 259748 172576 259754 172628
rect 56738 172508 56744 172560
rect 56796 172548 56802 172560
rect 67962 172548 67968 172560
rect 56796 172520 67968 172548
rect 56796 172508 56802 172520
rect 67962 172508 67968 172520
rect 68020 172508 68026 172560
rect 151590 172508 151596 172560
rect 151648 172548 151654 172560
rect 164470 172548 164476 172560
rect 151648 172520 164476 172548
rect 151648 172508 151654 172520
rect 164470 172508 164476 172520
rect 164528 172508 164534 172560
rect 236874 172508 236880 172560
rect 236932 172548 236938 172560
rect 250030 172548 250036 172560
rect 236932 172520 250036 172548
rect 236932 172508 236938 172520
rect 250030 172508 250036 172520
rect 250088 172508 250094 172560
rect 63546 172440 63552 172492
rect 63604 172480 63610 172492
rect 75230 172480 75236 172492
rect 63604 172452 75236 172480
rect 63604 172440 63610 172452
rect 75230 172440 75236 172452
rect 75288 172440 75294 172492
rect 153154 172440 153160 172492
rect 153212 172480 153218 172492
rect 167322 172480 167328 172492
rect 153212 172452 167328 172480
rect 153212 172440 153218 172452
rect 167322 172440 167328 172452
rect 167380 172440 167386 172492
rect 246902 172440 246908 172492
rect 246960 172480 246966 172492
rect 261162 172480 261168 172492
rect 246960 172452 261168 172480
rect 246960 172440 246966 172452
rect 261162 172440 261168 172452
rect 261220 172440 261226 172492
rect 62166 172372 62172 172424
rect 62224 172412 62230 172424
rect 74218 172412 74224 172424
rect 62224 172384 74224 172412
rect 62224 172372 62230 172384
rect 74218 172372 74224 172384
rect 74276 172372 74282 172424
rect 154534 172372 154540 172424
rect 154592 172412 154598 172424
rect 168702 172412 168708 172424
rect 154592 172384 168708 172412
rect 154592 172372 154598 172384
rect 168702 172372 168708 172384
rect 168760 172372 168766 172424
rect 248374 172372 248380 172424
rect 248432 172412 248438 172424
rect 262450 172412 262456 172424
rect 248432 172384 262456 172412
rect 248432 172372 248438 172384
rect 262450 172372 262456 172384
rect 262508 172372 262514 172424
rect 60694 172304 60700 172356
rect 60752 172344 60758 172356
rect 73114 172344 73120 172356
rect 60752 172316 73120 172344
rect 60752 172304 60758 172316
rect 73114 172304 73120 172316
rect 73172 172304 73178 172356
rect 154626 172304 154632 172356
rect 154684 172344 154690 172356
rect 170082 172344 170088 172356
rect 154684 172316 170088 172344
rect 154684 172304 154690 172316
rect 170082 172304 170088 172316
rect 170140 172304 170146 172356
rect 248558 172304 248564 172356
rect 248616 172344 248622 172356
rect 263830 172344 263836 172356
rect 248616 172316 263836 172344
rect 248616 172304 248622 172316
rect 263830 172304 263836 172316
rect 263888 172304 263894 172356
rect 245798 172236 245804 172288
rect 245856 172276 245862 172288
rect 256930 172276 256936 172288
rect 245856 172248 256936 172276
rect 245856 172236 245862 172248
rect 256930 172236 256936 172248
rect 256988 172236 256994 172288
rect 249018 172168 249024 172220
rect 249076 172208 249082 172220
rect 254909 172211 254967 172217
rect 254909 172208 254921 172211
rect 249076 172180 254921 172208
rect 249076 172168 249082 172180
rect 254909 172177 254921 172180
rect 254955 172177 254967 172211
rect 254909 172171 254967 172177
rect 247638 171896 247644 171948
rect 247696 171936 247702 171948
rect 248466 171936 248472 171948
rect 247696 171908 248472 171936
rect 247696 171896 247702 171908
rect 248466 171896 248472 171908
rect 248524 171896 248530 171948
rect 338534 171896 338540 171948
rect 338592 171936 338598 171948
rect 347274 171936 347280 171948
rect 338592 171908 347280 171936
rect 338592 171896 338598 171908
rect 347274 171896 347280 171908
rect 347332 171896 347338 171948
rect 251870 171760 251876 171812
rect 251928 171800 251934 171812
rect 258954 171800 258960 171812
rect 251928 171772 258960 171800
rect 251928 171760 251934 171772
rect 258954 171760 258960 171772
rect 259012 171760 259018 171812
rect 46710 171624 46716 171676
rect 46768 171664 46774 171676
rect 46894 171664 46900 171676
rect 46768 171636 46900 171664
rect 46768 171624 46774 171636
rect 46894 171624 46900 171636
rect 46952 171664 46958 171676
rect 72654 171664 72660 171676
rect 46952 171636 72660 171664
rect 46952 171624 46958 171636
rect 72654 171624 72660 171636
rect 72712 171624 72718 171676
rect 369722 170264 369728 170316
rect 369780 170304 369786 170316
rect 369906 170304 369912 170316
rect 369780 170276 369912 170304
rect 369780 170264 369786 170276
rect 369906 170264 369912 170276
rect 369964 170264 369970 170316
rect 79186 170196 79192 170248
rect 79244 170236 79250 170248
rect 123990 170236 123996 170248
rect 79244 170208 123996 170236
rect 79244 170196 79250 170208
rect 123990 170196 123996 170208
rect 124048 170196 124054 170248
rect 312038 170196 312044 170248
rect 312096 170236 312102 170248
rect 328414 170236 328420 170248
rect 312096 170208 328420 170236
rect 312096 170196 312102 170208
rect 328414 170196 328420 170208
rect 328472 170196 328478 170248
rect 123990 169516 123996 169568
rect 124048 169556 124054 169568
rect 140274 169556 140280 169568
rect 124048 169528 140280 169556
rect 124048 169516 124054 169528
rect 140274 169516 140280 169528
rect 140332 169516 140338 169568
rect 267234 169516 267240 169568
rect 267292 169556 267298 169568
rect 312038 169556 312044 169568
rect 267292 169528 312044 169556
rect 267292 169516 267298 169528
rect 312038 169516 312044 169528
rect 312096 169516 312102 169568
rect 73482 169420 73488 169432
rect 73443 169392 73488 169420
rect 73482 169380 73488 169392
rect 73540 169380 73546 169432
rect 132178 168904 132184 168956
rect 132236 168944 132242 168956
rect 140550 168944 140556 168956
rect 132236 168916 140556 168944
rect 132236 168904 132242 168916
rect 140550 168904 140556 168916
rect 140608 168904 140614 168956
rect 226018 168904 226024 168956
rect 226076 168944 226082 168956
rect 233470 168944 233476 168956
rect 226076 168916 233476 168944
rect 226076 168904 226082 168916
rect 233470 168904 233476 168916
rect 233528 168904 233534 168956
rect 46986 168836 46992 168888
rect 47044 168876 47050 168888
rect 49194 168876 49200 168888
rect 47044 168848 49200 168876
rect 47044 168836 47050 168848
rect 49194 168836 49200 168848
rect 49252 168876 49258 168888
rect 73485 168879 73543 168885
rect 73485 168876 73497 168879
rect 49252 168848 73497 168876
rect 49252 168836 49258 168848
rect 73485 168845 73497 168848
rect 73531 168845 73543 168879
rect 73485 168839 73543 168845
rect 222154 168564 222160 168616
rect 222212 168604 222218 168616
rect 369262 168604 369268 168616
rect 222212 168576 369268 168604
rect 222212 168564 222218 168576
rect 369262 168564 369268 168576
rect 369320 168564 369326 168616
rect 128130 168496 128136 168548
rect 128188 168536 128194 168548
rect 369170 168536 369176 168548
rect 128188 168508 369176 168536
rect 128188 168496 128194 168508
rect 369170 168496 369176 168508
rect 369228 168496 369234 168548
rect 361166 168156 361172 168208
rect 361224 168196 361230 168208
rect 423634 168196 423640 168208
rect 361224 168168 423640 168196
rect 361224 168156 361230 168168
rect 423634 168156 423640 168168
rect 423692 168156 423698 168208
rect 77254 167544 77260 167596
rect 77312 167584 77318 167596
rect 87190 167584 87196 167596
rect 77312 167556 87196 167584
rect 77312 167544 77318 167556
rect 87190 167544 87196 167556
rect 87248 167544 87254 167596
rect 132270 167544 132276 167596
rect 132328 167584 132334 167596
rect 140550 167584 140556 167596
rect 132328 167556 140556 167584
rect 132328 167544 132334 167556
rect 140550 167544 140556 167556
rect 140608 167544 140614 167596
rect 225926 167544 225932 167596
rect 225984 167584 225990 167596
rect 233470 167584 233476 167596
rect 225984 167556 233476 167584
rect 225984 167544 225990 167556
rect 233470 167544 233476 167556
rect 233528 167544 233534 167596
rect 110190 166796 110196 166848
rect 110248 166836 110254 166848
rect 112674 166836 112680 166848
rect 110248 166808 112680 166836
rect 110248 166796 110254 166808
rect 112674 166796 112680 166808
rect 112732 166796 112738 166848
rect 203846 166796 203852 166848
rect 203904 166836 203910 166848
rect 206514 166836 206520 166848
rect 203904 166808 206520 166836
rect 203904 166796 203910 166808
rect 206514 166796 206520 166808
rect 206572 166796 206578 166848
rect 217186 166796 217192 166848
rect 217244 166836 217250 166848
rect 225190 166836 225196 166848
rect 217244 166808 225196 166836
rect 217244 166796 217250 166808
rect 225190 166796 225196 166808
rect 225248 166796 225254 166848
rect 297870 166796 297876 166848
rect 297928 166836 297934 166848
rect 300354 166836 300360 166848
rect 297928 166808 300360 166836
rect 297928 166796 297934 166808
rect 300354 166796 300360 166808
rect 300412 166796 300418 166848
rect 311210 166796 311216 166848
rect 311268 166836 311274 166848
rect 319214 166836 319220 166848
rect 311268 166808 319220 166836
rect 311268 166796 311274 166808
rect 319214 166796 319220 166808
rect 319272 166796 319278 166848
rect 123530 166524 123536 166576
rect 123588 166564 123594 166576
rect 129234 166564 129240 166576
rect 123588 166536 129240 166564
rect 123588 166524 123594 166536
rect 129234 166524 129240 166536
rect 129292 166524 129298 166576
rect 284530 166252 284536 166304
rect 284588 166292 284594 166304
rect 285818 166292 285824 166304
rect 284588 166264 285824 166292
rect 284588 166252 284594 166264
rect 285818 166252 285824 166264
rect 285876 166252 285882 166304
rect 77254 166184 77260 166236
rect 77312 166224 77318 166236
rect 87098 166224 87104 166236
rect 77312 166196 87104 166224
rect 77312 166184 77318 166196
rect 87098 166184 87104 166196
rect 87156 166184 87162 166236
rect 132086 166184 132092 166236
rect 132144 166224 132150 166236
rect 140550 166224 140556 166236
rect 132144 166196 140556 166224
rect 132144 166184 132150 166196
rect 140550 166184 140556 166196
rect 140608 166184 140614 166236
rect 225834 166184 225840 166236
rect 225892 166224 225898 166236
rect 233470 166224 233476 166236
rect 225892 166196 233476 166224
rect 225892 166184 225898 166196
rect 233470 166184 233476 166196
rect 233528 166184 233534 166236
rect 361718 165436 361724 165488
rect 361776 165476 361782 165488
rect 420874 165476 420880 165488
rect 361776 165448 420880 165476
rect 361776 165436 361782 165448
rect 420874 165436 420880 165448
rect 420932 165436 420938 165488
rect 77254 164756 77260 164808
rect 77312 164796 77318 164808
rect 87282 164796 87288 164808
rect 77312 164768 87288 164796
rect 77312 164756 77318 164768
rect 87282 164756 87288 164768
rect 87340 164756 87346 164808
rect 132638 164756 132644 164808
rect 132696 164796 132702 164808
rect 139630 164796 139636 164808
rect 132696 164768 139636 164796
rect 132696 164756 132702 164768
rect 139630 164756 139636 164768
rect 139688 164756 139694 164808
rect 225650 164756 225656 164808
rect 225708 164796 225714 164808
rect 233470 164796 233476 164808
rect 225708 164768 233476 164796
rect 225708 164756 225714 164768
rect 233470 164756 233476 164768
rect 233528 164756 233534 164808
rect 131350 163464 131356 163516
rect 131408 163504 131414 163516
rect 137606 163504 137612 163516
rect 131408 163476 137612 163504
rect 131408 163464 131414 163476
rect 137606 163464 137612 163476
rect 137664 163464 137670 163516
rect 226294 163464 226300 163516
rect 226352 163504 226358 163516
rect 231446 163504 231452 163516
rect 226352 163476 231452 163504
rect 226352 163464 226358 163476
rect 231446 163464 231452 163476
rect 231504 163464 231510 163516
rect 321606 163464 321612 163516
rect 321664 163504 321670 163516
rect 327218 163504 327224 163516
rect 321664 163476 327224 163504
rect 321664 163464 321670 163476
rect 327218 163464 327224 163476
rect 327276 163464 327282 163516
rect 77254 163396 77260 163448
rect 77312 163436 77318 163448
rect 87190 163436 87196 163448
rect 77312 163408 87196 163436
rect 77312 163396 77318 163408
rect 87190 163396 87196 163408
rect 87248 163396 87254 163448
rect 131902 163396 131908 163448
rect 131960 163436 131966 163448
rect 139630 163436 139636 163448
rect 131960 163408 139636 163436
rect 131960 163396 131966 163408
rect 139630 163396 139636 163408
rect 139688 163396 139694 163448
rect 226386 163396 226392 163448
rect 226444 163436 226450 163448
rect 233470 163436 233476 163448
rect 226444 163408 233476 163436
rect 226444 163396 226450 163408
rect 233470 163396 233476 163408
rect 233528 163396 233534 163448
rect 272846 163396 272852 163448
rect 272904 163436 272910 163448
rect 274870 163436 274876 163448
rect 272904 163408 274876 163436
rect 272904 163396 272910 163408
rect 274870 163396 274876 163408
rect 274928 163396 274934 163448
rect 361718 162648 361724 162700
rect 361776 162688 361782 162700
rect 418206 162688 418212 162700
rect 361776 162660 418212 162688
rect 361776 162648 361782 162660
rect 418206 162648 418212 162660
rect 418264 162648 418270 162700
rect 321606 162376 321612 162428
rect 321664 162416 321670 162428
rect 327494 162416 327500 162428
rect 321664 162388 327500 162416
rect 321664 162376 321670 162388
rect 327494 162376 327500 162388
rect 327552 162376 327558 162428
rect 131994 162104 132000 162156
rect 132052 162144 132058 162156
rect 139538 162144 139544 162156
rect 132052 162116 139544 162144
rect 132052 162104 132058 162116
rect 139538 162104 139544 162116
rect 139596 162104 139602 162156
rect 226386 162104 226392 162156
rect 226444 162144 226450 162156
rect 233470 162144 233476 162156
rect 226444 162116 233476 162144
rect 226444 162104 226450 162116
rect 233470 162104 233476 162116
rect 233528 162104 233534 162156
rect 132362 162036 132368 162088
rect 132420 162076 132426 162088
rect 139630 162076 139636 162088
rect 132420 162048 139636 162076
rect 132420 162036 132426 162048
rect 139630 162036 139636 162048
rect 139688 162036 139694 162088
rect 226202 162036 226208 162088
rect 226260 162076 226266 162088
rect 234574 162076 234580 162088
rect 226260 162048 234580 162076
rect 226260 162036 226266 162048
rect 234574 162036 234580 162048
rect 234632 162036 234638 162088
rect 131994 161968 132000 162020
rect 132052 162008 132058 162020
rect 132270 162008 132276 162020
rect 132052 161980 132276 162008
rect 132052 161968 132058 161980
rect 132270 161968 132276 161980
rect 132328 161968 132334 162020
rect 222430 161560 222436 161612
rect 222488 161560 222494 161612
rect 321054 161560 321060 161612
rect 321112 161600 321118 161612
rect 327218 161600 327224 161612
rect 321112 161572 327224 161600
rect 321112 161560 321118 161572
rect 327218 161560 327224 161572
rect 327276 161560 327282 161612
rect 173302 161492 173308 161544
rect 173360 161532 173366 161544
rect 222448 161532 222476 161560
rect 173360 161504 222476 161532
rect 173360 161492 173366 161504
rect 321606 161424 321612 161476
rect 321664 161464 321670 161476
rect 328414 161464 328420 161476
rect 321664 161436 328420 161464
rect 321664 161424 321670 161436
rect 328414 161424 328420 161436
rect 328472 161424 328478 161476
rect 272938 161084 272944 161136
rect 272996 161124 273002 161136
rect 275146 161124 275152 161136
rect 272996 161096 275152 161124
rect 272996 161084 273002 161096
rect 275146 161084 275152 161096
rect 275204 161084 275210 161136
rect 131350 160676 131356 160728
rect 131408 160716 131414 160728
rect 140458 160716 140464 160728
rect 131408 160688 140464 160716
rect 131408 160676 131414 160688
rect 140458 160676 140464 160688
rect 140516 160676 140522 160728
rect 131442 160608 131448 160660
rect 131500 160648 131506 160660
rect 140826 160648 140832 160660
rect 131500 160620 140832 160648
rect 131500 160608 131506 160620
rect 140826 160608 140832 160620
rect 140884 160608 140890 160660
rect 174038 160608 174044 160660
rect 174096 160648 174102 160660
rect 176246 160648 176252 160660
rect 174096 160620 176252 160648
rect 174096 160608 174102 160620
rect 176246 160608 176252 160620
rect 176304 160608 176310 160660
rect 179006 160608 179012 160660
rect 179064 160648 179070 160660
rect 182318 160648 182324 160660
rect 179064 160620 182324 160648
rect 179064 160608 179070 160620
rect 182318 160608 182324 160620
rect 182376 160608 182382 160660
rect 226294 160608 226300 160660
rect 226352 160648 226358 160660
rect 234298 160648 234304 160660
rect 226352 160620 234304 160648
rect 226352 160608 226358 160620
rect 234298 160608 234304 160620
rect 234356 160608 234362 160660
rect 266590 160608 266596 160660
rect 266648 160648 266654 160660
rect 269994 160648 270000 160660
rect 266648 160620 270000 160648
rect 266648 160608 266654 160620
rect 269994 160608 270000 160620
rect 270052 160608 270058 160660
rect 77254 160540 77260 160592
rect 77312 160580 77318 160592
rect 87190 160580 87196 160592
rect 77312 160552 87196 160580
rect 77312 160540 77318 160552
rect 87190 160540 87196 160552
rect 87248 160540 87254 160592
rect 131350 159316 131356 159368
rect 131408 159356 131414 159368
rect 140550 159356 140556 159368
rect 131408 159328 140556 159356
rect 131408 159316 131414 159328
rect 140550 159316 140556 159328
rect 140608 159316 140614 159368
rect 173670 159316 173676 159368
rect 173728 159356 173734 159368
rect 181490 159356 181496 159368
rect 173728 159328 181496 159356
rect 173728 159316 173734 159328
rect 181490 159316 181496 159328
rect 181548 159316 181554 159368
rect 266590 159316 266596 159368
rect 266648 159356 266654 159368
rect 275698 159356 275704 159368
rect 266648 159328 275704 159356
rect 266648 159316 266654 159328
rect 275698 159316 275704 159328
rect 275756 159316 275762 159368
rect 320594 159316 320600 159368
rect 320652 159356 320658 159368
rect 327310 159356 327316 159368
rect 320652 159328 327316 159356
rect 320652 159316 320658 159328
rect 327310 159316 327316 159328
rect 327368 159316 327374 159368
rect 79278 159248 79284 159300
rect 79336 159288 79342 159300
rect 79336 159260 85764 159288
rect 79336 159248 79342 159260
rect 85736 159152 85764 159260
rect 131810 159248 131816 159300
rect 131868 159288 131874 159300
rect 139630 159288 139636 159300
rect 131868 159260 139636 159288
rect 131868 159248 131874 159260
rect 139630 159248 139636 159260
rect 139688 159248 139694 159300
rect 172750 159248 172756 159300
rect 172808 159288 172814 159300
rect 181674 159288 181680 159300
rect 172808 159260 181680 159288
rect 172808 159248 172814 159260
rect 181674 159248 181680 159260
rect 181732 159248 181738 159300
rect 226110 159248 226116 159300
rect 226168 159288 226174 159300
rect 228686 159288 228692 159300
rect 226168 159260 228692 159288
rect 226168 159248 226174 159260
rect 228686 159248 228692 159260
rect 228744 159248 228750 159300
rect 231354 159248 231360 159300
rect 231412 159288 231418 159300
rect 233470 159288 233476 159300
rect 231412 159260 233476 159288
rect 231412 159248 231418 159260
rect 233470 159248 233476 159260
rect 233528 159248 233534 159300
rect 272754 159248 272760 159300
rect 272812 159288 272818 159300
rect 275146 159288 275152 159300
rect 272812 159260 275152 159288
rect 272812 159248 272818 159260
rect 275146 159248 275152 159260
rect 275204 159248 275210 159300
rect 87282 159152 87288 159164
rect 85736 159124 87288 159152
rect 87282 159112 87288 159124
rect 87340 159112 87346 159164
rect 131902 159112 131908 159164
rect 131960 159152 131966 159164
rect 132086 159152 132092 159164
rect 131960 159124 132092 159152
rect 131960 159112 131966 159124
rect 132086 159112 132092 159124
rect 132144 159112 132150 159164
rect 81762 159044 81768 159096
rect 81820 159084 81826 159096
rect 87190 159084 87196 159096
rect 81820 159056 87196 159084
rect 81820 159044 81826 159056
rect 87190 159044 87196 159056
rect 87248 159044 87254 159096
rect 361718 158500 361724 158552
rect 361776 158540 361782 158552
rect 415538 158540 415544 158552
rect 361776 158512 415544 158540
rect 361776 158500 361782 158512
rect 415538 158500 415544 158512
rect 415596 158500 415602 158552
rect 321606 158160 321612 158212
rect 321664 158200 321670 158212
rect 327218 158200 327224 158212
rect 321664 158172 327224 158200
rect 321664 158160 321670 158172
rect 327218 158160 327224 158172
rect 327276 158160 327282 158212
rect 173670 158024 173676 158076
rect 173728 158064 173734 158076
rect 181858 158064 181864 158076
rect 173728 158036 181864 158064
rect 173728 158024 173734 158036
rect 181858 158024 181864 158036
rect 181916 158024 181922 158076
rect 178914 157956 178920 158008
rect 178972 157996 178978 158008
rect 181398 157996 181404 158008
rect 178972 157968 181404 157996
rect 178972 157956 178978 157968
rect 181398 157956 181404 157968
rect 181456 157956 181462 158008
rect 266590 157956 266596 158008
rect 266648 157996 266654 158008
rect 271374 157996 271380 158008
rect 266648 157968 271380 157996
rect 266648 157956 266654 157968
rect 271374 157956 271380 157968
rect 271432 157956 271438 158008
rect 321054 157956 321060 158008
rect 321112 157996 321118 158008
rect 327402 157996 327408 158008
rect 321112 157968 327408 157996
rect 321112 157956 321118 157968
rect 327402 157956 327408 157968
rect 327460 157956 327466 158008
rect 79738 157888 79744 157940
rect 79796 157928 79802 157940
rect 79796 157900 84476 157928
rect 79796 157888 79802 157900
rect 84448 157792 84476 157900
rect 132178 157888 132184 157940
rect 132236 157928 132242 157940
rect 138894 157928 138900 157940
rect 132236 157900 138900 157928
rect 132236 157888 132242 157900
rect 138894 157888 138900 157900
rect 138952 157888 138958 157940
rect 173486 157888 173492 157940
rect 173544 157928 173550 157940
rect 182318 157928 182324 157940
rect 173544 157900 182324 157928
rect 173544 157888 173550 157900
rect 182318 157888 182324 157900
rect 182376 157888 182382 157940
rect 266958 157888 266964 157940
rect 267016 157928 267022 157940
rect 274870 157928 274876 157940
rect 267016 157900 274876 157928
rect 267016 157888 267022 157900
rect 274870 157888 274876 157900
rect 274928 157888 274934 157940
rect 87190 157792 87196 157804
rect 84448 157764 87196 157792
rect 87190 157752 87196 157764
rect 87248 157752 87254 157804
rect 222798 157140 222804 157192
rect 222856 157180 222862 157192
rect 233470 157180 233476 157192
rect 222856 157152 233476 157180
rect 222856 157140 222862 157152
rect 233470 157140 233476 157152
rect 233528 157140 233534 157192
rect 321606 157140 321612 157192
rect 321664 157180 321670 157192
rect 327218 157180 327224 157192
rect 321664 157152 327224 157180
rect 321664 157140 321670 157152
rect 327218 157140 327224 157152
rect 327276 157140 327282 157192
rect 77254 156460 77260 156512
rect 77312 156500 77318 156512
rect 77312 156472 85212 156500
rect 77312 156460 77318 156472
rect 85184 156432 85212 156472
rect 173118 156460 173124 156512
rect 173176 156500 173182 156512
rect 173302 156500 173308 156512
rect 173176 156472 173308 156500
rect 173176 156460 173182 156472
rect 173302 156460 173308 156472
rect 173360 156460 173366 156512
rect 173670 156460 173676 156512
rect 173728 156500 173734 156512
rect 182318 156500 182324 156512
rect 173728 156472 182324 156500
rect 173728 156460 173734 156472
rect 182318 156460 182324 156472
rect 182376 156460 182382 156512
rect 369814 156500 369820 156512
rect 369775 156472 369820 156500
rect 369814 156460 369820 156472
rect 369872 156460 369878 156512
rect 87190 156432 87196 156444
rect 85184 156404 87196 156432
rect 87190 156392 87196 156404
rect 87248 156392 87254 156444
rect 173578 156392 173584 156444
rect 173636 156432 173642 156444
rect 182134 156432 182140 156444
rect 173636 156404 182140 156432
rect 173636 156392 173642 156404
rect 182134 156392 182140 156404
rect 182192 156392 182198 156444
rect 267418 156392 267424 156444
rect 267476 156432 267482 156444
rect 274870 156432 274876 156444
rect 267476 156404 274876 156432
rect 267476 156392 267482 156404
rect 274870 156392 274876 156404
rect 274928 156392 274934 156444
rect 267050 155780 267056 155832
rect 267108 155820 267114 155832
rect 267694 155820 267700 155832
rect 267108 155792 267700 155820
rect 267108 155780 267114 155792
rect 267694 155780 267700 155792
rect 267752 155780 267758 155832
rect 361718 155712 361724 155764
rect 361776 155752 361782 155764
rect 412870 155752 412876 155764
rect 361776 155724 412876 155752
rect 361776 155712 361782 155724
rect 412870 155712 412876 155724
rect 412928 155712 412934 155764
rect 321054 155372 321060 155424
rect 321112 155412 321118 155424
rect 327218 155412 327224 155424
rect 321112 155384 327224 155412
rect 321112 155372 321118 155384
rect 327218 155372 327224 155384
rect 327276 155372 327282 155424
rect 173854 155100 173860 155152
rect 173912 155140 173918 155152
rect 182318 155140 182324 155152
rect 173912 155112 182324 155140
rect 173912 155100 173918 155112
rect 182318 155100 182324 155112
rect 182376 155100 182382 155152
rect 267786 155100 267792 155152
rect 267844 155140 267850 155152
rect 274962 155140 274968 155152
rect 267844 155112 274968 155140
rect 267844 155100 267850 155112
rect 274962 155100 274968 155112
rect 275020 155100 275026 155152
rect 321606 155100 321612 155152
rect 321664 155140 321670 155152
rect 321664 155112 321836 155140
rect 321664 155100 321670 155112
rect 79738 155032 79744 155084
rect 79796 155072 79802 155084
rect 87190 155072 87196 155084
rect 79796 155044 87196 155072
rect 79796 155032 79802 155044
rect 87190 155032 87196 155044
rect 87248 155032 87254 155084
rect 137606 155032 137612 155084
rect 137664 155072 137670 155084
rect 139630 155072 139636 155084
rect 137664 155044 139636 155072
rect 137664 155032 137670 155044
rect 139630 155032 139636 155044
rect 139688 155032 139694 155084
rect 173394 155032 173400 155084
rect 173452 155032 173458 155084
rect 173578 155032 173584 155084
rect 173636 155072 173642 155084
rect 181766 155072 181772 155084
rect 173636 155044 181772 155072
rect 173636 155032 173642 155044
rect 181766 155032 181772 155044
rect 181824 155032 181830 155084
rect 231446 155032 231452 155084
rect 231504 155072 231510 155084
rect 233470 155072 233476 155084
rect 231504 155044 233476 155072
rect 231504 155032 231510 155044
rect 233470 155032 233476 155044
rect 233528 155032 233534 155084
rect 266682 155032 266688 155084
rect 266740 155072 266746 155084
rect 275054 155072 275060 155084
rect 266740 155044 275060 155072
rect 266740 155032 266746 155044
rect 275054 155032 275060 155044
rect 275112 155032 275118 155084
rect 321808 155072 321836 155112
rect 328414 155072 328420 155084
rect 321808 155044 328420 155072
rect 328414 155032 328420 155044
rect 328472 155032 328478 155084
rect 173412 155004 173440 155032
rect 182318 155004 182324 155016
rect 173412 154976 182324 155004
rect 182318 154964 182324 154976
rect 182376 154964 182382 155016
rect 267602 154964 267608 155016
rect 267660 155004 267666 155016
rect 274870 155004 274876 155016
rect 267660 154976 274876 155004
rect 267660 154964 267666 154976
rect 274870 154964 274876 154976
rect 274928 154964 274934 155016
rect 173394 154896 173400 154948
rect 173452 154936 173458 154948
rect 181306 154936 181312 154948
rect 173452 154908 181312 154936
rect 173452 154896 173458 154908
rect 181306 154896 181312 154908
rect 181364 154896 181370 154948
rect 266590 154896 266596 154948
rect 266648 154936 266654 154948
rect 272846 154936 272852 154948
rect 266648 154908 272852 154936
rect 266648 154896 266654 154908
rect 272846 154896 272852 154908
rect 272904 154896 272910 154948
rect 12670 154760 12676 154812
rect 12728 154800 12734 154812
rect 16258 154800 16264 154812
rect 12728 154772 16264 154800
rect 12728 154760 12734 154772
rect 16258 154760 16264 154772
rect 16316 154760 16322 154812
rect 81762 154352 81768 154404
rect 81820 154392 81826 154404
rect 87190 154392 87196 154404
rect 81820 154364 87196 154392
rect 81820 154352 81826 154364
rect 87190 154352 87196 154364
rect 87248 154352 87254 154404
rect 320870 153740 320876 153792
rect 320928 153780 320934 153792
rect 328414 153780 328420 153792
rect 320928 153752 328420 153780
rect 320928 153740 320934 153752
rect 328414 153740 328420 153752
rect 328472 153740 328478 153792
rect 172934 153672 172940 153724
rect 172992 153712 172998 153724
rect 181398 153712 181404 153724
rect 172992 153684 181404 153712
rect 172992 153672 172998 153684
rect 181398 153672 181404 153684
rect 181456 153672 181462 153724
rect 267142 153672 267148 153724
rect 267200 153712 267206 153724
rect 274962 153712 274968 153724
rect 267200 153684 274968 153712
rect 267200 153672 267206 153684
rect 274962 153672 274968 153684
rect 275020 153672 275026 153724
rect 369814 153712 369820 153724
rect 369775 153684 369820 153712
rect 369814 153672 369820 153684
rect 369872 153672 369878 153724
rect 173210 153604 173216 153656
rect 173268 153644 173274 153656
rect 182318 153644 182324 153656
rect 173268 153616 182324 153644
rect 173268 153604 173274 153616
rect 182318 153604 182324 153616
rect 182376 153604 182382 153656
rect 267510 153604 267516 153656
rect 267568 153644 267574 153656
rect 274870 153644 274876 153656
rect 267568 153616 274876 153644
rect 267568 153604 267574 153616
rect 274870 153604 274876 153616
rect 274928 153604 274934 153656
rect 266590 153536 266596 153588
rect 266648 153576 266654 153588
rect 272938 153576 272944 153588
rect 266648 153548 272944 153576
rect 266648 153536 266654 153548
rect 272938 153536 272944 153548
rect 272996 153536 273002 153588
rect 81762 152992 81768 153044
rect 81820 153032 81826 153044
rect 87190 153032 87196 153044
rect 81820 153004 87196 153032
rect 81820 152992 81826 153004
rect 87190 152992 87196 153004
rect 87248 152992 87254 153044
rect 321606 152448 321612 152500
rect 321664 152488 321670 152500
rect 328230 152488 328236 152500
rect 321664 152460 328236 152488
rect 321664 152448 321670 152460
rect 328230 152448 328236 152460
rect 328288 152448 328294 152500
rect 79738 152380 79744 152432
rect 79796 152420 79802 152432
rect 87190 152420 87196 152432
rect 79796 152392 87196 152420
rect 79796 152380 79802 152392
rect 87190 152380 87196 152392
rect 87248 152380 87254 152432
rect 173578 152380 173584 152432
rect 173636 152420 173642 152432
rect 180294 152420 180300 152432
rect 173636 152392 180300 152420
rect 173636 152380 173642 152392
rect 180294 152380 180300 152392
rect 180352 152380 180358 152432
rect 320502 152380 320508 152432
rect 320560 152420 320566 152432
rect 323170 152420 323176 152432
rect 320560 152392 323176 152420
rect 320560 152380 320566 152392
rect 323170 152380 323176 152392
rect 323228 152380 323234 152432
rect 173302 152312 173308 152364
rect 173360 152352 173366 152364
rect 182318 152352 182324 152364
rect 173360 152324 182324 152352
rect 173360 152312 173366 152324
rect 182318 152312 182324 152324
rect 182376 152312 182382 152364
rect 267878 152312 267884 152364
rect 267936 152352 267942 152364
rect 274870 152352 274876 152364
rect 267936 152324 274876 152352
rect 267936 152312 267942 152324
rect 274870 152312 274876 152324
rect 274928 152312 274934 152364
rect 173670 151672 173676 151684
rect 173631 151644 173676 151672
rect 173670 151632 173676 151644
rect 173728 151632 173734 151684
rect 320778 151360 320784 151412
rect 320836 151400 320842 151412
rect 323262 151400 323268 151412
rect 320836 151372 323268 151400
rect 320836 151360 320842 151372
rect 323262 151360 323268 151372
rect 323320 151360 323326 151412
rect 131350 150884 131356 150936
rect 131408 150924 131414 150936
rect 140642 150924 140648 150936
rect 131408 150896 140648 150924
rect 131408 150884 131414 150896
rect 140642 150884 140648 150896
rect 140700 150884 140706 150936
rect 173762 150884 173768 150936
rect 173820 150924 173826 150936
rect 182318 150924 182324 150936
rect 173820 150896 182324 150924
rect 173820 150884 173826 150896
rect 182318 150884 182324 150896
rect 182376 150884 182382 150936
rect 225742 150884 225748 150936
rect 225800 150924 225806 150936
rect 233470 150924 233476 150936
rect 225800 150896 233476 150924
rect 225800 150884 225806 150896
rect 233470 150884 233476 150896
rect 233528 150884 233534 150936
rect 266590 150884 266596 150936
rect 266648 150924 266654 150936
rect 275790 150924 275796 150936
rect 266648 150896 275796 150924
rect 266648 150884 266654 150896
rect 275790 150884 275796 150896
rect 275848 150884 275854 150936
rect 323170 150884 323176 150936
rect 323228 150924 323234 150936
rect 328414 150924 328420 150936
rect 323228 150896 328420 150924
rect 323228 150884 323234 150896
rect 328414 150884 328420 150896
rect 328472 150884 328478 150936
rect 176246 150816 176252 150868
rect 176304 150856 176310 150868
rect 182226 150856 182232 150868
rect 176304 150828 182232 150856
rect 176304 150816 176310 150828
rect 182226 150816 182232 150828
rect 182284 150816 182290 150868
rect 225558 150816 225564 150868
rect 225616 150856 225622 150868
rect 232734 150856 232740 150868
rect 225616 150828 232740 150856
rect 225616 150816 225622 150828
rect 232734 150816 232740 150828
rect 232792 150816 232798 150868
rect 267694 150816 267700 150868
rect 267752 150856 267758 150868
rect 274870 150856 274876 150868
rect 267752 150828 274876 150856
rect 267752 150816 267758 150828
rect 274870 150816 274876 150828
rect 274928 150816 274934 150868
rect 173578 150748 173584 150800
rect 173636 150788 173642 150800
rect 179006 150788 179012 150800
rect 173636 150760 179012 150788
rect 173636 150748 173642 150760
rect 179006 150748 179012 150760
rect 179064 150748 179070 150800
rect 269994 150748 270000 150800
rect 270052 150788 270058 150800
rect 274962 150788 274968 150800
rect 270052 150760 274968 150788
rect 270052 150748 270058 150760
rect 274962 150748 274968 150760
rect 275020 150748 275026 150800
rect 173673 150655 173731 150661
rect 173673 150621 173685 150655
rect 173719 150652 173731 150655
rect 173946 150652 173952 150664
rect 173719 150624 173952 150652
rect 173719 150621 173731 150624
rect 173673 150615 173731 150621
rect 173946 150612 173952 150624
rect 174004 150612 174010 150664
rect 80106 149592 80112 149644
rect 80164 149632 80170 149644
rect 87190 149632 87196 149644
rect 80164 149604 87196 149632
rect 80164 149592 80170 149604
rect 87190 149592 87196 149604
rect 87248 149592 87254 149644
rect 321606 149592 321612 149644
rect 321664 149632 321670 149644
rect 327218 149632 327224 149644
rect 321664 149604 327224 149632
rect 321664 149592 321670 149604
rect 327218 149592 327224 149604
rect 327276 149592 327282 149644
rect 81762 149524 81768 149576
rect 81820 149564 81826 149576
rect 88110 149564 88116 149576
rect 81820 149536 88116 149564
rect 81820 149524 81826 149536
rect 88110 149524 88116 149536
rect 88168 149524 88174 149576
rect 131350 149524 131356 149576
rect 131408 149564 131414 149576
rect 140734 149564 140740 149576
rect 131408 149536 140740 149564
rect 131408 149524 131414 149536
rect 140734 149524 140740 149536
rect 140792 149524 140798 149576
rect 225926 149524 225932 149576
rect 225984 149564 225990 149576
rect 234114 149564 234120 149576
rect 225984 149536 234120 149564
rect 225984 149524 225990 149536
rect 234114 149524 234120 149536
rect 234172 149524 234178 149576
rect 266590 149524 266596 149576
rect 266648 149564 266654 149576
rect 272754 149564 272760 149576
rect 266648 149536 272760 149564
rect 266648 149524 266654 149536
rect 272754 149524 272760 149536
rect 272812 149524 272818 149576
rect 323262 149524 323268 149576
rect 323320 149564 323326 149576
rect 328414 149564 328420 149576
rect 323320 149536 328420 149564
rect 323320 149524 323326 149536
rect 328414 149524 328420 149536
rect 328472 149524 328478 149576
rect 271374 149456 271380 149508
rect 271432 149496 271438 149508
rect 274870 149496 274876 149508
rect 271432 149468 274876 149496
rect 271432 149456 271438 149468
rect 274870 149456 274876 149468
rect 274928 149456 274934 149508
rect 228686 149388 228692 149440
rect 228744 149428 228750 149440
rect 233470 149428 233476 149440
rect 228744 149400 233476 149428
rect 228744 149388 228750 149400
rect 233470 149388 233476 149400
rect 233528 149388 233534 149440
rect 226294 149116 226300 149168
rect 226352 149156 226358 149168
rect 231354 149156 231360 149168
rect 226352 149128 231360 149156
rect 226352 149116 226358 149128
rect 231354 149116 231360 149128
rect 231412 149116 231418 149168
rect 321606 148368 321612 148420
rect 321664 148408 321670 148420
rect 328322 148408 328328 148420
rect 321664 148380 328328 148408
rect 321664 148368 321670 148380
rect 328322 148368 328328 148380
rect 328380 148368 328386 148420
rect 321054 148232 321060 148284
rect 321112 148272 321118 148284
rect 328506 148272 328512 148284
rect 321112 148244 328512 148272
rect 321112 148232 321118 148244
rect 328506 148232 328512 148244
rect 328564 148232 328570 148284
rect 173578 148164 173584 148216
rect 173636 148204 173642 148216
rect 178914 148204 178920 148216
rect 173636 148176 178920 148204
rect 173636 148164 173642 148176
rect 178914 148164 178920 148176
rect 178972 148164 178978 148216
rect 227214 148164 227220 148216
rect 227272 148204 227278 148216
rect 233470 148204 233476 148216
rect 227272 148176 233476 148204
rect 227272 148164 227278 148176
rect 233470 148164 233476 148176
rect 233528 148164 233534 148216
rect 321790 148164 321796 148216
rect 321848 148204 321854 148216
rect 328414 148204 328420 148216
rect 321848 148176 328420 148204
rect 321848 148164 321854 148176
rect 328414 148164 328420 148176
rect 328472 148164 328478 148216
rect 427314 148164 427320 148216
rect 427372 148204 427378 148216
rect 429430 148204 429436 148216
rect 427372 148176 429436 148204
rect 427372 148164 427378 148176
rect 429430 148164 429436 148176
rect 429488 148164 429494 148216
rect 79738 148096 79744 148148
rect 79796 148136 79802 148148
rect 87098 148136 87104 148148
rect 79796 148108 87104 148136
rect 79796 148096 79802 148108
rect 87098 148096 87104 148108
rect 87156 148096 87162 148148
rect 369814 146804 369820 146856
rect 369872 146804 369878 146856
rect 132546 146736 132552 146788
rect 132604 146776 132610 146788
rect 139630 146776 139636 146788
rect 132604 146748 139636 146776
rect 132604 146736 132610 146748
rect 139630 146736 139636 146748
rect 139688 146736 139694 146788
rect 226386 146736 226392 146788
rect 226444 146776 226450 146788
rect 233470 146776 233476 146788
rect 226444 146748 233476 146776
rect 226444 146736 226450 146748
rect 233470 146736 233476 146748
rect 233528 146736 233534 146788
rect 267878 146736 267884 146788
rect 267936 146776 267942 146788
rect 275514 146776 275520 146788
rect 267936 146748 275520 146776
rect 267936 146736 267942 146748
rect 275514 146736 275520 146748
rect 275572 146736 275578 146788
rect 369832 146720 369860 146804
rect 369814 146668 369820 146720
rect 369872 146668 369878 146720
rect 79738 145376 79744 145428
rect 79796 145416 79802 145428
rect 87190 145416 87196 145428
rect 79796 145388 87196 145416
rect 79796 145376 79802 145388
rect 87190 145376 87196 145388
rect 87248 145376 87254 145428
rect 91698 145376 91704 145428
rect 91756 145416 91762 145428
rect 128130 145416 128136 145428
rect 91756 145388 128136 145416
rect 91756 145376 91762 145388
rect 128130 145376 128136 145388
rect 128188 145376 128194 145428
rect 132270 145376 132276 145428
rect 132328 145416 132334 145428
rect 139630 145416 139636 145428
rect 132328 145388 139636 145416
rect 132328 145376 132334 145388
rect 139630 145376 139636 145388
rect 139688 145376 139694 145428
rect 185630 145376 185636 145428
rect 185688 145416 185694 145428
rect 222154 145416 222160 145428
rect 185688 145388 222160 145416
rect 185688 145376 185694 145388
rect 222154 145376 222160 145388
rect 222212 145376 222218 145428
rect 226110 145376 226116 145428
rect 226168 145416 226174 145428
rect 233470 145416 233476 145428
rect 226168 145388 233476 145416
rect 226168 145376 226174 145388
rect 233470 145376 233476 145388
rect 233528 145376 233534 145428
rect 266774 145376 266780 145428
rect 266832 145416 266838 145428
rect 275606 145416 275612 145428
rect 266832 145388 275612 145416
rect 266832 145376 266838 145388
rect 275606 145376 275612 145388
rect 275664 145376 275670 145428
rect 279654 145376 279660 145428
rect 279712 145416 279718 145428
rect 322894 145416 322900 145428
rect 279712 145388 322900 145416
rect 279712 145376 279718 145388
rect 322894 145376 322900 145388
rect 322952 145376 322958 145428
rect 116078 144832 116084 144884
rect 116136 144872 116142 144884
rect 128038 144872 128044 144884
rect 116136 144844 128044 144872
rect 116136 144832 116142 144844
rect 128038 144832 128044 144844
rect 128096 144832 128102 144884
rect 211022 144832 211028 144884
rect 211080 144872 211086 144884
rect 230986 144872 230992 144884
rect 211080 144844 230992 144872
rect 211080 144832 211086 144844
rect 230986 144832 230992 144844
rect 231044 144832 231050 144884
rect 103658 144764 103664 144816
rect 103716 144804 103722 144816
rect 124266 144804 124272 144816
rect 103716 144776 124272 144804
rect 103716 144764 103722 144776
rect 124266 144764 124272 144776
rect 124324 144764 124330 144816
rect 197498 144764 197504 144816
rect 197556 144804 197562 144816
rect 218290 144804 218296 144816
rect 197556 144776 218296 144804
rect 197556 144764 197562 144776
rect 218290 144764 218296 144776
rect 218348 144764 218354 144816
rect 292718 144764 292724 144816
rect 292776 144804 292782 144816
rect 312314 144804 312320 144816
rect 292776 144776 312320 144804
rect 292776 144764 292782 144776
rect 312314 144764 312320 144776
rect 312372 144764 312378 144816
rect 91238 144696 91244 144748
rect 91296 144736 91302 144748
rect 120678 144736 120684 144748
rect 91296 144708 120684 144736
rect 91296 144696 91302 144708
rect 120678 144696 120684 144708
rect 120736 144696 120742 144748
rect 185078 144696 185084 144748
rect 185136 144736 185142 144748
rect 214702 144736 214708 144748
rect 185136 144708 214708 144736
rect 185136 144696 185142 144708
rect 214702 144696 214708 144708
rect 214760 144696 214766 144748
rect 280298 144696 280304 144748
rect 280356 144736 280362 144748
rect 308726 144736 308732 144748
rect 280356 144708 308732 144736
rect 280356 144696 280362 144708
rect 308726 144696 308732 144708
rect 308784 144696 308790 144748
rect 216174 144356 216180 144408
rect 216232 144396 216238 144408
rect 221970 144396 221976 144408
rect 216232 144368 221976 144396
rect 216232 144356 216238 144368
rect 221970 144356 221976 144368
rect 222028 144356 222034 144408
rect 310014 144152 310020 144204
rect 310072 144192 310078 144204
rect 315994 144192 316000 144204
rect 310072 144164 316000 144192
rect 310072 144152 310078 144164
rect 315994 144152 316000 144164
rect 316052 144152 316058 144204
rect 79738 144016 79744 144068
rect 79796 144056 79802 144068
rect 87282 144056 87288 144068
rect 79796 144028 87288 144056
rect 79796 144016 79802 144028
rect 87282 144016 87288 144028
rect 87340 144016 87346 144068
rect 132362 144016 132368 144068
rect 132420 144056 132426 144068
rect 139630 144056 139636 144068
rect 132420 144028 139636 144056
rect 132420 144016 132426 144028
rect 139630 144016 139636 144028
rect 139688 144016 139694 144068
rect 226478 144016 226484 144068
rect 226536 144056 226542 144068
rect 233470 144056 233476 144068
rect 226536 144028 233476 144056
rect 226536 144016 226542 144028
rect 233470 144016 233476 144028
rect 233528 144016 233534 144068
rect 303850 143404 303856 143456
rect 303908 143444 303914 143456
rect 305046 143444 305052 143456
rect 303908 143416 305052 143444
rect 303908 143404 303914 143416
rect 305046 143404 305052 143416
rect 305104 143444 305110 143456
rect 324642 143444 324648 143456
rect 305104 143416 324648 143444
rect 305104 143404 305110 143416
rect 324642 143404 324648 143416
rect 324700 143404 324706 143456
rect 297778 143336 297784 143388
rect 297836 143376 297842 143388
rect 325378 143376 325384 143388
rect 297836 143348 325384 143376
rect 297836 143336 297842 143348
rect 325378 143336 325384 143348
rect 325436 143336 325442 143388
rect 193453 142835 193511 142841
rect 193453 142801 193465 142835
rect 193499 142832 193511 142835
rect 200166 142832 200172 142844
rect 193499 142804 200172 142832
rect 193499 142801 193511 142804
rect 193453 142795 193511 142801
rect 200166 142792 200172 142804
rect 200224 142832 200230 142844
rect 203021 142835 203079 142841
rect 203021 142832 203033 142835
rect 200224 142804 203033 142832
rect 200224 142792 200230 142804
rect 203021 142801 203033 142804
rect 203067 142801 203079 142835
rect 203021 142795 203079 142801
rect 186737 142359 186795 142365
rect 186737 142356 186749 142359
rect 176816 142328 186749 142356
rect 176816 142288 176844 142328
rect 186737 142325 186749 142328
rect 186783 142325 186795 142359
rect 186737 142319 186795 142325
rect 167800 142260 176844 142288
rect 203021 142291 203079 142297
rect 167800 142232 167828 142260
rect 203021 142257 203033 142291
rect 203067 142288 203079 142291
rect 203067 142260 205824 142288
rect 203067 142257 203079 142260
rect 203021 142251 203079 142257
rect 167782 142180 167788 142232
rect 167840 142180 167846 142232
rect 186737 142223 186795 142229
rect 186737 142189 186749 142223
rect 186783 142220 186795 142223
rect 193453 142223 193511 142229
rect 193453 142220 193465 142223
rect 186783 142192 193465 142220
rect 186783 142189 186795 142192
rect 186737 142183 186795 142189
rect 193453 142189 193465 142192
rect 193499 142189 193511 142223
rect 193453 142183 193511 142189
rect 205796 142084 205824 142260
rect 231354 142084 231360 142096
rect 205796 142056 231360 142084
rect 231354 142044 231360 142056
rect 231412 142044 231418 142096
rect 290970 142044 290976 142096
rect 291028 142084 291034 142096
rect 325930 142084 325936 142096
rect 291028 142056 325936 142084
rect 291028 142044 291034 142056
rect 325930 142044 325936 142056
rect 325988 142044 325994 142096
rect 127210 141976 127216 142028
rect 127268 142016 127274 142028
rect 140366 142016 140372 142028
rect 127268 141988 140372 142016
rect 127268 141976 127274 141988
rect 140366 141976 140372 141988
rect 140424 141976 140430 142028
rect 173578 141976 173584 142028
rect 173636 142016 173642 142028
rect 219670 142016 219676 142028
rect 173636 141988 219676 142016
rect 173636 141976 173642 141988
rect 219670 141976 219676 141988
rect 219728 142016 219734 142028
rect 233470 142016 233476 142028
rect 219728 141988 233476 142016
rect 219728 141976 219734 141988
rect 233470 141976 233476 141988
rect 233528 141976 233534 142028
rect 267326 141976 267332 142028
rect 267384 142016 267390 142028
rect 316270 142016 316276 142028
rect 267384 141988 316276 142016
rect 267384 141976 267390 141988
rect 316270 141976 316276 141988
rect 316328 141976 316334 142028
rect 360430 141976 360436 142028
rect 360488 142016 360494 142028
rect 361074 142016 361080 142028
rect 360488 141988 361080 142016
rect 360488 141976 360494 141988
rect 361074 141976 361080 141988
rect 361132 141976 361138 142028
rect 77254 141296 77260 141348
rect 77312 141336 77318 141348
rect 127210 141336 127216 141348
rect 77312 141308 127216 141336
rect 77312 141296 77318 141308
rect 127210 141296 127216 141308
rect 127268 141296 127274 141348
rect 136962 141296 136968 141348
rect 137020 141336 137026 141348
rect 150394 141336 150400 141348
rect 137020 141308 150400 141336
rect 137020 141296 137026 141308
rect 150394 141296 150400 141308
rect 150452 141336 150458 141348
rect 167782 141336 167788 141348
rect 150452 141308 167788 141336
rect 150452 141296 150458 141308
rect 167782 141296 167788 141308
rect 167840 141296 167846 141348
rect 316270 141296 316276 141348
rect 316328 141336 316334 141348
rect 328414 141336 328420 141348
rect 316328 141308 328420 141336
rect 316328 141296 316334 141308
rect 328414 141296 328420 141308
rect 328472 141296 328478 141348
rect 77714 141228 77720 141280
rect 77772 141268 77778 141280
rect 113410 141268 113416 141280
rect 77772 141240 113416 141268
rect 77772 141228 77778 141240
rect 113410 141228 113416 141240
rect 113468 141268 113474 141280
rect 114698 141268 114704 141280
rect 113468 141240 114704 141268
rect 113468 141228 113474 141240
rect 114698 141228 114704 141240
rect 114756 141228 114762 141280
rect 82314 140752 82320 140804
rect 82372 140792 82378 140804
rect 85813 140795 85871 140801
rect 85813 140792 85825 140795
rect 82372 140764 85825 140792
rect 82372 140752 82378 140764
rect 85813 140761 85825 140764
rect 85859 140761 85871 140795
rect 85813 140755 85871 140761
rect 85813 140659 85871 140665
rect 85813 140625 85825 140659
rect 85859 140656 85871 140659
rect 85859 140628 95424 140656
rect 85859 140625 85871 140628
rect 85813 140619 85871 140625
rect 95396 140588 95424 140628
rect 114698 140616 114704 140668
rect 114756 140656 114762 140668
rect 137606 140656 137612 140668
rect 114756 140628 137612 140656
rect 114756 140616 114762 140628
rect 137606 140616 137612 140628
rect 137664 140616 137670 140668
rect 102278 140588 102284 140600
rect 95396 140560 102284 140588
rect 102278 140548 102284 140560
rect 102336 140548 102342 140600
rect 102370 140548 102376 140600
rect 102428 140588 102434 140600
rect 137330 140588 137336 140600
rect 102428 140560 137336 140588
rect 102428 140548 102434 140560
rect 137330 140548 137336 140560
rect 137388 140548 137394 140600
rect 207894 140548 207900 140600
rect 207952 140588 207958 140600
rect 231262 140588 231268 140600
rect 207952 140560 231268 140588
rect 207952 140548 207958 140560
rect 231262 140548 231268 140560
rect 231320 140548 231326 140600
rect 302010 140548 302016 140600
rect 302068 140588 302074 140600
rect 324826 140588 324832 140600
rect 302068 140560 324832 140588
rect 302068 140548 302074 140560
rect 324826 140548 324832 140560
rect 324884 140548 324890 140600
rect 141838 139868 141844 139920
rect 141896 139908 141902 139920
rect 152602 139908 152608 139920
rect 141896 139880 152608 139908
rect 141896 139868 141902 139880
rect 152602 139868 152608 139880
rect 152660 139868 152666 139920
rect 157941 139911 157999 139917
rect 157941 139877 157953 139911
rect 157987 139908 157999 139911
rect 166126 139908 166132 139920
rect 157987 139880 166132 139908
rect 157987 139877 157999 139880
rect 157941 139871 157999 139877
rect 166126 139868 166132 139880
rect 166184 139868 166190 139920
rect 255921 139911 255979 139917
rect 255921 139877 255933 139911
rect 255967 139908 255979 139911
rect 260150 139908 260156 139920
rect 255967 139880 260156 139908
rect 255967 139877 255979 139880
rect 255921 139871 255979 139877
rect 260150 139868 260156 139880
rect 260208 139868 260214 139920
rect 70446 139840 70452 139852
rect 65680 139812 70452 139840
rect 64834 139732 64840 139784
rect 64892 139772 64898 139784
rect 65680 139772 65708 139812
rect 70446 139800 70452 139812
rect 70504 139800 70510 139852
rect 150486 139800 150492 139852
rect 150544 139840 150550 139852
rect 162262 139840 162268 139852
rect 150544 139812 162268 139840
rect 150544 139800 150550 139812
rect 162262 139800 162268 139812
rect 162320 139800 162326 139852
rect 239542 139800 239548 139852
rect 239600 139840 239606 139852
rect 322802 139840 322808 139852
rect 239600 139812 322808 139840
rect 239600 139800 239606 139812
rect 322802 139800 322808 139812
rect 322860 139800 322866 139852
rect 74218 139772 74224 139784
rect 64892 139744 65708 139772
rect 65772 139744 74224 139772
rect 64892 139732 64898 139744
rect 62258 139664 62264 139716
rect 62316 139704 62322 139716
rect 65772 139704 65800 139744
rect 74218 139732 74224 139744
rect 74276 139732 74282 139784
rect 151774 139732 151780 139784
rect 151832 139772 151838 139784
rect 164562 139772 164568 139784
rect 151832 139744 164568 139772
rect 151832 139732 151838 139744
rect 164562 139732 164568 139744
rect 164620 139732 164626 139784
rect 247086 139732 247092 139784
rect 247144 139772 247150 139784
rect 259230 139772 259236 139784
rect 247144 139744 259236 139772
rect 247144 139732 247150 139744
rect 259230 139732 259236 139744
rect 259288 139732 259294 139784
rect 73114 139704 73120 139716
rect 62316 139676 65800 139704
rect 65864 139676 73120 139704
rect 62316 139664 62322 139676
rect 59498 139596 59504 139648
rect 59556 139636 59562 139648
rect 59556 139608 60372 139636
rect 59556 139596 59562 139608
rect 57658 139528 57664 139580
rect 57716 139568 57722 139580
rect 60234 139568 60240 139580
rect 57716 139540 60240 139568
rect 57716 139528 57722 139540
rect 60234 139528 60240 139540
rect 60292 139528 60298 139580
rect 60344 139568 60372 139608
rect 60878 139596 60884 139648
rect 60936 139636 60942 139648
rect 65864 139636 65892 139676
rect 73114 139664 73120 139676
rect 73172 139664 73178 139716
rect 154718 139664 154724 139716
rect 154776 139704 154782 139716
rect 167322 139704 167328 139716
rect 154776 139676 167328 139704
rect 154776 139664 154782 139676
rect 167322 139664 167328 139676
rect 167380 139664 167386 139716
rect 244326 139664 244332 139716
rect 244384 139704 244390 139716
rect 256286 139704 256292 139716
rect 244384 139676 256292 139704
rect 244384 139664 244390 139676
rect 256286 139664 256292 139676
rect 256344 139664 256350 139716
rect 60936 139608 65892 139636
rect 60936 139596 60942 139608
rect 65938 139596 65944 139648
rect 65996 139636 66002 139648
rect 70538 139636 70544 139648
rect 65996 139608 70544 139636
rect 65996 139596 66002 139608
rect 70538 139596 70544 139608
rect 70596 139596 70602 139648
rect 153338 139596 153344 139648
rect 153396 139636 153402 139648
rect 157941 139639 157999 139645
rect 157941 139636 157953 139639
rect 153396 139608 157953 139636
rect 153396 139596 153402 139608
rect 157941 139605 157953 139608
rect 157987 139605 157999 139639
rect 163274 139636 163280 139648
rect 157941 139599 157999 139605
rect 158048 139608 163280 139636
rect 71090 139568 71096 139580
rect 60344 139540 71096 139568
rect 71090 139528 71096 139540
rect 71148 139528 71154 139580
rect 150578 139528 150584 139580
rect 150636 139568 150642 139580
rect 158048 139568 158076 139608
rect 163274 139596 163280 139608
rect 163332 139596 163338 139648
rect 242486 139596 242492 139648
rect 242544 139636 242550 139648
rect 249110 139636 249116 139648
rect 242544 139608 249116 139636
rect 242544 139596 242550 139608
rect 249110 139596 249116 139608
rect 249168 139596 249174 139648
rect 251318 139596 251324 139648
rect 251376 139636 251382 139648
rect 264106 139636 264112 139648
rect 251376 139608 264112 139636
rect 251376 139596 251382 139608
rect 264106 139596 264112 139608
rect 264164 139596 264170 139648
rect 150636 139540 158076 139568
rect 150636 139528 150642 139540
rect 158122 139528 158128 139580
rect 158180 139568 158186 139580
rect 158858 139568 158864 139580
rect 158180 139540 158864 139568
rect 158180 139528 158186 139540
rect 158858 139528 158864 139540
rect 158916 139528 158922 139580
rect 160974 139528 160980 139580
rect 161032 139568 161038 139580
rect 161618 139568 161624 139580
rect 161032 139540 161624 139568
rect 161032 139528 161038 139540
rect 161618 139528 161624 139540
rect 161676 139528 161682 139580
rect 161986 139528 161992 139580
rect 162044 139568 162050 139580
rect 162998 139568 163004 139580
rect 162044 139540 163004 139568
rect 162044 139528 162050 139540
rect 162998 139528 163004 139540
rect 163056 139528 163062 139580
rect 249846 139528 249852 139580
rect 249904 139568 249910 139580
rect 253066 139568 253072 139580
rect 249904 139540 253072 139568
rect 249904 139528 249910 139540
rect 253066 139528 253072 139540
rect 253124 139528 253130 139580
rect 254909 139571 254967 139577
rect 254909 139568 254921 139571
rect 253176 139540 254921 139568
rect 63638 139460 63644 139512
rect 63696 139500 63702 139512
rect 75230 139500 75236 139512
rect 63696 139472 75236 139500
rect 63696 139460 63702 139472
rect 75230 139460 75236 139472
rect 75288 139460 75294 139512
rect 151866 139460 151872 139512
rect 151924 139500 151930 139512
rect 151924 139472 156144 139500
rect 151924 139460 151930 139472
rect 58118 139392 58124 139444
rect 58176 139432 58182 139444
rect 70078 139432 70084 139444
rect 58176 139404 70084 139432
rect 58176 139392 58182 139404
rect 70078 139392 70084 139404
rect 70136 139392 70142 139444
rect 155178 139392 155184 139444
rect 155236 139432 155242 139444
rect 156006 139432 156012 139444
rect 155236 139404 156012 139432
rect 155236 139392 155242 139404
rect 156006 139392 156012 139404
rect 156064 139392 156070 139444
rect 156116 139432 156144 139472
rect 157386 139460 157392 139512
rect 157444 139500 157450 139512
rect 169990 139500 169996 139512
rect 157444 139472 169996 139500
rect 157444 139460 157450 139472
rect 169990 139460 169996 139472
rect 170048 139460 170054 139512
rect 249202 139460 249208 139512
rect 249260 139500 249266 139512
rect 252054 139500 252060 139512
rect 249260 139472 252060 139500
rect 249260 139460 249266 139472
rect 252054 139460 252060 139472
rect 252112 139460 252118 139512
rect 165206 139432 165212 139444
rect 156116 139404 165212 139432
rect 165206 139392 165212 139404
rect 165264 139392 165270 139444
rect 248558 139392 248564 139444
rect 248616 139432 248622 139444
rect 253176 139432 253204 139540
rect 254909 139537 254921 139540
rect 254955 139537 254967 139571
rect 254909 139531 254967 139537
rect 254998 139528 255004 139580
rect 255056 139568 255062 139580
rect 257482 139568 257488 139580
rect 255056 139540 257488 139568
rect 255056 139528 255062 139540
rect 257482 139528 257488 139540
rect 257540 139528 257546 139580
rect 333382 139528 333388 139580
rect 333440 139568 333446 139580
rect 334118 139568 334124 139580
rect 333440 139540 334124 139568
rect 333440 139528 333446 139540
rect 334118 139528 334124 139540
rect 334176 139528 334182 139580
rect 334394 139528 334400 139580
rect 334452 139568 334458 139580
rect 335498 139568 335504 139580
rect 334452 139540 335504 139568
rect 334452 139528 334458 139540
rect 335498 139528 335504 139540
rect 335556 139528 335562 139580
rect 253253 139503 253311 139509
rect 253253 139469 253265 139503
rect 253299 139500 253311 139503
rect 255921 139503 255979 139509
rect 255921 139500 255933 139503
rect 253299 139472 255933 139500
rect 253299 139469 253311 139472
rect 253253 139463 253311 139469
rect 255921 139469 255933 139472
rect 255967 139469 255979 139503
rect 255921 139463 255979 139469
rect 256010 139460 256016 139512
rect 256068 139500 256074 139512
rect 258678 139500 258684 139512
rect 256068 139472 258684 139500
rect 256068 139460 256074 139472
rect 258678 139460 258684 139472
rect 258736 139460 258742 139512
rect 248616 139404 253204 139432
rect 253345 139435 253403 139441
rect 248616 139392 248622 139404
rect 253345 139401 253357 139435
rect 253391 139432 253403 139435
rect 258310 139432 258316 139444
rect 253391 139404 258316 139432
rect 253391 139401 253403 139404
rect 253345 139395 253403 139401
rect 258310 139392 258316 139404
rect 258368 139392 258374 139444
rect 56738 139324 56744 139376
rect 56796 139364 56802 139376
rect 67962 139364 67968 139376
rect 56796 139336 67968 139364
rect 56796 139324 56802 139336
rect 67962 139324 67968 139336
rect 68020 139324 68026 139376
rect 154626 139324 154632 139376
rect 154684 139364 154690 139376
rect 168058 139364 168064 139376
rect 154684 139336 168064 139364
rect 154684 139324 154690 139336
rect 168058 139324 168064 139336
rect 168116 139324 168122 139376
rect 244418 139324 244424 139376
rect 244476 139364 244482 139376
rect 257298 139364 257304 139376
rect 244476 139336 257304 139364
rect 244476 139324 244482 139336
rect 257298 139324 257304 139336
rect 257356 139324 257362 139376
rect 55358 139256 55364 139308
rect 55416 139296 55422 139308
rect 66950 139296 66956 139308
rect 55416 139268 66956 139296
rect 55416 139256 55422 139268
rect 66950 139256 66956 139268
rect 67008 139256 67014 139308
rect 155914 139256 155920 139308
rect 155972 139296 155978 139308
rect 169070 139296 169076 139308
rect 155972 139268 169076 139296
rect 155972 139256 155978 139268
rect 169070 139256 169076 139268
rect 169128 139256 169134 139308
rect 241474 139256 241480 139308
rect 241532 139296 241538 139308
rect 249662 139296 249668 139308
rect 241532 139268 249668 139296
rect 241532 139256 241538 139268
rect 249662 139256 249668 139268
rect 249720 139256 249726 139308
rect 249846 139256 249852 139308
rect 249904 139296 249910 139308
rect 254817 139299 254875 139305
rect 254817 139296 254829 139299
rect 249904 139268 254829 139296
rect 249904 139256 249910 139268
rect 254817 139265 254829 139268
rect 254863 139265 254875 139299
rect 254817 139259 254875 139265
rect 254909 139299 254967 139305
rect 254909 139265 254921 139299
rect 254955 139296 254967 139299
rect 261162 139296 261168 139308
rect 254955 139268 261168 139296
rect 254955 139265 254967 139268
rect 254909 139259 254967 139265
rect 261162 139256 261168 139268
rect 261220 139256 261226 139308
rect 338534 139256 338540 139308
rect 338592 139296 338598 139308
rect 339546 139296 339552 139308
rect 338592 139268 339552 139296
rect 338592 139256 338598 139268
rect 339546 139256 339552 139268
rect 339604 139256 339610 139308
rect 60786 139188 60792 139240
rect 60844 139228 60850 139240
rect 72102 139228 72108 139240
rect 60844 139200 72108 139228
rect 60844 139188 60850 139200
rect 72102 139188 72108 139200
rect 72160 139188 72166 139240
rect 74310 139188 74316 139240
rect 74368 139228 74374 139240
rect 116170 139228 116176 139240
rect 74368 139200 116176 139228
rect 74368 139188 74374 139200
rect 116170 139188 116176 139200
rect 116228 139228 116234 139240
rect 136870 139228 136876 139240
rect 116228 139200 136876 139228
rect 116228 139188 116234 139200
rect 136870 139188 136876 139200
rect 136928 139188 136934 139240
rect 144598 139188 144604 139240
rect 144656 139228 144662 139240
rect 170634 139228 170640 139240
rect 144656 139200 170640 139228
rect 144656 139188 144662 139200
rect 170634 139188 170640 139200
rect 170692 139188 170698 139240
rect 238622 139188 238628 139240
rect 238680 139228 238686 139240
rect 264474 139228 264480 139240
rect 238680 139200 264480 139228
rect 238680 139188 238686 139200
rect 264474 139188 264480 139200
rect 264532 139188 264538 139240
rect 63822 139120 63828 139172
rect 63880 139160 63886 139172
rect 68606 139160 68612 139172
rect 63880 139132 68612 139160
rect 63880 139120 63886 139132
rect 68606 139120 68612 139132
rect 68664 139120 68670 139172
rect 249938 139120 249944 139172
rect 249996 139160 250002 139172
rect 254817 139163 254875 139169
rect 249996 139132 254768 139160
rect 249996 139120 250002 139132
rect 252146 139052 252152 139104
rect 252204 139092 252210 139104
rect 254170 139092 254176 139104
rect 252204 139064 254176 139092
rect 252204 139052 252210 139064
rect 254170 139052 254176 139064
rect 254228 139052 254234 139104
rect 254740 139092 254768 139132
rect 254817 139129 254829 139163
rect 254863 139160 254875 139163
rect 263094 139160 263100 139172
rect 254863 139132 263100 139160
rect 254863 139129 254875 139132
rect 254817 139123 254875 139129
rect 263094 139120 263100 139132
rect 263152 139120 263158 139172
rect 262082 139092 262088 139104
rect 254740 139064 262088 139092
rect 262082 139052 262088 139064
rect 262140 139052 262146 139104
rect 251134 138984 251140 139036
rect 251192 139024 251198 139036
rect 253986 139024 253992 139036
rect 251192 138996 253992 139024
rect 251192 138984 251198 138996
rect 253986 138984 253992 138996
rect 254044 138984 254050 139036
rect 247178 138916 247184 138968
rect 247236 138956 247242 138968
rect 253253 138959 253311 138965
rect 253253 138956 253265 138959
rect 247236 138928 253265 138956
rect 247236 138916 247242 138928
rect 253253 138925 253265 138928
rect 253299 138925 253311 138959
rect 253253 138919 253311 138925
rect 62810 138848 62816 138900
rect 62868 138888 62874 138900
rect 62868 138860 63132 138888
rect 62868 138848 62874 138860
rect 59682 138780 59688 138832
rect 59740 138820 59746 138832
rect 62994 138820 63000 138832
rect 59740 138792 63000 138820
rect 59740 138780 59746 138792
rect 62994 138780 63000 138792
rect 63052 138780 63058 138832
rect 63104 138820 63132 138860
rect 245798 138848 245804 138900
rect 245856 138888 245862 138900
rect 253345 138891 253403 138897
rect 253345 138888 253357 138891
rect 245856 138860 253357 138888
rect 245856 138848 245862 138860
rect 253345 138857 253357 138860
rect 253391 138857 253403 138891
rect 253345 138851 253403 138857
rect 340926 138848 340932 138900
rect 340984 138888 340990 138900
rect 340984 138860 341984 138888
rect 340984 138848 340990 138860
rect 67686 138820 67692 138832
rect 63104 138792 67692 138820
rect 67686 138780 67692 138792
rect 67744 138780 67750 138832
rect 253894 138780 253900 138832
rect 253952 138820 253958 138832
rect 256654 138820 256660 138832
rect 253952 138792 256660 138820
rect 253952 138780 253958 138792
rect 256654 138780 256660 138792
rect 256712 138780 256718 138832
rect 341018 138780 341024 138832
rect 341076 138820 341082 138832
rect 341757 138823 341815 138829
rect 341757 138820 341769 138823
rect 341076 138792 341769 138820
rect 341076 138780 341082 138792
rect 341757 138789 341769 138792
rect 341803 138789 341815 138823
rect 341956 138820 341984 138860
rect 345894 138848 345900 138900
rect 345952 138888 345958 138900
rect 349942 138888 349948 138900
rect 345952 138860 349948 138888
rect 345952 138848 345958 138860
rect 349942 138848 349948 138860
rect 350000 138848 350006 138900
rect 347918 138820 347924 138832
rect 341956 138792 347924 138820
rect 341757 138783 341815 138789
rect 347918 138780 347924 138792
rect 347976 138780 347982 138832
rect 61798 138712 61804 138764
rect 61856 138752 61862 138764
rect 65754 138752 65760 138764
rect 61856 138724 65760 138752
rect 61856 138712 61862 138724
rect 65754 138712 65760 138724
rect 65812 138712 65818 138764
rect 145242 138712 145248 138764
rect 145300 138752 145306 138764
rect 365214 138752 365220 138764
rect 145300 138724 365220 138752
rect 145300 138712 145306 138724
rect 365214 138712 365220 138724
rect 365272 138712 365278 138764
rect 58670 138644 58676 138696
rect 58728 138684 58734 138696
rect 63086 138684 63092 138696
rect 58728 138656 63092 138684
rect 58728 138644 58734 138656
rect 63086 138644 63092 138656
rect 63144 138644 63150 138696
rect 338074 138644 338080 138696
rect 338132 138684 338138 138696
rect 341662 138684 341668 138696
rect 338132 138656 341668 138684
rect 338132 138644 338138 138656
rect 341662 138644 341668 138656
rect 341720 138644 341726 138696
rect 341757 138687 341815 138693
rect 341757 138653 341769 138687
rect 341803 138684 341815 138687
rect 346814 138684 346820 138696
rect 341803 138656 346820 138684
rect 341803 138653 341815 138656
rect 341757 138647 341815 138653
rect 346814 138644 346820 138656
rect 346872 138644 346878 138696
rect 60694 138576 60700 138628
rect 60752 138616 60758 138628
rect 63178 138616 63184 138628
rect 60752 138588 63184 138616
rect 60752 138576 60758 138588
rect 63178 138576 63184 138588
rect 63236 138576 63242 138628
rect 252698 138576 252704 138628
rect 252756 138616 252762 138628
rect 254814 138616 254820 138628
rect 252756 138588 254820 138616
rect 252756 138576 252762 138588
rect 254814 138576 254820 138588
rect 254872 138576 254878 138628
rect 338258 138576 338264 138628
rect 338316 138616 338322 138628
rect 342674 138616 342680 138628
rect 338316 138588 342680 138616
rect 338316 138576 338322 138588
rect 342674 138576 342680 138588
rect 342732 138576 342738 138628
rect 344514 138576 344520 138628
rect 344572 138616 344578 138628
rect 345802 138616 345808 138628
rect 344572 138588 345808 138616
rect 344572 138576 344578 138588
rect 345802 138576 345808 138588
rect 345860 138576 345866 138628
rect 345986 138576 345992 138628
rect 346044 138616 346050 138628
rect 348930 138616 348936 138628
rect 346044 138588 348936 138616
rect 346044 138576 346050 138588
rect 348930 138576 348936 138588
rect 348988 138576 348994 138628
rect 287198 137828 287204 137880
rect 287256 137868 287262 137880
rect 324734 137868 324740 137880
rect 287256 137840 324740 137868
rect 287256 137828 287262 137840
rect 324734 137828 324740 137840
rect 324792 137828 324798 137880
rect 343962 137828 343968 137880
rect 344020 137868 344026 137880
rect 360890 137868 360896 137880
rect 344020 137840 360896 137868
rect 344020 137828 344026 137840
rect 360890 137828 360896 137840
rect 360948 137828 360954 137880
rect 325930 137148 325936 137200
rect 325988 137188 325994 137200
rect 326574 137188 326580 137200
rect 325988 137160 326580 137188
rect 325988 137148 325994 137160
rect 326574 137148 326580 137160
rect 326632 137188 326638 137200
rect 343962 137188 343968 137200
rect 326632 137160 343968 137188
rect 326632 137148 326638 137160
rect 343962 137148 343968 137160
rect 344020 137148 344026 137200
rect 74126 137080 74132 137132
rect 74184 137120 74190 137132
rect 74402 137120 74408 137132
rect 74184 137092 74408 137120
rect 74184 137080 74190 137092
rect 74402 137080 74408 137092
rect 74460 137080 74466 137132
rect 427498 137080 427504 137132
rect 427556 137120 427562 137132
rect 429430 137120 429436 137132
rect 427556 137092 429436 137120
rect 427556 137080 427562 137092
rect 429430 137080 429436 137092
rect 429488 137080 429494 137132
rect 210010 136400 210016 136452
rect 210068 136440 210074 136452
rect 216174 136440 216180 136452
rect 210068 136412 216180 136440
rect 210068 136400 210074 136412
rect 216174 136400 216180 136412
rect 216232 136400 216238 136452
rect 304034 136400 304040 136452
rect 304092 136440 304098 136452
rect 310014 136440 310020 136452
rect 304092 136412 310020 136440
rect 304092 136400 304098 136412
rect 310014 136400 310020 136412
rect 310072 136400 310078 136452
rect 291522 136264 291528 136316
rect 291580 136304 291586 136316
rect 292718 136304 292724 136316
rect 291580 136276 292724 136304
rect 291580 136264 291586 136276
rect 292718 136264 292724 136276
rect 292776 136264 292782 136316
rect 279102 136128 279108 136180
rect 279160 136168 279166 136180
rect 280298 136168 280304 136180
rect 279160 136140 280304 136168
rect 279160 136128 279166 136140
rect 280298 136128 280304 136140
rect 280356 136128 280362 136180
rect 346538 135040 346544 135092
rect 346596 135080 346602 135092
rect 360614 135080 360620 135092
rect 346596 135052 360620 135080
rect 346596 135040 346602 135052
rect 360614 135040 360620 135052
rect 360672 135040 360678 135092
rect 325378 134428 325384 134480
rect 325436 134468 325442 134480
rect 345710 134468 345716 134480
rect 325436 134440 345716 134468
rect 325436 134428 325442 134440
rect 345710 134428 345716 134440
rect 345768 134468 345774 134480
rect 346538 134468 346544 134480
rect 345768 134440 346544 134468
rect 345768 134428 345774 134440
rect 346538 134428 346544 134440
rect 346596 134428 346602 134480
rect 51586 134360 51592 134412
rect 51644 134400 51650 134412
rect 51862 134400 51868 134412
rect 51644 134372 51868 134400
rect 51644 134360 51650 134372
rect 51862 134360 51868 134372
rect 51920 134360 51926 134412
rect 236230 134400 236236 134412
rect 236191 134372 236236 134400
rect 236230 134360 236236 134372
rect 236288 134360 236294 134412
rect 357673 134403 357731 134409
rect 357673 134369 357685 134403
rect 357719 134400 357731 134403
rect 360706 134400 360712 134412
rect 357719 134372 360712 134400
rect 357719 134369 357731 134372
rect 357673 134363 357731 134369
rect 360706 134360 360712 134372
rect 360764 134360 360770 134412
rect 346538 133748 346544 133800
rect 346596 133788 346602 133800
rect 360522 133788 360528 133800
rect 346596 133760 360528 133788
rect 346596 133748 346602 133760
rect 360522 133748 360528 133760
rect 360580 133748 360586 133800
rect 283150 133680 283156 133732
rect 283208 133720 283214 133732
rect 324550 133720 324556 133732
rect 283208 133692 324556 133720
rect 283208 133680 283214 133692
rect 324550 133680 324556 133692
rect 324608 133680 324614 133732
rect 343318 133680 343324 133732
rect 343376 133720 343382 133732
rect 360982 133720 360988 133732
rect 343376 133692 360988 133720
rect 343376 133680 343382 133692
rect 360982 133680 360988 133692
rect 361040 133680 361046 133732
rect 324550 133068 324556 133120
rect 324608 133108 324614 133120
rect 343318 133108 343324 133120
rect 324608 133080 343324 133108
rect 324608 133068 324614 133080
rect 343318 133068 343324 133080
rect 343376 133068 343382 133120
rect 324826 133000 324832 133052
rect 324884 133040 324890 133052
rect 325470 133040 325476 133052
rect 324884 133012 325476 133040
rect 324884 133000 324890 133012
rect 325470 133000 325476 133012
rect 325528 133040 325534 133052
rect 346354 133040 346360 133052
rect 325528 133012 346360 133040
rect 325528 133000 325534 133012
rect 346354 133000 346360 133012
rect 346412 133040 346418 133052
rect 346538 133040 346544 133052
rect 346412 133012 346544 133040
rect 346412 133000 346418 133012
rect 346538 133000 346544 133012
rect 346596 133000 346602 133052
rect 13038 132932 13044 132984
rect 13096 132972 13102 132984
rect 16442 132972 16448 132984
rect 13096 132944 16448 132972
rect 13096 132932 13102 132944
rect 16442 132932 16448 132944
rect 16500 132932 16506 132984
rect 369630 132972 369636 132984
rect 369591 132944 369636 132972
rect 369630 132932 369636 132944
rect 369688 132932 369694 132984
rect 369538 132904 369544 132916
rect 369499 132876 369544 132904
rect 369538 132864 369544 132876
rect 369596 132864 369602 132916
rect 230986 132796 230992 132848
rect 231044 132836 231050 132848
rect 231446 132836 231452 132848
rect 231044 132808 231452 132836
rect 231044 132796 231050 132808
rect 231446 132796 231452 132808
rect 231504 132796 231510 132848
rect 136870 132320 136876 132372
rect 136928 132360 136934 132372
rect 137330 132360 137336 132372
rect 136928 132332 137336 132360
rect 136928 132320 136934 132332
rect 137330 132320 137336 132332
rect 137388 132320 137394 132372
rect 343962 132320 343968 132372
rect 344020 132360 344026 132372
rect 360798 132360 360804 132372
rect 344020 132332 360804 132360
rect 344020 132320 344026 132332
rect 360798 132320 360804 132332
rect 360856 132320 360862 132372
rect 324642 132252 324648 132304
rect 324700 132292 324706 132304
rect 346998 132292 347004 132304
rect 324700 132264 347004 132292
rect 324700 132252 324706 132264
rect 346998 132252 347004 132264
rect 347056 132252 347062 132304
rect 354910 132252 354916 132304
rect 354968 132292 354974 132304
rect 355830 132292 355836 132304
rect 354968 132264 355836 132292
rect 354968 132252 354974 132264
rect 355830 132252 355836 132264
rect 355888 132252 355894 132304
rect 339454 131708 339460 131760
rect 339512 131748 339518 131760
rect 339730 131748 339736 131760
rect 339512 131720 339736 131748
rect 339512 131708 339518 131720
rect 339730 131708 339736 131720
rect 339788 131708 339794 131760
rect 324734 131640 324740 131692
rect 324792 131680 324798 131692
rect 325562 131680 325568 131692
rect 324792 131652 325568 131680
rect 324792 131640 324798 131652
rect 325562 131640 325568 131652
rect 325620 131680 325626 131692
rect 343962 131680 343968 131692
rect 325620 131652 343968 131680
rect 325620 131640 325626 131652
rect 343962 131640 343968 131652
rect 344020 131640 344026 131692
rect 346998 131640 347004 131692
rect 347056 131680 347062 131692
rect 360430 131680 360436 131692
rect 347056 131652 360436 131680
rect 347056 131640 347062 131652
rect 360430 131640 360436 131652
rect 360488 131680 360494 131692
rect 361074 131680 361080 131692
rect 360488 131652 361080 131680
rect 360488 131640 360494 131652
rect 361074 131640 361080 131652
rect 361132 131640 361138 131692
rect 59682 131572 59688 131624
rect 59740 131612 59746 131624
rect 60786 131612 60792 131624
rect 59740 131584 60792 131612
rect 59740 131572 59746 131584
rect 60786 131572 60792 131584
rect 60844 131572 60850 131624
rect 245338 131572 245344 131624
rect 245396 131612 245402 131624
rect 245798 131612 245804 131624
rect 245396 131584 245804 131612
rect 245396 131572 245402 131584
rect 245798 131572 245804 131584
rect 245856 131572 245862 131624
rect 248006 131572 248012 131624
rect 248064 131612 248070 131624
rect 248558 131612 248564 131624
rect 248064 131584 248564 131612
rect 248064 131572 248070 131584
rect 248558 131572 248564 131584
rect 248616 131572 248622 131624
rect 250674 131572 250680 131624
rect 250732 131612 250738 131624
rect 251318 131612 251324 131624
rect 250732 131584 251324 131612
rect 250732 131572 250738 131584
rect 251318 131572 251324 131584
rect 251376 131572 251382 131624
rect 63178 131504 63184 131556
rect 63236 131544 63242 131556
rect 65938 131544 65944 131556
rect 63236 131516 65944 131544
rect 63236 131504 63242 131516
rect 65938 131504 65944 131516
rect 65996 131504 66002 131556
rect 339546 131504 339552 131556
rect 339604 131544 339610 131556
rect 350954 131544 350960 131556
rect 339604 131516 350960 131544
rect 339604 131504 339610 131516
rect 350954 131504 350960 131516
rect 351012 131504 351018 131556
rect 338166 131436 338172 131488
rect 338224 131476 338230 131488
rect 350402 131476 350408 131488
rect 338224 131448 350408 131476
rect 338224 131436 338230 131448
rect 350402 131436 350408 131448
rect 350460 131436 350466 131488
rect 161618 131368 161624 131420
rect 161676 131408 161682 131420
rect 163458 131408 163464 131420
rect 161676 131380 163464 131408
rect 161676 131368 161682 131380
rect 163458 131368 163464 131380
rect 163516 131368 163522 131420
rect 248466 131368 248472 131420
rect 248524 131408 248530 131420
rect 250950 131408 250956 131420
rect 248524 131380 250956 131408
rect 248524 131368 248530 131380
rect 250950 131368 250956 131380
rect 251008 131368 251014 131420
rect 342398 131368 342404 131420
rect 342456 131408 342462 131420
rect 345894 131408 345900 131420
rect 342456 131380 345900 131408
rect 342456 131368 342462 131380
rect 345894 131368 345900 131380
rect 345952 131368 345958 131420
rect 158766 131300 158772 131352
rect 158824 131340 158830 131352
rect 161710 131340 161716 131352
rect 158824 131312 161716 131340
rect 158824 131300 158830 131312
rect 161710 131300 161716 131312
rect 161768 131300 161774 131352
rect 231354 131300 231360 131352
rect 231412 131340 231418 131352
rect 322710 131340 322716 131352
rect 231412 131312 322716 131340
rect 231412 131300 231418 131312
rect 322710 131300 322716 131312
rect 322768 131300 322774 131352
rect 335498 131300 335504 131352
rect 335556 131340 335562 131352
rect 348562 131340 348568 131352
rect 335556 131312 348568 131340
rect 335556 131300 335562 131312
rect 348562 131300 348568 131312
rect 348620 131300 348626 131352
rect 258954 131232 258960 131284
rect 259012 131272 259018 131284
rect 368802 131272 368808 131284
rect 259012 131244 368808 131272
rect 259012 131232 259018 131244
rect 368802 131232 368808 131244
rect 368860 131232 368866 131284
rect 336878 131164 336884 131216
rect 336936 131204 336942 131216
rect 349758 131204 349764 131216
rect 336936 131176 349764 131204
rect 336936 131164 336942 131176
rect 349758 131164 349764 131176
rect 349816 131164 349822 131216
rect 334118 131096 334124 131148
rect 334176 131136 334182 131148
rect 348010 131136 348016 131148
rect 334176 131108 348016 131136
rect 334176 131096 334182 131108
rect 348010 131096 348016 131108
rect 348068 131096 348074 131148
rect 332738 131028 332744 131080
rect 332796 131068 332802 131080
rect 340009 131071 340067 131077
rect 340009 131068 340021 131071
rect 332796 131040 340021 131068
rect 332796 131028 332802 131040
rect 340009 131037 340021 131040
rect 340055 131037 340067 131071
rect 340009 131031 340067 131037
rect 340834 131028 340840 131080
rect 340892 131068 340898 131080
rect 352242 131068 352248 131080
rect 340892 131040 352248 131068
rect 340892 131028 340898 131040
rect 352242 131028 352248 131040
rect 352300 131028 352306 131080
rect 335406 130960 335412 131012
rect 335464 131000 335470 131012
rect 349390 131000 349396 131012
rect 335464 130972 349396 131000
rect 335464 130960 335470 130972
rect 349390 130960 349396 130972
rect 349448 130960 349454 131012
rect 57014 130892 57020 130944
rect 57072 130932 57078 130944
rect 68054 130932 68060 130944
rect 57072 130904 68060 130932
rect 57072 130892 57078 130904
rect 68054 130892 68060 130904
rect 68112 130892 68118 130944
rect 345253 130935 345311 130941
rect 345253 130901 345265 130935
rect 345299 130932 345311 130935
rect 361166 130932 361172 130944
rect 345299 130904 361172 130932
rect 345299 130901 345311 130904
rect 345253 130895 345311 130901
rect 361166 130892 361172 130904
rect 361224 130892 361230 130944
rect 340009 130867 340067 130873
rect 340009 130833 340021 130867
rect 340055 130864 340067 130867
rect 347274 130864 347280 130876
rect 340055 130836 347280 130864
rect 340055 130833 340067 130836
rect 340009 130827 340067 130833
rect 347274 130824 347280 130836
rect 347332 130824 347338 130876
rect 342490 130796 342496 130808
rect 337356 130768 342496 130796
rect 160238 130688 160244 130740
rect 160296 130728 160302 130740
rect 162630 130728 162636 130740
rect 160296 130700 162636 130728
rect 160296 130688 160302 130700
rect 162630 130688 162636 130700
rect 162688 130688 162694 130740
rect 246258 130552 246264 130604
rect 246316 130592 246322 130604
rect 247086 130592 247092 130604
rect 246316 130564 247092 130592
rect 246316 130552 246322 130564
rect 247086 130552 247092 130564
rect 247144 130552 247150 130604
rect 60234 130484 60240 130536
rect 60292 130524 60298 130536
rect 63270 130524 63276 130536
rect 60292 130496 63276 130524
rect 60292 130484 60298 130496
rect 63270 130484 63276 130496
rect 63328 130484 63334 130536
rect 156098 130484 156104 130536
rect 156156 130524 156162 130536
rect 159042 130524 159048 130536
rect 156156 130496 159048 130524
rect 156156 130484 156162 130496
rect 159042 130484 159048 130496
rect 159100 130484 159106 130536
rect 62994 130416 63000 130468
rect 63052 130456 63058 130468
rect 65018 130456 65024 130468
rect 63052 130428 65024 130456
rect 63052 130416 63058 130428
rect 65018 130416 65024 130428
rect 65076 130416 65082 130468
rect 156006 130416 156012 130468
rect 156064 130456 156070 130468
rect 158122 130456 158128 130468
rect 156064 130428 158128 130456
rect 156064 130416 156070 130428
rect 158122 130416 158128 130428
rect 158180 130416 158186 130468
rect 62350 130348 62356 130400
rect 62408 130388 62414 130400
rect 63638 130388 63644 130400
rect 62408 130360 63644 130388
rect 62408 130348 62414 130360
rect 63638 130348 63644 130360
rect 63696 130348 63702 130400
rect 154534 130348 154540 130400
rect 154592 130388 154598 130400
rect 157294 130388 157300 130400
rect 154592 130360 157300 130388
rect 154592 130348 154598 130360
rect 157294 130348 157300 130360
rect 157352 130348 157358 130400
rect 157478 130348 157484 130400
rect 157536 130388 157542 130400
rect 159962 130388 159968 130400
rect 157536 130360 159968 130388
rect 157536 130348 157542 130360
rect 159962 130348 159968 130360
rect 160020 130348 160026 130400
rect 325286 130348 325292 130400
rect 325344 130388 325350 130400
rect 337356 130388 337384 130768
rect 342490 130756 342496 130768
rect 342548 130796 342554 130808
rect 345253 130799 345311 130805
rect 345253 130796 345265 130799
rect 342548 130768 345265 130796
rect 342548 130756 342554 130768
rect 345253 130765 345265 130768
rect 345299 130765 345311 130799
rect 345253 130759 345311 130765
rect 339638 130688 339644 130740
rect 339696 130728 339702 130740
rect 351598 130728 351604 130740
rect 339696 130700 351604 130728
rect 339696 130688 339702 130700
rect 351598 130688 351604 130700
rect 351656 130688 351662 130740
rect 341754 130620 341760 130672
rect 341812 130660 341818 130672
rect 345986 130660 345992 130672
rect 341812 130632 345992 130660
rect 341812 130620 341818 130632
rect 345986 130620 345992 130632
rect 346044 130620 346050 130672
rect 339546 130552 339552 130604
rect 339604 130592 339610 130604
rect 344514 130592 344520 130604
rect 339604 130564 344520 130592
rect 339604 130552 339610 130564
rect 344514 130552 344520 130564
rect 344572 130552 344578 130604
rect 339362 130484 339368 130536
rect 339420 130524 339426 130536
rect 343870 130524 343876 130536
rect 339420 130496 343876 130524
rect 339420 130484 339426 130496
rect 343870 130484 343876 130496
rect 343928 130484 343934 130536
rect 338718 130416 338724 130468
rect 338776 130456 338782 130468
rect 342766 130456 342772 130468
rect 338776 130428 342772 130456
rect 338776 130416 338782 130428
rect 342766 130416 342772 130428
rect 342824 130416 342830 130468
rect 325344 130360 337384 130388
rect 325344 130348 325350 130360
rect 61430 130280 61436 130332
rect 61488 130320 61494 130332
rect 62258 130320 62264 130332
rect 61488 130292 62264 130320
rect 61488 130280 61494 130292
rect 62258 130280 62264 130292
rect 62316 130280 62322 130332
rect 63086 130280 63092 130332
rect 63144 130320 63150 130332
rect 64098 130320 64104 130332
rect 63144 130292 64104 130320
rect 63144 130280 63150 130292
rect 64098 130280 64104 130292
rect 64156 130280 64162 130332
rect 65754 130280 65760 130332
rect 65812 130320 65818 130332
rect 66766 130320 66772 130332
rect 65812 130292 66772 130320
rect 65812 130280 65818 130292
rect 66766 130280 66772 130292
rect 66824 130280 66830 130332
rect 149290 130280 149296 130332
rect 149348 130320 149354 130332
rect 150486 130320 150492 130332
rect 149348 130292 150492 130320
rect 149348 130280 149354 130292
rect 150486 130280 150492 130292
rect 150544 130280 150550 130332
rect 151038 130280 151044 130332
rect 151096 130320 151102 130332
rect 151774 130320 151780 130332
rect 151096 130292 151780 130320
rect 151096 130280 151102 130292
rect 151774 130280 151780 130292
rect 151832 130280 151838 130332
rect 153706 130280 153712 130332
rect 153764 130320 153770 130332
rect 154718 130320 154724 130332
rect 153764 130292 154724 130320
rect 153764 130280 153770 130292
rect 154718 130280 154724 130292
rect 154776 130280 154782 130332
rect 156374 130280 156380 130332
rect 156432 130320 156438 130332
rect 157386 130320 157392 130332
rect 156432 130292 157392 130320
rect 156432 130280 156438 130292
rect 157386 130280 157392 130292
rect 157444 130280 157450 130332
rect 158858 130280 158864 130332
rect 158916 130320 158922 130332
rect 160790 130320 160796 130332
rect 158916 130292 160796 130320
rect 158916 130280 158922 130292
rect 160790 130280 160796 130292
rect 160848 130280 160854 130332
rect 162998 130280 163004 130332
rect 163056 130320 163062 130332
rect 164378 130320 164384 130332
rect 163056 130292 164384 130320
rect 163056 130280 163062 130292
rect 164378 130280 164384 130292
rect 164436 130280 164442 130332
rect 243590 130280 243596 130332
rect 243648 130320 243654 130332
rect 244326 130320 244332 130332
rect 243648 130292 244332 130320
rect 243648 130280 243654 130292
rect 244326 130280 244332 130292
rect 244384 130280 244390 130332
rect 248926 130280 248932 130332
rect 248984 130320 248990 130332
rect 249938 130320 249944 130332
rect 248984 130292 249944 130320
rect 248984 130280 248990 130292
rect 249938 130280 249944 130292
rect 249996 130280 250002 130332
rect 254814 130280 254820 130332
rect 254872 130320 254878 130332
rect 255550 130320 255556 130332
rect 254872 130292 255556 130320
rect 254872 130280 254878 130292
rect 255550 130280 255556 130292
rect 255608 130280 255614 130332
rect 323170 130280 323176 130332
rect 323228 130320 323234 130332
rect 323228 130292 337476 130320
rect 323228 130280 323234 130292
rect 231262 130212 231268 130264
rect 231320 130252 231326 130264
rect 246442 130252 246448 130264
rect 231320 130224 246448 130252
rect 231320 130212 231326 130224
rect 246442 130212 246448 130224
rect 246500 130212 246506 130264
rect 337448 130252 337476 130292
rect 337522 130280 337528 130332
rect 337580 130320 337586 130332
rect 338074 130320 338080 130332
rect 337580 130292 338080 130320
rect 337580 130280 337586 130292
rect 338074 130280 338080 130292
rect 338132 130280 338138 130332
rect 338184 130292 340512 130320
rect 338184 130252 338212 130292
rect 337448 130224 338212 130252
rect 340484 130252 340512 130292
rect 340558 130280 340564 130332
rect 340616 130320 340622 130332
rect 341018 130320 341024 130332
rect 340616 130292 341024 130320
rect 340616 130280 340622 130292
rect 341018 130280 341024 130292
rect 341076 130280 341082 130332
rect 357673 130323 357731 130329
rect 357673 130320 357685 130323
rect 345222 130292 357685 130320
rect 344882 130252 344888 130264
rect 340484 130224 344888 130252
rect 344882 130212 344888 130224
rect 344940 130252 344946 130264
rect 345222 130252 345250 130292
rect 357673 130289 357685 130292
rect 357719 130289 357731 130323
rect 357673 130283 357731 130289
rect 344940 130224 345250 130252
rect 344940 130212 344946 130224
rect 73850 127492 73856 127544
rect 73908 127492 73914 127544
rect 74218 127492 74224 127544
rect 74276 127532 74282 127544
rect 74402 127532 74408 127544
rect 74276 127504 74408 127532
rect 74276 127492 74282 127504
rect 74402 127492 74408 127504
rect 74460 127492 74466 127544
rect 137054 127492 137060 127544
rect 137112 127532 137118 127544
rect 137238 127532 137244 127544
rect 137112 127504 137244 127532
rect 137112 127492 137118 127504
rect 137238 127492 137244 127504
rect 137296 127492 137302 127544
rect 73868 127396 73896 127492
rect 74034 127396 74040 127408
rect 73868 127368 74040 127396
rect 74034 127356 74040 127368
rect 74092 127356 74098 127408
rect 38798 126744 38804 126796
rect 38856 126784 38862 126796
rect 54070 126784 54076 126796
rect 38856 126756 54076 126784
rect 38856 126744 38862 126756
rect 54070 126744 54076 126756
rect 54128 126744 54134 126796
rect 357670 126744 357676 126796
rect 357728 126784 357734 126796
rect 405970 126784 405976 126796
rect 357728 126756 405976 126784
rect 357728 126744 357734 126756
rect 405970 126744 405976 126756
rect 406028 126744 406034 126796
rect 38246 126064 38252 126116
rect 38304 126104 38310 126116
rect 51218 126104 51224 126116
rect 38304 126076 51224 126104
rect 38304 126064 38310 126076
rect 51218 126064 51224 126076
rect 51276 126064 51282 126116
rect 356198 126064 356204 126116
rect 356256 126104 356262 126116
rect 405970 126104 405976 126116
rect 356256 126076 405976 126104
rect 356256 126064 356262 126076
rect 405970 126064 405976 126076
rect 406028 126064 406034 126116
rect 76886 125452 76892 125504
rect 76944 125492 76950 125504
rect 81670 125492 81676 125504
rect 76944 125464 81676 125492
rect 76944 125452 76950 125464
rect 81670 125452 81676 125464
rect 81728 125452 81734 125504
rect 169990 125384 169996 125436
rect 170048 125424 170054 125436
rect 170634 125424 170640 125436
rect 170048 125396 170640 125424
rect 170048 125384 170054 125396
rect 170634 125384 170640 125396
rect 170692 125424 170698 125436
rect 175510 125424 175516 125436
rect 170692 125396 175516 125424
rect 170692 125384 170698 125396
rect 175510 125384 175516 125396
rect 175568 125384 175574 125436
rect 263830 125248 263836 125300
rect 263888 125288 263894 125300
rect 264474 125288 264480 125300
rect 263888 125260 264480 125288
rect 263888 125248 263894 125260
rect 264474 125248 264480 125260
rect 264532 125288 264538 125300
rect 270362 125288 270368 125300
rect 264532 125260 270368 125288
rect 264532 125248 264538 125260
rect 270362 125248 270368 125260
rect 270420 125248 270426 125300
rect 76150 125044 76156 125096
rect 76208 125084 76214 125096
rect 76886 125084 76892 125096
rect 76208 125056 76892 125084
rect 76208 125044 76214 125056
rect 76886 125044 76892 125056
rect 76944 125044 76950 125096
rect 369538 124880 369544 124892
rect 369499 124852 369544 124880
rect 369538 124840 369544 124852
rect 369596 124840 369602 124892
rect 236230 124812 236236 124824
rect 236191 124784 236236 124812
rect 236230 124772 236236 124784
rect 236288 124772 236294 124824
rect 357673 124815 357731 124821
rect 357673 124781 357685 124815
rect 357719 124812 357731 124815
rect 360614 124812 360620 124824
rect 357719 124784 360620 124812
rect 357719 124781 357731 124784
rect 357673 124775 357731 124781
rect 360614 124772 360620 124784
rect 360672 124772 360678 124824
rect 74034 124744 74040 124756
rect 73995 124716 74040 124744
rect 74034 124704 74040 124716
rect 74092 124704 74098 124756
rect 369630 124676 369636 124688
rect 369591 124648 369636 124676
rect 369630 124636 369636 124648
rect 369688 124636 369694 124688
rect 38798 122596 38804 122648
rect 38856 122636 38862 122648
rect 53150 122636 53156 122648
rect 38856 122608 53156 122636
rect 38856 122596 38862 122608
rect 53150 122596 53156 122608
rect 53208 122596 53214 122648
rect 356290 122596 356296 122648
rect 356348 122636 356354 122648
rect 405970 122636 405976 122648
rect 356348 122608 405976 122636
rect 356348 122596 356354 122608
rect 405970 122596 405976 122608
rect 406028 122596 406034 122648
rect 137606 121984 137612 122036
rect 137664 122024 137670 122036
rect 144230 122024 144236 122036
rect 137664 121996 144236 122024
rect 137664 121984 137670 121996
rect 144230 121984 144236 121996
rect 144288 121984 144294 122036
rect 231446 121984 231452 122036
rect 231504 122024 231510 122036
rect 240370 122024 240376 122036
rect 231504 121996 240376 122024
rect 231504 121984 231510 121996
rect 240370 121984 240376 121996
rect 240428 121984 240434 122036
rect 325378 121984 325384 122036
rect 325436 122024 325442 122036
rect 334210 122024 334216 122036
rect 325436 121996 334216 122024
rect 325436 121984 325442 121996
rect 334210 121984 334216 121996
rect 334268 121984 334274 122036
rect 13222 121916 13228 121968
rect 13280 121956 13286 121968
rect 16534 121956 16540 121968
rect 13280 121928 16540 121956
rect 13280 121916 13286 121928
rect 16534 121916 16540 121928
rect 16592 121916 16598 121968
rect 38798 120556 38804 120608
rect 38856 120596 38862 120608
rect 52598 120596 52604 120608
rect 38856 120568 52604 120596
rect 38856 120556 38862 120568
rect 52598 120556 52604 120568
rect 52656 120556 52662 120608
rect 356198 120556 356204 120608
rect 356256 120596 356262 120608
rect 405970 120596 405976 120608
rect 356256 120568 405976 120596
rect 356256 120556 356262 120568
rect 405970 120556 405976 120568
rect 406028 120556 406034 120608
rect 324550 119876 324556 119928
rect 324608 119916 324614 119928
rect 326574 119916 326580 119928
rect 324608 119888 326580 119916
rect 324608 119876 324614 119888
rect 326574 119876 326580 119888
rect 326632 119876 326638 119928
rect 261162 117904 261168 117956
rect 261220 117944 261226 117956
rect 268614 117944 268620 117956
rect 261220 117916 268620 117944
rect 261220 117904 261226 117916
rect 268614 117904 268620 117916
rect 268672 117904 268678 117956
rect 167874 117836 167880 117888
rect 167932 117876 167938 117888
rect 174866 117876 174872 117888
rect 167932 117848 174872 117876
rect 167932 117836 167938 117848
rect 174866 117836 174872 117848
rect 174924 117836 174930 117888
rect 360338 117876 360344 117888
rect 360264 117848 360344 117876
rect 360264 117820 360292 117848
rect 360338 117836 360344 117848
rect 360396 117836 360402 117888
rect 360430 117836 360436 117888
rect 360488 117876 360494 117888
rect 360614 117876 360620 117888
rect 360488 117848 360620 117876
rect 360488 117836 360494 117848
rect 360614 117836 360620 117848
rect 360672 117836 360678 117888
rect 73482 117768 73488 117820
rect 73540 117808 73546 117820
rect 74218 117808 74224 117820
rect 73540 117780 74224 117808
rect 73540 117768 73546 117780
rect 74218 117768 74224 117780
rect 74276 117768 74282 117820
rect 360246 117768 360252 117820
rect 360304 117768 360310 117820
rect 74034 117740 74040 117752
rect 73995 117712 74040 117740
rect 74034 117700 74040 117712
rect 74092 117700 74098 117752
rect 38246 117088 38252 117140
rect 38304 117128 38310 117140
rect 54070 117128 54076 117140
rect 38304 117100 54076 117128
rect 38304 117088 38310 117100
rect 54070 117088 54076 117100
rect 54128 117088 54134 117140
rect 354910 117088 354916 117140
rect 354968 117128 354974 117140
rect 405970 117128 405976 117140
rect 354968 117100 405976 117128
rect 354968 117088 354974 117100
rect 405970 117088 405976 117100
rect 406028 117088 406034 117140
rect 38798 115048 38804 115100
rect 38856 115088 38862 115100
rect 51218 115088 51224 115100
rect 38856 115060 51224 115088
rect 38856 115048 38862 115060
rect 51218 115048 51224 115060
rect 51276 115048 51282 115100
rect 51681 115091 51739 115097
rect 51681 115057 51693 115091
rect 51727 115088 51739 115091
rect 51862 115088 51868 115100
rect 51727 115060 51868 115088
rect 51727 115057 51739 115060
rect 51681 115051 51739 115057
rect 51862 115048 51868 115060
rect 51920 115048 51926 115100
rect 74034 115048 74040 115100
rect 74092 115088 74098 115100
rect 74218 115088 74224 115100
rect 74092 115060 74224 115088
rect 74092 115048 74098 115060
rect 74218 115048 74224 115060
rect 74276 115048 74282 115100
rect 236230 115088 236236 115100
rect 236191 115060 236236 115088
rect 236230 115048 236236 115060
rect 236288 115048 236294 115100
rect 356198 115048 356204 115100
rect 356256 115088 356262 115100
rect 360249 115091 360307 115097
rect 360249 115088 360261 115091
rect 356256 115060 360261 115088
rect 356256 115048 356262 115060
rect 360249 115057 360261 115060
rect 360295 115057 360307 115091
rect 360249 115051 360307 115057
rect 360433 115091 360491 115097
rect 360433 115057 360445 115091
rect 360479 115088 360491 115091
rect 369817 115091 369875 115097
rect 369817 115088 369829 115091
rect 360479 115060 369829 115088
rect 360479 115057 360491 115060
rect 360433 115051 360491 115057
rect 369817 115057 369829 115060
rect 369863 115057 369875 115091
rect 405970 115088 405976 115100
rect 369817 115051 369875 115057
rect 370200 115060 405976 115088
rect 370001 115023 370059 115029
rect 370001 114989 370013 115023
rect 370047 115020 370059 115023
rect 370200 115020 370228 115060
rect 405970 115048 405976 115060
rect 406028 115048 406034 115100
rect 370047 114992 370228 115020
rect 370047 114989 370059 114992
rect 370001 114983 370059 114989
rect 38798 112940 38804 112992
rect 38856 112980 38862 112992
rect 52138 112980 52144 112992
rect 38856 112952 52144 112980
rect 38856 112940 38862 112952
rect 52138 112940 52144 112952
rect 52196 112940 52202 112992
rect 136870 112940 136876 112992
rect 136928 112980 136934 112992
rect 147358 112980 147364 112992
rect 136928 112952 147364 112980
rect 136928 112940 136934 112952
rect 147358 112940 147364 112952
rect 147416 112940 147422 112992
rect 355002 112940 355008 112992
rect 355060 112980 355066 112992
rect 405970 112980 405976 112992
rect 355060 112952 405976 112980
rect 355060 112940 355066 112952
rect 405970 112940 405976 112952
rect 406028 112940 406034 112992
rect 427406 112056 427412 112108
rect 427464 112096 427470 112108
rect 429430 112096 429436 112108
rect 427464 112068 429436 112096
rect 427464 112056 427470 112068
rect 429430 112056 429436 112068
rect 429488 112056 429494 112108
rect 12854 111512 12860 111564
rect 12912 111552 12918 111564
rect 16350 111552 16356 111564
rect 12912 111524 16356 111552
rect 12912 111512 12918 111524
rect 16350 111512 16356 111524
rect 16408 111512 16414 111564
rect 38246 110900 38252 110952
rect 38304 110940 38310 110952
rect 52598 110940 52604 110952
rect 38304 110912 52604 110940
rect 38304 110900 38310 110912
rect 52598 110900 52604 110912
rect 52656 110900 52662 110952
rect 136870 110900 136876 110952
rect 136928 110940 136934 110952
rect 145334 110940 145340 110952
rect 136928 110912 145340 110940
rect 136928 110900 136934 110912
rect 145334 110900 145340 110912
rect 145392 110900 145398 110952
rect 231630 110900 231636 110952
rect 231688 110940 231694 110952
rect 239082 110940 239088 110952
rect 231688 110912 239088 110940
rect 231688 110900 231694 110912
rect 239082 110900 239088 110912
rect 239140 110940 239146 110952
rect 240094 110940 240100 110952
rect 239140 110912 240100 110940
rect 239140 110900 239146 110912
rect 240094 110900 240100 110912
rect 240152 110900 240158 110952
rect 356198 110900 356204 110952
rect 356256 110940 356262 110952
rect 406062 110940 406068 110952
rect 356256 110912 406068 110940
rect 356256 110900 356262 110912
rect 406062 110900 406068 110912
rect 406120 110900 406126 110952
rect 74402 109472 74408 109524
rect 74460 109512 74466 109524
rect 81670 109512 81676 109524
rect 74460 109484 81676 109512
rect 74460 109472 74466 109484
rect 81670 109472 81676 109484
rect 81728 109472 81734 109524
rect 137698 108180 137704 108232
rect 137756 108220 137762 108232
rect 143954 108220 143960 108232
rect 137756 108192 143960 108220
rect 137756 108180 137762 108192
rect 143954 108180 143960 108192
rect 144012 108180 144018 108232
rect 231538 108180 231544 108232
rect 231596 108220 231602 108232
rect 240370 108220 240376 108232
rect 231596 108192 240376 108220
rect 231596 108180 231602 108192
rect 240370 108180 240376 108192
rect 240428 108180 240434 108232
rect 325470 108180 325476 108232
rect 325528 108220 325534 108232
rect 334210 108220 334216 108232
rect 325528 108192 334216 108220
rect 325528 108180 325534 108192
rect 334210 108180 334216 108192
rect 334268 108180 334274 108232
rect 51678 108016 51684 108028
rect 51639 107988 51684 108016
rect 51678 107976 51684 107988
rect 51736 107976 51742 108028
rect 38798 107432 38804 107484
rect 38856 107472 38862 107484
rect 51678 107472 51684 107484
rect 38856 107444 51684 107472
rect 38856 107432 38862 107444
rect 51678 107432 51684 107444
rect 51736 107432 51742 107484
rect 353530 107432 353536 107484
rect 353588 107472 353594 107484
rect 405970 107472 405976 107484
rect 353588 107444 405976 107472
rect 353588 107432 353594 107444
rect 405970 107432 405976 107444
rect 406028 107432 406034 107484
rect 13314 105460 13320 105512
rect 13372 105500 13378 105512
rect 18098 105500 18104 105512
rect 13372 105472 18104 105500
rect 13372 105460 13378 105472
rect 18098 105460 18104 105472
rect 18156 105460 18162 105512
rect 236230 105500 236236 105512
rect 236191 105472 236236 105500
rect 236230 105460 236236 105472
rect 236288 105460 236294 105512
rect 427682 105460 427688 105512
rect 427740 105500 427746 105512
rect 430074 105500 430080 105512
rect 427740 105472 430080 105500
rect 427740 105460 427746 105472
rect 430074 105460 430080 105472
rect 430132 105460 430138 105512
rect 38798 105392 38804 105444
rect 38856 105432 38862 105444
rect 52598 105432 52604 105444
rect 38856 105404 52604 105432
rect 38856 105392 38862 105404
rect 52598 105392 52604 105404
rect 52656 105392 52662 105444
rect 356198 105392 356204 105444
rect 356256 105432 356262 105444
rect 405970 105432 405976 105444
rect 356256 105404 405976 105432
rect 356256 105392 356262 105404
rect 405970 105392 405976 105404
rect 406028 105392 406034 105444
rect 352702 101924 352708 101976
rect 352760 101964 352766 101976
rect 405970 101964 405976 101976
rect 352760 101936 405976 101964
rect 352760 101924 352766 101936
rect 405970 101924 405976 101936
rect 406028 101924 406034 101976
rect 50022 101516 50028 101568
rect 50080 101556 50086 101568
rect 51310 101556 51316 101568
rect 50080 101528 51316 101556
rect 50080 101516 50086 101528
rect 51310 101516 51316 101528
rect 51368 101516 51374 101568
rect 38614 101312 38620 101364
rect 38672 101352 38678 101364
rect 50022 101352 50028 101364
rect 38672 101324 50028 101352
rect 38672 101312 38678 101324
rect 50022 101312 50028 101324
rect 50080 101312 50086 101364
rect 12854 100768 12860 100820
rect 12912 100808 12918 100820
rect 16166 100808 16172 100820
rect 12912 100780 16172 100808
rect 12912 100768 12918 100780
rect 16166 100768 16172 100780
rect 16224 100768 16230 100820
rect 38798 100564 38804 100616
rect 38856 100604 38862 100616
rect 52598 100604 52604 100616
rect 38856 100576 52604 100604
rect 38856 100564 38862 100576
rect 52598 100564 52604 100576
rect 52656 100564 52662 100616
rect 356198 100564 356204 100616
rect 356256 100604 356262 100616
rect 405970 100604 405976 100616
rect 356256 100576 405976 100604
rect 356256 100564 356262 100576
rect 405970 100564 405976 100576
rect 406028 100564 406034 100616
rect 13406 99884 13412 99936
rect 13464 99924 13470 99936
rect 17454 99924 17460 99936
rect 13464 99896 17460 99924
rect 13464 99884 13470 99896
rect 17454 99884 17460 99896
rect 17512 99884 17518 99936
rect 168242 98592 168248 98644
rect 168300 98632 168306 98644
rect 169254 98632 169260 98644
rect 168300 98604 169260 98632
rect 168300 98592 168306 98604
rect 169254 98592 169260 98604
rect 169312 98592 169318 98644
rect 427682 98524 427688 98576
rect 427740 98564 427746 98576
rect 429430 98564 429436 98576
rect 427740 98536 429436 98564
rect 427740 98524 427746 98536
rect 429430 98524 429436 98536
rect 429488 98524 429494 98576
rect 73942 98388 73948 98440
rect 74000 98428 74006 98440
rect 74218 98428 74224 98440
rect 74000 98400 74224 98428
rect 74000 98388 74006 98400
rect 74218 98388 74224 98400
rect 74276 98388 74282 98440
rect 38798 97776 38804 97828
rect 38856 97816 38862 97828
rect 49930 97816 49936 97828
rect 38856 97788 49936 97816
rect 38856 97776 38862 97788
rect 49930 97776 49936 97788
rect 49988 97776 49994 97828
rect 352794 97776 352800 97828
rect 352852 97816 352858 97828
rect 405970 97816 405976 97828
rect 352852 97788 405976 97816
rect 352852 97776 352858 97788
rect 405970 97776 405976 97788
rect 406028 97776 406034 97828
rect 13498 95804 13504 95856
rect 13556 95844 13562 95856
rect 18098 95844 18104 95856
rect 13556 95816 18104 95844
rect 13556 95804 13562 95816
rect 18098 95804 18104 95816
rect 18156 95804 18162 95856
rect 427222 95804 427228 95856
rect 427280 95844 427286 95856
rect 430166 95844 430172 95856
rect 427280 95816 430172 95844
rect 427280 95804 427286 95816
rect 430166 95804 430172 95816
rect 430224 95804 430230 95856
rect 38062 95736 38068 95788
rect 38120 95776 38126 95788
rect 52598 95776 52604 95788
rect 38120 95748 52604 95776
rect 38120 95736 38126 95748
rect 52598 95736 52604 95748
rect 52656 95736 52662 95788
rect 236230 95776 236236 95788
rect 236143 95748 236236 95776
rect 236230 95736 236236 95748
rect 236288 95776 236294 95788
rect 237242 95776 237248 95788
rect 236288 95748 237248 95776
rect 236288 95736 236294 95748
rect 237242 95736 237248 95748
rect 237300 95736 237306 95788
rect 356198 95736 356204 95788
rect 356256 95776 356262 95788
rect 405970 95776 405976 95788
rect 356256 95748 405976 95776
rect 356256 95736 356262 95748
rect 405970 95736 405976 95748
rect 406028 95736 406034 95788
rect 231814 94988 231820 95040
rect 231872 95028 231878 95040
rect 236233 95031 236291 95037
rect 236233 95028 236245 95031
rect 231872 95000 236245 95028
rect 231872 94988 231878 95000
rect 236233 94997 236245 95000
rect 236279 94997 236291 95031
rect 236233 94991 236291 94997
rect 325838 94648 325844 94700
rect 325896 94688 325902 94700
rect 330070 94688 330076 94700
rect 325896 94660 330076 94688
rect 325896 94648 325902 94660
rect 330070 94648 330076 94660
rect 330128 94648 330134 94700
rect 138158 94376 138164 94428
rect 138216 94416 138222 94428
rect 142390 94416 142396 94428
rect 138216 94388 142396 94416
rect 138216 94376 138222 94388
rect 142390 94376 142396 94388
rect 142448 94376 142454 94428
rect 232734 94376 232740 94428
rect 232792 94416 232798 94428
rect 240370 94416 240376 94428
rect 232792 94388 240376 94416
rect 232792 94376 232798 94388
rect 240370 94376 240376 94388
rect 240428 94376 240434 94428
rect 326666 94376 326672 94428
rect 326724 94416 326730 94428
rect 334210 94416 334216 94428
rect 326724 94388 334216 94416
rect 326724 94376 326730 94388
rect 334210 94376 334216 94388
rect 334268 94376 334274 94428
rect 72562 94308 72568 94360
rect 72620 94348 72626 94360
rect 73942 94348 73948 94360
rect 72620 94320 73948 94348
rect 72620 94308 72626 94320
rect 73942 94308 73948 94320
rect 74000 94308 74006 94360
rect 74678 94308 74684 94360
rect 74736 94348 74742 94360
rect 78174 94348 78180 94360
rect 74736 94320 78180 94348
rect 74736 94308 74742 94320
rect 78174 94308 78180 94320
rect 78232 94308 78238 94360
rect 73574 93832 73580 93884
rect 73632 93872 73638 93884
rect 73758 93872 73764 93884
rect 73632 93844 73764 93872
rect 73632 93832 73638 93844
rect 73758 93832 73764 93844
rect 73816 93832 73822 93884
rect 73390 93696 73396 93748
rect 73448 93736 73454 93748
rect 73574 93736 73580 93748
rect 73448 93708 73580 93736
rect 73448 93696 73454 93708
rect 73574 93696 73580 93708
rect 73632 93696 73638 93748
rect 74126 92948 74132 93000
rect 74184 92988 74190 93000
rect 81670 92988 81676 93000
rect 74184 92960 81676 92988
rect 74184 92948 74190 92960
rect 81670 92948 81676 92960
rect 81728 92948 81734 93000
rect 169254 92948 169260 93000
rect 169312 92988 169318 93000
rect 175510 92988 175516 93000
rect 169312 92960 175516 92988
rect 169312 92948 169318 92960
rect 175510 92948 175516 92960
rect 175568 92948 175574 93000
rect 263094 92948 263100 93000
rect 263152 92988 263158 93000
rect 270362 92988 270368 93000
rect 263152 92960 270368 92988
rect 263152 92948 263158 92960
rect 270362 92948 270368 92960
rect 270420 92948 270426 93000
rect 37602 92268 37608 92320
rect 37660 92308 37666 92320
rect 48550 92308 48556 92320
rect 37660 92280 48556 92308
rect 37660 92268 37666 92280
rect 48550 92268 48556 92280
rect 48608 92268 48614 92320
rect 352794 92268 352800 92320
rect 352852 92308 352858 92320
rect 405970 92308 405976 92320
rect 352852 92280 405976 92308
rect 352852 92268 352858 92280
rect 405970 92268 405976 92280
rect 406028 92268 406034 92320
rect 73850 91248 73856 91300
rect 73908 91288 73914 91300
rect 76794 91288 76800 91300
rect 73908 91260 76800 91288
rect 73908 91248 73914 91260
rect 76794 91248 76800 91260
rect 76852 91248 76858 91300
rect 17270 90268 17276 90280
rect 14068 90240 17276 90268
rect 13222 90160 13228 90212
rect 13280 90200 13286 90212
rect 14068 90200 14096 90240
rect 17270 90228 17276 90240
rect 17328 90228 17334 90280
rect 52598 90268 52604 90280
rect 48476 90240 52604 90268
rect 13280 90172 14096 90200
rect 13280 90160 13286 90172
rect 38798 90160 38804 90212
rect 38856 90200 38862 90212
rect 48476 90200 48504 90240
rect 52598 90228 52604 90240
rect 52656 90228 52662 90280
rect 38856 90172 48504 90200
rect 38856 90160 38862 90172
rect 356198 90160 356204 90212
rect 356256 90200 356262 90212
rect 405970 90200 405976 90212
rect 356256 90172 405976 90200
rect 356256 90160 356262 90172
rect 405970 90160 405976 90172
rect 406028 90160 406034 90212
rect 369722 88800 369728 88852
rect 369780 88840 369786 88852
rect 369906 88840 369912 88852
rect 369780 88812 369912 88840
rect 369780 88800 369786 88812
rect 369906 88800 369912 88812
rect 369964 88800 369970 88852
rect 251318 87508 251324 87560
rect 251376 87548 251382 87560
rect 260058 87548 260064 87560
rect 251376 87520 260064 87548
rect 251376 87508 251382 87520
rect 260058 87508 260064 87520
rect 260116 87508 260122 87560
rect 23894 87440 23900 87492
rect 23952 87480 23958 87492
rect 72562 87480 72568 87492
rect 23952 87452 72568 87480
rect 23952 87440 23958 87452
rect 72562 87440 72568 87452
rect 72620 87440 72626 87492
rect 154718 87480 154724 87492
rect 154677 87452 154724 87480
rect 154718 87440 154724 87452
rect 154776 87480 154782 87492
rect 172014 87480 172020 87492
rect 154776 87452 172020 87480
rect 154776 87440 154782 87452
rect 172014 87440 172020 87452
rect 172072 87440 172078 87492
rect 326574 87440 326580 87492
rect 326632 87480 326638 87492
rect 327218 87480 327224 87492
rect 326632 87452 327224 87480
rect 326632 87440 326638 87452
rect 327218 87440 327224 87452
rect 327276 87480 327282 87492
rect 412870 87480 412876 87492
rect 327276 87452 412876 87480
rect 327276 87440 327282 87452
rect 412870 87440 412876 87452
rect 412928 87440 412934 87492
rect 26562 87372 26568 87424
rect 26620 87412 26626 87424
rect 73666 87412 73672 87424
rect 26620 87384 73672 87412
rect 26620 87372 26626 87384
rect 73666 87372 73672 87384
rect 73724 87372 73730 87424
rect 243406 87372 243412 87424
rect 243464 87412 243470 87424
rect 250766 87412 250772 87424
rect 243464 87384 250772 87412
rect 243464 87372 243470 87384
rect 250766 87372 250772 87384
rect 250824 87372 250830 87424
rect 359694 87372 359700 87424
rect 359752 87412 359758 87424
rect 360154 87412 360160 87424
rect 359752 87384 360160 87412
rect 359752 87372 359758 87384
rect 360154 87372 360160 87384
rect 360212 87412 360218 87424
rect 423542 87412 423548 87424
rect 360212 87384 423548 87412
rect 360212 87372 360218 87384
rect 423542 87372 423548 87384
rect 423600 87372 423606 87424
rect 29230 87304 29236 87356
rect 29288 87344 29294 87356
rect 73758 87344 73764 87356
rect 29288 87316 73764 87344
rect 29288 87304 29294 87316
rect 73758 87304 73764 87316
rect 73816 87304 73822 87356
rect 149198 87304 149204 87356
rect 149256 87344 149262 87356
rect 156926 87344 156932 87356
rect 149256 87316 156932 87344
rect 149256 87304 149262 87316
rect 156926 87304 156932 87316
rect 156984 87304 156990 87356
rect 249018 87304 249024 87356
rect 249076 87344 249082 87356
rect 258954 87344 258960 87356
rect 249076 87316 258960 87344
rect 249076 87304 249082 87316
rect 258954 87304 258960 87316
rect 259012 87304 259018 87356
rect 344974 87304 344980 87356
rect 345032 87344 345038 87356
rect 363834 87344 363840 87356
rect 345032 87316 363840 87344
rect 345032 87304 345038 87316
rect 363834 87304 363840 87316
rect 363892 87304 363898 87356
rect 369998 87304 370004 87356
rect 370056 87344 370062 87356
rect 410202 87344 410208 87356
rect 370056 87316 410208 87344
rect 370056 87304 370062 87316
rect 410202 87304 410208 87316
rect 410260 87304 410266 87356
rect 31898 87236 31904 87288
rect 31956 87276 31962 87288
rect 73482 87276 73488 87288
rect 31956 87248 73488 87276
rect 31956 87236 31962 87248
rect 73482 87236 73488 87248
rect 73540 87236 73546 87288
rect 149750 87236 149756 87288
rect 149808 87276 149814 87288
rect 158950 87276 158956 87288
rect 149808 87248 158956 87276
rect 149808 87236 149814 87248
rect 158950 87236 158956 87248
rect 159008 87236 159014 87288
rect 341018 87236 341024 87288
rect 341076 87276 341082 87288
rect 352150 87276 352156 87288
rect 341076 87248 352156 87276
rect 341076 87236 341082 87248
rect 352150 87236 352156 87248
rect 352208 87236 352214 87288
rect 34566 87168 34572 87220
rect 34624 87208 34630 87220
rect 73574 87208 73580 87220
rect 34624 87180 73580 87208
rect 34624 87168 34630 87180
rect 73574 87168 73580 87180
rect 73632 87168 73638 87220
rect 151038 87168 151044 87220
rect 151096 87208 151102 87220
rect 161710 87208 161716 87220
rect 151096 87180 161716 87208
rect 151096 87168 151102 87180
rect 161710 87168 161716 87180
rect 161768 87168 161774 87220
rect 243958 87168 243964 87220
rect 244016 87208 244022 87220
rect 252974 87208 252980 87220
rect 244016 87180 252980 87208
rect 244016 87168 244022 87180
rect 252974 87168 252980 87180
rect 253032 87168 253038 87220
rect 344330 87168 344336 87220
rect 344388 87208 344394 87220
rect 347274 87208 347280 87220
rect 344388 87180 347280 87208
rect 344388 87168 344394 87180
rect 347274 87168 347280 87180
rect 347332 87168 347338 87220
rect 21226 87100 21232 87152
rect 21284 87140 21290 87152
rect 34658 87140 34664 87152
rect 21284 87112 34664 87140
rect 21284 87100 21290 87112
rect 34658 87100 34664 87112
rect 34716 87100 34722 87152
rect 64374 87100 64380 87152
rect 64432 87140 64438 87152
rect 65938 87140 65944 87152
rect 64432 87112 65944 87140
rect 64432 87100 64438 87112
rect 65938 87100 65944 87112
rect 65996 87100 66002 87152
rect 150394 87100 150400 87152
rect 150452 87140 150458 87152
rect 159594 87140 159600 87152
rect 150452 87112 159600 87140
rect 150452 87100 150458 87112
rect 159594 87100 159600 87112
rect 159652 87100 159658 87152
rect 243038 87100 243044 87152
rect 243096 87140 243102 87152
rect 255090 87140 255096 87152
rect 243096 87112 255096 87140
rect 243096 87100 243102 87112
rect 255090 87100 255096 87112
rect 255148 87100 255154 87152
rect 338074 87100 338080 87152
rect 338132 87140 338138 87152
rect 349574 87140 349580 87152
rect 338132 87112 349580 87140
rect 338132 87100 338138 87112
rect 349574 87100 349580 87112
rect 349632 87100 349638 87152
rect 150578 87032 150584 87084
rect 150636 87072 150642 87084
rect 162078 87072 162084 87084
rect 150636 87044 162084 87072
rect 150636 87032 150642 87044
rect 162078 87032 162084 87044
rect 162136 87032 162142 87084
rect 244418 87032 244424 87084
rect 244476 87072 244482 87084
rect 253526 87072 253532 87084
rect 244476 87044 253532 87072
rect 244476 87032 244482 87044
rect 253526 87032 253532 87044
rect 253584 87032 253590 87084
rect 334118 87032 334124 87084
rect 334176 87072 334182 87084
rect 346170 87072 346176 87084
rect 334176 87044 346176 87072
rect 334176 87032 334182 87044
rect 346170 87032 346176 87044
rect 346228 87032 346234 87084
rect 149198 86964 149204 87016
rect 149256 87004 149262 87016
rect 161434 87004 161440 87016
rect 149256 86976 161440 87004
rect 149256 86964 149262 86976
rect 161434 86964 161440 86976
rect 161492 86964 161498 87016
rect 241658 86964 241664 87016
rect 241716 87004 241722 87016
rect 254538 87004 254544 87016
rect 241716 86976 254544 87004
rect 241716 86964 241722 86976
rect 254538 86964 254544 86976
rect 254596 86964 254602 87016
rect 339638 86964 339644 87016
rect 339696 87004 339702 87016
rect 340745 87007 340803 87013
rect 339696 86976 340512 87004
rect 339696 86964 339702 86976
rect 56094 86896 56100 86948
rect 56152 86936 56158 86948
rect 65846 86936 65852 86948
rect 56152 86908 65852 86936
rect 56152 86896 56158 86908
rect 65846 86896 65852 86908
rect 65904 86896 65910 86948
rect 146438 86896 146444 86948
rect 146496 86936 146502 86948
rect 160238 86936 160244 86948
rect 146496 86908 160244 86936
rect 146496 86896 146502 86908
rect 160238 86896 160244 86908
rect 160296 86896 160302 86948
rect 245338 86896 245344 86948
rect 245396 86936 245402 86948
rect 255550 86936 255556 86948
rect 245396 86908 255556 86936
rect 245396 86896 245402 86908
rect 255550 86896 255556 86908
rect 255608 86896 255614 86948
rect 335406 86896 335412 86948
rect 335464 86936 335470 86948
rect 340377 86939 340435 86945
rect 340377 86936 340389 86939
rect 335464 86908 340389 86936
rect 335464 86896 335470 86908
rect 340377 86905 340389 86908
rect 340423 86905 340435 86939
rect 340484 86936 340512 86976
rect 340745 86973 340757 87007
rect 340791 87004 340803 87007
rect 348746 87004 348752 87016
rect 340791 86976 348752 87004
rect 340791 86973 340803 86976
rect 340745 86967 340803 86973
rect 348746 86964 348752 86976
rect 348804 86964 348810 87016
rect 351230 86936 351236 86948
rect 340484 86908 351236 86936
rect 340377 86899 340435 86905
rect 351230 86896 351236 86908
rect 351288 86896 351294 86948
rect 59682 86828 59688 86880
rect 59740 86868 59746 86880
rect 70722 86868 70728 86880
rect 59740 86840 70728 86868
rect 59740 86828 59746 86840
rect 70722 86828 70728 86840
rect 70780 86828 70786 86880
rect 147818 86828 147824 86880
rect 147876 86868 147882 86880
rect 160882 86868 160888 86880
rect 147876 86840 160888 86868
rect 147876 86828 147882 86840
rect 160882 86828 160888 86840
rect 160940 86828 160946 86880
rect 160974 86828 160980 86880
rect 161032 86868 161038 86880
rect 162722 86868 162728 86880
rect 161032 86840 162728 86868
rect 161032 86828 161038 86840
rect 162722 86828 162728 86840
rect 162780 86828 162786 86880
rect 240278 86828 240284 86880
rect 240336 86868 240342 86880
rect 254262 86868 254268 86880
rect 240336 86840 254268 86868
rect 240336 86828 240342 86840
rect 254262 86828 254268 86840
rect 254320 86828 254326 86880
rect 335498 86828 335504 86880
rect 335556 86868 335562 86880
rect 348010 86868 348016 86880
rect 335556 86840 348016 86868
rect 335556 86828 335562 86840
rect 348010 86828 348016 86840
rect 348068 86828 348074 86880
rect 57014 86760 57020 86812
rect 57072 86800 57078 86812
rect 67870 86800 67876 86812
rect 57072 86772 67876 86800
rect 57072 86760 57078 86772
rect 67870 86760 67876 86772
rect 67928 86760 67934 86812
rect 145058 86760 145064 86812
rect 145116 86800 145122 86812
rect 159318 86800 159324 86812
rect 145116 86772 159324 86800
rect 145116 86760 145122 86772
rect 159318 86760 159324 86772
rect 159376 86760 159382 86812
rect 238898 86760 238904 86812
rect 238956 86800 238962 86812
rect 253250 86800 253256 86812
rect 238956 86772 253256 86800
rect 238956 86760 238962 86772
rect 253250 86760 253256 86772
rect 253308 86760 253314 86812
rect 332738 86760 332744 86812
rect 332796 86800 332802 86812
rect 345434 86800 345440 86812
rect 332796 86772 345440 86800
rect 332796 86760 332802 86772
rect 345434 86760 345440 86772
rect 345492 86760 345498 86812
rect 153430 86692 153436 86744
rect 153488 86732 153494 86744
rect 154626 86732 154632 86744
rect 153488 86704 154632 86732
rect 153488 86692 153494 86704
rect 154626 86692 154632 86704
rect 154684 86692 154690 86744
rect 340377 86735 340435 86741
rect 340377 86701 340389 86735
rect 340423 86732 340435 86735
rect 346998 86732 347004 86744
rect 340423 86704 347004 86732
rect 340423 86701 340435 86704
rect 340377 86695 340435 86701
rect 346998 86692 347004 86704
rect 347056 86692 347062 86744
rect 336878 86624 336884 86676
rect 336936 86664 336942 86676
rect 340745 86667 340803 86673
rect 340745 86664 340757 86667
rect 336936 86636 340757 86664
rect 336936 86624 336942 86636
rect 340745 86633 340757 86636
rect 340791 86633 340803 86667
rect 340745 86627 340803 86633
rect 257574 86488 257580 86540
rect 257632 86528 257638 86540
rect 258402 86528 258408 86540
rect 257632 86500 258408 86528
rect 257632 86488 257638 86500
rect 258402 86488 258408 86500
rect 258460 86488 258466 86540
rect 156834 86284 156840 86336
rect 156892 86324 156898 86336
rect 163274 86324 163280 86336
rect 156892 86296 163280 86324
rect 156892 86284 156898 86296
rect 163274 86284 163280 86296
rect 163332 86284 163338 86336
rect 152234 86216 152240 86268
rect 152292 86256 152298 86268
rect 153338 86256 153344 86268
rect 152292 86228 153344 86256
rect 152292 86216 152298 86228
rect 153338 86216 153344 86228
rect 153396 86216 153402 86268
rect 250674 86216 250680 86268
rect 250732 86256 250738 86268
rect 256378 86256 256384 86268
rect 250732 86228 256384 86256
rect 250732 86216 250738 86228
rect 256378 86216 256384 86228
rect 256436 86216 256442 86268
rect 341662 86216 341668 86268
rect 341720 86256 341726 86268
rect 344606 86256 344612 86268
rect 341720 86228 344612 86256
rect 341720 86216 341726 86228
rect 344606 86216 344612 86228
rect 344664 86216 344670 86268
rect 61614 86148 61620 86200
rect 61672 86188 61678 86200
rect 63270 86188 63276 86200
rect 61672 86160 63276 86188
rect 61672 86148 61678 86160
rect 63270 86148 63276 86160
rect 63328 86148 63334 86200
rect 67134 86148 67140 86200
rect 67192 86188 67198 86200
rect 68606 86188 68612 86200
rect 67192 86160 68612 86188
rect 67192 86148 67198 86160
rect 68606 86148 68612 86160
rect 68664 86148 68670 86200
rect 253434 86148 253440 86200
rect 253492 86188 253498 86200
rect 257666 86188 257672 86200
rect 253492 86160 257672 86188
rect 253492 86148 253498 86160
rect 257666 86148 257672 86160
rect 257724 86148 257730 86200
rect 337614 86148 337620 86200
rect 337672 86188 337678 86200
rect 339086 86188 339092 86200
rect 337672 86160 339092 86188
rect 337672 86148 337678 86160
rect 339086 86148 339092 86160
rect 339144 86148 339150 86200
rect 340098 86148 340104 86200
rect 340156 86188 340162 86200
rect 341754 86188 341760 86200
rect 340156 86160 341760 86188
rect 340156 86148 340162 86160
rect 341754 86148 341760 86160
rect 341812 86148 341818 86200
rect 342398 86148 342404 86200
rect 342456 86188 342462 86200
rect 344698 86188 344704 86200
rect 342456 86160 344704 86188
rect 342456 86148 342462 86160
rect 344698 86148 344704 86160
rect 344756 86148 344762 86200
rect 61430 86080 61436 86132
rect 61488 86120 61494 86132
rect 62258 86120 62264 86132
rect 61488 86092 62264 86120
rect 61488 86080 61494 86092
rect 62258 86080 62264 86092
rect 62316 86080 62322 86132
rect 62350 86080 62356 86132
rect 62408 86120 62414 86132
rect 63638 86120 63644 86132
rect 62408 86092 63644 86120
rect 62408 86080 62414 86092
rect 63638 86080 63644 86092
rect 63696 86080 63702 86132
rect 65754 86080 65760 86132
rect 65812 86120 65818 86132
rect 66766 86120 66772 86132
rect 65812 86092 66772 86120
rect 65812 86080 65818 86092
rect 66766 86080 66772 86092
rect 66824 86080 66830 86132
rect 68514 86080 68520 86132
rect 68572 86120 68578 86132
rect 69434 86120 69440 86132
rect 68572 86092 69440 86120
rect 68572 86080 68578 86092
rect 69434 86080 69440 86092
rect 69492 86080 69498 86132
rect 246534 86080 246540 86132
rect 246592 86120 246598 86132
rect 247086 86120 247092 86132
rect 246592 86092 247092 86120
rect 246592 86080 246598 86092
rect 247086 86080 247092 86092
rect 247144 86080 247150 86132
rect 247730 86080 247736 86132
rect 247788 86120 247794 86132
rect 248558 86120 248564 86132
rect 247788 86092 248564 86120
rect 247788 86080 247794 86092
rect 248558 86080 248564 86092
rect 248616 86080 248622 86132
rect 254814 86080 254820 86132
rect 254872 86120 254878 86132
rect 255734 86120 255740 86132
rect 254872 86092 255740 86120
rect 254872 86080 254878 86092
rect 255734 86080 255740 86092
rect 255792 86080 255798 86132
rect 256194 86080 256200 86132
rect 256252 86120 256258 86132
rect 256930 86120 256936 86132
rect 256252 86092 256936 86120
rect 256252 86080 256258 86092
rect 256930 86080 256936 86092
rect 256988 86080 256994 86132
rect 338258 86080 338264 86132
rect 338316 86120 338322 86132
rect 338994 86120 339000 86132
rect 338316 86092 339000 86120
rect 338316 86080 338322 86092
rect 338994 86080 339000 86092
rect 339052 86080 339058 86132
rect 340926 86080 340932 86132
rect 340984 86120 340990 86132
rect 341846 86120 341852 86132
rect 340984 86092 341852 86120
rect 340984 86080 340990 86092
rect 341846 86080 341852 86092
rect 341904 86080 341910 86132
rect 343502 86080 343508 86132
rect 343560 86120 343566 86132
rect 344514 86120 344520 86132
rect 343560 86092 344520 86120
rect 343560 86080 343566 86092
rect 344514 86080 344520 86092
rect 344572 86080 344578 86132
rect 66674 86012 66680 86064
rect 66732 86052 66738 86064
rect 67318 86052 67324 86064
rect 66732 86024 67324 86052
rect 66732 86012 66738 86024
rect 67318 86012 67324 86024
rect 67376 86012 67382 86064
rect 230986 85876 230992 85928
rect 231044 85916 231050 85928
rect 232734 85916 232740 85928
rect 231044 85888 232740 85916
rect 231044 85876 231050 85888
rect 232734 85876 232740 85888
rect 232792 85876 232798 85928
rect 324550 85740 324556 85792
rect 324608 85780 324614 85792
rect 326666 85780 326672 85792
rect 324608 85752 326672 85780
rect 324608 85740 324614 85752
rect 326666 85740 326672 85752
rect 326724 85740 326730 85792
rect 138158 85468 138164 85520
rect 138216 85508 138222 85520
rect 144414 85508 144420 85520
rect 138216 85480 144420 85508
rect 138216 85468 138222 85480
rect 144414 85468 144420 85480
rect 144472 85468 144478 85520
rect 354910 84040 354916 84092
rect 354968 84080 354974 84092
rect 355830 84080 355836 84092
rect 354968 84052 355836 84080
rect 354968 84040 354974 84052
rect 355830 84040 355836 84052
rect 355888 84040 355894 84092
rect 88478 81932 88484 81984
rect 88536 81972 88542 81984
rect 182410 81972 182416 81984
rect 88536 81944 182416 81972
rect 88536 81932 88542 81944
rect 182410 81932 182416 81944
rect 182468 81972 182474 81984
rect 276250 81972 276256 81984
rect 182468 81944 276256 81972
rect 182468 81932 182474 81944
rect 276250 81932 276256 81944
rect 276308 81932 276314 81984
rect 95746 81864 95752 81916
rect 95804 81904 95810 81916
rect 176154 81904 176160 81916
rect 95804 81876 176160 81904
rect 95804 81864 95810 81876
rect 176154 81864 176160 81876
rect 176212 81904 176218 81916
rect 189494 81904 189500 81916
rect 176212 81876 189500 81904
rect 176212 81864 176218 81876
rect 189494 81864 189500 81876
rect 189552 81904 189558 81916
rect 283426 81904 283432 81916
rect 189552 81876 283432 81904
rect 189552 81864 189558 81876
rect 283426 81864 283432 81876
rect 283484 81864 283490 81916
rect 102922 81796 102928 81848
rect 102980 81836 102986 81848
rect 174774 81836 174780 81848
rect 102980 81808 174780 81836
rect 102980 81796 102986 81808
rect 174774 81796 174780 81808
rect 174832 81836 174838 81848
rect 196670 81836 196676 81848
rect 174832 81808 196676 81836
rect 174832 81796 174838 81808
rect 196670 81796 196676 81808
rect 196728 81836 196734 81848
rect 290326 81836 290332 81848
rect 196728 81808 290332 81836
rect 196728 81796 196734 81808
rect 290326 81796 290332 81808
rect 290384 81796 290390 81848
rect 285818 81320 285824 81372
rect 285876 81360 285882 81372
rect 297502 81360 297508 81372
rect 285876 81332 297508 81360
rect 285876 81320 285882 81332
rect 297502 81320 297508 81332
rect 297560 81320 297566 81372
rect 369906 81360 369912 81372
rect 369867 81332 369912 81360
rect 369906 81320 369912 81332
rect 369964 81320 369970 81372
rect 96758 81252 96764 81304
rect 96816 81292 96822 81304
rect 109822 81292 109828 81304
rect 96816 81264 109828 81292
rect 96816 81252 96822 81264
rect 109822 81252 109828 81264
rect 109880 81252 109886 81304
rect 190598 81252 190604 81304
rect 190656 81292 190662 81304
rect 203754 81292 203760 81304
rect 190656 81264 203760 81292
rect 190656 81252 190662 81264
rect 203754 81252 203760 81264
rect 203812 81252 203818 81304
rect 283426 81252 283432 81304
rect 283484 81292 283490 81304
rect 428050 81292 428056 81304
rect 283484 81264 428056 81292
rect 283484 81252 283490 81264
rect 428050 81252 428056 81264
rect 428108 81252 428114 81304
rect 129234 80572 129240 80624
rect 129292 80612 129298 80624
rect 131258 80612 131264 80624
rect 129292 80584 131264 80612
rect 129292 80572 129298 80584
rect 131258 80572 131264 80584
rect 131316 80572 131322 80624
rect 223074 80572 223080 80624
rect 223132 80612 223138 80624
rect 225190 80612 225196 80624
rect 223132 80584 225196 80612
rect 223132 80572 223138 80584
rect 225190 80572 225196 80584
rect 225248 80572 225254 80624
rect 316914 80572 316920 80624
rect 316972 80612 316978 80624
rect 319122 80612 319128 80624
rect 316972 80584 319128 80612
rect 316972 80572 316978 80584
rect 319122 80572 319128 80584
rect 319180 80572 319186 80624
rect 60234 79144 60240 79196
rect 60292 79184 60298 79196
rect 64374 79184 64380 79196
rect 60292 79156 64380 79184
rect 60292 79144 60298 79156
rect 64374 79144 64380 79156
rect 64432 79144 64438 79196
rect 153338 79144 153344 79196
rect 153396 79184 153402 79196
rect 156834 79184 156840 79196
rect 153396 79156 156840 79184
rect 153396 79144 153402 79156
rect 156834 79144 156840 79156
rect 156892 79144 156898 79196
rect 156926 79144 156932 79196
rect 156984 79184 156990 79196
rect 157570 79184 157576 79196
rect 156984 79156 157576 79184
rect 156984 79144 156990 79156
rect 157570 79144 157576 79156
rect 157628 79144 157634 79196
rect 159594 79144 159600 79196
rect 159652 79184 159658 79196
rect 160330 79184 160336 79196
rect 159652 79156 160336 79184
rect 159652 79144 159658 79156
rect 160330 79144 160336 79156
rect 160388 79144 160394 79196
rect 250766 79144 250772 79196
rect 250824 79184 250830 79196
rect 251410 79184 251416 79196
rect 250824 79156 251416 79184
rect 250824 79144 250830 79156
rect 251410 79144 251416 79156
rect 251468 79144 251474 79196
rect 253526 79144 253532 79196
rect 253584 79184 253590 79196
rect 254170 79184 254176 79196
rect 253584 79156 254176 79184
rect 253584 79144 253590 79156
rect 254170 79144 254176 79156
rect 254228 79144 254234 79196
rect 333382 79144 333388 79196
rect 333440 79184 333446 79196
rect 334118 79184 334124 79196
rect 333440 79156 334124 79184
rect 333440 79144 333446 79156
rect 334118 79144 334124 79156
rect 334176 79144 334182 79196
rect 334394 79144 334400 79196
rect 334452 79184 334458 79196
rect 335406 79184 335412 79196
rect 334452 79156 335412 79184
rect 334452 79144 334458 79156
rect 335406 79144 335412 79156
rect 335464 79144 335470 79196
rect 339546 79144 339552 79196
rect 339604 79184 339610 79196
rect 343778 79184 343784 79196
rect 339604 79156 343784 79184
rect 339604 79144 339610 79156
rect 343778 79144 343784 79156
rect 343836 79144 343842 79196
rect 344698 79144 344704 79196
rect 344756 79184 344762 79196
rect 344756 79156 346952 79184
rect 344756 79144 344762 79156
rect 59222 79076 59228 79128
rect 59280 79116 59286 79128
rect 63822 79116 63828 79128
rect 59280 79088 63828 79116
rect 59280 79076 59286 79088
rect 63822 79076 63828 79088
rect 63880 79076 63886 79128
rect 66674 79116 66680 79128
rect 63932 79088 66680 79116
rect 58210 78940 58216 78992
rect 58268 78980 58274 78992
rect 63730 78980 63736 78992
rect 58268 78952 63736 78980
rect 58268 78940 58274 78952
rect 63730 78940 63736 78952
rect 63788 78940 63794 78992
rect 62350 78872 62356 78924
rect 62408 78912 62414 78924
rect 63932 78912 63960 79088
rect 66674 79076 66680 79088
rect 66732 79076 66738 79128
rect 154534 79076 154540 79128
rect 154592 79116 154598 79128
rect 154718 79116 154724 79128
rect 154592 79088 154724 79116
rect 154592 79076 154598 79088
rect 154718 79076 154724 79088
rect 154776 79076 154782 79128
rect 250398 79076 250404 79128
rect 250456 79116 250462 79128
rect 257574 79116 257580 79128
rect 250456 79088 257580 79116
rect 250456 79076 250462 79088
rect 257574 79076 257580 79088
rect 257632 79076 257638 79128
rect 338994 79076 339000 79128
rect 339052 79116 339058 79128
rect 342674 79116 342680 79128
rect 339052 79088 342680 79116
rect 339052 79076 339058 79088
rect 342674 79076 342680 79088
rect 342732 79076 342738 79128
rect 344606 79076 344612 79128
rect 344664 79116 344670 79128
rect 346814 79116 346820 79128
rect 344664 79088 346820 79116
rect 344664 79076 344670 79088
rect 346814 79076 346820 79088
rect 346872 79076 346878 79128
rect 346924 79116 346952 79156
rect 347274 79144 347280 79196
rect 347332 79184 347338 79196
rect 349942 79184 349948 79196
rect 347332 79156 349948 79184
rect 347332 79144 347338 79156
rect 349942 79144 349948 79156
rect 350000 79144 350006 79196
rect 369262 79144 369268 79196
rect 369320 79184 369326 79196
rect 369814 79184 369820 79196
rect 369320 79156 369820 79184
rect 369320 79144 369326 79156
rect 369814 79144 369820 79156
rect 369872 79144 369878 79196
rect 347918 79116 347924 79128
rect 346924 79088 347924 79116
rect 347918 79076 347924 79088
rect 347976 79076 347982 79128
rect 337522 79008 337528 79060
rect 337580 79048 337586 79060
rect 338258 79048 338264 79060
rect 337580 79020 338264 79048
rect 337580 79008 337586 79020
rect 338258 79008 338264 79020
rect 338316 79008 338322 79060
rect 341846 79008 341852 79060
rect 341904 79048 341910 79060
rect 345802 79048 345808 79060
rect 341904 79020 345808 79048
rect 341904 79008 341910 79020
rect 345802 79008 345808 79020
rect 345860 79008 345866 79060
rect 151958 78980 151964 78992
rect 151884 78952 151964 78980
rect 62408 78884 63960 78912
rect 62408 78872 62414 78884
rect 64374 78872 64380 78924
rect 64432 78912 64438 78924
rect 68514 78912 68520 78924
rect 64432 78884 68520 78912
rect 64432 78872 64438 78884
rect 68514 78872 68520 78884
rect 68572 78872 68578 78924
rect 63638 78804 63644 78856
rect 63696 78844 63702 78856
rect 74770 78844 74776 78856
rect 63696 78816 74776 78844
rect 63696 78804 63702 78816
rect 74770 78804 74776 78816
rect 74828 78804 74834 78856
rect 62258 78736 62264 78788
rect 62316 78776 62322 78788
rect 65389 78779 65447 78785
rect 65389 78776 65401 78779
rect 62316 78748 65401 78776
rect 62316 78736 62322 78748
rect 65389 78745 65401 78748
rect 65435 78745 65447 78779
rect 65389 78739 65447 78745
rect 65478 78736 65484 78788
rect 65536 78776 65542 78788
rect 69342 78776 69348 78788
rect 65536 78748 69348 78776
rect 65536 78736 65542 78748
rect 69342 78736 69348 78748
rect 69400 78736 69406 78788
rect 151884 78776 151912 78952
rect 151958 78940 151964 78952
rect 152016 78940 152022 78992
rect 156098 78940 156104 78992
rect 156156 78980 156162 78992
rect 164470 78980 164476 78992
rect 156156 78952 164476 78980
rect 156156 78940 156162 78952
rect 164470 78940 164476 78952
rect 164528 78940 164534 78992
rect 341754 78940 341760 78992
rect 341812 78980 341818 78992
rect 344790 78980 344796 78992
rect 341812 78952 344796 78980
rect 341812 78940 341818 78952
rect 344790 78940 344796 78952
rect 344848 78940 344854 78992
rect 154718 78872 154724 78924
rect 154776 78912 154782 78924
rect 163182 78912 163188 78924
rect 154776 78884 163188 78912
rect 154776 78872 154782 78884
rect 163182 78872 163188 78884
rect 163240 78872 163246 78924
rect 247638 78872 247644 78924
rect 247696 78912 247702 78924
rect 256194 78912 256200 78924
rect 247696 78884 256200 78912
rect 247696 78872 247702 78884
rect 256194 78872 256200 78884
rect 256252 78872 256258 78924
rect 151958 78804 151964 78856
rect 152016 78844 152022 78856
rect 160974 78844 160980 78856
rect 152016 78816 160980 78844
rect 152016 78804 152022 78816
rect 160974 78804 160980 78816
rect 161032 78804 161038 78856
rect 244878 78804 244884 78856
rect 244936 78844 244942 78856
rect 254814 78844 254820 78856
rect 244936 78816 254820 78844
rect 244936 78804 244942 78816
rect 254814 78804 254820 78816
rect 254872 78804 254878 78856
rect 163090 78776 163096 78788
rect 151884 78748 163096 78776
rect 163090 78736 163096 78748
rect 163148 78736 163154 78788
rect 245798 78736 245804 78788
rect 245856 78776 245862 78788
rect 256930 78776 256936 78788
rect 245856 78748 256936 78776
rect 245856 78736 245862 78748
rect 256930 78736 256936 78748
rect 256988 78736 256994 78788
rect 339086 78736 339092 78788
rect 339144 78776 339150 78788
rect 341662 78776 341668 78788
rect 339144 78748 341668 78776
rect 339144 78736 339150 78748
rect 341662 78736 341668 78748
rect 341720 78736 341726 78788
rect 63362 78668 63368 78720
rect 63420 78708 63426 78720
rect 67134 78708 67140 78720
rect 63420 78680 67140 78708
rect 63420 78668 63426 78680
rect 67134 78668 67140 78680
rect 67192 78668 67198 78720
rect 153246 78668 153252 78720
rect 153304 78708 153310 78720
rect 164562 78708 164568 78720
rect 153304 78680 164568 78708
rect 153304 78668 153310 78680
rect 164562 78668 164568 78680
rect 164620 78668 164626 78720
rect 247086 78668 247092 78720
rect 247144 78708 247150 78720
rect 258402 78708 258408 78720
rect 247144 78680 258408 78708
rect 247144 78668 247150 78680
rect 258402 78668 258408 78680
rect 258460 78668 258466 78720
rect 60878 78600 60884 78652
rect 60936 78640 60942 78652
rect 72654 78640 72660 78652
rect 60936 78612 72660 78640
rect 60936 78600 60942 78612
rect 72654 78600 72660 78612
rect 72712 78600 72718 78652
rect 154626 78600 154632 78652
rect 154684 78640 154690 78652
rect 167322 78640 167328 78652
rect 154684 78612 167328 78640
rect 154684 78600 154690 78612
rect 167322 78600 167328 78612
rect 167380 78600 167386 78652
rect 248558 78600 248564 78652
rect 248616 78640 248622 78652
rect 261070 78640 261076 78652
rect 248616 78612 261076 78640
rect 248616 78600 248622 78612
rect 261070 78600 261076 78612
rect 261128 78600 261134 78652
rect 58118 78532 58124 78584
rect 58176 78572 58182 78584
rect 69618 78572 69624 78584
rect 58176 78544 69624 78572
rect 58176 78532 58182 78544
rect 69618 78532 69624 78544
rect 69676 78532 69682 78584
rect 153062 78532 153068 78584
rect 153120 78572 153126 78584
rect 165942 78572 165948 78584
rect 153120 78544 165948 78572
rect 153120 78532 153126 78544
rect 165942 78532 165948 78544
rect 166000 78532 166006 78584
rect 247178 78532 247184 78584
rect 247236 78572 247242 78584
rect 259690 78572 259696 78584
rect 247236 78544 259696 78572
rect 247236 78532 247242 78544
rect 259690 78532 259696 78544
rect 259748 78532 259754 78584
rect 344514 78532 344520 78584
rect 344572 78572 344578 78584
rect 348930 78572 348936 78584
rect 344572 78544 348936 78572
rect 344572 78532 344578 78544
rect 348930 78532 348936 78544
rect 348988 78532 348994 78584
rect 55358 78464 55364 78516
rect 55416 78504 55422 78516
rect 66490 78504 66496 78516
rect 55416 78476 66496 78504
rect 55416 78464 55422 78476
rect 66490 78464 66496 78476
rect 66548 78464 66554 78516
rect 154534 78464 154540 78516
rect 154592 78504 154598 78516
rect 168702 78504 168708 78516
rect 154592 78476 168708 78504
rect 154592 78464 154598 78476
rect 168702 78464 168708 78476
rect 168760 78464 168766 78516
rect 248466 78464 248472 78516
rect 248524 78504 248530 78516
rect 262450 78504 262456 78516
rect 248524 78476 262456 78504
rect 248524 78464 248530 78476
rect 262450 78464 262456 78476
rect 262508 78464 262514 78516
rect 338534 78464 338540 78516
rect 338592 78504 338598 78516
rect 349482 78504 349488 78516
rect 338592 78476 349488 78504
rect 338592 78464 338598 78476
rect 349482 78464 349488 78476
rect 349540 78464 349546 78516
rect 59498 78396 59504 78448
rect 59556 78436 59562 78448
rect 70630 78436 70636 78448
rect 59556 78408 70636 78436
rect 59556 78396 59562 78408
rect 70630 78396 70636 78408
rect 70688 78396 70694 78448
rect 65389 78371 65447 78377
rect 65389 78337 65401 78371
rect 65435 78368 65447 78371
rect 73758 78368 73764 78380
rect 65435 78340 73764 78368
rect 65435 78337 65447 78340
rect 65389 78331 65447 78337
rect 73758 78328 73764 78340
rect 73816 78328 73822 78380
rect 65846 78192 65852 78244
rect 65904 78232 65910 78244
rect 67502 78232 67508 78244
rect 65904 78204 67508 78232
rect 65904 78192 65910 78204
rect 67502 78192 67508 78204
rect 67560 78192 67566 78244
rect 246258 78124 246264 78176
rect 246316 78164 246322 78176
rect 250674 78164 250680 78176
rect 246316 78136 250680 78164
rect 246316 78124 246322 78136
rect 250674 78124 250680 78136
rect 250732 78124 250738 78176
rect 57198 78056 57204 78108
rect 57256 78096 57262 78108
rect 61614 78096 61620 78108
rect 57256 78068 61620 78096
rect 57256 78056 57262 78068
rect 61614 78056 61620 78068
rect 61672 78056 61678 78108
rect 61338 77988 61344 78040
rect 61396 78028 61402 78040
rect 65754 78028 65760 78040
rect 61396 78000 65760 78028
rect 61396 77988 61402 78000
rect 65754 77988 65760 78000
rect 65812 77988 65818 78040
rect 249018 77920 249024 77972
rect 249076 77960 249082 77972
rect 253434 77960 253440 77972
rect 249076 77932 253440 77960
rect 249076 77920 249082 77932
rect 253434 77920 253440 77932
rect 253492 77920 253498 77972
rect 75782 77852 75788 77904
rect 75840 77892 75846 77904
rect 76886 77892 76892 77904
rect 75840 77864 76892 77892
rect 75840 77852 75846 77864
rect 76886 77852 76892 77864
rect 76944 77852 76950 77904
rect 369906 76464 369912 76476
rect 369867 76436 369912 76464
rect 369906 76424 369912 76436
rect 369964 76424 369970 76476
rect 78910 76356 78916 76408
rect 78968 76396 78974 76408
rect 123990 76396 123996 76408
rect 78968 76368 123996 76396
rect 78968 76356 78974 76368
rect 123990 76356 123996 76368
rect 124048 76396 124054 76408
rect 139630 76396 139636 76408
rect 124048 76368 139636 76396
rect 124048 76356 124054 76368
rect 139630 76356 139636 76368
rect 139688 76356 139694 76408
rect 173854 76356 173860 76408
rect 173912 76396 173918 76408
rect 218014 76396 218020 76408
rect 173912 76368 218020 76396
rect 173912 76356 173918 76368
rect 218014 76356 218020 76368
rect 218072 76396 218078 76408
rect 233470 76396 233476 76408
rect 218072 76368 233476 76396
rect 218072 76356 218078 76368
rect 233470 76356 233476 76368
rect 233528 76356 233534 76408
rect 266590 76356 266596 76408
rect 266648 76396 266654 76408
rect 312038 76396 312044 76408
rect 266648 76368 312044 76396
rect 266648 76356 266654 76368
rect 312038 76356 312044 76368
rect 312096 76396 312102 76408
rect 328414 76396 328420 76408
rect 312096 76368 328420 76396
rect 312096 76356 312102 76368
rect 328414 76356 328420 76368
rect 328472 76356 328478 76408
rect 427406 76356 427412 76408
rect 427464 76396 427470 76408
rect 429430 76396 429436 76408
rect 427464 76368 429436 76396
rect 427464 76356 427470 76368
rect 429430 76356 429436 76368
rect 429488 76356 429494 76408
rect 155362 75512 155368 75524
rect 155323 75484 155368 75512
rect 155362 75472 155368 75484
rect 155420 75472 155426 75524
rect 249202 75444 249208 75456
rect 249163 75416 249208 75444
rect 249202 75404 249208 75416
rect 249260 75404 249266 75456
rect 78910 73704 78916 73756
rect 78968 73744 78974 73756
rect 87374 73744 87380 73756
rect 78968 73716 87380 73744
rect 78968 73704 78974 73716
rect 87374 73704 87380 73716
rect 87432 73704 87438 73756
rect 155365 73747 155423 73753
rect 155365 73713 155377 73747
rect 155411 73744 155423 73747
rect 170634 73744 170640 73756
rect 155411 73716 170640 73744
rect 155411 73713 155423 73716
rect 155365 73707 155423 73713
rect 170634 73704 170640 73716
rect 170692 73704 170698 73756
rect 249205 73747 249263 73753
rect 249205 73713 249217 73747
rect 249251 73744 249263 73747
rect 264474 73744 264480 73756
rect 249251 73716 264480 73744
rect 249251 73713 249263 73716
rect 249205 73707 249263 73713
rect 264474 73704 264480 73716
rect 264532 73704 264538 73756
rect 304862 73704 304868 73756
rect 304920 73744 304926 73756
rect 305046 73744 305052 73756
rect 304920 73716 305052 73744
rect 304920 73704 304926 73716
rect 305046 73704 305052 73716
rect 305104 73704 305110 73756
rect 110190 73432 110196 73484
rect 110248 73472 110254 73484
rect 116814 73472 116820 73484
rect 110248 73444 116820 73472
rect 110248 73432 110254 73444
rect 116814 73432 116820 73444
rect 116872 73432 116878 73484
rect 204122 72956 204128 73008
rect 204180 72996 204186 73008
rect 210930 72996 210936 73008
rect 204180 72968 210936 72996
rect 204180 72956 204186 72968
rect 210930 72956 210936 72968
rect 210988 72956 210994 73008
rect 217554 72956 217560 73008
rect 217612 72996 217618 73008
rect 223074 72996 223080 73008
rect 217612 72968 223080 72996
rect 217612 72956 217618 72968
rect 223074 72956 223080 72968
rect 223132 72956 223138 73008
rect 311210 72480 311216 72532
rect 311268 72520 311274 72532
rect 316914 72520 316920 72532
rect 311268 72492 316920 72520
rect 311268 72480 311274 72492
rect 316914 72480 316920 72492
rect 316972 72480 316978 72532
rect 78910 72344 78916 72396
rect 78968 72384 78974 72396
rect 87190 72384 87196 72396
rect 78968 72356 87196 72384
rect 78968 72344 78974 72356
rect 87190 72344 87196 72356
rect 87248 72344 87254 72396
rect 123530 72344 123536 72396
rect 123588 72384 123594 72396
rect 129234 72384 129240 72396
rect 123588 72356 129240 72384
rect 123588 72344 123594 72356
rect 129234 72344 129240 72356
rect 129292 72344 129298 72396
rect 173486 72344 173492 72396
rect 173544 72384 173550 72396
rect 178270 72384 178276 72396
rect 173544 72356 178276 72384
rect 173544 72344 173550 72356
rect 178270 72344 178276 72356
rect 178328 72344 178334 72396
rect 230158 72344 230164 72396
rect 230216 72384 230222 72396
rect 233470 72384 233476 72396
rect 230216 72356 233476 72384
rect 230216 72344 230222 72356
rect 233470 72344 233476 72356
rect 233528 72344 233534 72396
rect 266590 72344 266596 72396
rect 266648 72384 266654 72396
rect 274962 72384 274968 72396
rect 266648 72356 274968 72384
rect 266648 72344 266654 72356
rect 274962 72344 274968 72356
rect 275020 72344 275026 72396
rect 284530 72344 284536 72396
rect 284588 72384 284594 72396
rect 285818 72384 285824 72396
rect 284588 72356 285824 72384
rect 284588 72344 284594 72356
rect 285818 72344 285824 72356
rect 285876 72344 285882 72396
rect 297870 72344 297876 72396
rect 297928 72384 297934 72396
rect 304862 72384 304868 72396
rect 297928 72356 304868 72384
rect 297928 72344 297934 72356
rect 304862 72344 304868 72356
rect 304920 72344 304926 72396
rect 173486 71732 173492 71784
rect 173544 71772 173550 71784
rect 178362 71772 178368 71784
rect 173544 71744 178368 71772
rect 173544 71732 173550 71744
rect 178362 71732 178368 71744
rect 178420 71732 178426 71784
rect 78910 70984 78916 71036
rect 78968 71024 78974 71036
rect 85718 71024 85724 71036
rect 78968 70996 85724 71024
rect 78968 70984 78974 70996
rect 85718 70984 85724 70996
rect 85776 70984 85782 71036
rect 173302 70984 173308 71036
rect 173360 71024 173366 71036
rect 180846 71024 180852 71036
rect 173360 70996 180852 71024
rect 173360 70984 173366 70996
rect 180846 70984 180852 70996
rect 180904 70984 180910 71036
rect 266682 70984 266688 71036
rect 266740 71024 266746 71036
rect 274778 71024 274784 71036
rect 266740 70996 274784 71024
rect 266740 70984 266746 70996
rect 274778 70984 274784 70996
rect 274836 70984 274842 71036
rect 266590 70916 266596 70968
rect 266648 70956 266654 70968
rect 274686 70956 274692 70968
rect 266648 70928 274692 70956
rect 266648 70916 266654 70928
rect 274686 70916 274692 70928
rect 274744 70916 274750 70968
rect 173302 70032 173308 70084
rect 173360 70072 173366 70084
rect 178454 70072 178460 70084
rect 173360 70044 178460 70072
rect 173360 70032 173366 70044
rect 178454 70032 178460 70044
rect 178512 70032 178518 70084
rect 78910 69556 78916 69608
rect 78968 69596 78974 69608
rect 84890 69596 84896 69608
rect 78968 69568 84896 69596
rect 78968 69556 78974 69568
rect 84890 69556 84896 69568
rect 84948 69556 84954 69608
rect 229882 69556 229888 69608
rect 229940 69596 229946 69608
rect 233562 69596 233568 69608
rect 229940 69568 233568 69596
rect 229940 69556 229946 69568
rect 233562 69556 233568 69568
rect 233620 69556 233626 69608
rect 266590 69556 266596 69608
rect 266648 69596 266654 69608
rect 270546 69596 270552 69608
rect 266648 69568 270552 69596
rect 266648 69556 266654 69568
rect 270546 69556 270552 69568
rect 270604 69556 270610 69608
rect 131442 69488 131448 69540
rect 131500 69528 131506 69540
rect 139630 69528 139636 69540
rect 131500 69500 139636 69528
rect 131500 69488 131506 69500
rect 139630 69488 139636 69500
rect 139688 69488 139694 69540
rect 172934 69488 172940 69540
rect 172992 69528 172998 69540
rect 182318 69528 182324 69540
rect 172992 69500 182324 69528
rect 172992 69488 172998 69500
rect 182318 69488 182324 69500
rect 182376 69488 182382 69540
rect 226294 69488 226300 69540
rect 226352 69528 226358 69540
rect 233930 69528 233936 69540
rect 226352 69500 233936 69528
rect 226352 69488 226358 69500
rect 233930 69488 233936 69500
rect 233988 69488 233994 69540
rect 267418 69488 267424 69540
rect 267476 69528 267482 69540
rect 274870 69528 274876 69540
rect 267476 69500 274876 69528
rect 267476 69488 267482 69500
rect 274870 69488 274876 69500
rect 274928 69488 274934 69540
rect 369722 69488 369728 69540
rect 369780 69528 369786 69540
rect 369906 69528 369912 69540
rect 369780 69500 369912 69528
rect 369780 69488 369786 69500
rect 369906 69488 369912 69500
rect 369964 69488 369970 69540
rect 131350 69420 131356 69472
rect 131408 69460 131414 69472
rect 139814 69460 139820 69472
rect 131408 69432 139820 69460
rect 131408 69420 131414 69432
rect 139814 69420 139820 69432
rect 139872 69420 139878 69472
rect 178270 69420 178276 69472
rect 178328 69460 178334 69472
rect 181674 69460 181680 69472
rect 178328 69432 181680 69460
rect 178328 69420 178334 69432
rect 181674 69420 181680 69432
rect 181732 69420 181738 69472
rect 226386 69420 226392 69472
rect 226444 69460 226450 69472
rect 230158 69460 230164 69472
rect 226444 69432 230164 69460
rect 226444 69420 226450 69432
rect 230158 69420 230164 69432
rect 230216 69420 230222 69472
rect 321606 68536 321612 68588
rect 321664 68576 321670 68588
rect 327034 68576 327040 68588
rect 321664 68548 327040 68576
rect 321664 68536 321670 68548
rect 327034 68536 327040 68548
rect 327092 68536 327098 68588
rect 321606 68332 321612 68384
rect 321664 68372 321670 68384
rect 327862 68372 327868 68384
rect 321664 68344 327868 68372
rect 321664 68332 321670 68344
rect 327862 68332 327868 68344
rect 327920 68332 327926 68384
rect 78910 68196 78916 68248
rect 78968 68236 78974 68248
rect 85626 68236 85632 68248
rect 78968 68208 85632 68236
rect 78968 68196 78974 68208
rect 85626 68196 85632 68208
rect 85684 68196 85690 68248
rect 136686 68196 136692 68248
rect 136744 68236 136750 68248
rect 139630 68236 139636 68248
rect 136744 68208 139636 68236
rect 136744 68196 136750 68208
rect 139630 68196 139636 68208
rect 139688 68196 139694 68248
rect 173118 68196 173124 68248
rect 173176 68236 173182 68248
rect 178270 68236 178276 68248
rect 173176 68208 178276 68236
rect 173176 68196 173182 68208
rect 178270 68196 178276 68208
rect 178328 68196 178334 68248
rect 266590 68196 266596 68248
rect 266648 68236 266654 68248
rect 272662 68236 272668 68248
rect 266648 68208 272668 68236
rect 266648 68196 266654 68208
rect 272662 68196 272668 68208
rect 272720 68196 272726 68248
rect 85718 68128 85724 68180
rect 85776 68168 85782 68180
rect 87190 68168 87196 68180
rect 85776 68140 87196 68168
rect 85776 68128 85782 68140
rect 87190 68128 87196 68140
rect 87248 68128 87254 68180
rect 132362 68128 132368 68180
rect 132420 68168 132426 68180
rect 139722 68168 139728 68180
rect 132420 68140 139728 68168
rect 132420 68128 132426 68140
rect 139722 68128 139728 68140
rect 139780 68128 139786 68180
rect 178362 68128 178368 68180
rect 178420 68168 178426 68180
rect 181398 68168 181404 68180
rect 178420 68140 181404 68168
rect 178420 68128 178426 68140
rect 181398 68128 181404 68140
rect 181456 68128 181462 68180
rect 226294 68128 226300 68180
rect 226352 68168 226358 68180
rect 233470 68168 233476 68180
rect 226352 68140 233476 68168
rect 226352 68128 226358 68140
rect 233470 68128 233476 68140
rect 233528 68128 233534 68180
rect 79554 67516 79560 67568
rect 79612 67556 79618 67568
rect 129418 67556 129424 67568
rect 79612 67528 129424 67556
rect 79612 67516 79618 67528
rect 129418 67516 129424 67528
rect 129476 67516 129482 67568
rect 173394 67516 173400 67568
rect 173452 67556 173458 67568
rect 223442 67556 223448 67568
rect 173452 67528 223448 67556
rect 173452 67516 173458 67528
rect 223442 67516 223448 67528
rect 223500 67516 223506 67568
rect 267234 67516 267240 67568
rect 267292 67556 267298 67568
rect 317558 67556 317564 67568
rect 267292 67528 317564 67556
rect 267292 67516 267298 67528
rect 317558 67516 317564 67528
rect 317616 67516 317622 67568
rect 320502 67176 320508 67228
rect 320560 67216 320566 67228
rect 327126 67216 327132 67228
rect 320560 67188 327132 67216
rect 320560 67176 320566 67188
rect 327126 67176 327132 67188
rect 327184 67176 327190 67228
rect 78910 67040 78916 67092
rect 78968 67080 78974 67092
rect 81670 67080 81676 67092
rect 78968 67052 81676 67080
rect 78968 67040 78974 67052
rect 81670 67040 81676 67052
rect 81728 67040 81734 67092
rect 78910 66904 78916 66956
rect 78968 66944 78974 66956
rect 85166 66944 85172 66956
rect 78968 66916 85172 66944
rect 78968 66904 78974 66916
rect 85166 66904 85172 66916
rect 85224 66904 85230 66956
rect 174038 66904 174044 66956
rect 174096 66944 174102 66956
rect 179098 66944 179104 66956
rect 174096 66916 179104 66944
rect 174096 66904 174102 66916
rect 179098 66904 179104 66916
rect 179156 66904 179162 66956
rect 136778 66836 136784 66888
rect 136836 66876 136842 66888
rect 139722 66876 139728 66888
rect 136836 66848 139728 66876
rect 136836 66836 136842 66848
rect 139722 66836 139728 66848
rect 139780 66836 139786 66888
rect 266682 66836 266688 66888
rect 266740 66876 266746 66888
rect 272478 66876 272484 66888
rect 266740 66848 272484 66876
rect 266740 66836 266746 66848
rect 272478 66836 272484 66848
rect 272536 66836 272542 66888
rect 321054 66836 321060 66888
rect 321112 66876 321118 66888
rect 328414 66876 328420 66888
rect 321112 66848 328420 66876
rect 321112 66836 321118 66848
rect 328414 66836 328420 66848
rect 328472 66836 328478 66888
rect 136134 66768 136140 66820
rect 136192 66808 136198 66820
rect 139630 66808 139636 66820
rect 136192 66780 139636 66808
rect 136192 66768 136198 66780
rect 139630 66768 139636 66780
rect 139688 66768 139694 66820
rect 173670 66768 173676 66820
rect 173728 66808 173734 66820
rect 175602 66808 175608 66820
rect 173728 66780 175608 66808
rect 173728 66768 173734 66780
rect 175602 66768 175608 66780
rect 175660 66768 175666 66820
rect 230066 66768 230072 66820
rect 230124 66808 230130 66820
rect 233470 66808 233476 66820
rect 230124 66780 233476 66808
rect 230124 66768 230130 66780
rect 233470 66768 233476 66780
rect 233528 66768 233534 66820
rect 266590 66768 266596 66820
rect 266648 66808 266654 66820
rect 272754 66808 272760 66820
rect 266648 66780 272760 66808
rect 266648 66768 266654 66780
rect 272754 66768 272760 66780
rect 272812 66768 272818 66820
rect 369262 66768 369268 66820
rect 369320 66808 369326 66820
rect 369814 66808 369820 66820
rect 369320 66780 369820 66808
rect 369320 66768 369326 66780
rect 369814 66768 369820 66780
rect 369872 66768 369878 66820
rect 80290 66700 80296 66752
rect 80348 66740 80354 66752
rect 87190 66740 87196 66752
rect 80348 66712 87196 66740
rect 80348 66700 80354 66712
rect 87190 66700 87196 66712
rect 87248 66700 87254 66752
rect 129418 66740 129424 66752
rect 129379 66712 129424 66740
rect 129418 66700 129424 66712
rect 129476 66700 129482 66752
rect 132362 66700 132368 66752
rect 132420 66740 132426 66752
rect 139906 66740 139912 66752
rect 132420 66712 139912 66740
rect 132420 66700 132426 66712
rect 139906 66700 139912 66712
rect 139964 66700 139970 66752
rect 226294 66700 226300 66752
rect 226352 66740 226358 66752
rect 233746 66740 233752 66752
rect 226352 66712 233752 66740
rect 226352 66700 226358 66712
rect 233746 66700 233752 66712
rect 233804 66700 233810 66752
rect 270546 66700 270552 66752
rect 270604 66740 270610 66752
rect 274870 66740 274876 66752
rect 270604 66712 274876 66740
rect 270604 66700 270610 66712
rect 274870 66700 274876 66712
rect 274928 66700 274934 66752
rect 84890 66632 84896 66684
rect 84948 66672 84954 66684
rect 87282 66672 87288 66684
rect 84948 66644 87288 66672
rect 84948 66632 84954 66644
rect 87282 66632 87288 66644
rect 87340 66632 87346 66684
rect 131350 66632 131356 66684
rect 131408 66672 131414 66684
rect 139998 66672 140004 66684
rect 131408 66644 140004 66672
rect 131408 66632 131414 66644
rect 139998 66632 140004 66644
rect 140056 66632 140062 66684
rect 226294 66360 226300 66412
rect 226352 66400 226358 66412
rect 229882 66400 229888 66412
rect 226352 66372 229888 66400
rect 226352 66360 226358 66372
rect 229882 66360 229888 66372
rect 229940 66360 229946 66412
rect 178454 66156 178460 66208
rect 178512 66196 178518 66208
rect 181766 66196 181772 66208
rect 178512 66168 181772 66196
rect 178512 66156 178518 66168
rect 181766 66156 181772 66168
rect 181824 66156 181830 66208
rect 321606 65816 321612 65868
rect 321664 65856 321670 65868
rect 326942 65856 326948 65868
rect 321664 65828 326948 65856
rect 321664 65816 321670 65828
rect 326942 65816 326948 65828
rect 327000 65816 327006 65868
rect 174038 65680 174044 65732
rect 174096 65720 174102 65732
rect 178730 65720 178736 65732
rect 174096 65692 178736 65720
rect 174096 65680 174102 65692
rect 178730 65680 178736 65692
rect 178788 65680 178794 65732
rect 321422 65680 321428 65732
rect 321480 65720 321486 65732
rect 326850 65720 326856 65732
rect 321480 65692 326856 65720
rect 321480 65680 321486 65692
rect 326850 65680 326856 65692
rect 326908 65680 326914 65732
rect 78910 65408 78916 65460
rect 78968 65448 78974 65460
rect 84430 65448 84436 65460
rect 78968 65420 84436 65448
rect 78968 65408 78974 65420
rect 84430 65408 84436 65420
rect 84488 65408 84494 65460
rect 229422 65408 229428 65460
rect 229480 65448 229486 65460
rect 233470 65448 233476 65460
rect 229480 65420 233476 65448
rect 229480 65408 229486 65420
rect 233470 65408 233476 65420
rect 233528 65408 233534 65460
rect 266590 65408 266596 65460
rect 266648 65448 266654 65460
rect 274962 65448 274968 65460
rect 266648 65420 274968 65448
rect 266648 65408 266654 65420
rect 274962 65408 274968 65420
rect 275020 65408 275026 65460
rect 321698 65408 321704 65460
rect 321756 65448 321762 65460
rect 328414 65448 328420 65460
rect 321756 65420 328420 65448
rect 321756 65408 321762 65420
rect 328414 65408 328420 65420
rect 328472 65408 328478 65460
rect 81670 65340 81676 65392
rect 81728 65380 81734 65392
rect 87190 65380 87196 65392
rect 81728 65352 87196 65380
rect 81728 65340 81734 65352
rect 87190 65340 87196 65352
rect 87248 65340 87254 65392
rect 131442 65340 131448 65392
rect 131500 65380 131506 65392
rect 136778 65380 136784 65392
rect 131500 65352 136784 65380
rect 131500 65340 131506 65352
rect 136778 65340 136784 65352
rect 136836 65340 136842 65392
rect 178270 65340 178276 65392
rect 178328 65380 178334 65392
rect 182318 65380 182324 65392
rect 178328 65352 182324 65380
rect 178328 65340 178334 65352
rect 182318 65340 182324 65352
rect 182376 65340 182382 65392
rect 225926 65340 225932 65392
rect 225984 65380 225990 65392
rect 233562 65380 233568 65392
rect 225984 65352 233568 65380
rect 225984 65340 225990 65352
rect 233562 65340 233568 65352
rect 233620 65340 233626 65392
rect 272478 65340 272484 65392
rect 272536 65380 272542 65392
rect 274870 65380 274876 65392
rect 272536 65352 274876 65380
rect 272536 65340 272542 65352
rect 274870 65340 274876 65352
rect 274928 65340 274934 65392
rect 85626 65272 85632 65324
rect 85684 65312 85690 65324
rect 87282 65312 87288 65324
rect 85684 65284 87288 65312
rect 85684 65272 85690 65284
rect 87282 65272 87288 65284
rect 87340 65272 87346 65324
rect 131350 65272 131356 65324
rect 131408 65312 131414 65324
rect 136686 65312 136692 65324
rect 131408 65284 136692 65312
rect 131408 65272 131414 65284
rect 136686 65272 136692 65284
rect 136744 65272 136750 65324
rect 175602 65272 175608 65324
rect 175660 65312 175666 65324
rect 181582 65312 181588 65324
rect 175660 65284 181588 65312
rect 175660 65272 175666 65284
rect 181582 65272 181588 65284
rect 181640 65272 181646 65324
rect 226202 65272 226208 65324
rect 226260 65312 226266 65324
rect 233654 65312 233660 65324
rect 226260 65284 233660 65312
rect 226260 65272 226266 65284
rect 233654 65272 233660 65284
rect 233712 65272 233718 65324
rect 272662 65272 272668 65324
rect 272720 65312 272726 65324
rect 275054 65312 275060 65324
rect 272720 65284 275060 65312
rect 272720 65272 272726 65284
rect 275054 65272 275060 65284
rect 275112 65272 275118 65324
rect 321422 65068 321428 65120
rect 321480 65108 321486 65120
rect 327678 65108 327684 65120
rect 321480 65080 327684 65108
rect 321480 65068 321486 65080
rect 327678 65068 327684 65080
rect 327736 65068 327742 65120
rect 321606 64728 321612 64780
rect 321664 64768 321670 64780
rect 327034 64768 327040 64780
rect 321664 64740 327040 64768
rect 321664 64728 321670 64740
rect 327034 64728 327040 64740
rect 327092 64728 327098 64780
rect 173118 64524 173124 64576
rect 173176 64564 173182 64576
rect 176062 64564 176068 64576
rect 173176 64536 176068 64564
rect 173176 64524 173182 64536
rect 176062 64524 176068 64536
rect 176120 64524 176126 64576
rect 78910 64456 78916 64508
rect 78968 64496 78974 64508
rect 81670 64496 81676 64508
rect 78968 64468 81676 64496
rect 78968 64456 78974 64468
rect 81670 64456 81676 64468
rect 81728 64456 81734 64508
rect 266590 64048 266596 64100
rect 266648 64088 266654 64100
rect 273030 64088 273036 64100
rect 266648 64060 273036 64088
rect 266648 64048 266654 64060
rect 273030 64048 273036 64060
rect 273088 64048 273094 64100
rect 132362 63980 132368 64032
rect 132420 64020 132426 64032
rect 136134 64020 136140 64032
rect 132420 63992 136140 64020
rect 132420 63980 132426 63992
rect 136134 63980 136140 63992
rect 136192 63980 136198 64032
rect 179098 63980 179104 64032
rect 179156 64020 179162 64032
rect 182318 64020 182324 64032
rect 179156 63992 182324 64020
rect 179156 63980 179162 63992
rect 182318 63980 182324 63992
rect 182376 63980 182382 64032
rect 225742 63980 225748 64032
rect 225800 64020 225806 64032
rect 230066 64020 230072 64032
rect 225800 63992 230072 64020
rect 225800 63980 225806 63992
rect 230066 63980 230072 63992
rect 230124 63980 230130 64032
rect 85166 63572 85172 63624
rect 85224 63612 85230 63624
rect 87190 63612 87196 63624
rect 85224 63584 87196 63612
rect 85224 63572 85230 63584
rect 87190 63572 87196 63584
rect 87248 63572 87254 63624
rect 272754 63572 272760 63624
rect 272812 63612 272818 63624
rect 274870 63612 274876 63624
rect 272812 63584 274876 63612
rect 272812 63572 272818 63584
rect 274870 63572 274876 63584
rect 274928 63572 274934 63624
rect 78910 62960 78916 63012
rect 78968 63000 78974 63012
rect 81762 63000 81768 63012
rect 78968 62972 81768 63000
rect 78968 62960 78974 62972
rect 81762 62960 81768 62972
rect 81820 62960 81826 63012
rect 174038 62688 174044 62740
rect 174096 62728 174102 62740
rect 178270 62728 178276 62740
rect 174096 62700 178276 62728
rect 174096 62688 174102 62700
rect 178270 62688 178276 62700
rect 178328 62688 178334 62740
rect 266682 62688 266688 62740
rect 266740 62728 266746 62740
rect 272754 62728 272760 62740
rect 266740 62700 272760 62728
rect 266740 62688 266746 62700
rect 272754 62688 272760 62700
rect 272812 62688 272818 62740
rect 78910 62620 78916 62672
rect 78968 62660 78974 62672
rect 87374 62660 87380 62672
rect 78968 62632 87380 62660
rect 78968 62620 78974 62632
rect 87374 62620 87380 62632
rect 87432 62620 87438 62672
rect 173486 62620 173492 62672
rect 173544 62660 173550 62672
rect 175602 62660 175608 62672
rect 173544 62632 175608 62660
rect 173544 62620 173550 62632
rect 175602 62620 175608 62632
rect 175660 62620 175666 62672
rect 230158 62620 230164 62672
rect 230216 62660 230222 62672
rect 233470 62660 233476 62672
rect 230216 62632 233476 62660
rect 230216 62620 230222 62632
rect 233470 62620 233476 62632
rect 233528 62620 233534 62672
rect 266590 62620 266596 62672
rect 266648 62660 266654 62672
rect 275054 62660 275060 62672
rect 266648 62632 275060 62660
rect 266648 62620 266654 62632
rect 275054 62620 275060 62632
rect 275112 62620 275118 62672
rect 81670 62552 81676 62604
rect 81728 62592 81734 62604
rect 87190 62592 87196 62604
rect 81728 62564 87196 62592
rect 81728 62552 81734 62564
rect 87190 62552 87196 62564
rect 87248 62552 87254 62604
rect 131718 62552 131724 62604
rect 131776 62592 131782 62604
rect 139630 62592 139636 62604
rect 131776 62564 139636 62592
rect 131776 62552 131782 62564
rect 139630 62552 139636 62564
rect 139688 62552 139694 62604
rect 176062 62552 176068 62604
rect 176120 62592 176126 62604
rect 181582 62592 181588 62604
rect 176120 62564 181588 62592
rect 176120 62552 176126 62564
rect 181582 62552 181588 62564
rect 181640 62552 181646 62604
rect 225926 62552 225932 62604
rect 225984 62592 225990 62604
rect 234574 62592 234580 62604
rect 225984 62564 234580 62592
rect 225984 62552 225990 62564
rect 234574 62552 234580 62564
rect 234632 62552 234638 62604
rect 273030 62552 273036 62604
rect 273088 62592 273094 62604
rect 274870 62592 274876 62604
rect 273088 62564 274876 62592
rect 273088 62552 273094 62564
rect 274870 62552 274876 62564
rect 274928 62552 274934 62604
rect 84430 62484 84436 62536
rect 84488 62524 84494 62536
rect 87282 62524 87288 62536
rect 84488 62496 87288 62524
rect 84488 62484 84494 62496
rect 87282 62484 87288 62496
rect 87340 62484 87346 62536
rect 131350 62484 131356 62536
rect 131408 62524 131414 62536
rect 139906 62524 139912 62536
rect 131408 62496 139912 62524
rect 131408 62484 131414 62496
rect 139906 62484 139912 62496
rect 139964 62484 139970 62536
rect 178730 62484 178736 62536
rect 178788 62524 178794 62536
rect 182318 62524 182324 62536
rect 178788 62496 182324 62524
rect 178788 62484 178794 62496
rect 182318 62484 182324 62496
rect 182376 62484 182382 62536
rect 226294 62348 226300 62400
rect 226352 62388 226358 62400
rect 229422 62388 229428 62400
rect 226352 62360 229428 62388
rect 226352 62348 226358 62360
rect 229422 62348 229428 62360
rect 229480 62348 229486 62400
rect 321238 62348 321244 62400
rect 321296 62388 321302 62400
rect 327310 62388 327316 62400
rect 321296 62360 327316 62388
rect 321296 62348 321302 62360
rect 327310 62348 327316 62360
rect 327368 62348 327374 62400
rect 173118 61600 173124 61652
rect 173176 61640 173182 61652
rect 175510 61640 175516 61652
rect 173176 61612 175516 61640
rect 173176 61600 173182 61612
rect 175510 61600 175516 61612
rect 175568 61600 175574 61652
rect 78910 61328 78916 61380
rect 78968 61368 78974 61380
rect 81670 61368 81676 61380
rect 78968 61340 81676 61368
rect 78968 61328 78974 61340
rect 81670 61328 81676 61340
rect 81728 61328 81734 61380
rect 266590 61260 266596 61312
rect 266648 61300 266654 61312
rect 272662 61300 272668 61312
rect 266648 61272 272668 61300
rect 266648 61260 266654 61272
rect 272662 61260 272668 61272
rect 272720 61260 272726 61312
rect 321054 61260 321060 61312
rect 321112 61300 321118 61312
rect 328506 61300 328512 61312
rect 321112 61272 328512 61300
rect 321112 61260 321118 61272
rect 328506 61260 328512 61272
rect 328564 61260 328570 61312
rect 81762 61192 81768 61244
rect 81820 61232 81826 61244
rect 87190 61232 87196 61244
rect 81820 61204 87196 61232
rect 81820 61192 81826 61204
rect 87190 61192 87196 61204
rect 87248 61192 87254 61244
rect 131350 61192 131356 61244
rect 131408 61232 131414 61244
rect 139722 61232 139728 61244
rect 131408 61204 139728 61232
rect 131408 61192 131414 61204
rect 139722 61192 139728 61204
rect 139780 61192 139786 61244
rect 175602 61192 175608 61244
rect 175660 61232 175666 61244
rect 181214 61232 181220 61244
rect 175660 61204 181220 61232
rect 175660 61192 175666 61204
rect 181214 61192 181220 61204
rect 181272 61192 181278 61244
rect 272754 61192 272760 61244
rect 272812 61232 272818 61244
rect 274870 61232 274876 61244
rect 272812 61204 274876 61232
rect 272812 61192 272818 61204
rect 274870 61192 274876 61204
rect 274928 61192 274934 61244
rect 226294 61056 226300 61108
rect 226352 61096 226358 61108
rect 230158 61096 230164 61108
rect 226352 61068 230164 61096
rect 226352 61056 226358 61068
rect 230158 61056 230164 61068
rect 230216 61056 230222 61108
rect 320870 60988 320876 61040
rect 320928 61028 320934 61040
rect 328046 61028 328052 61040
rect 320928 61000 328052 61028
rect 320928 60988 320934 61000
rect 328046 60988 328052 61000
rect 328104 60988 328110 61040
rect 78910 59900 78916 59952
rect 78968 59940 78974 59952
rect 85718 59940 85724 59952
rect 78968 59912 85724 59940
rect 78968 59900 78974 59912
rect 85718 59900 85724 59912
rect 85776 59900 85782 59952
rect 136778 59900 136784 59952
rect 136836 59940 136842 59952
rect 139722 59940 139728 59952
rect 136836 59912 139728 59940
rect 136836 59900 136842 59912
rect 139722 59900 139728 59912
rect 139780 59900 139786 59952
rect 173486 59900 173492 59952
rect 173544 59940 173550 59952
rect 175602 59940 175608 59952
rect 173544 59912 175608 59940
rect 173544 59900 173550 59912
rect 175602 59900 175608 59912
rect 175660 59900 175666 59952
rect 266590 59900 266596 59952
rect 266648 59940 266654 59952
rect 274962 59940 274968 59952
rect 266648 59912 274968 59940
rect 266648 59900 266654 59912
rect 274962 59900 274968 59912
rect 275020 59900 275026 59952
rect 369722 59900 369728 59952
rect 369780 59940 369786 59952
rect 369998 59940 370004 59952
rect 369780 59912 370004 59940
rect 369780 59900 369786 59912
rect 369998 59900 370004 59912
rect 370056 59900 370062 59952
rect 81670 59832 81676 59884
rect 81728 59872 81734 59884
rect 87190 59872 87196 59884
rect 81728 59844 87196 59872
rect 81728 59832 81734 59844
rect 87190 59832 87196 59844
rect 87248 59832 87254 59884
rect 132638 59832 132644 59884
rect 132696 59872 132702 59884
rect 139814 59872 139820 59884
rect 132696 59844 139820 59872
rect 132696 59832 132702 59844
rect 139814 59832 139820 59844
rect 139872 59832 139878 59884
rect 175510 59832 175516 59884
rect 175568 59872 175574 59884
rect 181582 59872 181588 59884
rect 175568 59844 181588 59872
rect 175568 59832 175574 59844
rect 181582 59832 181588 59844
rect 181640 59832 181646 59884
rect 226110 59832 226116 59884
rect 226168 59872 226174 59884
rect 233562 59872 233568 59884
rect 226168 59844 233568 59872
rect 226168 59832 226174 59844
rect 233562 59832 233568 59844
rect 233620 59832 233626 59884
rect 272662 59832 272668 59884
rect 272720 59872 272726 59884
rect 274870 59872 274876 59884
rect 272720 59844 274876 59872
rect 272720 59832 272726 59844
rect 274870 59832 274876 59844
rect 274928 59832 274934 59884
rect 369262 59832 369268 59884
rect 369320 59872 369326 59884
rect 369814 59872 369820 59884
rect 369320 59844 369820 59872
rect 369320 59832 369326 59844
rect 369814 59832 369820 59844
rect 369872 59832 369878 59884
rect 132546 59764 132552 59816
rect 132604 59804 132610 59816
rect 139630 59804 139636 59816
rect 132604 59776 139636 59804
rect 132604 59764 132610 59776
rect 139630 59764 139636 59776
rect 139688 59764 139694 59816
rect 178270 59764 178276 59816
rect 178328 59804 178334 59816
rect 182318 59804 182324 59816
rect 178328 59776 182324 59804
rect 178328 59764 178334 59776
rect 182318 59764 182324 59776
rect 182376 59764 182382 59816
rect 226294 59764 226300 59816
rect 226352 59804 226358 59816
rect 233470 59804 233476 59816
rect 226352 59776 233476 59804
rect 226352 59764 226358 59776
rect 233470 59764 233476 59776
rect 233528 59764 233534 59816
rect 321606 58744 321612 58796
rect 321664 58784 321670 58796
rect 328322 58784 328328 58796
rect 321664 58756 328328 58784
rect 321664 58744 321670 58756
rect 328322 58744 328328 58756
rect 328380 58744 328386 58796
rect 135490 58608 135496 58660
rect 135548 58648 135554 58660
rect 139722 58648 139728 58660
rect 135548 58620 139728 58648
rect 135548 58608 135554 58620
rect 139722 58608 139728 58620
rect 139780 58608 139786 58660
rect 230342 58608 230348 58660
rect 230400 58648 230406 58660
rect 233562 58648 233568 58660
rect 230400 58620 233568 58648
rect 230400 58608 230406 58620
rect 233562 58608 233568 58620
rect 233620 58608 233626 58660
rect 266590 58608 266596 58660
rect 266648 58648 266654 58660
rect 272570 58648 272576 58660
rect 266648 58620 272576 58648
rect 266648 58608 266654 58620
rect 272570 58608 272576 58620
rect 272628 58608 272634 58660
rect 136410 58540 136416 58592
rect 136468 58580 136474 58592
rect 139630 58580 139636 58592
rect 136468 58552 139636 58580
rect 136468 58540 136474 58552
rect 139630 58540 139636 58552
rect 139688 58540 139694 58592
rect 230618 58540 230624 58592
rect 230676 58580 230682 58592
rect 233470 58580 233476 58592
rect 230676 58552 233476 58580
rect 230676 58540 230682 58552
rect 233470 58540 233476 58552
rect 233528 58540 233534 58592
rect 266682 58540 266688 58592
rect 266740 58580 266746 58592
rect 272754 58580 272760 58592
rect 266740 58552 272760 58580
rect 266740 58540 266746 58552
rect 272754 58540 272760 58552
rect 272812 58540 272818 58592
rect 85718 58472 85724 58524
rect 85776 58512 85782 58524
rect 87190 58512 87196 58524
rect 85776 58484 87196 58512
rect 85776 58472 85782 58484
rect 87190 58472 87196 58484
rect 87248 58472 87254 58524
rect 132638 58472 132644 58524
rect 132696 58512 132702 58524
rect 136778 58512 136784 58524
rect 132696 58484 136784 58512
rect 132696 58472 132702 58484
rect 136778 58472 136784 58484
rect 136836 58472 136842 58524
rect 175602 58472 175608 58524
rect 175660 58512 175666 58524
rect 182318 58512 182324 58524
rect 175660 58484 182324 58512
rect 175660 58472 175666 58484
rect 182318 58472 182324 58484
rect 182376 58472 182382 58524
rect 226294 58472 226300 58524
rect 226352 58512 226358 58524
rect 233654 58512 233660 58524
rect 226352 58484 233660 58512
rect 226352 58472 226358 58484
rect 233654 58472 233660 58484
rect 233712 58472 233718 58524
rect 173486 57384 173492 57436
rect 173544 57424 173550 57436
rect 176246 57424 176252 57436
rect 173544 57396 176252 57424
rect 173544 57384 173550 57396
rect 176246 57384 176252 57396
rect 176304 57384 176310 57436
rect 320870 57180 320876 57232
rect 320928 57220 320934 57232
rect 328414 57220 328420 57232
rect 320928 57192 328420 57220
rect 320928 57180 320934 57192
rect 328414 57180 328420 57192
rect 328472 57180 328478 57232
rect 78910 57112 78916 57164
rect 78968 57152 78974 57164
rect 87374 57152 87380 57164
rect 78968 57124 87380 57152
rect 78968 57112 78974 57124
rect 87374 57112 87380 57124
rect 87432 57112 87438 57164
rect 129421 57155 129479 57161
rect 129421 57121 129433 57155
rect 129467 57152 129479 57155
rect 129510 57152 129516 57164
rect 129467 57124 129516 57152
rect 129467 57121 129479 57124
rect 129421 57115 129479 57121
rect 129510 57112 129516 57124
rect 129568 57112 129574 57164
rect 266590 57112 266596 57164
rect 266648 57152 266654 57164
rect 274962 57152 274968 57164
rect 266648 57124 274968 57152
rect 266648 57112 266654 57124
rect 274962 57112 274968 57124
rect 275020 57112 275026 57164
rect 80382 57044 80388 57096
rect 80440 57084 80446 57096
rect 87190 57084 87196 57096
rect 80440 57056 87196 57084
rect 80440 57044 80446 57056
rect 87190 57044 87196 57056
rect 87248 57044 87254 57096
rect 132638 57044 132644 57096
rect 132696 57084 132702 57096
rect 135490 57084 135496 57096
rect 132696 57056 135496 57084
rect 132696 57044 132702 57056
rect 135490 57044 135496 57056
rect 135548 57044 135554 57096
rect 272754 57044 272760 57096
rect 272812 57084 272818 57096
rect 274870 57084 274876 57096
rect 272812 57056 274876 57084
rect 272812 57044 272818 57056
rect 274870 57044 274876 57056
rect 274928 57044 274934 57096
rect 80290 56976 80296 57028
rect 80348 57016 80354 57028
rect 87282 57016 87288 57028
rect 80348 56988 87288 57016
rect 80348 56976 80354 56988
rect 87282 56976 87288 56988
rect 87340 56976 87346 57028
rect 132546 56976 132552 57028
rect 132604 57016 132610 57028
rect 136410 57016 136416 57028
rect 132604 56988 136416 57016
rect 132604 56976 132610 56988
rect 136410 56976 136416 56988
rect 136468 56976 136474 57028
rect 272570 56976 272576 57028
rect 272628 57016 272634 57028
rect 275054 57016 275060 57028
rect 272628 56988 275060 57016
rect 272628 56976 272634 56988
rect 275054 56976 275060 56988
rect 275112 56976 275118 57028
rect 226294 56908 226300 56960
rect 226352 56948 226358 56960
rect 230342 56948 230348 56960
rect 226352 56920 230348 56948
rect 226352 56908 226358 56920
rect 230342 56908 230348 56920
rect 230400 56908 230406 56960
rect 225374 56636 225380 56688
rect 225432 56676 225438 56688
rect 230618 56676 230624 56688
rect 225432 56648 230624 56676
rect 225432 56636 225438 56648
rect 230618 56636 230624 56648
rect 230676 56636 230682 56688
rect 174130 56568 174136 56620
rect 174188 56608 174194 56620
rect 181766 56608 181772 56620
rect 174188 56580 181772 56608
rect 174188 56568 174194 56580
rect 181766 56568 181772 56580
rect 181824 56568 181830 56620
rect 174222 56432 174228 56484
rect 174280 56472 174286 56484
rect 182318 56472 182324 56484
rect 174280 56444 182324 56472
rect 174280 56432 174286 56444
rect 182318 56432 182324 56444
rect 182376 56432 182382 56484
rect 321606 56296 321612 56348
rect 321664 56336 321670 56348
rect 327678 56336 327684 56348
rect 321664 56308 327684 56336
rect 321664 56296 321670 56308
rect 327678 56296 327684 56308
rect 327736 56296 327742 56348
rect 321054 56024 321060 56076
rect 321112 56064 321118 56076
rect 328506 56064 328512 56076
rect 321112 56036 328512 56064
rect 321112 56024 321118 56036
rect 328506 56024 328512 56036
rect 328564 56024 328570 56076
rect 78910 55752 78916 55804
rect 78968 55792 78974 55804
rect 81670 55792 81676 55804
rect 78968 55764 81676 55792
rect 78968 55752 78974 55764
rect 81670 55752 81676 55764
rect 81728 55752 81734 55804
rect 172750 55752 172756 55804
rect 172808 55792 172814 55804
rect 176798 55792 176804 55804
rect 172808 55764 176804 55792
rect 172808 55752 172814 55764
rect 176798 55752 176804 55764
rect 176856 55752 176862 55804
rect 266590 55752 266596 55804
rect 266648 55792 266654 55804
rect 273398 55792 273404 55804
rect 266648 55764 273404 55792
rect 266648 55752 266654 55764
rect 273398 55752 273404 55764
rect 273456 55752 273462 55804
rect 324550 55752 324556 55804
rect 324608 55792 324614 55804
rect 327494 55792 327500 55804
rect 324608 55764 327500 55792
rect 324608 55752 324614 55764
rect 327494 55752 327500 55764
rect 327552 55752 327558 55804
rect 132638 55684 132644 55736
rect 132696 55724 132702 55736
rect 139630 55724 139636 55736
rect 132696 55696 139636 55724
rect 132696 55684 132702 55696
rect 139630 55684 139636 55696
rect 139688 55684 139694 55736
rect 176246 55684 176252 55736
rect 176304 55724 176310 55736
rect 181674 55724 181680 55736
rect 176304 55696 181680 55724
rect 176304 55684 176310 55696
rect 181674 55684 181680 55696
rect 181732 55684 181738 55736
rect 225374 55684 225380 55736
rect 225432 55724 225438 55736
rect 233470 55724 233476 55736
rect 225432 55696 233476 55724
rect 225432 55684 225438 55696
rect 233470 55684 233476 55696
rect 233528 55684 233534 55736
rect 134202 55112 134208 55124
rect 134036 55084 134208 55112
rect 134036 55053 134064 55084
rect 134202 55072 134208 55084
rect 134260 55072 134266 55124
rect 369722 55072 369728 55124
rect 369780 55112 369786 55124
rect 369998 55112 370004 55124
rect 369780 55084 370004 55112
rect 369780 55072 369786 55084
rect 369998 55072 370004 55084
rect 370056 55072 370062 55124
rect 134021 55047 134079 55053
rect 134021 55013 134033 55047
rect 134067 55013 134079 55047
rect 134021 55007 134079 55013
rect 223442 55004 223448 55056
rect 223500 55044 223506 55056
rect 233470 55044 233476 55056
rect 223500 55016 233476 55044
rect 223500 55004 223506 55016
rect 233470 55004 233476 55016
rect 233528 55004 233534 55056
rect 317466 55004 317472 55056
rect 317524 55044 317530 55056
rect 328506 55044 328512 55056
rect 317524 55016 328512 55044
rect 317524 55004 317530 55016
rect 328506 55004 328512 55016
rect 328564 55004 328570 55056
rect 358498 55004 358504 55056
rect 358556 55044 358562 55056
rect 389410 55044 389416 55056
rect 358556 55016 389416 55044
rect 358556 55004 358562 55016
rect 389410 55004 389416 55016
rect 389468 55004 389474 55056
rect 321606 54936 321612 54988
rect 321664 54976 321670 54988
rect 328322 54976 328328 54988
rect 321664 54948 328328 54976
rect 321664 54936 321670 54948
rect 328322 54936 328328 54948
rect 328380 54936 328386 54988
rect 129510 54868 129516 54920
rect 129568 54908 129574 54920
rect 134021 54911 134079 54917
rect 134021 54908 134033 54911
rect 129568 54880 134033 54908
rect 129568 54868 129574 54880
rect 134021 54877 134033 54880
rect 134067 54877 134079 54911
rect 134021 54871 134079 54877
rect 78910 54392 78916 54444
rect 78968 54432 78974 54444
rect 87282 54432 87288 54444
rect 78968 54404 87288 54432
rect 78968 54392 78974 54404
rect 87282 54392 87288 54404
rect 87340 54392 87346 54444
rect 134110 54392 134116 54444
rect 134168 54432 134174 54444
rect 139630 54432 139636 54444
rect 134168 54404 139636 54432
rect 134168 54392 134174 54404
rect 139630 54392 139636 54404
rect 139688 54392 139694 54444
rect 174038 54392 174044 54444
rect 174096 54432 174102 54444
rect 233470 54432 233476 54444
rect 174096 54404 181076 54432
rect 174096 54392 174102 54404
rect 81670 54324 81676 54376
rect 81728 54364 81734 54376
rect 87190 54364 87196 54376
rect 81728 54336 87196 54364
rect 81728 54324 81734 54336
rect 87190 54324 87196 54336
rect 87248 54324 87254 54376
rect 132638 54324 132644 54376
rect 132696 54364 132702 54376
rect 139538 54364 139544 54376
rect 132696 54336 139544 54364
rect 132696 54324 132702 54336
rect 139538 54324 139544 54336
rect 139596 54324 139602 54376
rect 181048 54296 181076 54404
rect 223736 54404 233476 54432
rect 223534 54324 223540 54376
rect 223592 54364 223598 54376
rect 223736 54364 223764 54404
rect 233470 54392 233476 54404
rect 233528 54392 233534 54444
rect 266590 54392 266596 54444
rect 266648 54432 266654 54444
rect 317466 54432 317472 54444
rect 266648 54404 275560 54432
rect 266648 54392 266654 54404
rect 223592 54336 223764 54364
rect 223592 54324 223598 54336
rect 226294 54324 226300 54376
rect 226352 54364 226358 54376
rect 234390 54364 234396 54376
rect 226352 54336 234396 54364
rect 226352 54324 226358 54336
rect 234390 54324 234396 54336
rect 234448 54324 234454 54376
rect 273398 54324 273404 54376
rect 273456 54364 273462 54376
rect 274870 54364 274876 54376
rect 273456 54336 274876 54364
rect 273456 54324 273462 54336
rect 274870 54324 274876 54336
rect 274928 54324 274934 54376
rect 223552 54296 223580 54324
rect 181048 54268 223580 54296
rect 275532 54296 275560 54404
rect 316748 54404 317472 54432
rect 316748 54296 316776 54404
rect 317466 54392 317472 54404
rect 317524 54432 317530 54444
rect 328414 54432 328420 54444
rect 317524 54404 328420 54432
rect 317524 54392 317530 54404
rect 328414 54392 328420 54404
rect 328472 54392 328478 54444
rect 320962 54324 320968 54376
rect 321020 54364 321026 54376
rect 324550 54364 324556 54376
rect 321020 54336 324556 54364
rect 321020 54324 321026 54336
rect 324550 54324 324556 54336
rect 324608 54324 324614 54376
rect 275532 54268 316776 54296
rect 176798 54188 176804 54240
rect 176856 54228 176862 54240
rect 182318 54228 182324 54240
rect 176856 54200 182324 54228
rect 176856 54188 176862 54200
rect 182318 54188 182324 54200
rect 182376 54188 182382 54240
rect 78910 53712 78916 53764
rect 78968 53752 78974 53764
rect 118194 53752 118200 53764
rect 78968 53724 118200 53752
rect 78968 53712 78974 53724
rect 118194 53712 118200 53724
rect 118252 53752 118258 53764
rect 139630 53752 139636 53764
rect 118252 53724 139636 53752
rect 118252 53712 118258 53724
rect 139630 53712 139636 53724
rect 139688 53712 139694 53764
rect 87282 53644 87288 53696
rect 87340 53684 87346 53696
rect 128682 53684 128688 53696
rect 87340 53656 128688 53684
rect 87340 53644 87346 53656
rect 128682 53644 128688 53656
rect 128740 53684 128746 53696
rect 134110 53684 134116 53696
rect 128740 53656 134116 53684
rect 128740 53644 128746 53656
rect 134110 53644 134116 53656
rect 134168 53644 134174 53696
rect 174038 53644 174044 53696
rect 174096 53684 174102 53696
rect 212034 53684 212040 53696
rect 174096 53656 212040 53684
rect 174096 53644 174102 53656
rect 212034 53644 212040 53656
rect 212092 53684 212098 53696
rect 233470 53684 233476 53696
rect 212092 53656 233476 53684
rect 212092 53644 212098 53656
rect 233470 53644 233476 53656
rect 233528 53644 233534 53696
rect 266590 53644 266596 53696
rect 266648 53684 266654 53696
rect 306978 53684 306984 53696
rect 266648 53656 306984 53684
rect 266648 53644 266654 53656
rect 306978 53644 306984 53656
rect 307036 53684 307042 53696
rect 328414 53684 328420 53696
rect 307036 53656 328420 53684
rect 307036 53644 307042 53656
rect 328414 53644 328420 53656
rect 328472 53644 328478 53696
rect 129050 52284 129056 52336
rect 129108 52324 129114 52336
rect 129510 52324 129516 52336
rect 129108 52296 129516 52324
rect 129108 52284 129114 52296
rect 129510 52284 129516 52296
rect 129568 52284 129574 52336
rect 91238 51536 91244 51588
rect 91296 51576 91302 51588
rect 134754 51576 134760 51588
rect 91296 51548 134760 51576
rect 91296 51536 91302 51548
rect 134754 51536 134760 51548
rect 134812 51536 134818 51588
rect 184986 51536 184992 51588
rect 185044 51576 185050 51588
rect 228594 51576 228600 51588
rect 185044 51548 228600 51576
rect 185044 51536 185050 51548
rect 228594 51536 228600 51548
rect 228652 51536 228658 51588
rect 279010 51536 279016 51588
rect 279068 51576 279074 51588
rect 323814 51576 323820 51588
rect 279068 51548 323820 51576
rect 279068 51536 279074 51548
rect 323814 51536 323820 51548
rect 323872 51536 323878 51588
rect 427590 51536 427596 51588
rect 427648 51576 427654 51588
rect 429798 51576 429804 51588
rect 427648 51548 429804 51576
rect 427648 51536 427654 51548
rect 429798 51536 429804 51548
rect 429856 51536 429862 51588
rect 78174 51468 78180 51520
rect 78232 51508 78238 51520
rect 93630 51508 93636 51520
rect 78232 51480 93636 51508
rect 78232 51468 78238 51480
rect 93630 51468 93636 51480
rect 93688 51468 93694 51520
rect 170174 51468 170180 51520
rect 170232 51508 170238 51520
rect 170634 51508 170640 51520
rect 170232 51480 170640 51508
rect 170232 51468 170238 51480
rect 170634 51468 170640 51480
rect 170692 51508 170698 51520
rect 189678 51508 189684 51520
rect 170692 51480 189684 51508
rect 170692 51468 170698 51480
rect 189678 51468 189684 51480
rect 189736 51468 189742 51520
rect 111938 51128 111944 51180
rect 111996 51168 112002 51180
rect 121230 51168 121236 51180
rect 111996 51140 121236 51168
rect 111996 51128 112002 51140
rect 121230 51128 121236 51140
rect 121288 51128 121294 51180
rect 205778 51128 205784 51180
rect 205836 51168 205842 51180
rect 215530 51168 215536 51180
rect 205836 51140 215536 51168
rect 205836 51128 205842 51140
rect 215530 51128 215536 51140
rect 215588 51128 215594 51180
rect 299618 51128 299624 51180
rect 299676 51168 299682 51180
rect 309554 51168 309560 51180
rect 299676 51140 309560 51168
rect 299676 51128 299682 51140
rect 309554 51128 309560 51140
rect 309612 51128 309618 51180
rect 106418 51060 106424 51112
rect 106476 51100 106482 51112
rect 118930 51100 118936 51112
rect 106476 51072 118936 51100
rect 106476 51060 106482 51072
rect 118930 51060 118936 51072
rect 118988 51060 118994 51112
rect 200258 51060 200264 51112
rect 200316 51100 200322 51112
rect 213230 51100 213236 51112
rect 200316 51072 213236 51100
rect 200316 51060 200322 51072
rect 213230 51060 213236 51072
rect 213288 51060 213294 51112
rect 294098 51060 294104 51112
rect 294156 51100 294162 51112
rect 307254 51100 307260 51112
rect 294156 51072 307260 51100
rect 294156 51060 294162 51072
rect 307254 51060 307260 51072
rect 307312 51060 307318 51112
rect 102278 50992 102284 51044
rect 102336 51032 102342 51044
rect 116538 51032 116544 51044
rect 102336 51004 116544 51032
rect 102336 50992 102342 51004
rect 116538 50992 116544 51004
rect 116596 50992 116602 51044
rect 196118 50992 196124 51044
rect 196176 51032 196182 51044
rect 210838 51032 210844 51044
rect 196176 51004 210844 51032
rect 196176 50992 196182 51004
rect 210838 50992 210844 51004
rect 210896 50992 210902 51044
rect 289958 50992 289964 51044
rect 290016 51032 290022 51044
rect 304862 51032 304868 51044
rect 290016 51004 304868 51032
rect 290016 50992 290022 51004
rect 304862 50992 304868 51004
rect 304920 50992 304926 51044
rect 96761 50967 96819 50973
rect 96761 50933 96773 50967
rect 96807 50964 96819 50967
rect 114146 50964 114152 50976
rect 96807 50936 114152 50964
rect 96807 50933 96819 50936
rect 96761 50927 96819 50933
rect 114146 50924 114152 50936
rect 114204 50924 114210 50976
rect 122334 50924 122340 50976
rect 122392 50964 122398 50976
rect 125922 50964 125928 50976
rect 122392 50936 125928 50964
rect 122392 50924 122398 50936
rect 125922 50924 125928 50936
rect 125980 50924 125986 50976
rect 190598 50924 190604 50976
rect 190656 50964 190662 50976
rect 208446 50964 208452 50976
rect 190656 50936 208452 50964
rect 190656 50924 190662 50936
rect 208446 50924 208452 50936
rect 208504 50924 208510 50976
rect 284438 50924 284444 50976
rect 284496 50964 284502 50976
rect 302470 50964 302476 50976
rect 284496 50936 302476 50964
rect 284496 50924 284502 50936
rect 302470 50924 302476 50936
rect 302528 50924 302534 50976
rect 91238 50856 91244 50908
rect 91296 50896 91302 50908
rect 112030 50896 112036 50908
rect 91296 50868 112036 50896
rect 91296 50856 91302 50868
rect 112030 50856 112036 50868
rect 112088 50856 112094 50908
rect 116078 50856 116084 50908
rect 116136 50896 116142 50908
rect 123622 50896 123628 50908
rect 116136 50868 123628 50896
rect 116136 50856 116142 50868
rect 123622 50856 123628 50868
rect 123680 50856 123686 50908
rect 185078 50856 185084 50908
rect 185136 50896 185142 50908
rect 206146 50896 206152 50908
rect 185136 50868 206152 50896
rect 185136 50856 185142 50868
rect 206146 50856 206152 50868
rect 206204 50856 206210 50908
rect 280298 50856 280304 50908
rect 280356 50896 280362 50908
rect 300170 50896 300176 50908
rect 280356 50868 300176 50896
rect 280356 50856 280362 50868
rect 300170 50856 300176 50868
rect 300228 50856 300234 50908
rect 305138 50856 305144 50908
rect 305196 50896 305202 50908
rect 311946 50896 311952 50908
rect 305196 50868 311952 50896
rect 305196 50856 305202 50868
rect 311946 50856 311952 50868
rect 312004 50856 312010 50908
rect 216174 50652 216180 50704
rect 216232 50692 216238 50704
rect 220222 50692 220228 50704
rect 216232 50664 220228 50692
rect 216232 50652 216238 50664
rect 220222 50652 220228 50664
rect 220280 50652 220286 50704
rect 211298 50380 211304 50432
rect 211356 50420 211362 50432
rect 217922 50420 217928 50432
rect 211356 50392 217928 50420
rect 211356 50380 211362 50392
rect 217922 50380 217928 50392
rect 217980 50380 217986 50432
rect 310014 50380 310020 50432
rect 310072 50420 310078 50432
rect 314246 50420 314252 50432
rect 310072 50392 314252 50420
rect 310072 50380 310078 50392
rect 314246 50380 314252 50392
rect 314304 50380 314310 50432
rect 79002 50312 79008 50364
rect 79060 50352 79066 50364
rect 108626 50352 108632 50364
rect 79060 50324 108632 50352
rect 79060 50312 79066 50324
rect 108626 50312 108632 50324
rect 108684 50352 108690 50364
rect 139722 50352 139728 50364
rect 108684 50324 139728 50352
rect 108684 50312 108690 50324
rect 139722 50312 139728 50324
rect 139780 50312 139786 50364
rect 173946 50312 173952 50364
rect 174004 50352 174010 50364
rect 202558 50352 202564 50364
rect 174004 50324 202564 50352
rect 174004 50312 174010 50324
rect 202558 50312 202564 50324
rect 202616 50352 202622 50364
rect 233562 50352 233568 50364
rect 202616 50324 233568 50352
rect 202616 50312 202622 50324
rect 233562 50312 233568 50324
rect 233620 50312 233626 50364
rect 266682 50312 266688 50364
rect 266740 50352 266746 50364
rect 296582 50352 296588 50364
rect 266740 50324 296588 50352
rect 266740 50312 266746 50324
rect 296582 50312 296588 50324
rect 296640 50352 296646 50364
rect 327678 50352 327684 50364
rect 296640 50324 327684 50352
rect 296640 50312 296646 50324
rect 327678 50312 327684 50324
rect 327736 50312 327742 50364
rect 78910 50244 78916 50296
rect 78968 50284 78974 50296
rect 103566 50284 103572 50296
rect 78968 50256 103572 50284
rect 78968 50244 78974 50256
rect 103566 50244 103572 50256
rect 103624 50284 103630 50296
rect 139630 50284 139636 50296
rect 103624 50256 139636 50284
rect 103624 50244 103630 50256
rect 139630 50244 139636 50256
rect 139688 50244 139694 50296
rect 174038 50244 174044 50296
rect 174096 50284 174102 50296
rect 197498 50284 197504 50296
rect 174096 50256 197504 50284
rect 174096 50244 174102 50256
rect 197498 50244 197504 50256
rect 197556 50284 197562 50296
rect 233470 50284 233476 50296
rect 197556 50256 233476 50284
rect 197556 50244 197562 50256
rect 233470 50244 233476 50256
rect 233528 50244 233534 50296
rect 266590 50244 266596 50296
rect 266648 50284 266654 50296
rect 291522 50284 291528 50296
rect 266648 50256 291528 50284
rect 266648 50244 266654 50256
rect 291522 50244 291528 50256
rect 291580 50284 291586 50296
rect 328414 50284 328420 50296
rect 291580 50256 328420 50284
rect 291580 50244 291586 50256
rect 328414 50244 328420 50256
rect 328472 50244 328478 50296
rect 288302 50176 288308 50228
rect 288360 50216 288366 50228
rect 327218 50216 327224 50228
rect 288360 50188 327224 50216
rect 288360 50176 288366 50188
rect 327218 50176 327224 50188
rect 327276 50176 327282 50228
rect 274962 49564 274968 49616
rect 275020 49604 275026 49616
rect 275606 49604 275612 49616
rect 275020 49576 275612 49604
rect 275020 49564 275026 49576
rect 275606 49564 275612 49576
rect 275664 49604 275670 49616
rect 288302 49604 288308 49616
rect 275664 49576 288308 49604
rect 275664 49564 275670 49576
rect 288302 49564 288308 49576
rect 288360 49564 288366 49616
rect 87466 49496 87472 49548
rect 87524 49536 87530 49548
rect 88386 49536 88392 49548
rect 87524 49508 88392 49536
rect 87524 49496 87530 49508
rect 88386 49496 88392 49508
rect 88444 49536 88450 49548
rect 102370 49536 102376 49548
rect 88444 49508 102376 49536
rect 88444 49496 88450 49508
rect 102370 49496 102376 49508
rect 102428 49496 102434 49548
rect 181858 49496 181864 49548
rect 181916 49536 181922 49548
rect 194370 49536 194376 49548
rect 181916 49508 194376 49536
rect 181916 49496 181922 49508
rect 194370 49496 194376 49508
rect 194428 49496 194434 49548
rect 275054 49496 275060 49548
rect 275112 49536 275118 49548
rect 275882 49536 275888 49548
rect 275112 49508 275888 49536
rect 275112 49496 275118 49508
rect 275882 49496 275888 49508
rect 275940 49536 275946 49548
rect 297778 49536 297784 49548
rect 275940 49508 297784 49536
rect 275940 49496 275946 49508
rect 297778 49496 297784 49508
rect 297836 49536 297842 49548
rect 357305 49539 357363 49545
rect 357305 49536 357317 49539
rect 297836 49508 357317 49536
rect 297836 49496 297842 49508
rect 357305 49505 357317 49508
rect 357351 49505 357363 49539
rect 357305 49499 357363 49505
rect 78910 48884 78916 48936
rect 78968 48924 78974 48936
rect 98598 48924 98604 48936
rect 78968 48896 98604 48924
rect 78968 48884 78974 48896
rect 98598 48884 98604 48896
rect 98656 48924 98662 48936
rect 140550 48924 140556 48936
rect 98656 48896 140556 48924
rect 98656 48884 98662 48896
rect 140550 48884 140556 48896
rect 140608 48884 140614 48936
rect 173302 48884 173308 48936
rect 173360 48924 173366 48936
rect 192530 48924 192536 48936
rect 173360 48896 192536 48924
rect 173360 48884 173366 48896
rect 192530 48884 192536 48896
rect 192588 48924 192594 48936
rect 233470 48924 233476 48936
rect 192588 48896 233476 48924
rect 192588 48884 192594 48896
rect 233470 48884 233476 48896
rect 233528 48884 233534 48936
rect 266590 48884 266596 48936
rect 266648 48924 266654 48936
rect 286554 48924 286560 48936
rect 266648 48896 286560 48924
rect 266648 48884 266654 48896
rect 286554 48884 286560 48896
rect 286612 48924 286618 48936
rect 328506 48924 328512 48936
rect 286612 48896 328512 48924
rect 286612 48884 286618 48896
rect 328506 48884 328512 48896
rect 328564 48884 328570 48936
rect 357305 48927 357363 48933
rect 357305 48893 357317 48927
rect 357351 48924 357363 48927
rect 359694 48924 359700 48936
rect 357351 48896 359700 48924
rect 357351 48893 357363 48896
rect 357305 48887 357363 48893
rect 359694 48884 359700 48896
rect 359752 48884 359758 48936
rect 96758 48516 96764 48528
rect 96719 48488 96764 48516
rect 96758 48476 96764 48488
rect 96816 48476 96822 48528
rect 182226 48136 182232 48188
rect 182284 48176 182290 48188
rect 196670 48176 196676 48188
rect 182284 48148 196676 48176
rect 182284 48136 182290 48148
rect 196670 48136 196676 48148
rect 196728 48136 196734 48188
rect 275790 48136 275796 48188
rect 275848 48176 275854 48188
rect 276066 48176 276072 48188
rect 275848 48148 276072 48176
rect 275848 48136 275854 48148
rect 276066 48136 276072 48148
rect 276124 48176 276130 48188
rect 290694 48176 290700 48188
rect 276124 48148 290700 48176
rect 276124 48136 276130 48148
rect 290694 48136 290700 48148
rect 290752 48136 290758 48188
rect 357302 48176 357308 48188
rect 357263 48148 357308 48176
rect 357302 48136 357308 48148
rect 357360 48136 357366 48188
rect 124453 47771 124511 47777
rect 124453 47737 124465 47771
rect 124499 47768 124511 47771
rect 134021 47771 134079 47777
rect 134021 47768 134033 47771
rect 124499 47740 134033 47768
rect 124499 47737 124511 47740
rect 124453 47731 124511 47737
rect 134021 47737 134033 47740
rect 134067 47737 134079 47771
rect 134021 47731 134079 47737
rect 109365 47703 109423 47709
rect 109365 47669 109377 47703
rect 109411 47700 109423 47703
rect 139998 47700 140004 47712
rect 109411 47672 118792 47700
rect 109411 47669 109423 47672
rect 109365 47663 109423 47669
rect 105041 47635 105099 47641
rect 105041 47601 105053 47635
rect 105087 47632 105099 47635
rect 109181 47635 109239 47641
rect 109181 47632 109193 47635
rect 105087 47604 109193 47632
rect 105087 47601 105099 47604
rect 105041 47595 105099 47601
rect 109181 47601 109193 47604
rect 109227 47601 109239 47635
rect 118764 47632 118792 47672
rect 138176 47672 140004 47700
rect 124453 47635 124511 47641
rect 124453 47632 124465 47635
rect 118764 47604 124465 47632
rect 109181 47595 109239 47601
rect 124453 47601 124465 47604
rect 124499 47601 124511 47635
rect 124453 47595 124511 47601
rect 134021 47635 134079 47641
rect 134021 47601 134033 47635
rect 134067 47632 134079 47635
rect 138176 47632 138204 47672
rect 139998 47660 140004 47672
rect 140056 47660 140062 47712
rect 134067 47604 138204 47632
rect 134067 47601 134079 47604
rect 134021 47595 134079 47601
rect 95105 47567 95163 47573
rect 95105 47533 95117 47567
rect 95151 47564 95163 47567
rect 95473 47567 95531 47573
rect 95473 47564 95485 47567
rect 95151 47536 95485 47564
rect 95151 47533 95163 47536
rect 95105 47527 95163 47533
rect 95473 47533 95485 47536
rect 95519 47533 95531 47567
rect 95473 47527 95531 47533
rect 142850 47524 142856 47576
rect 142908 47564 142914 47576
rect 159502 47564 159508 47576
rect 142908 47536 159508 47564
rect 142908 47524 142914 47536
rect 159502 47524 159508 47536
rect 159560 47524 159566 47576
rect 100438 47456 100444 47508
rect 100496 47496 100502 47508
rect 100898 47496 100904 47508
rect 100496 47468 100904 47496
rect 100496 47456 100502 47468
rect 100898 47456 100904 47468
rect 100956 47496 100962 47508
rect 156834 47496 156840 47508
rect 100956 47468 156840 47496
rect 100956 47456 100962 47468
rect 156834 47456 156840 47468
rect 156892 47496 156898 47508
rect 167598 47496 167604 47508
rect 156892 47468 167604 47496
rect 156892 47456 156898 47468
rect 167598 47456 167604 47468
rect 167656 47456 167662 47508
rect 174038 47456 174044 47508
rect 174096 47496 174102 47508
rect 187562 47496 187568 47508
rect 174096 47468 187568 47496
rect 174096 47456 174102 47468
rect 187562 47456 187568 47468
rect 187620 47496 187626 47508
rect 233470 47496 233476 47508
rect 187620 47468 233476 47496
rect 187620 47456 187626 47468
rect 233470 47456 233476 47468
rect 233528 47456 233534 47508
rect 266590 47456 266596 47508
rect 266648 47496 266654 47508
rect 281586 47496 281592 47508
rect 266648 47468 281592 47496
rect 266648 47456 266654 47468
rect 281586 47456 281592 47468
rect 281644 47496 281650 47508
rect 328046 47496 328052 47508
rect 281644 47468 328052 47496
rect 281644 47456 281650 47468
rect 328046 47456 328052 47468
rect 328104 47456 328110 47508
rect 369262 47456 369268 47508
rect 369320 47496 369326 47508
rect 369814 47496 369820 47508
rect 369320 47468 369820 47496
rect 369320 47456 369326 47468
rect 369814 47456 369820 47468
rect 369872 47456 369878 47508
rect 13038 47388 13044 47440
rect 13096 47428 13102 47440
rect 16534 47428 16540 47440
rect 13096 47400 16540 47428
rect 13096 47388 13102 47400
rect 16534 47388 16540 47400
rect 16592 47388 16598 47440
rect 60694 47388 60700 47440
rect 60752 47428 60758 47440
rect 72562 47428 72568 47440
rect 60752 47400 72568 47428
rect 60752 47388 60758 47400
rect 72562 47388 72568 47400
rect 72620 47428 72626 47440
rect 73298 47428 73304 47440
rect 72620 47400 73304 47428
rect 72620 47388 72626 47400
rect 73298 47388 73304 47400
rect 73356 47388 73362 47440
rect 95473 47431 95531 47437
rect 95473 47397 95485 47431
rect 95519 47428 95531 47431
rect 105041 47431 105099 47437
rect 105041 47428 105053 47431
rect 95519 47400 105053 47428
rect 95519 47397 95531 47400
rect 95473 47391 95531 47397
rect 105041 47397 105053 47400
rect 105087 47397 105099 47431
rect 105041 47391 105099 47397
rect 294190 47388 294196 47440
rect 294248 47428 294254 47440
rect 295478 47428 295484 47440
rect 294248 47400 295484 47428
rect 294248 47388 294254 47400
rect 295478 47388 295484 47400
rect 295536 47428 295542 47440
rect 353622 47428 353628 47440
rect 295536 47400 353628 47428
rect 295536 47388 295542 47400
rect 353622 47388 353628 47400
rect 353680 47428 353686 47440
rect 419770 47428 419776 47440
rect 353680 47400 419776 47428
rect 353680 47388 353686 47400
rect 419770 47388 419776 47400
rect 419828 47388 419834 47440
rect 285910 47320 285916 47372
rect 285968 47360 285974 47372
rect 339638 47360 339644 47372
rect 285968 47332 339644 47360
rect 285968 47320 285974 47332
rect 339638 47320 339644 47332
rect 339696 47320 339702 47372
rect 87098 47184 87104 47236
rect 87156 47224 87162 47236
rect 93630 47224 93636 47236
rect 87156 47196 93636 47224
rect 87156 47184 87162 47196
rect 93630 47184 93636 47196
rect 93688 47224 93694 47236
rect 95105 47227 95163 47233
rect 95105 47224 95117 47227
rect 93688 47196 95117 47224
rect 93688 47184 93694 47196
rect 95105 47193 95117 47196
rect 95151 47193 95163 47227
rect 95105 47187 95163 47193
rect 86089 46819 86147 46825
rect 86089 46785 86101 46819
rect 86135 46816 86147 46819
rect 88018 46816 88024 46828
rect 86135 46788 88024 46816
rect 86135 46785 86147 46788
rect 86089 46779 86147 46785
rect 88018 46776 88024 46788
rect 88076 46816 88082 46828
rect 100898 46816 100904 46828
rect 88076 46788 100904 46816
rect 88076 46776 88082 46788
rect 100898 46776 100904 46788
rect 100956 46776 100962 46828
rect 74678 46708 74684 46760
rect 74736 46748 74742 46760
rect 87190 46748 87196 46760
rect 74736 46720 87196 46748
rect 74736 46708 74742 46720
rect 87190 46708 87196 46720
rect 87248 46708 87254 46760
rect 275882 46708 275888 46760
rect 275940 46748 275946 46760
rect 294190 46748 294196 46760
rect 275940 46720 294196 46748
rect 275940 46708 275946 46720
rect 294190 46708 294196 46720
rect 294248 46708 294254 46760
rect 71182 46164 71188 46216
rect 71240 46204 71246 46216
rect 74310 46204 74316 46216
rect 71240 46176 74316 46204
rect 71240 46164 71246 46176
rect 74310 46164 74316 46176
rect 74368 46204 74374 46216
rect 88202 46204 88208 46216
rect 74368 46176 88208 46204
rect 74368 46164 74374 46176
rect 88202 46164 88208 46176
rect 88260 46204 88266 46216
rect 106602 46204 106608 46216
rect 88260 46176 106608 46204
rect 88260 46164 88266 46176
rect 106602 46164 106608 46176
rect 106660 46164 106666 46216
rect 73298 46096 73304 46148
rect 73356 46136 73362 46148
rect 86089 46139 86147 46145
rect 86089 46136 86101 46139
rect 73356 46108 86101 46136
rect 73356 46096 73362 46108
rect 86089 46105 86101 46108
rect 86135 46105 86147 46139
rect 86089 46099 86147 46105
rect 87190 46096 87196 46148
rect 87248 46136 87254 46148
rect 88110 46136 88116 46148
rect 87248 46108 88116 46136
rect 87248 46096 87254 46108
rect 88110 46096 88116 46108
rect 88168 46136 88174 46148
rect 109454 46136 109460 46148
rect 88168 46108 109460 46136
rect 88168 46096 88174 46108
rect 109454 46096 109460 46108
rect 109512 46096 109518 46148
rect 50206 46028 50212 46080
rect 50264 46068 50270 46080
rect 369538 46068 369544 46080
rect 50264 46040 369544 46068
rect 50264 46028 50270 46040
rect 369538 46028 369544 46040
rect 369596 46028 369602 46080
rect 53702 45960 53708 46012
rect 53760 46000 53766 46012
rect 95470 46000 95476 46012
rect 53760 45972 95476 46000
rect 53760 45960 53766 45972
rect 95470 45960 95476 45972
rect 95528 45960 95534 46012
rect 144690 45960 144696 46012
rect 144748 46000 144754 46012
rect 369722 46000 369728 46012
rect 144748 45972 369728 46000
rect 144748 45960 144754 45972
rect 369722 45960 369728 45972
rect 369780 45960 369786 46012
rect 57198 45892 57204 45944
rect 57256 45932 57262 45944
rect 98046 45932 98052 45944
rect 57256 45904 98052 45932
rect 57256 45892 57262 45904
rect 98046 45892 98052 45904
rect 98104 45932 98110 45944
rect 153430 45932 153436 45944
rect 98104 45904 153436 45932
rect 98104 45892 98110 45904
rect 153430 45892 153436 45904
rect 153488 45892 153494 45944
rect 238622 45892 238628 45944
rect 238680 45932 238686 45944
rect 322618 45932 322624 45944
rect 238680 45904 322624 45932
rect 238680 45892 238686 45904
rect 322618 45892 322624 45904
rect 322676 45892 322682 45944
rect 338350 45892 338356 45944
rect 338408 45932 338414 45944
rect 343134 45932 343140 45944
rect 338408 45904 343140 45932
rect 338408 45892 338414 45904
rect 343134 45892 343140 45904
rect 343192 45892 343198 45944
rect 350126 45892 350132 45944
rect 350184 45932 350190 45944
rect 417010 45932 417016 45944
rect 350184 45904 417016 45932
rect 350184 45892 350190 45904
rect 417010 45892 417016 45904
rect 417068 45892 417074 45944
rect 95470 45824 95476 45876
rect 95528 45864 95534 45876
rect 95746 45864 95752 45876
rect 95528 45836 95752 45864
rect 95528 45824 95534 45836
rect 95746 45824 95752 45836
rect 95804 45864 95810 45876
rect 150578 45864 150584 45876
rect 95804 45836 150584 45864
rect 95804 45824 95810 45836
rect 150578 45824 150584 45836
rect 150636 45864 150642 45876
rect 170174 45864 170180 45876
rect 150636 45836 170180 45864
rect 150636 45824 150642 45836
rect 170174 45824 170180 45836
rect 170232 45824 170238 45876
rect 256930 45824 256936 45876
rect 256988 45864 256994 45876
rect 263186 45864 263192 45876
rect 256988 45836 263192 45864
rect 256988 45824 256994 45836
rect 263186 45824 263192 45836
rect 263244 45824 263250 45876
rect 283702 45824 283708 45876
rect 283760 45864 283766 45876
rect 336142 45864 336148 45876
rect 283760 45836 336148 45864
rect 283760 45824 283766 45836
rect 336142 45824 336148 45836
rect 336200 45824 336206 45876
rect 332646 45756 332652 45808
rect 332704 45796 332710 45808
rect 369814 45796 369820 45808
rect 332704 45768 369820 45796
rect 332704 45756 332710 45768
rect 369814 45756 369820 45768
rect 369872 45756 369878 45808
rect 182042 45416 182048 45468
rect 182100 45456 182106 45468
rect 201454 45456 201460 45468
rect 182100 45428 201460 45456
rect 182100 45416 182106 45428
rect 201454 45416 201460 45428
rect 201512 45416 201518 45468
rect 339638 45416 339644 45468
rect 339696 45456 339702 45468
rect 350770 45456 350776 45468
rect 339696 45428 350776 45456
rect 339696 45416 339702 45428
rect 350770 45416 350776 45428
rect 350828 45416 350834 45468
rect 168886 45348 168892 45400
rect 168944 45388 168950 45400
rect 181950 45388 181956 45400
rect 168944 45360 181956 45388
rect 168944 45348 168950 45360
rect 181950 45348 181956 45360
rect 182008 45388 182014 45400
rect 203754 45388 203760 45400
rect 182008 45360 203760 45388
rect 182008 45348 182014 45360
rect 203754 45348 203760 45360
rect 203812 45348 203818 45400
rect 275974 45348 275980 45400
rect 276032 45388 276038 45400
rect 293086 45388 293092 45400
rect 276032 45360 293092 45388
rect 276032 45348 276038 45360
rect 293086 45348 293092 45360
rect 293144 45388 293150 45400
rect 324550 45388 324556 45400
rect 293144 45360 324556 45388
rect 293144 45348 293150 45360
rect 324550 45348 324556 45360
rect 324608 45388 324614 45400
rect 350126 45388 350132 45400
rect 324608 45360 350132 45388
rect 324608 45348 324614 45360
rect 350126 45348 350132 45360
rect 350184 45348 350190 45400
rect 169714 44736 169720 44788
rect 169772 44776 169778 44788
rect 182042 44776 182048 44788
rect 169772 44748 182048 44776
rect 169772 44736 169778 44748
rect 182042 44736 182048 44748
rect 182100 44736 182106 44788
rect 263186 44736 263192 44788
rect 263244 44776 263250 44788
rect 275974 44776 275980 44788
rect 263244 44748 275980 44776
rect 263244 44736 263250 44748
rect 275974 44736 275980 44748
rect 276032 44736 276038 44788
rect 101358 37732 101364 37784
rect 101416 37772 101422 37784
rect 102278 37772 102284 37784
rect 101416 37744 102284 37772
rect 101416 37732 101422 37744
rect 102278 37732 102284 37744
rect 102336 37732 102342 37784
rect 210010 37732 210016 37784
rect 210068 37772 210074 37784
rect 211298 37772 211304 37784
rect 210068 37744 211304 37772
rect 210068 37732 210074 37744
rect 211298 37732 211304 37744
rect 211356 37732 211362 37784
rect 289038 37732 289044 37784
rect 289096 37772 289102 37784
rect 289958 37772 289964 37784
rect 289096 37744 289964 37772
rect 289096 37732 289102 37744
rect 289958 37732 289964 37744
rect 290016 37732 290022 37784
rect 304034 37732 304040 37784
rect 304092 37772 304098 37784
rect 305138 37772 305144 37784
rect 304092 37744 305144 37772
rect 304092 37732 304098 37744
rect 305138 37732 305144 37744
rect 305196 37732 305202 37784
rect 309094 37732 309100 37784
rect 309152 37772 309158 37784
rect 310014 37772 310020 37784
rect 309152 37744 310020 37772
rect 309152 37732 309158 37744
rect 310014 37732 310020 37744
rect 310072 37732 310078 37784
rect 126382 37596 126388 37648
rect 126440 37636 126446 37648
rect 128590 37636 128596 37648
rect 126440 37608 128596 37636
rect 126440 37596 126446 37608
rect 128590 37596 128596 37608
rect 128648 37596 128654 37648
rect 96390 37460 96396 37512
rect 96448 37500 96454 37512
rect 96758 37500 96764 37512
rect 96448 37472 96764 37500
rect 96448 37460 96454 37472
rect 96758 37460 96764 37472
rect 96816 37460 96822 37512
rect 195014 37392 195020 37444
rect 195072 37432 195078 37444
rect 196118 37432 196124 37444
rect 195072 37404 196124 37432
rect 195072 37392 195078 37404
rect 196118 37392 196124 37404
rect 196176 37392 196182 37444
rect 215070 37392 215076 37444
rect 215128 37432 215134 37444
rect 216174 37432 216180 37444
rect 215128 37404 216180 37432
rect 215128 37392 215134 37404
rect 216174 37392 216180 37404
rect 216232 37392 216238 37444
rect 220038 37392 220044 37444
rect 220096 37432 220102 37444
rect 222430 37432 222436 37444
rect 220096 37404 222436 37432
rect 220096 37392 220102 37404
rect 222430 37392 222436 37404
rect 222488 37392 222494 37444
rect 279102 37324 279108 37376
rect 279160 37364 279166 37376
rect 280298 37364 280304 37376
rect 279160 37336 280304 37364
rect 279160 37324 279166 37336
rect 280298 37324 280304 37336
rect 280356 37324 280362 37376
rect 121414 37256 121420 37308
rect 121472 37296 121478 37308
rect 122334 37296 122340 37308
rect 121472 37268 122340 37296
rect 121472 37256 121478 37268
rect 122334 37256 122340 37268
rect 122392 37256 122398 37308
rect 217554 37052 217560 37104
rect 217612 37092 217618 37104
rect 223534 37092 223540 37104
rect 217612 37064 223540 37092
rect 217612 37052 217618 37064
rect 223534 37052 223540 37064
rect 223592 37052 223598 37104
rect 123898 36712 123904 36764
rect 123956 36752 123962 36764
rect 128682 36752 128688 36764
rect 123956 36724 128688 36752
rect 123956 36712 123962 36724
rect 128682 36712 128688 36724
rect 128740 36712 128746 36764
rect 111386 36644 111392 36696
rect 111444 36684 111450 36696
rect 111938 36684 111944 36696
rect 111444 36656 111944 36684
rect 111444 36644 111450 36656
rect 111938 36644 111944 36656
rect 111996 36644 112002 36696
rect 311578 36508 311584 36560
rect 311636 36548 311642 36560
rect 317466 36548 317472 36560
rect 311636 36520 317472 36548
rect 311636 36508 311642 36520
rect 317466 36508 317472 36520
rect 317524 36508 317530 36560
rect 314062 36440 314068 36492
rect 314120 36480 314126 36492
rect 316270 36480 316276 36492
rect 314120 36452 316276 36480
rect 314120 36440 314126 36452
rect 316270 36440 316276 36452
rect 316328 36440 316334 36492
rect 12854 36304 12860 36356
rect 12912 36344 12918 36356
rect 16442 36344 16448 36356
rect 12912 36316 16448 36344
rect 12912 36304 12918 36316
rect 16442 36304 16448 36316
rect 16500 36304 16506 36356
rect 276158 33040 276164 33092
rect 276216 33080 276222 33092
rect 369630 33080 369636 33092
rect 276216 33052 369636 33080
rect 276216 33040 276222 33052
rect 369630 33040 369636 33052
rect 369688 33040 369694 33092
rect 182318 32972 182324 33024
rect 182376 33012 182382 33024
rect 369446 33012 369452 33024
rect 182376 32984 369452 33012
rect 182376 32972 182382 32984
rect 369446 32972 369452 32984
rect 369504 32972 369510 33024
rect 88478 32904 88484 32956
rect 88536 32944 88542 32956
rect 369170 32944 369176 32956
rect 88536 32916 369176 32944
rect 88536 32904 88542 32916
rect 369170 32904 369176 32916
rect 369228 32904 369234 32956
rect 427498 28076 427504 28128
rect 427556 28116 427562 28128
rect 429430 28116 429436 28128
rect 427556 28088 429436 28116
rect 427556 28076 427562 28088
rect 429430 28076 429436 28088
rect 429488 28076 429494 28128
rect 12670 24948 12676 25000
rect 12728 24988 12734 25000
rect 16258 24988 16264 25000
rect 12728 24960 16264 24988
rect 12728 24948 12734 24960
rect 16258 24948 16264 24960
rect 16316 24948 16322 25000
rect 185170 17060 185176 17112
rect 185228 17100 185234 17112
rect 186366 17100 186372 17112
rect 185228 17072 186372 17100
rect 185228 17060 185234 17072
rect 186366 17060 186372 17072
rect 186424 17060 186430 17112
rect 191334 17060 191340 17112
rect 191392 17100 191398 17112
rect 192070 17100 192076 17112
rect 191392 17072 192076 17100
rect 191392 17060 191398 17072
rect 192070 17060 192076 17072
rect 192128 17060 192134 17112
rect 288670 17060 288676 17112
rect 288728 17100 288734 17112
rect 290326 17100 290332 17112
rect 288728 17072 290332 17100
rect 288728 17060 288734 17072
rect 290326 17060 290332 17072
rect 290384 17060 290390 17112
rect 194554 16992 194560 17044
rect 194612 17032 194618 17044
rect 196302 17032 196308 17044
rect 194612 17004 196308 17032
rect 194612 16992 194618 17004
rect 196302 16992 196308 17004
rect 196360 16992 196366 17044
rect 92618 16788 92624 16840
rect 92676 16828 92682 16840
rect 105130 16828 105136 16840
rect 92676 16800 105136 16828
rect 92676 16788 92682 16800
rect 105130 16788 105136 16800
rect 105188 16788 105194 16840
rect 80750 16720 80756 16772
rect 80808 16760 80814 16772
rect 102370 16760 102376 16772
rect 80808 16732 102376 16760
rect 80808 16720 80814 16732
rect 102370 16720 102376 16732
rect 102428 16720 102434 16772
rect 285358 16720 285364 16772
rect 285416 16760 285422 16772
rect 299710 16760 299716 16772
rect 285416 16732 299716 16760
rect 285416 16720 285422 16732
rect 299710 16720 299716 16732
rect 299768 16720 299774 16772
rect 67870 16652 67876 16704
rect 67928 16692 67934 16704
rect 107062 16692 107068 16704
rect 67928 16664 107068 16692
rect 67928 16652 67934 16664
rect 107062 16652 107068 16664
rect 107120 16652 107126 16704
rect 170910 16652 170916 16704
rect 170968 16692 170974 16704
rect 201362 16692 201368 16704
rect 170968 16664 201368 16692
rect 170968 16652 170974 16664
rect 201362 16652 201368 16664
rect 201420 16652 201426 16704
rect 273950 16652 273956 16704
rect 274008 16692 274014 16704
rect 295386 16692 295392 16704
rect 274008 16664 295392 16692
rect 274008 16652 274014 16664
rect 295386 16652 295392 16664
rect 295444 16652 295450 16704
rect 54990 16584 54996 16636
rect 55048 16624 55054 16636
rect 112030 16624 112036 16636
rect 55048 16596 112036 16624
rect 55048 16584 55054 16596
rect 112030 16584 112036 16596
rect 112088 16584 112094 16636
rect 158030 16584 158036 16636
rect 158088 16624 158094 16636
rect 206330 16624 206336 16636
rect 158088 16596 206336 16624
rect 158088 16584 158094 16596
rect 206330 16584 206336 16596
rect 206388 16584 206394 16636
rect 261070 16584 261076 16636
rect 261128 16624 261134 16636
rect 300354 16624 300360 16636
rect 261128 16596 300360 16624
rect 261128 16584 261134 16596
rect 300354 16584 300360 16596
rect 300412 16584 300418 16636
rect 29230 16516 29236 16568
rect 29288 16556 29294 16568
rect 122058 16556 122064 16568
rect 29288 16528 122064 16556
rect 29288 16516 29294 16528
rect 122058 16516 122064 16528
rect 122116 16516 122122 16568
rect 145150 16516 145156 16568
rect 145208 16556 145214 16568
rect 211298 16556 211304 16568
rect 145208 16528 211304 16556
rect 145208 16516 145214 16528
rect 211298 16516 211304 16528
rect 211356 16516 211362 16568
rect 248190 16516 248196 16568
rect 248248 16556 248254 16568
rect 305322 16556 305328 16568
rect 248248 16528 305328 16556
rect 248248 16516 248254 16528
rect 305322 16516 305328 16528
rect 305380 16516 305386 16568
rect 42110 16448 42116 16500
rect 42168 16488 42174 16500
rect 116998 16488 117004 16500
rect 42168 16460 117004 16488
rect 42168 16448 42174 16460
rect 116998 16448 117004 16460
rect 117056 16448 117062 16500
rect 119390 16448 119396 16500
rect 119448 16488 119454 16500
rect 221326 16488 221332 16500
rect 119448 16460 221332 16488
rect 119448 16448 119454 16460
rect 221326 16448 221332 16460
rect 221384 16448 221390 16500
rect 235310 16448 235316 16500
rect 235368 16488 235374 16500
rect 310382 16488 310388 16500
rect 235368 16460 310388 16488
rect 235368 16448 235374 16460
rect 310382 16448 310388 16460
rect 310440 16448 310446 16500
rect 16350 16380 16356 16432
rect 16408 16420 16414 16432
rect 127210 16420 127216 16432
rect 16408 16392 127216 16420
rect 16408 16380 16414 16392
rect 127210 16380 127216 16392
rect 127268 16380 127274 16432
rect 132270 16380 132276 16432
rect 132328 16420 132334 16432
rect 216358 16420 216364 16432
rect 132328 16392 216364 16420
rect 132328 16380 132334 16392
rect 216358 16380 216364 16392
rect 216416 16380 216422 16432
rect 222430 16380 222436 16432
rect 222488 16420 222494 16432
rect 315350 16420 315356 16432
rect 222488 16392 315356 16420
rect 222488 16380 222494 16392
rect 315350 16380 315356 16392
rect 315408 16380 315414 16432
rect 95470 16040 95476 16092
rect 95528 16080 95534 16092
rect 97034 16080 97040 16092
rect 95528 16052 97040 16080
rect 95528 16040 95534 16052
rect 97034 16040 97040 16052
rect 97092 16040 97098 16092
rect 427314 15292 427320 15344
rect 427372 15332 427378 15344
rect 429430 15332 429436 15344
rect 427372 15304 429436 15332
rect 427372 15292 427378 15304
rect 429430 15292 429436 15304
rect 429488 15292 429494 15344
rect 12670 14204 12676 14256
rect 12728 14244 12734 14256
rect 16074 14244 16080 14256
rect 12728 14216 16080 14244
rect 12728 14204 12734 14216
rect 16074 14204 16080 14216
rect 16132 14204 16138 14256
rect 93630 12572 93636 12624
rect 93688 12612 93694 12624
rect 95470 12612 95476 12624
rect 93688 12584 95476 12612
rect 93688 12572 93694 12584
rect 95470 12572 95476 12584
rect 95528 12572 95534 12624
rect 286830 12368 286836 12420
rect 286888 12408 286894 12420
rect 288670 12408 288676 12420
rect 286888 12380 288676 12408
rect 286888 12368 286894 12380
rect 288670 12368 288676 12380
rect 288728 12368 288734 12420
rect 325286 12368 325292 12420
rect 325344 12408 325350 12420
rect 364110 12408 364116 12420
rect 325344 12380 364116 12408
rect 325344 12368 325350 12380
rect 364110 12368 364116 12380
rect 364168 12368 364174 12420
rect 376990 12368 376996 12420
rect 377048 12408 377054 12420
rect 378278 12408 378284 12420
rect 377048 12380 378284 12408
rect 377048 12368 377054 12380
rect 378278 12368 378284 12380
rect 378336 12368 378342 12420
rect 105130 12300 105136 12352
rect 105188 12340 105194 12352
rect 106510 12340 106516 12352
rect 105188 12312 106516 12340
rect 105188 12300 105194 12312
rect 106510 12300 106516 12312
rect 106568 12300 106574 12352
rect 183790 12300 183796 12352
rect 183848 12340 183854 12352
rect 194554 12340 194560 12352
rect 183848 12312 194560 12340
rect 183848 12300 183854 12312
rect 194554 12300 194560 12312
rect 194612 12300 194618 12352
rect 362454 12300 362460 12352
rect 362512 12340 362518 12352
rect 402750 12340 402756 12352
rect 362512 12312 402756 12340
rect 362512 12300 362518 12312
rect 402750 12300 402756 12312
rect 402808 12300 402814 12352
rect 185170 12232 185176 12284
rect 185228 12272 185234 12284
rect 209550 12272 209556 12284
rect 185228 12244 209556 12272
rect 185228 12232 185234 12244
rect 209550 12232 209556 12244
rect 209608 12232 209614 12284
rect 280390 12232 280396 12284
rect 280448 12272 280454 12284
rect 312590 12272 312596 12284
rect 280448 12244 312596 12272
rect 280448 12232 280454 12244
rect 312590 12232 312596 12244
rect 312648 12232 312654 12284
rect 322526 12232 322532 12284
rect 322584 12272 322590 12284
rect 415630 12272 415636 12284
rect 322584 12244 415636 12272
rect 322584 12232 322590 12244
rect 415630 12232 415636 12244
rect 415688 12232 415694 12284
rect 192070 12096 192076 12148
rect 192128 12136 192134 12148
rect 196670 12136 196676 12148
rect 192128 12108 196676 12136
rect 192128 12096 192134 12108
rect 196670 12096 196676 12108
rect 196728 12096 196734 12148
rect 350770 9376 350776 9428
rect 350828 9416 350834 9428
rect 351230 9416 351236 9428
rect 350828 9388 351236 9416
rect 350828 9376 350834 9388
rect 351230 9376 351236 9388
rect 351288 9376 351294 9428
rect 389410 9376 389416 9428
rect 389468 9416 389474 9428
rect 389870 9416 389876 9428
rect 389468 9388 389876 9416
rect 389468 9376 389474 9388
rect 389870 9376 389876 9388
rect 389928 9376 389934 9428
rect 428050 9376 428056 9428
rect 428108 9416 428114 9428
rect 428510 9416 428516 9428
rect 428108 9388 428516 9416
rect 428108 9376 428114 9388
rect 428510 9376 428516 9388
rect 428568 9376 428574 9428
<< via1 >>
rect 395120 395183 395172 395192
rect 395120 395149 395129 395183
rect 395129 395149 395163 395183
rect 395163 395149 395172 395183
rect 395120 395140 395172 395149
rect 22336 393780 22388 393832
rect 23164 393780 23216 393832
rect 48556 393780 48608 393832
rect 49660 393780 49712 393832
rect 128596 393780 128648 393832
rect 129424 393780 129476 393832
rect 154816 393780 154868 393832
rect 155920 393780 155972 393832
rect 234856 393780 234908 393832
rect 235684 393780 235736 393832
rect 261076 393780 261128 393832
rect 262180 393780 262232 393832
rect 279660 393168 279712 393220
rect 315356 393168 315408 393220
rect 102836 393100 102888 393152
rect 108908 393100 108960 393152
rect 314620 393100 314672 393152
rect 421616 393100 421668 393152
rect 284444 392488 284496 392540
rect 288768 392488 288820 392540
rect 13136 391060 13188 391112
rect 87196 391060 87248 391112
rect 299624 389700 299676 389752
rect 429436 389700 429488 389752
rect 108908 389428 108960 389480
rect 111300 389428 111352 389480
rect 195296 389156 195348 389208
rect 208636 389156 208688 389208
rect 76156 389088 76208 389140
rect 116268 389088 116320 389140
rect 182416 389088 182468 389140
rect 200356 389088 200408 389140
rect 48556 389020 48608 389072
rect 121328 389020 121380 389072
rect 154816 389020 154868 389072
rect 205324 389020 205376 389072
rect 261076 389020 261128 389072
rect 288952 389020 289004 389072
rect 22336 388952 22388 389004
rect 126296 388952 126348 389004
rect 128596 388952 128648 389004
rect 210292 388952 210344 389004
rect 234856 388952 234908 389004
rect 294196 388952 294248 389004
rect 91336 388680 91388 388732
rect 358504 388680 358556 388732
rect 13504 388612 13556 388664
rect 96304 388612 96356 388664
rect 13320 388544 13372 388596
rect 106332 388544 106384 388596
rect 13688 388476 13740 388528
rect 185360 388476 185412 388528
rect 190328 388476 190380 388528
rect 223080 388476 223132 388528
rect 304592 388476 304644 388528
rect 322532 388476 322584 388528
rect 13596 388408 13648 388460
rect 215352 388408 215404 388460
rect 220320 388408 220372 388460
rect 362460 388408 362512 388460
rect 13412 388340 13464 388392
rect 101272 388340 101324 388392
rect 309284 388340 309336 388392
rect 315632 388340 315684 388392
rect 395212 385552 395264 385604
rect 315816 378616 315868 378668
rect 429436 378616 429488 378668
rect 131816 371748 131868 371800
rect 134760 371748 134812 371800
rect 225840 371748 225892 371800
rect 265860 371748 265912 371800
rect 320140 371748 320192 371800
rect 323820 371748 323872 371800
rect 189040 368552 189092 368604
rect 190696 368552 190748 368604
rect 209004 368552 209056 368604
rect 210016 368552 210068 368604
rect 219032 368552 219084 368604
rect 220320 368552 220372 368604
rect 277544 368280 277596 368332
rect 280396 368280 280448 368332
rect 89864 367668 89916 367720
rect 92532 367668 92584 367720
rect 90048 367600 90100 367652
rect 91336 367600 91388 367652
rect 99984 367600 100036 367652
rect 100904 367600 100956 367652
rect 110012 367600 110064 367652
rect 112036 367600 112088 367652
rect 114980 367600 115032 367652
rect 116176 367600 116228 367652
rect 125008 367600 125060 367652
rect 126480 367600 126532 367652
rect 184072 367600 184124 367652
rect 185084 367600 185136 367652
rect 185268 367600 185320 367652
rect 186556 367600 186608 367652
rect 199068 367600 199120 367652
rect 200264 367600 200316 367652
rect 204036 367600 204088 367652
rect 205876 367600 205928 367652
rect 278372 367600 278424 367652
rect 280488 367600 280540 367652
rect 293368 367600 293420 367652
rect 294288 367600 294340 367652
rect 298244 367600 298296 367652
rect 299716 367600 299768 367652
rect 303304 367600 303356 367652
rect 305236 367600 305288 367652
rect 308364 367600 308416 367652
rect 309284 367600 309336 367652
rect 223080 367532 223132 367584
rect 429436 367532 429488 367584
rect 395304 366351 395356 366360
rect 395304 366317 395313 366351
rect 395313 366317 395347 366351
rect 395347 366317 395356 366351
rect 395304 366308 395356 366317
rect 395212 364948 395264 365000
rect 91336 363452 91388 363504
rect 92072 363452 92124 363504
rect 116176 363452 116228 363504
rect 116820 363452 116872 363504
rect 210016 363452 210068 363504
rect 210844 363452 210896 363504
rect 395304 363495 395356 363504
rect 395304 363461 395313 363495
rect 395313 363461 395347 363495
rect 395347 363461 395356 363495
rect 395304 363452 395356 363461
rect 53708 359780 53760 359832
rect 76984 359780 77036 359832
rect 50212 359712 50264 359764
rect 76800 359712 76852 359764
rect 64196 359644 64248 359696
rect 76064 359644 76116 359696
rect 60700 359576 60752 359628
rect 75880 359576 75932 359628
rect 57204 359508 57256 359560
rect 75788 359508 75840 359560
rect 67692 359372 67744 359424
rect 75972 359372 76024 359424
rect 80204 357876 80256 357928
rect 127216 357876 127268 357928
rect 139636 357876 139688 357928
rect 174044 357876 174096 357928
rect 221056 357876 221108 357928
rect 233476 357876 233528 357928
rect 266596 357876 266648 357928
rect 314896 357876 314948 357928
rect 328420 357876 328472 357928
rect 75880 357604 75932 357656
rect 76156 357604 76208 357656
rect 75788 357536 75840 357588
rect 71464 357468 71516 357520
rect 75880 357468 75932 357520
rect 74776 357400 74828 357452
rect 76892 357400 76944 357452
rect 80204 356516 80256 356568
rect 121696 356516 121748 356568
rect 139636 356516 139688 356568
rect 173492 356516 173544 356568
rect 215536 356516 215588 356568
rect 233476 356516 233528 356568
rect 266596 356516 266648 356568
rect 309376 356516 309428 356568
rect 328328 356516 328380 356568
rect 80204 355156 80256 355208
rect 117556 355156 117608 355208
rect 118016 355156 118068 355208
rect 120224 355156 120276 355208
rect 122064 355156 122116 355208
rect 139636 355156 139688 355208
rect 174044 355156 174096 355208
rect 211396 355156 211448 355208
rect 212684 355156 212736 355208
rect 214064 355156 214116 355208
rect 216364 355156 216416 355208
rect 233476 355156 233528 355208
rect 266596 355156 266648 355208
rect 305328 355156 305380 355208
rect 328420 355156 328472 355208
rect 79284 355088 79336 355140
rect 105044 355088 105096 355140
rect 107068 355088 107120 355140
rect 95384 355020 95436 355072
rect 97040 355020 97092 355072
rect 100904 355020 100956 355072
rect 102376 355020 102428 355072
rect 112128 354884 112180 354936
rect 139728 355088 139780 355140
rect 173768 355088 173820 355140
rect 205968 355088 206020 355140
rect 233568 355088 233620 355140
rect 266688 355088 266740 355140
rect 299808 355088 299860 355140
rect 328512 355088 328564 355140
rect 126480 355020 126532 355072
rect 127216 355020 127268 355072
rect 185084 355020 185136 355072
rect 186372 355020 186424 355072
rect 194744 355020 194796 355072
rect 196308 355020 196360 355072
rect 220320 355020 220372 355072
rect 221332 355020 221384 355072
rect 283064 355020 283116 355072
rect 285364 355020 285416 355072
rect 288584 355020 288636 355072
rect 290332 355020 290384 355072
rect 309284 355020 309336 355072
rect 310388 355020 310440 355072
rect 313424 355020 313476 355072
rect 315356 355020 315408 355072
rect 118016 354952 118068 355004
rect 212684 354952 212736 355004
rect 200264 354000 200316 354052
rect 201368 354000 201420 354052
rect 76248 353907 76300 353916
rect 76248 353873 76257 353907
rect 76257 353873 76291 353907
rect 76291 353873 76300 353907
rect 76248 353864 76300 353873
rect 196216 353864 196268 353916
rect 196492 353864 196544 353916
rect 390704 353864 390756 353916
rect 429436 353864 429488 353916
rect 80204 353796 80256 353848
rect 106516 353796 106568 353848
rect 139636 353796 139688 353848
rect 174044 353796 174096 353848
rect 200356 353796 200408 353848
rect 233476 353796 233528 353848
rect 266596 353796 266648 353848
rect 294196 353796 294248 353848
rect 328052 353796 328104 353848
rect 80204 352368 80256 352420
rect 102652 352368 102704 352420
rect 139636 352368 139688 352420
rect 174044 352368 174096 352420
rect 196216 352368 196268 352420
rect 233476 352368 233528 352420
rect 266596 352368 266648 352420
rect 290056 352368 290108 352420
rect 328512 352368 328564 352420
rect 191248 351867 191300 351876
rect 191248 351833 191257 351867
rect 191257 351833 191291 351867
rect 191291 351833 191300 351867
rect 191248 351824 191300 351833
rect 284536 351595 284588 351604
rect 284536 351561 284545 351595
rect 284545 351561 284579 351595
rect 284579 351561 284588 351595
rect 284536 351552 284588 351561
rect 96764 351527 96816 351536
rect 96764 351493 96773 351527
rect 96773 351493 96807 351527
rect 96807 351493 96816 351527
rect 96764 351484 96816 351493
rect 226300 351280 226352 351332
rect 231636 351280 231688 351332
rect 131816 351076 131868 351128
rect 139452 351076 139504 351128
rect 272024 351076 272076 351128
rect 274876 351076 274928 351128
rect 320600 351076 320652 351128
rect 328144 351076 328196 351128
rect 79836 351008 79888 351060
rect 89864 351008 89916 351060
rect 139636 351008 139688 351060
rect 173860 351008 173912 351060
rect 185268 351008 185320 351060
rect 233568 351008 233620 351060
rect 266688 351008 266740 351060
rect 277544 351008 277596 351060
rect 327868 351008 327920 351060
rect 80204 350328 80256 350380
rect 139728 350328 139780 350380
rect 173676 350328 173728 350380
rect 233476 350328 233528 350380
rect 266596 350328 266648 350380
rect 327500 350328 327552 350380
rect 131816 349716 131868 349768
rect 139544 349716 139596 349768
rect 271932 349716 271984 349768
rect 274876 349716 274928 349768
rect 321612 349716 321664 349768
rect 328328 349716 328380 349768
rect 76064 349648 76116 349700
rect 172848 349648 172900 349700
rect 182324 349648 182376 349700
rect 231636 349648 231688 349700
rect 233476 349648 233528 349700
rect 266596 349648 266648 349700
rect 272024 349648 272076 349700
rect 78916 348900 78968 348952
rect 87104 348900 87156 348952
rect 321704 348424 321756 348476
rect 327224 348424 327276 348476
rect 131816 348356 131868 348408
rect 137244 348356 137296 348408
rect 226484 348356 226536 348408
rect 232004 348356 232056 348408
rect 131908 348288 131960 348340
rect 137520 348288 137572 348340
rect 226392 348288 226444 348340
rect 231636 348288 231688 348340
rect 321612 348288 321664 348340
rect 327132 348288 327184 348340
rect 226576 348220 226628 348272
rect 233476 348220 233528 348272
rect 266596 348220 266648 348272
rect 271932 348220 271984 348272
rect 174044 347948 174096 348000
rect 180760 347948 180812 348000
rect 78916 347336 78968 347388
rect 87012 347336 87064 347388
rect 132184 346928 132236 346980
rect 139728 346928 139780 346980
rect 226392 346928 226444 346980
rect 228600 346928 228652 346980
rect 321060 346928 321112 346980
rect 323176 346928 323228 346980
rect 137520 346860 137572 346912
rect 139636 346860 139688 346912
rect 174044 346860 174096 346912
rect 180944 346860 180996 346912
rect 232004 346860 232056 346912
rect 233476 346860 233528 346912
rect 266596 346860 266648 346912
rect 274876 346860 274928 346912
rect 137244 346792 137296 346844
rect 139820 346792 139872 346844
rect 231636 346792 231688 346844
rect 233568 346792 233620 346844
rect 266688 346792 266740 346844
rect 274968 346792 275020 346844
rect 173124 346248 173176 346300
rect 180852 346248 180904 346300
rect 78916 346180 78968 346232
rect 87104 346180 87156 346232
rect 79008 345976 79060 346028
rect 86920 345976 86972 346028
rect 131816 345636 131868 345688
rect 134116 345636 134168 345688
rect 226484 345636 226536 345688
rect 228048 345636 228100 345688
rect 320416 345636 320468 345688
rect 323268 345636 323320 345688
rect 85816 345568 85868 345620
rect 87932 345568 87984 345620
rect 131908 345568 131960 345620
rect 139636 345568 139688 345620
rect 173032 345568 173084 345620
rect 182324 345568 182376 345620
rect 226392 345568 226444 345620
rect 234580 345568 234632 345620
rect 320508 345568 320560 345620
rect 327040 345568 327092 345620
rect 395396 345568 395448 345620
rect 228600 345500 228652 345552
rect 233476 345500 233528 345552
rect 266596 345500 266648 345552
rect 275060 345500 275112 345552
rect 323176 345500 323228 345552
rect 328052 345500 328104 345552
rect 173308 345160 173360 345212
rect 180760 345160 180812 345212
rect 85908 344616 85960 344668
rect 87472 344616 87524 344668
rect 226024 344616 226076 344668
rect 228508 344616 228560 344668
rect 321060 344616 321112 344668
rect 323176 344616 323228 344668
rect 78916 344412 78968 344464
rect 87012 344412 87064 344464
rect 321612 344344 321664 344396
rect 326856 344344 326908 344396
rect 131816 344208 131868 344260
rect 138164 344208 138216 344260
rect 226392 344208 226444 344260
rect 227956 344208 228008 344260
rect 132368 344140 132420 344192
rect 139728 344140 139780 344192
rect 172940 344140 172992 344192
rect 182324 344140 182376 344192
rect 228048 344072 228100 344124
rect 233476 344072 233528 344124
rect 266596 344072 266648 344124
rect 274968 344072 275020 344124
rect 323268 344072 323320 344124
rect 328512 344072 328564 344124
rect 173676 343732 173728 343784
rect 180852 343732 180904 343784
rect 78916 342916 78968 342968
rect 85816 342916 85868 342968
rect 321612 342848 321664 342900
rect 327132 342848 327184 342900
rect 131816 342780 131868 342832
rect 139820 342780 139872 342832
rect 173676 342780 173728 342832
rect 181404 342780 181456 342832
rect 226392 342780 226444 342832
rect 233660 342780 233712 342832
rect 78916 342712 78968 342764
rect 88116 342712 88168 342764
rect 134116 342712 134168 342764
rect 139636 342712 139688 342764
rect 228508 342712 228560 342764
rect 233476 342712 233528 342764
rect 266688 342712 266740 342764
rect 274876 342712 274928 342764
rect 323176 342712 323228 342764
rect 328052 342712 328104 342764
rect 266596 342644 266648 342696
rect 275244 342644 275296 342696
rect 172756 342236 172808 342288
rect 180944 342236 180996 342288
rect 78916 341488 78968 341540
rect 85908 341488 85960 341540
rect 131908 341488 131960 341540
rect 139728 341488 139780 341540
rect 226484 341488 226536 341540
rect 233568 341488 233620 341540
rect 321612 341488 321664 341540
rect 327040 341488 327092 341540
rect 131816 341420 131868 341472
rect 139912 341420 139964 341472
rect 226392 341420 226444 341472
rect 233752 341420 233804 341472
rect 321060 341420 321112 341472
rect 327224 341420 327276 341472
rect 394844 341420 394896 341472
rect 429436 341420 429488 341472
rect 78916 341352 78968 341404
rect 88484 341352 88536 341404
rect 138164 341352 138216 341404
rect 139636 341352 139688 341404
rect 227956 341352 228008 341404
rect 233476 341352 233528 341404
rect 266596 341352 266648 341404
rect 275060 341352 275112 341404
rect 76064 340060 76116 340112
rect 76248 340060 76300 340112
rect 85724 340060 85776 340112
rect 87564 340060 87616 340112
rect 131816 340060 131868 340112
rect 137336 340060 137388 340112
rect 173492 340060 173544 340112
rect 181404 340060 181456 340112
rect 226392 340060 226444 340112
rect 231912 340060 231964 340112
rect 272024 340060 272076 340112
rect 275060 340060 275112 340112
rect 320600 340060 320652 340112
rect 326948 340060 327000 340112
rect 78916 339992 78968 340044
rect 87380 339992 87432 340044
rect 266596 339992 266648 340044
rect 274968 339992 275020 340044
rect 226484 338768 226536 338820
rect 233660 338768 233712 338820
rect 321612 338768 321664 338820
rect 326672 338768 326724 338820
rect 131816 338700 131868 338752
rect 136140 338700 136192 338752
rect 173308 338700 173360 338752
rect 181588 338700 181640 338752
rect 84988 338632 85040 338684
rect 87380 338632 87432 338684
rect 131908 338632 131960 338684
rect 139636 338632 139688 338684
rect 173400 338632 173452 338684
rect 182324 338632 182376 338684
rect 225932 338632 225984 338684
rect 230808 338632 230860 338684
rect 321244 338632 321296 338684
rect 327132 338632 327184 338684
rect 80204 338564 80256 338616
rect 87472 338564 87524 338616
rect 173952 338564 174004 338616
rect 181772 338564 181824 338616
rect 266688 338564 266740 338616
rect 274876 338564 274928 338616
rect 78916 338496 78968 338548
rect 87288 338496 87340 338548
rect 174044 338496 174096 338548
rect 182140 338496 182192 338548
rect 266596 338496 266648 338548
rect 275152 338496 275204 338548
rect 131816 337272 131868 337324
rect 136232 337272 136284 337324
rect 225932 337272 225984 337324
rect 230716 337272 230768 337324
rect 271472 337272 271524 337324
rect 274876 337272 274928 337324
rect 321612 337272 321664 337324
rect 327040 337272 327092 337324
rect 137336 337204 137388 337256
rect 139728 337204 139780 337256
rect 231912 337204 231964 337256
rect 233476 337204 233528 337256
rect 266596 337204 266648 337256
rect 272024 337204 272076 337256
rect 80204 336048 80256 336100
rect 85724 336048 85776 336100
rect 321428 336048 321480 336100
rect 327316 336048 327368 336100
rect 131908 335980 131960 336032
rect 138072 335980 138124 336032
rect 85816 335912 85868 335964
rect 87840 335912 87892 335964
rect 131816 335912 131868 335964
rect 138164 335912 138216 335964
rect 172848 335912 172900 335964
rect 181588 335912 181640 335964
rect 225932 335912 225984 335964
rect 230900 335912 230952 335964
rect 321612 335912 321664 335964
rect 327224 335912 327276 335964
rect 395212 335912 395264 335964
rect 395304 335912 395356 335964
rect 230808 335844 230860 335896
rect 233476 335844 233528 335896
rect 266596 335844 266648 335896
rect 275060 335844 275112 335896
rect 80204 335096 80256 335148
rect 84988 335096 85040 335148
rect 75972 334756 76024 334808
rect 75880 334688 75932 334740
rect 76064 334688 76116 334740
rect 75972 334527 76024 334536
rect 75972 334493 75981 334527
rect 75981 334493 76015 334527
rect 76015 334493 76024 334527
rect 75972 334484 76024 334493
rect 76064 334484 76116 334536
rect 108264 334416 108316 334468
rect 131632 334416 131684 334468
rect 136140 334416 136192 334468
rect 139636 334416 139688 334468
rect 212316 334416 212368 334468
rect 230716 334416 230768 334468
rect 233476 334416 233528 334468
rect 266596 334416 266648 334468
rect 275612 334416 275664 334468
rect 75880 334348 75932 334400
rect 104860 334348 104912 334400
rect 131724 334348 131776 334400
rect 266688 334348 266740 334400
rect 271472 334348 271524 334400
rect 75972 334280 76024 334332
rect 76984 334280 77036 334332
rect 98236 334280 98288 334332
rect 111392 334280 111444 334332
rect 131540 334280 131592 334332
rect 80204 334212 80256 334264
rect 87840 334212 87892 334264
rect 114796 334212 114848 334264
rect 131448 334212 131500 334264
rect 136232 334212 136284 334264
rect 139636 334212 139688 334264
rect 225288 334212 225340 334264
rect 231360 334212 231412 334264
rect 78916 334144 78968 334196
rect 88024 334144 88076 334196
rect 118200 334144 118252 334196
rect 131356 334144 131408 334196
rect 131632 334144 131684 334196
rect 136968 334144 137020 334196
rect 116084 334008 116136 334060
rect 127860 334008 127912 334060
rect 131540 334076 131592 334128
rect 137060 334076 137112 334128
rect 137244 334008 137296 334060
rect 103664 333940 103716 333992
rect 124548 333940 124600 333992
rect 131448 333940 131500 333992
rect 137152 333940 137204 333992
rect 211304 333940 211356 333992
rect 221884 333940 221936 333992
rect 305144 333940 305196 333992
rect 316184 333940 316236 333992
rect 91244 333872 91296 333924
rect 121236 333872 121288 333924
rect 131724 333872 131776 333924
rect 137520 333872 137572 333924
rect 197504 333872 197556 333924
rect 218572 333872 218624 333924
rect 292724 333872 292776 333924
rect 312872 333872 312924 333924
rect 98236 333804 98288 333856
rect 137980 333804 138032 333856
rect 185084 333804 185136 333856
rect 215628 333804 215680 333856
rect 280304 333804 280356 333856
rect 309560 333804 309612 333856
rect 91888 333736 91940 333788
rect 134852 333736 134904 333788
rect 185912 333736 185964 333788
rect 228600 333736 228652 333788
rect 279568 333736 279620 333788
rect 322624 333736 322676 333788
rect 173308 333464 173360 333516
rect 180392 333464 180444 333516
rect 80204 333056 80256 333108
rect 87380 333056 87432 333108
rect 138072 333056 138124 333108
rect 139636 333056 139688 333108
rect 230900 333056 230952 333108
rect 233476 333056 233528 333108
rect 266596 333056 266648 333108
rect 274876 333056 274928 333108
rect 319312 331764 319364 331816
rect 325384 331764 325436 331816
rect 76892 331696 76944 331748
rect 118200 331696 118252 331748
rect 138164 331696 138216 331748
rect 139636 331696 139688 331748
rect 173676 331696 173728 331748
rect 180944 331696 180996 331748
rect 198700 331696 198752 331748
rect 114796 331628 114848 331680
rect 111392 331560 111444 331612
rect 226576 331696 226628 331748
rect 233476 331696 233528 331748
rect 266596 331696 266648 331748
rect 274968 331696 275020 331748
rect 299532 331696 299584 331748
rect 319220 331696 319272 331748
rect 225564 331560 225616 331612
rect 230808 331560 230860 331612
rect 80204 330608 80256 330660
rect 85816 330608 85868 330660
rect 319404 330472 319456 330524
rect 325568 330472 325620 330524
rect 319220 330404 319272 330456
rect 324648 330404 324700 330456
rect 305236 330336 305288 330388
rect 306248 330336 306300 330388
rect 319036 330336 319088 330388
rect 325752 330336 325804 330388
rect 75512 330175 75564 330184
rect 75512 330141 75521 330175
rect 75521 330141 75555 330175
rect 75555 330141 75564 330175
rect 75512 330132 75564 330141
rect 75420 330107 75472 330116
rect 75420 330073 75429 330107
rect 75429 330073 75463 330107
rect 75463 330073 75472 330107
rect 75420 330064 75472 330073
rect 158220 329180 158272 329232
rect 137520 329044 137572 329096
rect 158220 329044 158272 329096
rect 198884 329112 198936 329164
rect 172112 329044 172164 329096
rect 222528 329044 222580 329096
rect 233476 329044 233528 329096
rect 266596 329044 266648 329096
rect 316552 329044 316604 329096
rect 328420 329044 328472 329096
rect 78916 328976 78968 329028
rect 128504 328976 128556 329028
rect 140372 328976 140424 329028
rect 231360 328976 231412 329028
rect 255556 328976 255608 329028
rect 305236 328976 305288 329028
rect 325200 328976 325252 329028
rect 429436 328976 429488 329028
rect 208728 328908 208780 328960
rect 225196 328908 225248 328960
rect 231084 328908 231136 328960
rect 302476 328908 302528 328960
rect 303120 328908 303172 328960
rect 319128 328908 319180 328960
rect 325660 328908 325712 328960
rect 342496 327616 342548 327668
rect 346452 327616 346504 327668
rect 395120 327616 395172 327668
rect 395212 327616 395264 327668
rect 76064 327548 76116 327600
rect 100996 327548 101048 327600
rect 156288 327548 156340 327600
rect 156840 327548 156892 327600
rect 194836 327548 194888 327600
rect 241480 327548 241532 327600
rect 252888 327548 252940 327600
rect 254820 327548 254872 327600
rect 302476 327548 302528 327600
rect 339920 327548 339972 327600
rect 356020 327548 356072 327600
rect 65484 327480 65536 327532
rect 69440 327480 69492 327532
rect 137704 327480 137756 327532
rect 137980 327480 138032 327532
rect 155920 327480 155972 327532
rect 238628 327480 238680 327532
rect 249944 327480 249996 327532
rect 250036 327480 250088 327532
rect 250772 327480 250824 327532
rect 288676 327480 288728 327532
rect 289964 327480 290016 327532
rect 337160 327480 337212 327532
rect 352800 327480 352852 327532
rect 66864 327412 66916 327464
rect 70636 327412 70688 327464
rect 154816 327412 154868 327464
rect 59228 327344 59280 327396
rect 63644 327344 63696 327396
rect 66312 327344 66364 327396
rect 67508 327344 67560 327396
rect 69072 327344 69124 327396
rect 72660 327344 72712 327396
rect 151964 327344 152016 327396
rect 165212 327344 165264 327396
rect 192076 327412 192128 327464
rect 232004 327412 232056 327464
rect 248656 327412 248708 327464
rect 248748 327412 248800 327464
rect 249852 327412 249904 327464
rect 285916 327412 285968 327464
rect 338632 327412 338684 327464
rect 353628 327412 353680 327464
rect 238996 327344 239048 327396
rect 239916 327344 239968 327396
rect 244424 327344 244476 327396
rect 246908 327344 246960 327396
rect 281776 327344 281828 327396
rect 282236 327344 282288 327396
rect 332928 327344 332980 327396
rect 333664 327344 333716 327396
rect 334216 327344 334268 327396
rect 335228 327344 335280 327396
rect 341484 327344 341536 327396
rect 357584 327344 357636 327396
rect 60240 327276 60292 327328
rect 65024 327276 65076 327328
rect 66496 327276 66548 327328
rect 68520 327276 68572 327328
rect 151320 327276 151372 327328
rect 163188 327276 163240 327328
rect 245344 327276 245396 327328
rect 247920 327276 247972 327328
rect 68428 327208 68480 327260
rect 71648 327208 71700 327260
rect 149388 327208 149440 327260
rect 163280 327208 163332 327260
rect 247368 327208 247420 327260
rect 261168 327276 261220 327328
rect 339552 327276 339604 327328
rect 351972 327276 352024 327328
rect 258408 327208 258460 327260
rect 344796 327208 344848 327260
rect 358320 327208 358372 327260
rect 62356 327140 62408 327192
rect 66588 327140 66640 327192
rect 154172 327140 154224 327192
rect 168064 327140 168116 327192
rect 247184 327140 247236 327192
rect 258960 327140 259012 327192
rect 342404 327140 342456 327192
rect 355560 327140 355612 327192
rect 150768 327072 150820 327124
rect 164568 327072 164620 327124
rect 194836 327072 194888 327124
rect 232096 327072 232148 327124
rect 250036 327072 250088 327124
rect 250128 327072 250180 327124
rect 264020 327072 264072 327124
rect 289964 327072 290016 327124
rect 325292 327072 325344 327124
rect 341208 327072 341260 327124
rect 358412 327072 358464 327124
rect 64380 327004 64432 327056
rect 69164 327004 69216 327056
rect 153252 327004 153304 327056
rect 165120 327004 165172 327056
rect 233476 327004 233528 327056
rect 248656 327004 248708 327056
rect 248748 327004 248800 327056
rect 263100 327004 263152 327056
rect 285916 327004 285968 327056
rect 324556 327004 324608 327056
rect 339920 327004 339972 327056
rect 356756 327004 356808 327056
rect 137612 326936 137664 326988
rect 154816 326936 154868 326988
rect 154908 326936 154960 326988
rect 187936 326936 187988 326988
rect 230716 326936 230768 326988
rect 232004 326936 232056 326988
rect 244608 326936 244660 326988
rect 248288 326936 248340 326988
rect 268620 326936 268672 326988
rect 282236 326936 282288 326988
rect 325476 326936 325528 326988
rect 338540 326936 338592 326988
rect 355192 326936 355244 326988
rect 100996 326868 101048 326920
rect 136876 326868 136928 326920
rect 154264 326868 154316 326920
rect 326580 326868 326632 326920
rect 335688 326868 335740 326920
rect 336792 326868 336844 326920
rect 354364 326868 354416 326920
rect 363840 326868 363892 326920
rect 153528 326800 153580 326852
rect 167328 326800 167380 326852
rect 243136 326800 243188 326852
rect 57204 326732 57256 326784
rect 62264 326732 62316 326784
rect 152056 326732 152108 326784
rect 166132 326732 166184 326784
rect 239548 326732 239600 326784
rect 74316 326664 74368 326716
rect 76892 326664 76944 326716
rect 144604 326664 144656 326716
rect 155552 326664 155604 326716
rect 156196 326664 156248 326716
rect 169996 326664 170048 326716
rect 241940 326664 241992 326716
rect 242768 326664 242820 326716
rect 245896 326732 245948 326784
rect 250036 326664 250088 326716
rect 255464 326800 255516 326852
rect 256292 326800 256344 326852
rect 256936 326800 256988 326852
rect 262088 326800 262140 326852
rect 340840 326800 340892 326852
rect 260156 326732 260208 326784
rect 341576 326732 341628 326784
rect 354180 326732 354232 326784
rect 257304 326664 257356 326716
rect 343968 326664 344020 326716
rect 356940 326664 356992 326716
rect 63368 326596 63420 326648
rect 66772 326596 66824 326648
rect 145524 326596 145576 326648
rect 157576 326596 157628 326648
rect 169076 326596 169128 326648
rect 246356 326596 246408 326648
rect 258224 326596 258276 326648
rect 343232 326596 343284 326648
rect 355652 326596 355704 326648
rect 58216 326528 58268 326580
rect 62448 326528 62500 326580
rect 150400 326528 150452 326580
rect 161624 326528 161676 326580
rect 337068 326528 337120 326580
rect 14700 326392 14752 326444
rect 148468 326460 148520 326512
rect 160244 326460 160296 326512
rect 248840 326460 248892 326512
rect 345624 326460 345676 326512
rect 61344 326392 61396 326444
rect 66404 326392 66456 326444
rect 147916 326392 147968 326444
rect 148744 326392 148796 326444
rect 152332 326392 152384 326444
rect 163096 326392 163148 326444
rect 74040 326324 74092 326376
rect 76064 326324 76116 326376
rect 145156 326324 145208 326376
rect 145892 326324 145944 326376
rect 147456 326324 147508 326376
rect 156932 326324 156984 326376
rect 242492 326324 242544 326376
rect 250220 326324 250272 326376
rect 75788 326256 75840 326308
rect 76984 326256 77036 326308
rect 136876 326256 136928 326308
rect 156288 326256 156340 326308
rect 161532 326256 161584 326308
rect 162268 326256 162320 326308
rect 254912 326256 254964 326308
rect 259236 326256 259288 326308
rect 137704 326231 137756 326240
rect 137704 326197 137713 326231
rect 137713 326197 137747 326231
rect 137747 326197 137756 326231
rect 137704 326188 137756 326197
rect 352892 325168 352944 325220
rect 325292 324828 325344 324880
rect 343876 324828 343928 324880
rect 347188 324828 347240 324880
rect 210016 323468 210068 323520
rect 211304 323468 211356 323520
rect 279108 323468 279160 323520
rect 280304 323468 280356 323520
rect 291528 323468 291580 323520
rect 292724 323468 292776 323520
rect 304040 323468 304092 323520
rect 305144 323468 305196 323520
rect 324740 323468 324792 323520
rect 325752 323468 325804 323520
rect 347004 323468 347056 323520
rect 351236 323468 351288 323520
rect 344336 323400 344388 323452
rect 348016 323400 348068 323452
rect 325568 322108 325620 322160
rect 344336 322108 344388 322160
rect 346452 322040 346504 322092
rect 350408 322040 350460 322092
rect 395120 320748 395172 320800
rect 395212 320748 395264 320800
rect 324832 320680 324884 320732
rect 325660 320680 325712 320732
rect 346452 320680 346504 320732
rect 62264 320612 62316 320664
rect 63276 320612 63328 320664
rect 248932 320612 248984 320664
rect 256936 320612 256988 320664
rect 337160 320612 337212 320664
rect 337528 320612 337580 320664
rect 339276 320612 339328 320664
rect 339552 320612 339604 320664
rect 339920 320612 339972 320664
rect 340564 320612 340616 320664
rect 58768 320476 58820 320528
rect 66864 320544 66916 320596
rect 248748 320544 248800 320596
rect 249208 320544 249260 320596
rect 346084 320544 346136 320596
rect 349396 320544 349448 320596
rect 63644 320476 63696 320528
rect 65024 320476 65076 320528
rect 336976 320476 337028 320528
rect 351604 320476 351656 320528
rect 60608 320408 60660 320460
rect 69072 320408 69124 320460
rect 338356 320408 338408 320460
rect 352248 320408 352300 320460
rect 59688 320340 59740 320392
rect 68428 320340 68480 320392
rect 247920 320340 247972 320392
rect 257120 320340 257172 320392
rect 335596 320340 335648 320392
rect 350684 320340 350736 320392
rect 57020 320272 57072 320324
rect 66496 320272 66548 320324
rect 243136 320272 243188 320324
rect 243780 320272 243832 320324
rect 245896 320272 245948 320324
rect 246448 320272 246500 320324
rect 334216 320272 334268 320324
rect 349764 320272 349816 320324
rect 56100 320204 56152 320256
rect 66312 320204 66364 320256
rect 156932 320204 156984 320256
rect 159968 320204 160020 320256
rect 246908 320204 246960 320256
rect 256292 320204 256344 320256
rect 332836 320204 332888 320256
rect 348016 320204 348068 320256
rect 62356 320136 62408 320188
rect 74776 320136 74828 320188
rect 246264 320136 246316 320188
rect 254912 320136 254964 320188
rect 331456 320136 331508 320188
rect 347280 320136 347332 320188
rect 61436 320068 61488 320120
rect 73396 320068 73448 320120
rect 149296 320068 149348 320120
rect 161532 320068 161584 320120
rect 243596 320068 243648 320120
rect 255464 320068 255516 320120
rect 335688 320068 335740 320120
rect 350960 320068 351012 320120
rect 55272 320000 55324 320052
rect 66680 320000 66732 320052
rect 147916 320000 147968 320052
rect 57940 319932 57992 319984
rect 69348 319932 69400 319984
rect 62448 319864 62500 319916
rect 64104 319864 64156 319916
rect 145156 319864 145208 319916
rect 238996 320000 239048 320052
rect 252796 320000 252848 320052
rect 334308 320000 334360 320052
rect 349396 320000 349448 320052
rect 241940 319932 241992 319984
rect 255556 319932 255608 319984
rect 332928 319932 332980 319984
rect 348568 319932 348620 319984
rect 66772 319796 66824 319848
rect 68612 319796 68664 319848
rect 161716 319864 161768 319916
rect 250220 319864 250272 319916
rect 254452 319864 254504 319916
rect 159048 319728 159100 319780
rect 250036 319728 250088 319780
rect 251784 319728 251836 319780
rect 338540 319592 338592 319644
rect 339552 319592 339604 319644
rect 249944 319456 249996 319508
rect 250956 319456 251008 319508
rect 65116 319320 65168 319372
rect 65944 319320 65996 319372
rect 152056 319320 152108 319372
rect 152792 319320 152844 319372
rect 155552 319320 155604 319372
rect 157300 319320 157352 319372
rect 161624 319320 161676 319372
rect 162636 319320 162688 319372
rect 325384 319320 325436 319372
rect 341208 319320 341260 319372
rect 341760 319320 341812 319372
rect 345164 319320 345216 319372
rect 348108 319320 348160 319372
rect 163096 318504 163148 318556
rect 164108 318504 164160 318556
rect 231084 317892 231136 317944
rect 231360 317892 231412 317944
rect 246172 317892 246224 317944
rect 254820 317892 254872 317944
rect 137796 316600 137848 316652
rect 325476 316600 325528 316652
rect 343048 316600 343100 316652
rect 429436 316600 429488 316652
rect 38804 315852 38856 315904
rect 55088 315852 55140 315904
rect 357676 315852 357728 315904
rect 358320 315852 358372 315904
rect 405976 315852 406028 315904
rect 352892 315172 352944 315224
rect 353076 315172 353128 315224
rect 38436 313744 38488 313796
rect 51592 313744 51644 313796
rect 356204 313744 356256 313796
rect 405976 313744 406028 313796
rect 76984 313540 77036 313592
rect 81676 313540 81728 313592
rect 165120 313064 165172 313116
rect 175516 313064 175568 313116
rect 258960 313064 259012 313116
rect 270276 313064 270328 313116
rect 76156 312452 76208 312504
rect 76984 312452 77036 312504
rect 137796 311092 137848 311144
rect 136968 310820 137020 310872
rect 395028 311024 395080 311076
rect 395212 311024 395264 311076
rect 38804 310276 38856 310328
rect 54076 310276 54128 310328
rect 356940 310276 356992 310328
rect 405976 310276 406028 310328
rect 137704 309664 137756 309716
rect 145524 309664 145576 309716
rect 231452 309664 231504 309716
rect 240652 309664 240704 309716
rect 325384 309664 325436 309716
rect 334216 309664 334268 309716
rect 356296 309664 356348 309716
rect 356940 309664 356992 309716
rect 38804 308236 38856 308288
rect 51224 308236 51276 308288
rect 136416 308236 136468 308288
rect 136968 308236 137020 308288
rect 356204 308236 356256 308288
rect 405976 308236 406028 308288
rect 352708 306876 352760 306928
rect 352892 306876 352944 306928
rect 38804 306196 38856 306248
rect 54076 306196 54128 306248
rect 354916 306196 354968 306248
rect 355652 306196 355704 306248
rect 406068 306196 406120 306248
rect 73396 305380 73448 305432
rect 75512 305380 75564 305432
rect 38620 304088 38672 304140
rect 51868 304156 51920 304208
rect 232096 304156 232148 304208
rect 232740 304156 232792 304208
rect 356204 304088 356256 304140
rect 405976 304088 406028 304140
rect 232004 301368 232056 301420
rect 233476 301368 233528 301420
rect 234120 301368 234172 301420
rect 38804 300620 38856 300672
rect 50304 300620 50356 300672
rect 355560 300620 355612 300672
rect 405976 300620 406028 300672
rect 355008 300008 355060 300060
rect 355560 300008 355612 300060
rect 136416 298648 136468 298700
rect 136876 298648 136928 298700
rect 38252 298580 38304 298632
rect 51684 298580 51736 298632
rect 356204 298580 356256 298632
rect 405976 298580 406028 298632
rect 74224 297152 74276 297204
rect 81676 297152 81728 297204
rect 167880 297152 167932 297204
rect 175516 297152 175568 297204
rect 261720 297152 261772 297204
rect 269356 297152 269408 297204
rect 137796 295860 137848 295912
rect 145432 295860 145484 295912
rect 231544 295860 231596 295912
rect 240928 295860 240980 295912
rect 325476 295860 325528 295912
rect 334216 295860 334268 295912
rect 353536 295792 353588 295844
rect 354180 295792 354232 295844
rect 38804 295112 38856 295164
rect 51316 295112 51368 295164
rect 353536 295112 353588 295164
rect 405976 295112 406028 295164
rect 38436 293752 38488 293804
rect 52604 293752 52656 293804
rect 356204 293752 356256 293804
rect 405976 293752 406028 293804
rect 427872 293208 427924 293260
rect 428792 293208 428844 293260
rect 427688 293140 427740 293192
rect 429896 293140 429948 293192
rect 352708 291755 352760 291764
rect 352708 291721 352717 291755
rect 352717 291721 352751 291755
rect 352751 291721 352760 291755
rect 352708 291712 352760 291721
rect 395028 291712 395080 291764
rect 395212 291712 395264 291764
rect 38528 291644 38580 291696
rect 50028 291644 50080 291696
rect 50028 291236 50080 291288
rect 51500 291236 51552 291288
rect 405976 290964 406028 291016
rect 230716 289060 230768 289112
rect 236052 289060 236104 289112
rect 38528 288924 38580 288976
rect 54536 288992 54588 289044
rect 356204 288924 356256 288976
rect 405976 288924 406028 288976
rect 395120 288899 395172 288908
rect 395120 288865 395129 288899
rect 395129 288865 395163 288899
rect 395163 288865 395172 288899
rect 395120 288856 395172 288865
rect 261720 286544 261772 286596
rect 266596 286544 266648 286596
rect 168064 286204 168116 286256
rect 172756 286204 172808 286256
rect 38528 285456 38580 285508
rect 49936 285456 49988 285508
rect 353720 285456 353772 285508
rect 405976 285456 406028 285508
rect 427964 283552 428016 283604
rect 429436 283552 429488 283604
rect 141660 283484 141712 283536
rect 145616 283484 145668 283536
rect 231820 283484 231872 283536
rect 240928 283484 240980 283536
rect 325200 283484 325252 283536
rect 334216 283484 334268 283536
rect 38528 283416 38580 283468
rect 52052 283416 52104 283468
rect 356204 283416 356256 283468
rect 405976 283416 406028 283468
rect 231636 282804 231688 282856
rect 236236 282804 236288 282856
rect 324556 282736 324608 282788
rect 330076 282736 330128 282788
rect 136876 282328 136928 282380
rect 142396 282328 142448 282380
rect 143040 282328 143092 282380
rect 236236 282056 236288 282108
rect 236880 282056 236932 282108
rect 395304 282056 395356 282108
rect 74132 280628 74184 280680
rect 81676 280628 81728 280680
rect 172756 280628 172808 280680
rect 175792 280628 175844 280680
rect 266596 280628 266648 280680
rect 270276 280628 270328 280680
rect 38068 279948 38120 280000
rect 48556 279948 48608 280000
rect 13596 279336 13648 279388
rect 18104 279336 18156 279388
rect 352984 279379 353036 279388
rect 352984 279345 352993 279379
rect 352993 279345 353027 279379
rect 353027 279345 353036 279379
rect 352984 279336 353036 279345
rect 38620 279268 38672 279320
rect 52604 279268 52656 279320
rect 356204 279268 356256 279320
rect 405976 279268 406028 279320
rect 395120 279200 395172 279252
rect 395304 279200 395356 279252
rect 51500 277908 51552 277960
rect 51684 277908 51736 277960
rect 137520 275120 137572 275172
rect 155920 275120 155972 275172
rect 234120 275120 234172 275172
rect 249116 275120 249168 275172
rect 138624 275052 138676 275104
rect 155276 275052 155328 275104
rect 339644 274984 339696 275036
rect 351236 274984 351288 275036
rect 149756 274916 149808 274968
rect 160520 274916 160572 274968
rect 337620 274916 337672 274968
rect 339092 274916 339144 274968
rect 341024 274916 341076 274968
rect 352156 274916 352208 274968
rect 151964 274848 152016 274900
rect 153436 274780 153488 274832
rect 154540 274780 154592 274832
rect 162728 274848 162780 274900
rect 247920 274848 247972 274900
rect 249576 274848 249628 274900
rect 338264 274848 338316 274900
rect 349580 274848 349632 274900
rect 163280 274780 163332 274832
rect 244056 274780 244108 274832
rect 254452 274780 254504 274832
rect 334124 274780 334176 274832
rect 346176 274780 346228 274832
rect 63092 274712 63144 274764
rect 65024 274712 65076 274764
rect 151044 274712 151096 274764
rect 151780 274712 151832 274764
rect 152240 274712 152292 274764
rect 153344 274712 153396 274764
rect 154080 274712 154132 274764
rect 154632 274712 154684 274764
rect 162084 274712 162136 274764
rect 243044 274712 243096 274764
rect 255740 274712 255792 274764
rect 336884 274712 336936 274764
rect 348752 274712 348804 274764
rect 34572 274644 34624 274696
rect 47084 274644 47136 274696
rect 59688 274644 59740 274696
rect 60884 274644 60936 274696
rect 147824 274644 147876 274696
rect 161440 274644 161492 274696
rect 240284 274644 240336 274696
rect 254544 274644 254596 274696
rect 335412 274644 335464 274696
rect 347004 274644 347056 274696
rect 29236 274576 29288 274628
rect 46624 274576 46676 274628
rect 62356 274576 62408 274628
rect 63552 274576 63604 274628
rect 65024 274576 65076 274628
rect 68612 274576 68664 274628
rect 145064 274576 145116 274628
rect 160244 274576 160296 274628
rect 241664 274576 241716 274628
rect 255096 274576 255148 274628
rect 256200 274576 256252 274628
rect 256936 274576 256988 274628
rect 335504 274576 335556 274628
rect 348108 274576 348160 274628
rect 26568 274508 26620 274560
rect 46532 274508 46584 274560
rect 146444 274508 146496 274560
rect 160888 274508 160940 274560
rect 238904 274508 238956 274560
rect 254268 274508 254320 274560
rect 332744 274508 332796 274560
rect 345348 274508 345400 274560
rect 23900 274440 23952 274492
rect 46440 274440 46492 274492
rect 57020 274440 57072 274492
rect 67140 274440 67192 274492
rect 143684 274440 143736 274492
rect 159324 274440 159376 274492
rect 159600 274440 159652 274492
rect 164568 274440 164620 274492
rect 237524 274440 237576 274492
rect 149204 274372 149256 274424
rect 149112 274304 149164 274356
rect 156840 274304 156892 274356
rect 245344 274304 245396 274356
rect 245804 274304 245856 274356
rect 247736 274440 247788 274492
rect 248564 274440 248616 274492
rect 345164 274440 345216 274492
rect 365312 274440 365364 274492
rect 369912 274440 369964 274492
rect 410208 274440 410260 274492
rect 253440 274304 253492 274356
rect 150492 274236 150544 274288
rect 341760 274236 341812 274288
rect 344612 274236 344664 274288
rect 254820 274168 254872 274220
rect 258316 274168 258368 274220
rect 249024 274032 249076 274084
rect 249944 274032 249996 274084
rect 60240 273964 60292 274016
rect 63276 273964 63328 274016
rect 250680 273964 250732 274016
rect 256384 273964 256436 274016
rect 344336 273964 344388 274016
rect 347372 273964 347424 274016
rect 63000 273896 63052 273948
rect 65944 273896 65996 273948
rect 246540 273896 246592 273948
rect 247184 273896 247236 273948
rect 253440 273896 253492 273948
rect 257580 273896 257632 273948
rect 343508 273896 343560 273948
rect 347280 273896 347332 273948
rect 61620 273828 61672 273880
rect 64104 273828 64156 273880
rect 66404 273828 66456 273880
rect 70360 273828 70412 273880
rect 234120 273828 234172 273880
rect 234764 273828 234816 273880
rect 243504 273828 243556 273880
rect 250772 273828 250824 273880
rect 339276 273828 339328 273880
rect 341852 273828 341904 273880
rect 342404 273828 342456 273880
rect 344520 273828 344572 273880
rect 21232 273760 21284 273812
rect 22244 273760 22296 273812
rect 61436 273760 61488 273812
rect 62264 273760 62316 273812
rect 63644 273760 63696 273812
rect 67692 273760 67744 273812
rect 162360 273760 162412 273812
rect 163924 273760 163976 273812
rect 338172 273760 338224 273812
rect 339000 273760 339052 273812
rect 340104 273760 340156 273812
rect 340932 273760 340984 273812
rect 348660 273760 348712 273812
rect 350408 273760 350460 273812
rect 13044 273692 13096 273744
rect 31904 273692 31956 273744
rect 138072 273692 138124 273744
rect 141660 273692 141712 273744
rect 247276 273692 247328 273744
rect 252152 273692 252204 273744
rect 31904 273012 31956 273064
rect 46716 273012 46768 273064
rect 51500 272468 51552 272520
rect 352800 272400 352852 272452
rect 352984 272400 353036 272452
rect 51408 269723 51460 269732
rect 51408 269689 51417 269723
rect 51417 269689 51451 269723
rect 51451 269689 51460 269723
rect 51408 269680 51460 269689
rect 88392 269612 88444 269664
rect 182416 269612 182468 269664
rect 276440 269612 276492 269664
rect 290700 269612 290752 269664
rect 395396 269612 395448 269664
rect 427596 269612 427648 269664
rect 429436 269612 429488 269664
rect 102652 269544 102704 269596
rect 196676 269544 196728 269596
rect 197504 269544 197556 269596
rect 189500 269476 189552 269528
rect 283524 269476 283576 269528
rect 127768 269340 127820 269392
rect 131172 269340 131224 269392
rect 95568 269000 95620 269052
rect 109736 269000 109788 269052
rect 189316 269000 189368 269052
rect 203760 269000 203812 269052
rect 284536 269000 284588 269052
rect 297784 269000 297836 269052
rect 95476 268932 95528 268984
rect 174872 268932 174924 268984
rect 189500 268932 189552 268984
rect 197504 268932 197556 268984
rect 264480 268932 264532 268984
rect 290700 268932 290752 268984
rect 114796 268524 114848 268576
rect 116912 268524 116964 268576
rect 209924 268252 209976 268304
rect 210936 268252 210988 268304
rect 303764 268252 303816 268304
rect 304960 268252 305012 268304
rect 51316 267844 51368 267896
rect 52052 267844 52104 267896
rect 354916 267844 354968 267896
rect 355836 267844 355888 267896
rect 333388 266824 333440 266876
rect 334124 266824 334176 266876
rect 334400 266824 334452 266876
rect 335412 266824 335464 266876
rect 337528 266824 337580 266876
rect 338264 266824 338316 266876
rect 347280 266824 347332 266876
rect 348936 266824 348988 266876
rect 64840 266756 64892 266808
rect 69348 266756 69400 266808
rect 245712 266756 245764 266808
rect 344520 266756 344572 266808
rect 347924 266756 347976 266808
rect 59504 266688 59556 266740
rect 71096 266688 71148 266740
rect 153252 266688 153304 266740
rect 162360 266688 162412 266740
rect 246264 266688 246316 266740
rect 256200 266688 256252 266740
rect 60884 266620 60936 266672
rect 72108 266620 72160 266672
rect 150584 266620 150636 266672
rect 161716 266620 161768 266672
rect 245804 266620 245856 266672
rect 256936 266620 256988 266672
rect 62264 266552 62316 266604
rect 74224 266552 74276 266604
rect 244424 266552 244476 266604
rect 255556 266552 255608 266604
rect 57664 266484 57716 266536
rect 60240 266484 60292 266536
rect 143040 266484 143092 266536
rect 155736 266484 155788 266536
rect 247644 266484 247696 266536
rect 253440 266484 253492 266536
rect 56744 266416 56796 266468
rect 67968 266416 68020 266468
rect 153344 266416 153396 266468
rect 165948 266416 166000 266468
rect 247184 266416 247236 266468
rect 259696 266484 259748 266536
rect 344612 266484 344664 266536
rect 346820 266484 346872 266536
rect 258316 266416 258368 266468
rect 341852 266416 341904 266468
rect 343784 266416 343836 266468
rect 55364 266348 55416 266400
rect 66956 266348 67008 266400
rect 151872 266348 151924 266400
rect 164568 266348 164620 266400
rect 236880 266348 236932 266400
rect 250036 266348 250088 266400
rect 58124 266280 58176 266332
rect 70084 266280 70136 266332
rect 153160 266280 153212 266332
rect 167328 266280 167380 266332
rect 247092 266280 247144 266332
rect 250772 266280 250824 266332
rect 252796 266280 252848 266332
rect 60792 266212 60844 266264
rect 73120 266212 73172 266264
rect 154540 266212 154592 266264
rect 168708 266212 168760 266264
rect 248564 266212 248616 266264
rect 262456 266280 262508 266332
rect 347372 266280 347424 266332
rect 349948 266280 350000 266332
rect 261076 266212 261128 266264
rect 340840 266212 340892 266264
rect 345808 266212 345860 266264
rect 63552 266144 63604 266196
rect 75236 266144 75288 266196
rect 154632 266144 154684 266196
rect 170088 266144 170140 266196
rect 244884 266144 244936 266196
rect 250680 266144 250732 266196
rect 151780 266076 151832 266128
rect 163096 266076 163148 266128
rect 248472 266076 248524 266128
rect 263836 266144 263888 266196
rect 338540 266144 338592 266196
rect 348660 266144 348712 266196
rect 61804 265872 61856 265924
rect 66588 265872 66640 265924
rect 59688 265736 59740 265788
rect 63092 265736 63144 265788
rect 251876 265736 251928 265788
rect 258960 265736 259012 265788
rect 58676 265668 58728 265720
rect 61620 265668 61672 265720
rect 157852 265668 157904 265720
rect 165120 265668 165172 265720
rect 339000 265668 339052 265720
rect 342680 265668 342732 265720
rect 60700 265600 60752 265652
rect 63000 265600 63052 265652
rect 154724 265600 154776 265652
rect 159600 265600 159652 265652
rect 249024 265600 249076 265652
rect 254820 265600 254872 265652
rect 340932 265600 340984 265652
rect 344796 265600 344848 265652
rect 62816 265532 62868 265584
rect 63644 265532 63696 265584
rect 63828 265532 63880 265584
rect 65024 265532 65076 265584
rect 67140 265532 67192 265584
rect 68980 265532 69032 265584
rect 156840 265532 156892 265584
rect 158956 265532 159008 265584
rect 339092 265532 339144 265584
rect 341668 265532 341720 265584
rect 77260 264036 77312 264088
rect 123260 264036 123312 264088
rect 124364 264036 124416 264088
rect 310756 264036 310808 264088
rect 312044 264036 312096 264088
rect 327316 264036 327368 264088
rect 154448 263560 154500 263612
rect 73856 263467 73908 263476
rect 73856 263433 73865 263467
rect 73865 263433 73899 263467
rect 73899 263433 73908 263467
rect 73856 263424 73908 263433
rect 74040 263424 74092 263476
rect 124364 263424 124416 263476
rect 140280 263424 140332 263476
rect 267240 263560 267292 263612
rect 310756 263560 310808 263612
rect 358412 263560 358464 263612
rect 249944 263492 249996 263544
rect 358412 263424 358464 263476
rect 369544 263356 369596 263408
rect 225932 262880 225984 262932
rect 233476 262880 233528 262932
rect 132092 262744 132144 262796
rect 139820 262744 139872 262796
rect 13320 262676 13372 262728
rect 372856 262676 372908 262728
rect 13412 262608 13464 262660
rect 381136 262608 381188 262660
rect 13504 262540 13556 262592
rect 385276 262540 385328 262592
rect 47084 262472 47136 262524
rect 49200 262472 49252 262524
rect 228600 262268 228652 262320
rect 369728 262268 369780 262320
rect 360436 261996 360488 262048
rect 360804 261996 360856 262048
rect 422536 261996 422588 262048
rect 79744 261384 79796 261436
rect 87196 261384 87248 261436
rect 132000 261384 132052 261436
rect 140372 261384 140424 261436
rect 225840 261384 225892 261436
rect 233476 261384 233528 261436
rect 95568 261316 95620 261368
rect 96212 261316 96264 261368
rect 203852 261248 203904 261300
rect 209924 261248 209976 261300
rect 297876 261248 297928 261300
rect 303764 261248 303816 261300
rect 189316 260840 189368 260892
rect 190512 260840 190564 260892
rect 217192 260636 217244 260688
rect 225196 260636 225248 260688
rect 311216 260636 311268 260688
rect 319220 260636 319272 260688
rect 123536 260568 123588 260620
rect 127768 260568 127820 260620
rect 110196 260432 110248 260484
rect 114796 260432 114848 260484
rect 79744 260024 79796 260076
rect 85080 260024 85132 260076
rect 132368 260024 132420 260076
rect 140372 260024 140424 260076
rect 226300 260024 226352 260076
rect 233476 260024 233528 260076
rect 360528 259276 360580 259328
rect 419776 259276 419828 259328
rect 79744 258664 79796 258716
rect 84436 258664 84488 258716
rect 132644 258596 132696 258648
rect 140556 258596 140608 258648
rect 226208 258596 226260 258648
rect 233476 258596 233528 258648
rect 324556 258596 324608 258648
rect 328420 258596 328472 258648
rect 321244 258392 321296 258444
rect 327224 258392 327276 258444
rect 131356 257304 131408 257356
rect 135128 257304 135180 257356
rect 132276 257236 132328 257288
rect 140556 257236 140608 257288
rect 179196 257236 179248 257288
rect 182324 257236 182376 257288
rect 226116 257236 226168 257288
rect 233476 257236 233528 257288
rect 267148 257236 267200 257288
rect 274876 257236 274928 257288
rect 321060 257168 321112 257220
rect 326764 257168 326816 257220
rect 360620 257168 360672 257220
rect 417016 257168 417068 257220
rect 85080 256828 85132 256880
rect 87196 256828 87248 256880
rect 131724 256488 131776 256540
rect 132368 256488 132420 256540
rect 225656 256488 225708 256540
rect 226300 256488 226352 256540
rect 181036 256080 181088 256132
rect 181680 256080 181732 256132
rect 136232 255944 136284 255996
rect 140556 255944 140608 255996
rect 174044 255944 174096 255996
rect 181036 255944 181088 255996
rect 229980 255944 230032 255996
rect 233476 255944 233528 255996
rect 79744 255876 79796 255928
rect 87380 255876 87432 255928
rect 132368 255876 132420 255928
rect 139544 255876 139596 255928
rect 178276 255876 178328 255928
rect 182324 255876 182376 255928
rect 226300 255876 226352 255928
rect 233568 255876 233620 255928
rect 266596 255876 266648 255928
rect 275704 255876 275756 255928
rect 80296 255808 80348 255860
rect 87196 255808 87248 255860
rect 320692 255808 320744 255860
rect 327224 255808 327276 255860
rect 84436 255740 84488 255792
rect 87288 255740 87340 255792
rect 320876 255604 320928 255656
rect 324556 255604 324608 255656
rect 173124 255536 173176 255588
rect 222712 255536 222764 255588
rect 226300 254584 226352 254636
rect 234120 254584 234172 254636
rect 131448 254516 131500 254568
rect 135036 254516 135088 254568
rect 173308 254516 173360 254568
rect 182324 254516 182376 254568
rect 225564 254516 225616 254568
rect 234304 254516 234356 254568
rect 131356 254448 131408 254500
rect 134944 254448 134996 254500
rect 137520 254448 137572 254500
rect 140556 254448 140608 254500
rect 173768 254448 173820 254500
rect 176160 254448 176212 254500
rect 176252 254448 176304 254500
rect 181588 254448 181640 254500
rect 266596 254448 266648 254500
rect 272760 254448 272812 254500
rect 321612 253632 321664 253684
rect 328052 253632 328104 253684
rect 172940 253224 172992 253276
rect 174780 253224 174832 253276
rect 266596 253156 266648 253208
rect 274232 253156 274284 253208
rect 79744 253088 79796 253140
rect 131356 253088 131408 253140
rect 138900 253088 138952 253140
rect 178920 253088 178972 253140
rect 181772 253088 181824 253140
rect 225380 253088 225432 253140
rect 230072 253088 230124 253140
rect 231452 253088 231504 253140
rect 234212 253088 234264 253140
rect 267884 253088 267936 253140
rect 274876 253088 274928 253140
rect 267424 253020 267476 253072
rect 267700 253020 267752 253072
rect 321612 253020 321664 253072
rect 328420 253020 328472 253072
rect 361172 253020 361224 253072
rect 414256 253020 414308 253072
rect 87288 252952 87340 253004
rect 79836 252884 79888 252936
rect 87196 252884 87248 252936
rect 321612 252000 321664 252052
rect 327224 252000 327276 252052
rect 173676 251864 173728 251916
rect 180300 251864 180352 251916
rect 131356 251796 131408 251848
rect 136324 251796 136376 251848
rect 179012 251796 179064 251848
rect 181588 251796 181640 251848
rect 79744 251728 79796 251780
rect 173584 251728 173636 251780
rect 181772 251728 181824 251780
rect 225748 251728 225800 251780
rect 234120 251728 234172 251780
rect 266596 251728 266648 251780
rect 272852 251728 272904 251780
rect 87196 251660 87248 251712
rect 13136 251456 13188 251508
rect 17552 251456 17604 251508
rect 222804 250980 222856 251032
rect 233476 250980 233528 251032
rect 320600 250572 320652 250624
rect 327132 250572 327184 250624
rect 79744 250368 79796 250420
rect 173676 250300 173728 250352
rect 182324 250300 182376 250352
rect 87196 250232 87248 250284
rect 135128 250232 135180 250284
rect 140556 250232 140608 250284
rect 173400 250232 173452 250284
rect 181496 250232 181548 250284
rect 226392 250232 226444 250284
rect 233476 250232 233528 250284
rect 267516 250232 267568 250284
rect 274876 250232 274928 250284
rect 361448 250232 361500 250284
rect 412876 250232 412928 250284
rect 77260 249552 77312 249604
rect 87196 249552 87248 249604
rect 321060 249484 321112 249536
rect 327224 249484 327276 249536
rect 173308 249416 173360 249468
rect 179196 249416 179248 249468
rect 321612 249076 321664 249128
rect 328420 249076 328472 249128
rect 132000 248940 132052 248992
rect 136140 248940 136192 248992
rect 174044 248940 174096 248992
rect 182232 248940 182284 248992
rect 225380 248940 225432 248992
rect 227312 248940 227364 248992
rect 173492 248872 173544 248924
rect 181956 248872 182008 248924
rect 267608 248872 267660 248924
rect 274968 248872 275020 248924
rect 173768 248804 173820 248856
rect 181864 248804 181916 248856
rect 267700 248804 267752 248856
rect 274876 248804 274928 248856
rect 266596 248736 266648 248788
rect 275060 248736 275112 248788
rect 77260 248192 77312 248244
rect 87196 248192 87248 248244
rect 173308 247852 173360 247904
rect 178276 247852 178328 247904
rect 321612 247648 321664 247700
rect 328420 247648 328472 247700
rect 77260 247512 77312 247564
rect 88484 247512 88536 247564
rect 173860 247512 173912 247564
rect 182324 247512 182376 247564
rect 266596 247512 266648 247564
rect 275888 247512 275940 247564
rect 321796 247512 321848 247564
rect 328420 247512 328472 247564
rect 267700 247444 267752 247496
rect 274876 247444 274928 247496
rect 135036 247308 135088 247360
rect 140648 247308 140700 247360
rect 173676 246900 173728 246952
rect 176252 246900 176304 246952
rect 321244 246220 321296 246272
rect 78916 246152 78968 246204
rect 87196 246152 87248 246204
rect 134944 246152 134996 246204
rect 140556 246152 140608 246204
rect 173952 246152 174004 246204
rect 181680 246152 181732 246204
rect 267792 246152 267844 246204
rect 274876 246152 274928 246204
rect 327868 246152 327920 246204
rect 427504 246152 427556 246204
rect 429436 246152 429488 246204
rect 131356 246084 131408 246136
rect 136232 246084 136284 246136
rect 266596 246084 266648 246136
rect 274416 246084 274468 246136
rect 225380 245472 225432 245524
rect 229980 245472 230032 245524
rect 321704 244860 321756 244912
rect 323176 244860 323228 244912
rect 80204 244792 80256 244844
rect 87196 244792 87248 244844
rect 321612 244792 321664 244844
rect 78916 244724 78968 244776
rect 87288 244724 87340 244776
rect 131356 244724 131408 244776
rect 137520 244724 137572 244776
rect 225564 244724 225616 244776
rect 232740 244724 232792 244776
rect 272760 244724 272812 244776
rect 274876 244724 274928 244776
rect 327868 244724 327920 244776
rect 176160 244656 176212 244708
rect 182048 244656 182100 244708
rect 230072 244656 230124 244708
rect 233568 244656 233620 244708
rect 173308 244384 173360 244436
rect 178920 244384 178972 244436
rect 321612 243432 321664 243484
rect 327040 243432 327092 243484
rect 136324 243364 136376 243416
rect 140648 243364 140700 243416
rect 174780 243364 174832 243416
rect 181036 243364 181088 243416
rect 226392 243364 226444 243416
rect 232832 243364 232884 243416
rect 272852 243364 272904 243416
rect 275796 243364 275848 243416
rect 323176 243364 323228 243416
rect 327868 243364 327920 243416
rect 132644 243296 132696 243348
rect 140464 243296 140516 243348
rect 267884 243228 267936 243280
rect 274324 243228 274376 243280
rect 131908 243160 131960 243212
rect 140556 243160 140608 243212
rect 226300 243092 226352 243144
rect 231452 243092 231504 243144
rect 172940 242752 172992 242804
rect 179012 242752 179064 242804
rect 321612 242208 321664 242260
rect 327224 242208 327276 242260
rect 79008 242140 79060 242192
rect 87288 242140 87340 242192
rect 79100 242072 79152 242124
rect 87196 242072 87248 242124
rect 320508 242072 320560 242124
rect 327132 242072 327184 242124
rect 123076 241596 123128 241648
rect 124318 241596 124370 241648
rect 78916 240576 78968 240628
rect 87380 240576 87432 240628
rect 133380 240576 133432 240628
rect 140556 240576 140608 240628
rect 227220 240576 227272 240628
rect 233476 240576 233528 240628
rect 267884 240576 267936 240628
rect 275612 240576 275664 240628
rect 389876 240576 389928 240628
rect 390704 240576 390756 240628
rect 393832 240576 393884 240628
rect 394844 240576 394896 240628
rect 13320 240508 13372 240560
rect 17460 240508 17512 240560
rect 368624 239896 368676 239948
rect 377824 239896 377876 239948
rect 314896 239828 314948 239880
rect 316092 239828 316144 239880
rect 185636 239284 185688 239336
rect 186464 239284 186516 239336
rect 279660 239284 279712 239336
rect 280304 239284 280356 239336
rect 132184 239216 132236 239268
rect 140556 239216 140608 239268
rect 226024 239216 226076 239268
rect 233476 239216 233528 239268
rect 267884 239216 267936 239268
rect 275520 239216 275572 239268
rect 136140 239148 136192 239200
rect 140188 239148 140240 239200
rect 227312 239148 227364 239200
rect 233568 239148 233620 239200
rect 267516 239148 267568 239200
rect 274140 239148 274192 239200
rect 136968 238604 137020 238656
rect 142396 238604 142448 238656
rect 142764 238604 142816 238656
rect 294196 238604 294248 238656
rect 325200 238604 325252 238656
rect 200172 238536 200224 238588
rect 230900 238536 230952 238588
rect 286928 238536 286980 238588
rect 325568 238536 325620 238588
rect 127860 237176 127912 237228
rect 140372 237176 140424 237228
rect 172940 237176 172992 237228
rect 219768 237176 219820 237228
rect 233476 237176 233528 237228
rect 267332 237176 267384 237228
rect 316276 237176 316328 237228
rect 78916 236564 78968 236616
rect 127860 236564 127912 236616
rect 128136 236564 128188 236616
rect 316276 236564 316328 236616
rect 328420 236564 328472 236616
rect 297692 236292 297744 236344
rect 262548 236156 262600 236208
rect 203760 235816 203812 235868
rect 230808 235816 230860 235868
rect 232004 235816 232056 235868
rect 297692 235816 297744 235868
rect 325384 235816 325436 235868
rect 136968 235204 137020 235256
rect 137152 235204 137204 235256
rect 148652 235204 148704 235256
rect 150676 235204 150728 235256
rect 149204 235136 149256 235188
rect 196492 235136 196544 235188
rect 232004 235136 232056 235188
rect 244976 235136 245028 235188
rect 262548 235136 262600 235188
rect 363840 235068 363892 235120
rect 368716 235068 368768 235120
rect 46900 234388 46952 234440
rect 73488 234388 73540 234440
rect 113508 234456 113560 234508
rect 137336 234456 137388 234508
rect 139268 234456 139320 234508
rect 74408 234388 74460 234440
rect 117096 234388 117148 234440
rect 137704 234388 137756 234440
rect 207256 234388 207308 234440
rect 231176 234388 231228 234440
rect 231820 234388 231872 234440
rect 302016 234388 302068 234440
rect 324556 234388 324608 234440
rect 346544 234388 346596 234440
rect 360528 234388 360580 234440
rect 221056 233776 221108 233828
rect 222160 233776 222212 233828
rect 324556 233776 324608 233828
rect 324740 233776 324792 233828
rect 345440 233776 345492 233828
rect 346544 233776 346596 233828
rect 138164 233708 138216 233760
rect 146812 233708 146864 233760
rect 150584 233708 150636 233760
rect 162268 233708 162320 233760
rect 234764 233708 234816 233760
rect 241480 233708 241532 233760
rect 248932 233708 248984 233760
rect 262088 233708 262140 233760
rect 268620 233708 268672 233760
rect 368900 233708 368952 233760
rect 427412 233708 427464 233760
rect 429804 233708 429856 233760
rect 62264 233640 62316 233692
rect 74224 233640 74276 233692
rect 157484 233640 157536 233692
rect 169996 233640 170048 233692
rect 246264 233640 246316 233692
rect 259236 233640 259288 233692
rect 322624 233640 322676 233692
rect 368716 233640 368768 233692
rect 55364 233164 55416 233216
rect 66956 233572 67008 233624
rect 160980 233572 161032 233624
rect 163188 233572 163240 233624
rect 244424 233572 244476 233624
rect 256292 233572 256344 233624
rect 323820 233572 323872 233624
rect 368808 233572 368860 233624
rect 62816 233504 62868 233556
rect 65852 233504 65904 233556
rect 153344 233504 153396 233556
rect 166132 233504 166184 233556
rect 248012 233504 248064 233556
rect 261168 233504 261220 233556
rect 64840 233436 64892 233488
rect 67232 233436 67284 233488
rect 151964 233436 152016 233488
rect 165212 233436 165264 233488
rect 250680 233436 250732 233488
rect 264020 233436 264072 233488
rect 63828 233368 63880 233420
rect 67140 233368 67192 233420
rect 154724 233368 154776 233420
rect 167236 233368 167288 233420
rect 61804 233300 61856 233352
rect 65760 233300 65812 233352
rect 56744 233232 56796 233284
rect 67968 233232 68020 233284
rect 63644 233164 63696 233216
rect 75236 233300 75288 233352
rect 150492 233300 150544 233352
rect 231452 233300 231504 233352
rect 234764 233300 234816 233352
rect 249852 233300 249904 233352
rect 263100 233300 263152 233352
rect 341024 233300 341076 233352
rect 346820 233300 346872 233352
rect 151872 233232 151924 233284
rect 164568 233232 164620 233284
rect 231728 233232 231780 233284
rect 243044 233232 243096 233284
rect 245344 233232 245396 233284
rect 258408 233232 258460 233284
rect 154632 233164 154684 233216
rect 168064 233164 168116 233216
rect 231636 233164 231688 233216
rect 242124 233164 242176 233216
rect 244332 233164 244384 233216
rect 257304 233164 257356 233216
rect 58124 233096 58176 233148
rect 70084 233096 70136 233148
rect 144604 233096 144656 233148
rect 165120 233096 165172 233148
rect 238628 233096 238680 233148
rect 258960 233096 259012 233148
rect 60792 233028 60844 233080
rect 72108 233028 72160 233080
rect 74132 233028 74184 233080
rect 75144 233028 75196 233080
rect 105136 233028 105188 233080
rect 137152 233028 137204 233080
rect 145248 233028 145300 233080
rect 352892 233028 352944 233080
rect 340932 232960 340984 233012
rect 347924 232960 347976 233012
rect 60884 232892 60936 232944
rect 73120 232892 73172 232944
rect 163280 232892 163332 232944
rect 247092 232892 247144 232944
rect 260156 232892 260208 232944
rect 59504 232824 59556 232876
rect 71096 232824 71148 232876
rect 156012 232824 156064 232876
rect 169076 232824 169128 232876
rect 160060 232756 160112 232808
rect 161808 232756 161860 232808
rect 58676 232620 58728 232672
rect 63184 232620 63236 232672
rect 156104 232620 156156 232672
rect 158220 232620 158272 232672
rect 57664 232552 57716 232604
rect 61620 232552 61672 232604
rect 157116 232552 157168 232604
rect 159048 232552 159100 232604
rect 59688 232484 59740 232536
rect 63000 232484 63052 232536
rect 65944 232484 65996 232536
rect 68520 232484 68572 232536
rect 155184 232484 155236 232536
rect 157576 232484 157628 232536
rect 158128 232484 158180 232536
rect 160336 232484 160388 232536
rect 248288 232484 248340 232536
rect 250128 232484 250180 232536
rect 339000 232484 339052 232536
rect 341668 232484 341720 232536
rect 342864 232484 342916 232536
rect 345808 232484 345860 232536
rect 346728 232484 346780 232536
rect 349948 232484 350000 232536
rect 60700 232416 60752 232468
rect 63092 232416 63144 232468
rect 67324 232416 67376 232468
rect 68980 232416 69032 232468
rect 154264 232416 154316 232468
rect 156380 232416 156432 232468
rect 158864 232416 158916 232468
rect 160980 232416 161032 232468
rect 161992 232416 162044 232468
rect 163004 232416 163056 232468
rect 239548 232416 239600 232468
rect 240284 232416 240336 232468
rect 249944 232416 249996 232468
rect 252888 232416 252940 232468
rect 333388 232416 333440 232468
rect 334124 232416 334176 232468
rect 334400 232416 334452 232468
rect 335412 232416 335464 232468
rect 338540 232416 338592 232468
rect 339644 232416 339696 232468
rect 342956 232416 343008 232468
rect 344796 232416 344848 232468
rect 346636 232416 346688 232468
rect 348936 232416 348988 232468
rect 134852 232348 134904 232400
rect 368900 232348 368952 232400
rect 265860 232280 265912 232332
rect 368716 232280 368768 232332
rect 326580 232212 326632 232264
rect 368808 232212 368860 232264
rect 354916 232008 354968 232060
rect 355836 232008 355888 232060
rect 239640 231668 239692 231720
rect 324648 231668 324700 231720
rect 345164 231668 345216 231720
rect 360712 231668 360764 231720
rect 370004 231464 370056 231516
rect 369912 231260 369964 231312
rect 222620 230988 222672 231040
rect 222804 230988 222856 231040
rect 325568 230988 325620 231040
rect 343968 230988 344020 231040
rect 345164 230988 345216 231040
rect 12860 230920 12912 230972
rect 16172 230920 16224 230972
rect 47084 230920 47136 230972
rect 368900 230920 368952 230972
rect 76800 230852 76852 230904
rect 368716 230852 368768 230904
rect 134760 230784 134812 230836
rect 368808 230784 368860 230836
rect 115992 230376 116044 230428
rect 127216 230376 127268 230428
rect 210016 230376 210068 230428
rect 221056 230376 221108 230428
rect 304040 230376 304092 230428
rect 314896 230376 314948 230428
rect 103480 230308 103532 230360
rect 123076 230308 123128 230360
rect 197504 230308 197556 230360
rect 218296 230308 218348 230360
rect 291528 230308 291580 230360
rect 312136 230308 312188 230360
rect 339644 230308 339696 230360
rect 91060 230240 91112 230292
rect 120316 230240 120368 230292
rect 185084 230240 185136 230292
rect 214156 230240 214208 230292
rect 279108 230240 279160 230292
rect 307996 230240 308048 230292
rect 343784 230240 343836 230292
rect 360804 230240 360856 230292
rect 324648 229628 324700 229680
rect 325476 229628 325528 229680
rect 343048 229628 343100 229680
rect 343784 229628 343836 229680
rect 22244 229560 22296 229612
rect 368716 229560 368768 229612
rect 74040 228404 74092 228456
rect 368716 228404 368768 228456
rect 47084 228336 47136 228388
rect 368808 228336 368860 228388
rect 34020 228268 34072 228320
rect 368716 228268 368768 228320
rect 305144 227656 305196 227708
rect 322992 227656 323044 227708
rect 347004 227656 347056 227708
rect 360436 227656 360488 227708
rect 222436 227588 222488 227640
rect 222620 227588 222672 227640
rect 280304 227588 280356 227640
rect 353076 227588 353128 227640
rect 186464 227520 186516 227572
rect 369084 227520 369136 227572
rect 322992 226976 323044 227028
rect 347004 226976 347056 227028
rect 76800 226908 76852 226960
rect 368808 226908 368860 226960
rect 34572 226840 34624 226892
rect 368716 226840 368768 226892
rect 240284 226228 240336 226280
rect 353260 226228 353312 226280
rect 231360 226160 231412 226212
rect 353168 226160 353220 226212
rect 137612 226092 137664 226144
rect 353352 226092 353404 226144
rect 324556 225684 324608 225736
rect 325384 225684 325436 225736
rect 345716 225684 345768 225736
rect 172020 225616 172072 225668
rect 368808 225616 368860 225668
rect 137520 225548 137572 225600
rect 368716 225548 368768 225600
rect 134760 225480 134812 225532
rect 368900 225480 368952 225532
rect 251232 225412 251284 225464
rect 253992 225412 254044 225464
rect 255004 225412 255056 225464
rect 257488 225412 257540 225464
rect 338356 225412 338408 225464
rect 62356 225344 62408 225396
rect 63644 225344 63696 225396
rect 249208 225344 249260 225396
rect 252152 225344 252204 225396
rect 252244 225344 252296 225396
rect 254820 225344 254872 225396
rect 256016 225344 256068 225396
rect 258408 225344 258460 225396
rect 337160 225344 337212 225396
rect 339000 225344 339052 225396
rect 340196 225344 340248 225396
rect 341024 225344 341076 225396
rect 341392 225412 341444 225464
rect 346636 225412 346688 225464
rect 56100 225276 56152 225328
rect 56744 225276 56796 225328
rect 59688 225276 59740 225328
rect 60792 225276 60844 225328
rect 61436 225276 61488 225328
rect 62264 225276 62316 225328
rect 63184 225276 63236 225328
rect 64104 225276 64156 225328
rect 65760 225276 65812 225328
rect 66772 225276 66824 225328
rect 68520 225276 68572 225328
rect 70360 225276 70412 225328
rect 153712 225276 153764 225328
rect 154724 225276 154776 225328
rect 155460 225276 155512 225328
rect 156104 225276 156156 225328
rect 156380 225276 156432 225328
rect 157484 225276 157536 225328
rect 228600 225276 228652 225328
rect 61620 225208 61672 225260
rect 63276 225208 63328 225260
rect 65852 225208 65904 225260
rect 67692 225208 67744 225260
rect 254084 225208 254136 225260
rect 256660 225208 256712 225260
rect 339552 225208 339604 225260
rect 342036 225344 342088 225396
rect 346728 225344 346780 225396
rect 368716 225276 368768 225328
rect 343508 225208 343560 225260
rect 351604 225208 351656 225260
rect 151044 225140 151096 225192
rect 151872 225140 151924 225192
rect 163004 225140 163056 225192
rect 164384 225140 164436 225192
rect 252612 225140 252664 225192
rect 255740 225140 255792 225192
rect 339000 225140 339052 225192
rect 342956 225140 343008 225192
rect 63092 225072 63144 225124
rect 65944 225072 65996 225124
rect 335412 225072 335464 225124
rect 348568 225072 348620 225124
rect 58768 225004 58820 225056
rect 59504 225004 59556 225056
rect 337712 225004 337764 225056
rect 342588 225004 342640 225056
rect 342680 225004 342732 225056
rect 352248 225140 352300 225192
rect 63000 224936 63052 224988
rect 65024 224936 65076 224988
rect 334124 224936 334176 224988
rect 348016 224936 348068 224988
rect 335504 224868 335556 224920
rect 349396 224868 349448 224920
rect 149296 224800 149348 224852
rect 150584 224800 150636 224852
rect 332744 224800 332796 224852
rect 340840 224800 340892 224852
rect 341300 224800 341352 224852
rect 57020 224732 57072 224784
rect 67324 224732 67376 224784
rect 342864 224732 342916 224784
rect 343048 224732 343100 224784
rect 360620 224732 360672 224784
rect 338264 224596 338316 224648
rect 350684 224596 350736 224648
rect 67232 224528 67284 224580
rect 69440 224528 69492 224580
rect 339644 224528 339696 224580
rect 336884 224460 336936 224512
rect 349764 224460 349816 224512
rect 347280 224392 347332 224444
rect 160980 224324 161032 224376
rect 161716 224324 161768 224376
rect 325660 224324 325712 224376
rect 343048 224324 343100 224376
rect 67140 224256 67192 224308
rect 68612 224256 68664 224308
rect 325384 224256 325436 224308
rect 325752 224256 325804 224308
rect 344244 224256 344296 224308
rect 158220 224188 158272 224240
rect 159048 224188 159100 224240
rect 325200 224188 325252 224240
rect 325844 224188 325896 224240
rect 345164 224188 345216 224240
rect 243596 224120 243648 224172
rect 244424 224120 244476 224172
rect 322624 224120 322676 224172
rect 368808 224120 368860 224172
rect 369084 223712 369136 223764
rect 369360 223712 369412 223764
rect 351282 223032 351334 223084
rect 363840 222896 363892 222948
rect 368900 222896 368952 222948
rect 323820 222828 323872 222880
rect 368716 222828 368768 222880
rect 322716 222760 322768 222812
rect 368808 222760 368860 222812
rect 250128 222692 250180 222744
rect 250956 222692 251008 222744
rect 34572 221740 34624 221792
rect 34940 221740 34992 221792
rect 34020 221672 34072 221724
rect 34756 221672 34808 221724
rect 361080 221468 361132 221520
rect 368900 221468 368952 221520
rect 325200 221400 325252 221452
rect 368808 221400 368860 221452
rect 322900 221332 322952 221384
rect 368716 221332 368768 221384
rect 325292 220584 325344 220636
rect 353444 220584 353496 220636
rect 34664 220516 34716 220568
rect 34940 220516 34992 220568
rect 325384 220516 325436 220568
rect 368808 220516 368860 220568
rect 34756 220448 34808 220500
rect 322808 220448 322860 220500
rect 368716 220448 368768 220500
rect 38068 219904 38120 219956
rect 51868 219972 51920 220024
rect 359700 219972 359752 220024
rect 368900 219972 368952 220024
rect 76156 219496 76208 219548
rect 81676 219496 81728 219548
rect 369084 219471 369136 219480
rect 369084 219437 369093 219471
rect 369093 219437 369127 219471
rect 369127 219437 369136 219471
rect 369084 219428 369136 219437
rect 13044 219360 13096 219412
rect 16356 219360 16408 219412
rect 368900 219360 368952 219412
rect 369268 219360 369320 219412
rect 369360 219403 369412 219412
rect 369360 219369 369369 219403
rect 369369 219369 369403 219403
rect 369403 219369 369412 219403
rect 369360 219360 369412 219369
rect 165120 219224 165172 219276
rect 179288 219224 179340 219276
rect 258960 219224 259012 219276
rect 272944 219224 272996 219276
rect 368992 218952 369044 219004
rect 369176 218952 369228 219004
rect 365220 218680 365272 218732
rect 368808 218680 368860 218732
rect 352800 218612 352852 218664
rect 368716 218612 368768 218664
rect 394844 218612 394896 218664
rect 405976 218612 406028 218664
rect 352892 218476 352944 218528
rect 368808 218476 368860 218528
rect 352984 217184 353036 217236
rect 368716 217184 368768 217236
rect 38528 217116 38580 217168
rect 53248 217116 53300 217168
rect 353352 217116 353404 217168
rect 368808 217116 368860 217168
rect 358412 217048 358464 217100
rect 368716 217048 368768 217100
rect 369084 216887 369136 216896
rect 369084 216853 369093 216887
rect 369093 216853 369127 216887
rect 369127 216853 369136 216887
rect 369084 216844 369136 216853
rect 369084 216708 369136 216760
rect 137612 215824 137664 215876
rect 145156 215824 145208 215876
rect 231360 215824 231412 215876
rect 240928 215824 240980 215876
rect 325292 215824 325344 215876
rect 334216 215824 334268 215876
rect 353168 215756 353220 215808
rect 368992 215756 369044 215808
rect 353260 215688 353312 215740
rect 368716 215688 368768 215740
rect 358320 215620 358372 215672
rect 368808 215620 368860 215672
rect 369820 214532 369872 214584
rect 38528 214396 38580 214448
rect 51684 214464 51736 214516
rect 74224 214464 74276 214516
rect 74408 214464 74460 214516
rect 353076 214396 353128 214448
rect 368716 214396 368768 214448
rect 368992 214439 369044 214448
rect 368992 214405 369001 214439
rect 369001 214405 369035 214439
rect 369035 214405 369044 214439
rect 368992 214396 369044 214405
rect 361172 214260 361224 214312
rect 368900 214260 368952 214312
rect 356204 214056 356256 214108
rect 405976 214056 406028 214108
rect 355100 213988 355152 214040
rect 394844 213988 394896 214040
rect 365312 213920 365364 213972
rect 368900 213920 368952 213972
rect 34848 213895 34900 213904
rect 34848 213861 34857 213895
rect 34857 213861 34891 213895
rect 34891 213861 34900 213895
rect 34848 213852 34900 213861
rect 353444 213036 353496 213088
rect 368716 213036 368768 213088
rect 262364 211744 262416 211796
rect 268620 211744 268672 211796
rect 167972 211676 168024 211728
rect 174780 211676 174832 211728
rect 369912 211608 369964 211660
rect 370740 211608 370792 211660
rect 38712 210928 38764 210980
rect 54076 210928 54128 210980
rect 354916 210928 354968 210980
rect 405976 210928 406028 210980
rect 378284 210316 378336 210368
rect 383896 210316 383948 210368
rect 369176 209840 369228 209892
rect 369820 209840 369872 209892
rect 174780 209636 174832 209688
rect 178920 209636 178972 209688
rect 38528 209568 38580 209620
rect 51408 209568 51460 209620
rect 356020 209568 356072 209620
rect 405976 209568 406028 209620
rect 368992 209500 369044 209552
rect 369268 209500 369320 209552
rect 427320 208820 427372 208872
rect 429620 208820 429672 208872
rect 13044 208140 13096 208192
rect 16448 208140 16500 208192
rect 268620 207460 268672 207512
rect 272944 207460 272996 207512
rect 34848 206891 34900 206900
rect 34848 206857 34857 206891
rect 34857 206857 34891 206891
rect 34891 206857 34900 206891
rect 34848 206848 34900 206857
rect 38528 206780 38580 206832
rect 51408 206780 51460 206832
rect 355008 206780 355060 206832
rect 405976 206780 406028 206832
rect 38528 204740 38580 204792
rect 51408 204740 51460 204792
rect 136876 204740 136928 204792
rect 145340 204740 145392 204792
rect 232004 204740 232056 204792
rect 239640 204740 239692 204792
rect 356204 204740 356256 204792
rect 406068 204740 406120 204792
rect 34848 204715 34900 204724
rect 34848 204681 34857 204715
rect 34857 204681 34891 204715
rect 34891 204681 34900 204715
rect 34848 204672 34900 204681
rect 368992 204672 369044 204724
rect 369176 204672 369228 204724
rect 74316 203312 74368 203364
rect 81676 203312 81728 203364
rect 137796 202020 137848 202072
rect 145432 202020 145484 202072
rect 231452 202020 231504 202072
rect 240652 202020 240704 202072
rect 325476 202020 325528 202072
rect 334216 202020 334268 202072
rect 38528 201272 38580 201324
rect 51500 201272 51552 201324
rect 353536 201272 353588 201324
rect 405976 201272 406028 201324
rect 368900 199912 368952 199964
rect 369176 199912 369228 199964
rect 427136 199708 427188 199760
rect 428792 199708 428844 199760
rect 369820 199479 369872 199488
rect 369820 199445 369829 199479
rect 369829 199445 369863 199479
rect 369863 199445 369872 199479
rect 369820 199436 369872 199445
rect 13320 199300 13372 199352
rect 17644 199300 17696 199352
rect 38528 199232 38580 199284
rect 51776 199232 51828 199284
rect 355928 199232 355980 199284
rect 405976 199232 406028 199284
rect 13044 197736 13096 197788
rect 16264 197736 16316 197788
rect 427688 196512 427740 196564
rect 429528 196512 429580 196564
rect 38528 195764 38580 195816
rect 51316 195764 51368 195816
rect 352708 195764 352760 195816
rect 405976 195764 406028 195816
rect 369912 195220 369964 195272
rect 368992 195152 369044 195204
rect 369360 195152 369412 195204
rect 369728 195152 369780 195204
rect 38804 195084 38856 195136
rect 51316 195084 51368 195136
rect 356204 195084 356256 195136
rect 406068 195084 406120 195136
rect 230808 194472 230860 194524
rect 235316 194472 235368 194524
rect 369912 192364 369964 192416
rect 369912 192228 369964 192280
rect 38804 191616 38856 191668
rect 49936 191616 49988 191668
rect 352892 191616 352944 191668
rect 405976 191616 406028 191668
rect 426860 189848 426912 189900
rect 429344 189848 429396 189900
rect 13412 189644 13464 189696
rect 17092 189644 17144 189696
rect 38068 189576 38120 189628
rect 51776 189576 51828 189628
rect 355192 189576 355244 189628
rect 405976 189576 406028 189628
rect 324556 188896 324608 188948
rect 330076 188896 330128 188948
rect 232004 188760 232056 188812
rect 236236 188760 236288 188812
rect 137796 188284 137848 188336
rect 142396 188284 142448 188336
rect 143040 188284 143092 188336
rect 236236 188284 236288 188336
rect 236880 188284 236932 188336
rect 138900 188216 138952 188268
rect 145616 188216 145668 188268
rect 232740 188216 232792 188268
rect 240928 188216 240980 188268
rect 326580 188216 326632 188268
rect 334216 188216 334268 188268
rect 75420 186788 75472 186840
rect 81676 186788 81728 186840
rect 169260 186788 169312 186840
rect 178920 186788 178972 186840
rect 263100 186788 263152 186840
rect 272944 186788 272996 186840
rect 13044 186652 13096 186704
rect 16080 186652 16132 186704
rect 38068 186108 38120 186160
rect 48556 186108 48608 186160
rect 352800 186108 352852 186160
rect 405976 186108 406028 186160
rect 369084 185428 369136 185480
rect 369728 185428 369780 185480
rect 38804 184000 38856 184052
rect 51408 184000 51460 184052
rect 356204 184000 356256 184052
rect 405976 184000 406028 184052
rect 34388 183184 34440 183236
rect 34940 183184 34992 183236
rect 369820 182751 369872 182760
rect 369820 182717 369829 182751
rect 369829 182717 369863 182751
rect 369863 182717 369872 182751
rect 369820 182708 369872 182717
rect 34572 182640 34624 182692
rect 34756 182640 34808 182692
rect 261076 182028 261128 182080
rect 267516 182028 267568 182080
rect 21600 181280 21652 181332
rect 34388 181280 34440 181332
rect 59688 181280 59740 181332
rect 60884 181280 60936 181332
rect 61436 181280 61488 181332
rect 62172 181280 62224 181332
rect 245344 181280 245396 181332
rect 245804 181280 245856 181332
rect 247736 181280 247788 181332
rect 248380 181280 248432 181332
rect 337620 181280 337672 181332
rect 341116 181280 341168 181332
rect 344980 181280 345032 181332
rect 359700 181280 359752 181332
rect 370740 181280 370792 181332
rect 410208 181280 410260 181332
rect 60792 181212 60844 181264
rect 65024 181212 65076 181264
rect 338264 181212 338316 181264
rect 341760 181212 341812 181264
rect 343508 181212 343560 181264
rect 59412 181144 59464 181196
rect 64104 181144 64156 181196
rect 149756 181144 149808 181196
rect 159600 181144 159652 181196
rect 344336 181144 344388 181196
rect 347280 181212 347332 181264
rect 350408 181212 350460 181264
rect 348108 181144 348160 181196
rect 149204 181076 149256 181128
rect 158956 181076 159008 181128
rect 248472 181076 248524 181128
rect 257580 181076 257632 181128
rect 339644 181076 339696 181128
rect 351236 181076 351288 181128
rect 151964 181008 152016 181060
rect 163280 181008 163332 181060
rect 243504 181008 243556 181060
rect 252796 181008 252848 181060
rect 334124 181008 334176 181060
rect 346176 181008 346228 181060
rect 66404 180940 66456 180992
rect 70360 180940 70412 180992
rect 150308 180940 150360 180992
rect 162728 180940 162780 180992
rect 244056 180940 244108 180992
rect 253440 180940 253492 180992
rect 335504 180940 335556 180992
rect 347004 180940 347056 180992
rect 34664 180872 34716 180924
rect 46992 180872 47044 180924
rect 62356 180872 62408 180924
rect 63552 180872 63604 180924
rect 147824 180872 147876 180924
rect 161440 180872 161492 180924
rect 241664 180872 241716 180924
rect 255096 180872 255148 180924
rect 336884 180872 336936 180924
rect 348752 180872 348804 180924
rect 31812 180804 31864 180856
rect 46716 180804 46768 180856
rect 64932 180804 64984 180856
rect 68612 180804 68664 180856
rect 149204 180804 149256 180856
rect 162084 180804 162136 180856
rect 243044 180804 243096 180856
rect 255740 180804 255792 180856
rect 338264 180804 338316 180856
rect 349580 180804 349632 180856
rect 29512 180736 29564 180788
rect 46624 180736 46676 180788
rect 65024 180736 65076 180788
rect 69440 180736 69492 180788
rect 145064 180736 145116 180788
rect 160244 180736 160296 180788
rect 240284 180736 240336 180788
rect 254544 180736 254596 180788
rect 340932 180736 340984 180788
rect 349396 180736 349448 180788
rect 26936 180668 26988 180720
rect 46532 180668 46584 180720
rect 146444 180668 146496 180720
rect 160888 180668 160940 180720
rect 237524 180668 237576 180720
rect 253532 180668 253584 180720
rect 332744 180668 332796 180720
rect 345440 180668 345492 180720
rect 24176 180600 24228 180652
rect 46440 180600 46492 180652
rect 57020 180600 57072 180652
rect 67140 180600 67192 180652
rect 143684 180600 143736 180652
rect 159324 180600 159376 180652
rect 238904 180600 238956 180652
rect 254176 180600 254228 180652
rect 335412 180600 335464 180652
rect 348016 180600 348068 180652
rect 254820 180532 254872 180584
rect 256936 180532 256988 180584
rect 352156 180532 352208 180584
rect 340104 180328 340156 180380
rect 341024 180328 341076 180380
rect 341668 180192 341720 180244
rect 345992 180192 346044 180244
rect 60608 180124 60660 180176
rect 65944 180124 65996 180176
rect 63276 180056 63328 180108
rect 57848 179988 57900 180040
rect 62264 179988 62316 180040
rect 66772 179988 66824 180040
rect 340840 179988 340892 180040
rect 345256 179988 345308 180040
rect 63644 179920 63696 179972
rect 67692 179920 67744 179972
rect 152240 179920 152292 179972
rect 153252 179920 153304 179972
rect 153436 179920 153488 179972
rect 154632 179920 154684 179972
rect 342404 179920 342456 179972
rect 345900 179920 345952 179972
rect 230992 179716 231044 179768
rect 232740 179716 232792 179768
rect 324556 179444 324608 179496
rect 326580 179444 326632 179496
rect 273864 178492 273916 178544
rect 276256 178492 276308 178544
rect 369084 175840 369136 175892
rect 369912 175840 369964 175892
rect 13044 175772 13096 175824
rect 16080 175772 16132 175824
rect 88392 175772 88444 175824
rect 182416 175772 182468 175824
rect 182968 175772 183020 175824
rect 276440 175772 276492 175824
rect 95476 175704 95528 175756
rect 174872 175704 174924 175756
rect 189316 175704 189368 175756
rect 189500 175704 189552 175756
rect 283524 175704 283576 175756
rect 196676 175636 196728 175688
rect 264480 175636 264532 175688
rect 290700 175636 290752 175688
rect 96764 175160 96816 175212
rect 109736 175160 109788 175212
rect 112680 175160 112732 175212
rect 116912 175160 116964 175212
rect 174872 175160 174924 175212
rect 176160 175160 176212 175212
rect 189316 175160 189368 175212
rect 190604 175160 190656 175212
rect 203760 175160 203812 175212
rect 102652 175092 102704 175144
rect 174780 175092 174832 175144
rect 196676 175092 196728 175144
rect 285824 175092 285876 175144
rect 297784 175092 297836 175144
rect 354916 175092 354968 175144
rect 355836 175092 355888 175144
rect 206520 174752 206572 174804
rect 210936 174752 210988 174804
rect 129240 174412 129292 174464
rect 131172 174412 131224 174464
rect 300360 174412 300412 174464
rect 304960 174412 305012 174464
rect 57848 172984 57900 173036
rect 58124 172984 58176 173036
rect 58676 172984 58728 173036
rect 59412 172984 59464 173036
rect 59688 172984 59740 173036
rect 60792 172984 60844 173036
rect 62816 172984 62868 173036
rect 63644 172984 63696 173036
rect 63828 172984 63880 173036
rect 64932 172984 64984 173036
rect 67140 172984 67192 173036
rect 68980 172984 69032 173036
rect 153160 172984 153212 173036
rect 153344 172984 153396 173036
rect 159600 172984 159652 173036
rect 160336 172984 160388 173036
rect 253440 172984 253492 173036
rect 254176 172984 254228 173036
rect 333388 172984 333440 173036
rect 334124 172984 334176 173036
rect 341760 172984 341812 173036
rect 342680 172984 342732 173036
rect 345992 172984 346044 173036
rect 346820 172984 346872 173036
rect 427596 172984 427648 173036
rect 429896 172984 429948 173036
rect 154724 172916 154776 172968
rect 164660 172916 164712 172968
rect 246264 172916 246316 172968
rect 254820 172916 254872 172968
rect 258684 172916 258736 172968
rect 341024 172916 341076 172968
rect 344796 172916 344848 172968
rect 345900 172916 345952 172968
rect 347924 172916 347976 172968
rect 153344 172848 153396 172900
rect 163924 172848 163976 172900
rect 244884 172848 244936 172900
rect 256752 172848 256804 172900
rect 334400 172848 334452 172900
rect 335504 172848 335556 172900
rect 339552 172848 339604 172900
rect 343784 172848 343836 172900
rect 59504 172780 59556 172832
rect 71096 172780 71148 172832
rect 150400 172780 150452 172832
rect 161716 172780 161768 172832
rect 60884 172712 60936 172764
rect 72108 172712 72160 172764
rect 151320 172712 151372 172764
rect 163096 172712 163148 172764
rect 244424 172712 244476 172764
rect 255556 172712 255608 172764
rect 57940 172644 57992 172696
rect 70084 172644 70136 172696
rect 143040 172644 143092 172696
rect 155736 172644 155788 172696
rect 157852 172644 157904 172696
rect 165120 172644 165172 172696
rect 245528 172644 245580 172696
rect 258316 172644 258368 172696
rect 55364 172576 55416 172628
rect 66956 172576 67008 172628
rect 153252 172576 153304 172628
rect 165856 172576 165908 172628
rect 246816 172576 246868 172628
rect 259696 172576 259748 172628
rect 56744 172508 56796 172560
rect 67968 172508 68020 172560
rect 151596 172508 151648 172560
rect 164476 172508 164528 172560
rect 236880 172508 236932 172560
rect 250036 172508 250088 172560
rect 63552 172440 63604 172492
rect 75236 172440 75288 172492
rect 153160 172440 153212 172492
rect 167328 172440 167380 172492
rect 246908 172440 246960 172492
rect 261168 172440 261220 172492
rect 62172 172372 62224 172424
rect 74224 172372 74276 172424
rect 154540 172372 154592 172424
rect 168708 172372 168760 172424
rect 248380 172372 248432 172424
rect 262456 172372 262508 172424
rect 60700 172304 60752 172356
rect 73120 172304 73172 172356
rect 154632 172304 154684 172356
rect 170088 172304 170140 172356
rect 248564 172304 248616 172356
rect 263836 172304 263888 172356
rect 245804 172236 245856 172288
rect 256936 172236 256988 172288
rect 249024 172168 249076 172220
rect 247644 171896 247696 171948
rect 248472 171896 248524 171948
rect 338540 171896 338592 171948
rect 347280 171896 347332 171948
rect 251876 171760 251928 171812
rect 258960 171760 259012 171812
rect 46716 171624 46768 171676
rect 46900 171624 46952 171676
rect 72660 171624 72712 171676
rect 369728 170264 369780 170316
rect 369912 170264 369964 170316
rect 79192 170196 79244 170248
rect 123996 170196 124048 170248
rect 312044 170196 312096 170248
rect 328420 170196 328472 170248
rect 123996 169516 124048 169568
rect 140280 169516 140332 169568
rect 267240 169516 267292 169568
rect 312044 169516 312096 169568
rect 73488 169423 73540 169432
rect 73488 169389 73497 169423
rect 73497 169389 73531 169423
rect 73531 169389 73540 169423
rect 73488 169380 73540 169389
rect 132184 168904 132236 168956
rect 140556 168904 140608 168956
rect 226024 168904 226076 168956
rect 233476 168904 233528 168956
rect 46992 168836 47044 168888
rect 49200 168836 49252 168888
rect 222160 168564 222212 168616
rect 369268 168564 369320 168616
rect 128136 168496 128188 168548
rect 369176 168496 369228 168548
rect 361172 168156 361224 168208
rect 423640 168156 423692 168208
rect 77260 167544 77312 167596
rect 87196 167544 87248 167596
rect 132276 167544 132328 167596
rect 140556 167544 140608 167596
rect 225932 167544 225984 167596
rect 233476 167544 233528 167596
rect 110196 166796 110248 166848
rect 112680 166796 112732 166848
rect 203852 166796 203904 166848
rect 206520 166796 206572 166848
rect 217192 166796 217244 166848
rect 225196 166796 225248 166848
rect 297876 166796 297928 166848
rect 300360 166796 300412 166848
rect 311216 166796 311268 166848
rect 319220 166796 319272 166848
rect 123536 166524 123588 166576
rect 129240 166524 129292 166576
rect 284536 166252 284588 166304
rect 285824 166252 285876 166304
rect 77260 166184 77312 166236
rect 87104 166184 87156 166236
rect 132092 166184 132144 166236
rect 140556 166184 140608 166236
rect 225840 166184 225892 166236
rect 233476 166184 233528 166236
rect 361724 165436 361776 165488
rect 420880 165436 420932 165488
rect 77260 164756 77312 164808
rect 87288 164756 87340 164808
rect 132644 164756 132696 164808
rect 139636 164756 139688 164808
rect 225656 164756 225708 164808
rect 233476 164756 233528 164808
rect 131356 163464 131408 163516
rect 137612 163464 137664 163516
rect 226300 163464 226352 163516
rect 231452 163464 231504 163516
rect 321612 163464 321664 163516
rect 327224 163464 327276 163516
rect 77260 163396 77312 163448
rect 87196 163396 87248 163448
rect 131908 163396 131960 163448
rect 139636 163396 139688 163448
rect 226392 163396 226444 163448
rect 233476 163396 233528 163448
rect 272852 163396 272904 163448
rect 274876 163396 274928 163448
rect 361724 162648 361776 162700
rect 418212 162648 418264 162700
rect 321612 162376 321664 162428
rect 327500 162376 327552 162428
rect 132000 162104 132052 162156
rect 139544 162104 139596 162156
rect 226392 162104 226444 162156
rect 233476 162104 233528 162156
rect 132368 162036 132420 162088
rect 139636 162036 139688 162088
rect 226208 162036 226260 162088
rect 234580 162036 234632 162088
rect 132000 161968 132052 162020
rect 132276 161968 132328 162020
rect 222436 161560 222488 161612
rect 321060 161560 321112 161612
rect 327224 161560 327276 161612
rect 173308 161492 173360 161544
rect 321612 161424 321664 161476
rect 328420 161424 328472 161476
rect 272944 161084 272996 161136
rect 275152 161084 275204 161136
rect 131356 160676 131408 160728
rect 140464 160676 140516 160728
rect 131448 160608 131500 160660
rect 140832 160608 140884 160660
rect 174044 160608 174096 160660
rect 176252 160608 176304 160660
rect 179012 160608 179064 160660
rect 182324 160608 182376 160660
rect 226300 160608 226352 160660
rect 234304 160608 234356 160660
rect 266596 160608 266648 160660
rect 270000 160608 270052 160660
rect 77260 160540 77312 160592
rect 87196 160540 87248 160592
rect 131356 159316 131408 159368
rect 140556 159316 140608 159368
rect 173676 159316 173728 159368
rect 181496 159316 181548 159368
rect 266596 159316 266648 159368
rect 275704 159316 275756 159368
rect 320600 159316 320652 159368
rect 327316 159316 327368 159368
rect 79284 159248 79336 159300
rect 131816 159248 131868 159300
rect 139636 159248 139688 159300
rect 172756 159248 172808 159300
rect 181680 159248 181732 159300
rect 226116 159248 226168 159300
rect 228692 159248 228744 159300
rect 231360 159248 231412 159300
rect 233476 159248 233528 159300
rect 272760 159248 272812 159300
rect 275152 159248 275204 159300
rect 87288 159112 87340 159164
rect 131908 159112 131960 159164
rect 132092 159112 132144 159164
rect 81768 159044 81820 159096
rect 87196 159044 87248 159096
rect 361724 158500 361776 158552
rect 415544 158500 415596 158552
rect 321612 158160 321664 158212
rect 327224 158160 327276 158212
rect 173676 158024 173728 158076
rect 181864 158024 181916 158076
rect 178920 157956 178972 158008
rect 181404 157956 181456 158008
rect 266596 157956 266648 158008
rect 271380 157956 271432 158008
rect 321060 157956 321112 158008
rect 327408 157956 327460 158008
rect 79744 157888 79796 157940
rect 132184 157888 132236 157940
rect 138900 157888 138952 157940
rect 173492 157888 173544 157940
rect 182324 157888 182376 157940
rect 266964 157888 267016 157940
rect 274876 157888 274928 157940
rect 87196 157752 87248 157804
rect 222804 157140 222856 157192
rect 233476 157140 233528 157192
rect 321612 157140 321664 157192
rect 327224 157140 327276 157192
rect 77260 156460 77312 156512
rect 173124 156460 173176 156512
rect 173308 156460 173360 156512
rect 173676 156460 173728 156512
rect 182324 156460 182376 156512
rect 369820 156503 369872 156512
rect 369820 156469 369829 156503
rect 369829 156469 369863 156503
rect 369863 156469 369872 156503
rect 369820 156460 369872 156469
rect 87196 156392 87248 156444
rect 173584 156392 173636 156444
rect 182140 156392 182192 156444
rect 267424 156392 267476 156444
rect 274876 156392 274928 156444
rect 267056 155780 267108 155832
rect 267700 155780 267752 155832
rect 361724 155712 361776 155764
rect 412876 155712 412928 155764
rect 321060 155372 321112 155424
rect 327224 155372 327276 155424
rect 173860 155100 173912 155152
rect 182324 155100 182376 155152
rect 267792 155100 267844 155152
rect 274968 155100 275020 155152
rect 321612 155100 321664 155152
rect 79744 155032 79796 155084
rect 87196 155032 87248 155084
rect 137612 155032 137664 155084
rect 139636 155032 139688 155084
rect 173400 155032 173452 155084
rect 173584 155032 173636 155084
rect 181772 155032 181824 155084
rect 231452 155032 231504 155084
rect 233476 155032 233528 155084
rect 266688 155032 266740 155084
rect 275060 155032 275112 155084
rect 328420 155032 328472 155084
rect 182324 154964 182376 155016
rect 267608 154964 267660 155016
rect 274876 154964 274928 155016
rect 173400 154896 173452 154948
rect 181312 154896 181364 154948
rect 266596 154896 266648 154948
rect 272852 154896 272904 154948
rect 12676 154760 12728 154812
rect 16264 154760 16316 154812
rect 81768 154352 81820 154404
rect 87196 154352 87248 154404
rect 320876 153740 320928 153792
rect 328420 153740 328472 153792
rect 172940 153672 172992 153724
rect 181404 153672 181456 153724
rect 267148 153672 267200 153724
rect 274968 153672 275020 153724
rect 369820 153715 369872 153724
rect 369820 153681 369829 153715
rect 369829 153681 369863 153715
rect 369863 153681 369872 153715
rect 369820 153672 369872 153681
rect 173216 153604 173268 153656
rect 182324 153604 182376 153656
rect 267516 153604 267568 153656
rect 274876 153604 274928 153656
rect 266596 153536 266648 153588
rect 272944 153536 272996 153588
rect 81768 152992 81820 153044
rect 87196 152992 87248 153044
rect 321612 152448 321664 152500
rect 328236 152448 328288 152500
rect 79744 152380 79796 152432
rect 87196 152380 87248 152432
rect 173584 152380 173636 152432
rect 180300 152380 180352 152432
rect 320508 152380 320560 152432
rect 323176 152380 323228 152432
rect 173308 152312 173360 152364
rect 182324 152312 182376 152364
rect 267884 152312 267936 152364
rect 274876 152312 274928 152364
rect 173676 151675 173728 151684
rect 173676 151641 173685 151675
rect 173685 151641 173719 151675
rect 173719 151641 173728 151675
rect 173676 151632 173728 151641
rect 320784 151360 320836 151412
rect 323268 151360 323320 151412
rect 131356 150884 131408 150936
rect 140648 150884 140700 150936
rect 173768 150884 173820 150936
rect 182324 150884 182376 150936
rect 225748 150884 225800 150936
rect 233476 150884 233528 150936
rect 266596 150884 266648 150936
rect 275796 150884 275848 150936
rect 323176 150884 323228 150936
rect 328420 150884 328472 150936
rect 176252 150816 176304 150868
rect 182232 150816 182284 150868
rect 225564 150816 225616 150868
rect 232740 150816 232792 150868
rect 267700 150816 267752 150868
rect 274876 150816 274928 150868
rect 173584 150748 173636 150800
rect 179012 150748 179064 150800
rect 270000 150748 270052 150800
rect 274968 150748 275020 150800
rect 173952 150612 174004 150664
rect 80112 149592 80164 149644
rect 87196 149592 87248 149644
rect 321612 149592 321664 149644
rect 327224 149592 327276 149644
rect 81768 149524 81820 149576
rect 88116 149524 88168 149576
rect 131356 149524 131408 149576
rect 140740 149524 140792 149576
rect 225932 149524 225984 149576
rect 234120 149524 234172 149576
rect 266596 149524 266648 149576
rect 272760 149524 272812 149576
rect 323268 149524 323320 149576
rect 328420 149524 328472 149576
rect 271380 149456 271432 149508
rect 274876 149456 274928 149508
rect 228692 149388 228744 149440
rect 233476 149388 233528 149440
rect 226300 149116 226352 149168
rect 231360 149116 231412 149168
rect 321612 148368 321664 148420
rect 328328 148368 328380 148420
rect 321060 148232 321112 148284
rect 328512 148232 328564 148284
rect 173584 148164 173636 148216
rect 178920 148164 178972 148216
rect 227220 148164 227272 148216
rect 233476 148164 233528 148216
rect 321796 148164 321848 148216
rect 328420 148164 328472 148216
rect 427320 148164 427372 148216
rect 429436 148164 429488 148216
rect 79744 148096 79796 148148
rect 87104 148096 87156 148148
rect 369820 146804 369872 146856
rect 132552 146736 132604 146788
rect 139636 146736 139688 146788
rect 226392 146736 226444 146788
rect 233476 146736 233528 146788
rect 267884 146736 267936 146788
rect 275520 146736 275572 146788
rect 369820 146668 369872 146720
rect 79744 145376 79796 145428
rect 87196 145376 87248 145428
rect 91704 145376 91756 145428
rect 128136 145376 128188 145428
rect 132276 145376 132328 145428
rect 139636 145376 139688 145428
rect 185636 145376 185688 145428
rect 222160 145376 222212 145428
rect 226116 145376 226168 145428
rect 233476 145376 233528 145428
rect 266780 145376 266832 145428
rect 275612 145376 275664 145428
rect 279660 145376 279712 145428
rect 322900 145376 322952 145428
rect 116084 144832 116136 144884
rect 128044 144832 128096 144884
rect 211028 144832 211080 144884
rect 230992 144832 231044 144884
rect 103664 144764 103716 144816
rect 124272 144764 124324 144816
rect 197504 144764 197556 144816
rect 218296 144764 218348 144816
rect 292724 144764 292776 144816
rect 312320 144764 312372 144816
rect 91244 144696 91296 144748
rect 120684 144696 120736 144748
rect 185084 144696 185136 144748
rect 214708 144696 214760 144748
rect 280304 144696 280356 144748
rect 308732 144696 308784 144748
rect 216180 144356 216232 144408
rect 221976 144356 222028 144408
rect 310020 144152 310072 144204
rect 316000 144152 316052 144204
rect 79744 144016 79796 144068
rect 87288 144016 87340 144068
rect 132368 144016 132420 144068
rect 139636 144016 139688 144068
rect 226484 144016 226536 144068
rect 233476 144016 233528 144068
rect 303856 143404 303908 143456
rect 305052 143404 305104 143456
rect 324648 143404 324700 143456
rect 297784 143336 297836 143388
rect 325384 143336 325436 143388
rect 200172 142792 200224 142844
rect 167788 142180 167840 142232
rect 231360 142044 231412 142096
rect 290976 142044 291028 142096
rect 325936 142044 325988 142096
rect 127216 141976 127268 142028
rect 140372 141976 140424 142028
rect 173584 141976 173636 142028
rect 219676 141976 219728 142028
rect 233476 141976 233528 142028
rect 267332 141976 267384 142028
rect 316276 141976 316328 142028
rect 360436 141976 360488 142028
rect 361080 141976 361132 142028
rect 77260 141296 77312 141348
rect 127216 141296 127268 141348
rect 136968 141296 137020 141348
rect 150400 141296 150452 141348
rect 167788 141296 167840 141348
rect 316276 141296 316328 141348
rect 328420 141296 328472 141348
rect 77720 141228 77772 141280
rect 113416 141228 113468 141280
rect 114704 141228 114756 141280
rect 82320 140752 82372 140804
rect 114704 140616 114756 140668
rect 137612 140616 137664 140668
rect 102284 140548 102336 140600
rect 102376 140548 102428 140600
rect 137336 140548 137388 140600
rect 207900 140548 207952 140600
rect 231268 140548 231320 140600
rect 302016 140548 302068 140600
rect 324832 140548 324884 140600
rect 141844 139868 141896 139920
rect 152608 139868 152660 139920
rect 166132 139868 166184 139920
rect 260156 139868 260208 139920
rect 64840 139732 64892 139784
rect 70452 139800 70504 139852
rect 150492 139800 150544 139852
rect 162268 139800 162320 139852
rect 239548 139800 239600 139852
rect 322808 139800 322860 139852
rect 62264 139664 62316 139716
rect 74224 139732 74276 139784
rect 151780 139732 151832 139784
rect 164568 139732 164620 139784
rect 247092 139732 247144 139784
rect 259236 139732 259288 139784
rect 59504 139596 59556 139648
rect 57664 139528 57716 139580
rect 60240 139528 60292 139580
rect 60884 139596 60936 139648
rect 73120 139664 73172 139716
rect 154724 139664 154776 139716
rect 167328 139664 167380 139716
rect 244332 139664 244384 139716
rect 256292 139664 256344 139716
rect 65944 139596 65996 139648
rect 70544 139596 70596 139648
rect 153344 139596 153396 139648
rect 71096 139528 71148 139580
rect 150584 139528 150636 139580
rect 163280 139596 163332 139648
rect 242492 139596 242544 139648
rect 249116 139596 249168 139648
rect 251324 139596 251376 139648
rect 264112 139596 264164 139648
rect 158128 139528 158180 139580
rect 158864 139528 158916 139580
rect 160980 139528 161032 139580
rect 161624 139528 161676 139580
rect 161992 139528 162044 139580
rect 163004 139528 163056 139580
rect 249852 139528 249904 139580
rect 253072 139528 253124 139580
rect 63644 139460 63696 139512
rect 75236 139460 75288 139512
rect 151872 139460 151924 139512
rect 58124 139392 58176 139444
rect 70084 139392 70136 139444
rect 155184 139392 155236 139444
rect 156012 139392 156064 139444
rect 157392 139460 157444 139512
rect 169996 139460 170048 139512
rect 249208 139460 249260 139512
rect 252060 139460 252112 139512
rect 165212 139392 165264 139444
rect 248564 139392 248616 139444
rect 255004 139528 255056 139580
rect 257488 139528 257540 139580
rect 333388 139528 333440 139580
rect 334124 139528 334176 139580
rect 334400 139528 334452 139580
rect 335504 139528 335556 139580
rect 256016 139460 256068 139512
rect 258684 139460 258736 139512
rect 258316 139392 258368 139444
rect 56744 139324 56796 139376
rect 67968 139324 68020 139376
rect 154632 139324 154684 139376
rect 168064 139324 168116 139376
rect 244424 139324 244476 139376
rect 257304 139324 257356 139376
rect 55364 139256 55416 139308
rect 66956 139256 67008 139308
rect 155920 139256 155972 139308
rect 169076 139256 169128 139308
rect 241480 139256 241532 139308
rect 249668 139256 249720 139308
rect 249852 139256 249904 139308
rect 261168 139256 261220 139308
rect 338540 139256 338592 139308
rect 339552 139256 339604 139308
rect 60792 139188 60844 139240
rect 72108 139188 72160 139240
rect 74316 139188 74368 139240
rect 116176 139188 116228 139240
rect 136876 139188 136928 139240
rect 144604 139188 144656 139240
rect 170640 139188 170692 139240
rect 238628 139188 238680 139240
rect 264480 139188 264532 139240
rect 63828 139120 63880 139172
rect 68612 139120 68664 139172
rect 249944 139120 249996 139172
rect 252152 139052 252204 139104
rect 254176 139052 254228 139104
rect 263100 139120 263152 139172
rect 262088 139052 262140 139104
rect 251140 138984 251192 139036
rect 253992 138984 254044 139036
rect 247184 138916 247236 138968
rect 62816 138848 62868 138900
rect 59688 138780 59740 138832
rect 63000 138780 63052 138832
rect 245804 138848 245856 138900
rect 340932 138848 340984 138900
rect 67692 138780 67744 138832
rect 253900 138780 253952 138832
rect 256660 138780 256712 138832
rect 341024 138780 341076 138832
rect 345900 138848 345952 138900
rect 349948 138848 350000 138900
rect 347924 138780 347976 138832
rect 61804 138712 61856 138764
rect 65760 138712 65812 138764
rect 145248 138712 145300 138764
rect 365220 138712 365272 138764
rect 58676 138644 58728 138696
rect 63092 138644 63144 138696
rect 338080 138644 338132 138696
rect 341668 138644 341720 138696
rect 346820 138644 346872 138696
rect 60700 138576 60752 138628
rect 63184 138576 63236 138628
rect 252704 138576 252756 138628
rect 254820 138576 254872 138628
rect 338264 138576 338316 138628
rect 342680 138576 342732 138628
rect 344520 138576 344572 138628
rect 345808 138576 345860 138628
rect 345992 138576 346044 138628
rect 348936 138576 348988 138628
rect 287204 137828 287256 137880
rect 324740 137828 324792 137880
rect 343968 137828 344020 137880
rect 360896 137828 360948 137880
rect 325936 137148 325988 137200
rect 326580 137148 326632 137200
rect 343968 137148 344020 137200
rect 74132 137080 74184 137132
rect 74408 137080 74460 137132
rect 427504 137080 427556 137132
rect 429436 137080 429488 137132
rect 210016 136400 210068 136452
rect 216180 136400 216232 136452
rect 304040 136400 304092 136452
rect 310020 136400 310072 136452
rect 291528 136264 291580 136316
rect 292724 136264 292776 136316
rect 279108 136128 279160 136180
rect 280304 136128 280356 136180
rect 346544 135040 346596 135092
rect 360620 135040 360672 135092
rect 325384 134428 325436 134480
rect 345716 134428 345768 134480
rect 346544 134428 346596 134480
rect 51592 134360 51644 134412
rect 51868 134360 51920 134412
rect 236236 134403 236288 134412
rect 236236 134369 236245 134403
rect 236245 134369 236279 134403
rect 236279 134369 236288 134403
rect 236236 134360 236288 134369
rect 360712 134360 360764 134412
rect 346544 133748 346596 133800
rect 360528 133748 360580 133800
rect 283156 133680 283208 133732
rect 324556 133680 324608 133732
rect 343324 133680 343376 133732
rect 360988 133680 361040 133732
rect 324556 133068 324608 133120
rect 343324 133068 343376 133120
rect 324832 133000 324884 133052
rect 325476 133000 325528 133052
rect 346360 133000 346412 133052
rect 346544 133000 346596 133052
rect 13044 132932 13096 132984
rect 16448 132932 16500 132984
rect 369636 132975 369688 132984
rect 369636 132941 369645 132975
rect 369645 132941 369679 132975
rect 369679 132941 369688 132975
rect 369636 132932 369688 132941
rect 369544 132907 369596 132916
rect 369544 132873 369553 132907
rect 369553 132873 369587 132907
rect 369587 132873 369596 132907
rect 369544 132864 369596 132873
rect 230992 132796 231044 132848
rect 231452 132796 231504 132848
rect 136876 132320 136928 132372
rect 137336 132320 137388 132372
rect 343968 132320 344020 132372
rect 360804 132320 360856 132372
rect 324648 132252 324700 132304
rect 347004 132252 347056 132304
rect 354916 132252 354968 132304
rect 355836 132252 355888 132304
rect 339460 131708 339512 131760
rect 339736 131708 339788 131760
rect 324740 131640 324792 131692
rect 325568 131640 325620 131692
rect 343968 131640 344020 131692
rect 347004 131640 347056 131692
rect 360436 131640 360488 131692
rect 361080 131640 361132 131692
rect 59688 131572 59740 131624
rect 60792 131572 60844 131624
rect 245344 131572 245396 131624
rect 245804 131572 245856 131624
rect 248012 131572 248064 131624
rect 248564 131572 248616 131624
rect 250680 131572 250732 131624
rect 251324 131572 251376 131624
rect 63184 131504 63236 131556
rect 65944 131504 65996 131556
rect 339552 131504 339604 131556
rect 350960 131504 351012 131556
rect 338172 131436 338224 131488
rect 350408 131436 350460 131488
rect 161624 131368 161676 131420
rect 163464 131368 163516 131420
rect 248472 131368 248524 131420
rect 250956 131368 251008 131420
rect 342404 131368 342456 131420
rect 345900 131368 345952 131420
rect 158772 131300 158824 131352
rect 161716 131300 161768 131352
rect 231360 131300 231412 131352
rect 322716 131300 322768 131352
rect 335504 131300 335556 131352
rect 348568 131300 348620 131352
rect 258960 131232 259012 131284
rect 368808 131232 368860 131284
rect 336884 131164 336936 131216
rect 349764 131164 349816 131216
rect 334124 131096 334176 131148
rect 348016 131096 348068 131148
rect 332744 131028 332796 131080
rect 340840 131028 340892 131080
rect 352248 131028 352300 131080
rect 335412 130960 335464 131012
rect 349396 130960 349448 131012
rect 57020 130892 57072 130944
rect 68060 130892 68112 130944
rect 361172 130892 361224 130944
rect 347280 130824 347332 130876
rect 160244 130688 160296 130740
rect 162636 130688 162688 130740
rect 246264 130552 246316 130604
rect 247092 130552 247144 130604
rect 60240 130484 60292 130536
rect 63276 130484 63328 130536
rect 156104 130484 156156 130536
rect 159048 130484 159100 130536
rect 63000 130416 63052 130468
rect 65024 130416 65076 130468
rect 156012 130416 156064 130468
rect 158128 130416 158180 130468
rect 62356 130348 62408 130400
rect 63644 130348 63696 130400
rect 154540 130348 154592 130400
rect 157300 130348 157352 130400
rect 157484 130348 157536 130400
rect 159968 130348 160020 130400
rect 325292 130348 325344 130400
rect 342496 130756 342548 130808
rect 339644 130688 339696 130740
rect 351604 130688 351656 130740
rect 341760 130620 341812 130672
rect 345992 130620 346044 130672
rect 339552 130552 339604 130604
rect 344520 130552 344572 130604
rect 339368 130484 339420 130536
rect 343876 130484 343928 130536
rect 338724 130416 338776 130468
rect 342772 130416 342824 130468
rect 61436 130280 61488 130332
rect 62264 130280 62316 130332
rect 63092 130280 63144 130332
rect 64104 130280 64156 130332
rect 65760 130280 65812 130332
rect 66772 130280 66824 130332
rect 149296 130280 149348 130332
rect 150492 130280 150544 130332
rect 151044 130280 151096 130332
rect 151780 130280 151832 130332
rect 153712 130280 153764 130332
rect 154724 130280 154776 130332
rect 156380 130280 156432 130332
rect 157392 130280 157444 130332
rect 158864 130280 158916 130332
rect 160796 130280 160848 130332
rect 163004 130280 163056 130332
rect 164384 130280 164436 130332
rect 243596 130280 243648 130332
rect 244332 130280 244384 130332
rect 248932 130280 248984 130332
rect 249944 130280 249996 130332
rect 254820 130280 254872 130332
rect 255556 130280 255608 130332
rect 323176 130280 323228 130332
rect 231268 130212 231320 130264
rect 246448 130212 246500 130264
rect 337528 130280 337580 130332
rect 338080 130280 338132 130332
rect 340564 130280 340616 130332
rect 341024 130280 341076 130332
rect 344888 130212 344940 130264
rect 73856 127492 73908 127544
rect 74224 127492 74276 127544
rect 74408 127492 74460 127544
rect 137060 127492 137112 127544
rect 137244 127492 137296 127544
rect 74040 127356 74092 127408
rect 38804 126744 38856 126796
rect 54076 126744 54128 126796
rect 357676 126744 357728 126796
rect 405976 126744 406028 126796
rect 38252 126064 38304 126116
rect 51224 126064 51276 126116
rect 356204 126064 356256 126116
rect 405976 126064 406028 126116
rect 76892 125452 76944 125504
rect 81676 125452 81728 125504
rect 169996 125384 170048 125436
rect 170640 125384 170692 125436
rect 175516 125384 175568 125436
rect 263836 125248 263888 125300
rect 264480 125248 264532 125300
rect 270368 125248 270420 125300
rect 76156 125044 76208 125096
rect 76892 125044 76944 125096
rect 369544 124883 369596 124892
rect 369544 124849 369553 124883
rect 369553 124849 369587 124883
rect 369587 124849 369596 124883
rect 369544 124840 369596 124849
rect 236236 124815 236288 124824
rect 236236 124781 236245 124815
rect 236245 124781 236279 124815
rect 236279 124781 236288 124815
rect 236236 124772 236288 124781
rect 360620 124772 360672 124824
rect 74040 124747 74092 124756
rect 74040 124713 74049 124747
rect 74049 124713 74083 124747
rect 74083 124713 74092 124747
rect 74040 124704 74092 124713
rect 369636 124679 369688 124688
rect 369636 124645 369645 124679
rect 369645 124645 369679 124679
rect 369679 124645 369688 124679
rect 369636 124636 369688 124645
rect 38804 122596 38856 122648
rect 53156 122596 53208 122648
rect 356296 122596 356348 122648
rect 405976 122596 406028 122648
rect 137612 121984 137664 122036
rect 144236 121984 144288 122036
rect 231452 121984 231504 122036
rect 240376 121984 240428 122036
rect 325384 121984 325436 122036
rect 334216 121984 334268 122036
rect 13228 121916 13280 121968
rect 16540 121916 16592 121968
rect 38804 120556 38856 120608
rect 52604 120556 52656 120608
rect 356204 120556 356256 120608
rect 405976 120556 406028 120608
rect 324556 119876 324608 119928
rect 326580 119876 326632 119928
rect 261168 117904 261220 117956
rect 268620 117904 268672 117956
rect 167880 117836 167932 117888
rect 174872 117836 174924 117888
rect 360344 117836 360396 117888
rect 360436 117836 360488 117888
rect 360620 117836 360672 117888
rect 73488 117768 73540 117820
rect 74224 117768 74276 117820
rect 360252 117768 360304 117820
rect 74040 117743 74092 117752
rect 74040 117709 74049 117743
rect 74049 117709 74083 117743
rect 74083 117709 74092 117743
rect 74040 117700 74092 117709
rect 38252 117088 38304 117140
rect 54076 117088 54128 117140
rect 354916 117088 354968 117140
rect 405976 117088 406028 117140
rect 38804 115048 38856 115100
rect 51224 115048 51276 115100
rect 51868 115048 51920 115100
rect 74040 115048 74092 115100
rect 74224 115048 74276 115100
rect 236236 115091 236288 115100
rect 236236 115057 236245 115091
rect 236245 115057 236279 115091
rect 236279 115057 236288 115091
rect 236236 115048 236288 115057
rect 356204 115048 356256 115100
rect 405976 115048 406028 115100
rect 38804 112940 38856 112992
rect 52144 112940 52196 112992
rect 136876 112940 136928 112992
rect 147364 112940 147416 112992
rect 355008 112940 355060 112992
rect 405976 112940 406028 112992
rect 427412 112056 427464 112108
rect 429436 112056 429488 112108
rect 12860 111512 12912 111564
rect 16356 111512 16408 111564
rect 38252 110900 38304 110952
rect 52604 110900 52656 110952
rect 136876 110900 136928 110952
rect 145340 110900 145392 110952
rect 231636 110900 231688 110952
rect 239088 110900 239140 110952
rect 240100 110900 240152 110952
rect 356204 110900 356256 110952
rect 406068 110900 406120 110952
rect 74408 109472 74460 109524
rect 81676 109472 81728 109524
rect 137704 108180 137756 108232
rect 143960 108180 144012 108232
rect 231544 108180 231596 108232
rect 240376 108180 240428 108232
rect 325476 108180 325528 108232
rect 334216 108180 334268 108232
rect 51684 108019 51736 108028
rect 51684 107985 51693 108019
rect 51693 107985 51727 108019
rect 51727 107985 51736 108019
rect 51684 107976 51736 107985
rect 38804 107432 38856 107484
rect 51684 107432 51736 107484
rect 353536 107432 353588 107484
rect 405976 107432 406028 107484
rect 13320 105460 13372 105512
rect 18104 105460 18156 105512
rect 236236 105503 236288 105512
rect 236236 105469 236245 105503
rect 236245 105469 236279 105503
rect 236279 105469 236288 105503
rect 236236 105460 236288 105469
rect 427688 105460 427740 105512
rect 430080 105460 430132 105512
rect 38804 105392 38856 105444
rect 52604 105392 52656 105444
rect 356204 105392 356256 105444
rect 405976 105392 406028 105444
rect 352708 101924 352760 101976
rect 405976 101924 406028 101976
rect 50028 101516 50080 101568
rect 51316 101516 51368 101568
rect 38620 101312 38672 101364
rect 50028 101312 50080 101364
rect 12860 100768 12912 100820
rect 16172 100768 16224 100820
rect 38804 100564 38856 100616
rect 52604 100564 52656 100616
rect 356204 100564 356256 100616
rect 405976 100564 406028 100616
rect 13412 99884 13464 99936
rect 17460 99884 17512 99936
rect 168248 98592 168300 98644
rect 169260 98592 169312 98644
rect 427688 98524 427740 98576
rect 429436 98524 429488 98576
rect 73948 98388 74000 98440
rect 74224 98388 74276 98440
rect 38804 97776 38856 97828
rect 49936 97776 49988 97828
rect 352800 97776 352852 97828
rect 405976 97776 406028 97828
rect 13504 95804 13556 95856
rect 18104 95804 18156 95856
rect 427228 95804 427280 95856
rect 430172 95804 430224 95856
rect 38068 95736 38120 95788
rect 52604 95736 52656 95788
rect 236236 95779 236288 95788
rect 236236 95745 236245 95779
rect 236245 95745 236279 95779
rect 236279 95745 236288 95779
rect 236236 95736 236288 95745
rect 237248 95736 237300 95788
rect 356204 95736 356256 95788
rect 405976 95736 406028 95788
rect 231820 94988 231872 95040
rect 325844 94648 325896 94700
rect 330076 94648 330128 94700
rect 138164 94376 138216 94428
rect 142396 94376 142448 94428
rect 232740 94376 232792 94428
rect 240376 94376 240428 94428
rect 326672 94376 326724 94428
rect 334216 94376 334268 94428
rect 72568 94308 72620 94360
rect 73948 94308 74000 94360
rect 74684 94308 74736 94360
rect 78180 94308 78232 94360
rect 73580 93832 73632 93884
rect 73764 93832 73816 93884
rect 73396 93696 73448 93748
rect 73580 93696 73632 93748
rect 74132 92948 74184 93000
rect 81676 92948 81728 93000
rect 169260 92948 169312 93000
rect 175516 92948 175568 93000
rect 263100 92948 263152 93000
rect 270368 92948 270420 93000
rect 37608 92268 37660 92320
rect 48556 92268 48608 92320
rect 352800 92268 352852 92320
rect 405976 92268 406028 92320
rect 73856 91248 73908 91300
rect 76800 91248 76852 91300
rect 13228 90160 13280 90212
rect 17276 90228 17328 90280
rect 38804 90160 38856 90212
rect 52604 90228 52656 90280
rect 356204 90160 356256 90212
rect 405976 90160 406028 90212
rect 369728 88800 369780 88852
rect 369912 88800 369964 88852
rect 251324 87508 251376 87560
rect 260064 87508 260116 87560
rect 23900 87440 23952 87492
rect 72568 87440 72620 87492
rect 154724 87440 154776 87492
rect 172020 87440 172072 87492
rect 326580 87440 326632 87492
rect 327224 87440 327276 87492
rect 412876 87440 412928 87492
rect 26568 87372 26620 87424
rect 73672 87372 73724 87424
rect 243412 87372 243464 87424
rect 250772 87372 250824 87424
rect 359700 87372 359752 87424
rect 360160 87372 360212 87424
rect 423548 87372 423600 87424
rect 29236 87304 29288 87356
rect 73764 87304 73816 87356
rect 149204 87304 149256 87356
rect 156932 87304 156984 87356
rect 249024 87304 249076 87356
rect 258960 87304 259012 87356
rect 344980 87304 345032 87356
rect 363840 87304 363892 87356
rect 370004 87304 370056 87356
rect 410208 87304 410260 87356
rect 31904 87236 31956 87288
rect 73488 87236 73540 87288
rect 149756 87236 149808 87288
rect 158956 87236 159008 87288
rect 341024 87236 341076 87288
rect 352156 87236 352208 87288
rect 34572 87168 34624 87220
rect 73580 87168 73632 87220
rect 151044 87168 151096 87220
rect 161716 87168 161768 87220
rect 243964 87168 244016 87220
rect 252980 87168 253032 87220
rect 344336 87168 344388 87220
rect 347280 87168 347332 87220
rect 21232 87100 21284 87152
rect 34664 87100 34716 87152
rect 64380 87100 64432 87152
rect 65944 87100 65996 87152
rect 150400 87100 150452 87152
rect 159600 87100 159652 87152
rect 243044 87100 243096 87152
rect 255096 87100 255148 87152
rect 338080 87100 338132 87152
rect 349580 87100 349632 87152
rect 150584 87032 150636 87084
rect 162084 87032 162136 87084
rect 244424 87032 244476 87084
rect 253532 87032 253584 87084
rect 334124 87032 334176 87084
rect 346176 87032 346228 87084
rect 149204 86964 149256 87016
rect 161440 86964 161492 87016
rect 241664 86964 241716 87016
rect 254544 86964 254596 87016
rect 339644 86964 339696 87016
rect 56100 86896 56152 86948
rect 65852 86896 65904 86948
rect 146444 86896 146496 86948
rect 160244 86896 160296 86948
rect 245344 86896 245396 86948
rect 255556 86896 255608 86948
rect 335412 86896 335464 86948
rect 348752 86964 348804 87016
rect 351236 86896 351288 86948
rect 59688 86828 59740 86880
rect 70728 86828 70780 86880
rect 147824 86828 147876 86880
rect 160888 86828 160940 86880
rect 160980 86828 161032 86880
rect 162728 86828 162780 86880
rect 240284 86828 240336 86880
rect 254268 86828 254320 86880
rect 335504 86828 335556 86880
rect 348016 86828 348068 86880
rect 57020 86760 57072 86812
rect 67876 86760 67928 86812
rect 145064 86760 145116 86812
rect 159324 86760 159376 86812
rect 238904 86760 238956 86812
rect 253256 86760 253308 86812
rect 332744 86760 332796 86812
rect 345440 86760 345492 86812
rect 153436 86692 153488 86744
rect 154632 86692 154684 86744
rect 347004 86692 347056 86744
rect 336884 86624 336936 86676
rect 257580 86488 257632 86540
rect 258408 86488 258460 86540
rect 156840 86284 156892 86336
rect 163280 86284 163332 86336
rect 152240 86216 152292 86268
rect 153344 86216 153396 86268
rect 250680 86216 250732 86268
rect 256384 86216 256436 86268
rect 341668 86216 341720 86268
rect 344612 86216 344664 86268
rect 61620 86148 61672 86200
rect 63276 86148 63328 86200
rect 67140 86148 67192 86200
rect 68612 86148 68664 86200
rect 253440 86148 253492 86200
rect 257672 86148 257724 86200
rect 337620 86148 337672 86200
rect 339092 86148 339144 86200
rect 340104 86148 340156 86200
rect 341760 86148 341812 86200
rect 342404 86148 342456 86200
rect 344704 86148 344756 86200
rect 61436 86080 61488 86132
rect 62264 86080 62316 86132
rect 62356 86080 62408 86132
rect 63644 86080 63696 86132
rect 65760 86080 65812 86132
rect 66772 86080 66824 86132
rect 68520 86080 68572 86132
rect 69440 86080 69492 86132
rect 246540 86080 246592 86132
rect 247092 86080 247144 86132
rect 247736 86080 247788 86132
rect 248564 86080 248616 86132
rect 254820 86080 254872 86132
rect 255740 86080 255792 86132
rect 256200 86080 256252 86132
rect 256936 86080 256988 86132
rect 338264 86080 338316 86132
rect 339000 86080 339052 86132
rect 340932 86080 340984 86132
rect 341852 86080 341904 86132
rect 343508 86080 343560 86132
rect 344520 86080 344572 86132
rect 66680 86012 66732 86064
rect 67324 86012 67376 86064
rect 230992 85876 231044 85928
rect 232740 85876 232792 85928
rect 324556 85740 324608 85792
rect 326672 85740 326724 85792
rect 138164 85468 138216 85520
rect 144420 85468 144472 85520
rect 354916 84040 354968 84092
rect 355836 84040 355888 84092
rect 88484 81932 88536 81984
rect 182416 81932 182468 81984
rect 276256 81932 276308 81984
rect 95752 81864 95804 81916
rect 176160 81864 176212 81916
rect 189500 81864 189552 81916
rect 283432 81864 283484 81916
rect 102928 81796 102980 81848
rect 174780 81796 174832 81848
rect 196676 81796 196728 81848
rect 290332 81796 290384 81848
rect 285824 81320 285876 81372
rect 297508 81320 297560 81372
rect 369912 81363 369964 81372
rect 369912 81329 369921 81363
rect 369921 81329 369955 81363
rect 369955 81329 369964 81363
rect 369912 81320 369964 81329
rect 96764 81252 96816 81304
rect 109828 81252 109880 81304
rect 190604 81252 190656 81304
rect 203760 81252 203812 81304
rect 283432 81252 283484 81304
rect 428056 81252 428108 81304
rect 129240 80572 129292 80624
rect 131264 80572 131316 80624
rect 223080 80572 223132 80624
rect 225196 80572 225248 80624
rect 316920 80572 316972 80624
rect 319128 80572 319180 80624
rect 60240 79144 60292 79196
rect 64380 79144 64432 79196
rect 153344 79144 153396 79196
rect 156840 79144 156892 79196
rect 156932 79144 156984 79196
rect 157576 79144 157628 79196
rect 159600 79144 159652 79196
rect 160336 79144 160388 79196
rect 250772 79144 250824 79196
rect 251416 79144 251468 79196
rect 253532 79144 253584 79196
rect 254176 79144 254228 79196
rect 333388 79144 333440 79196
rect 334124 79144 334176 79196
rect 334400 79144 334452 79196
rect 335412 79144 335464 79196
rect 339552 79144 339604 79196
rect 343784 79144 343836 79196
rect 344704 79144 344756 79196
rect 59228 79076 59280 79128
rect 63828 79076 63880 79128
rect 58216 78940 58268 78992
rect 63736 78940 63788 78992
rect 62356 78872 62408 78924
rect 66680 79076 66732 79128
rect 154540 79076 154592 79128
rect 154724 79076 154776 79128
rect 250404 79076 250456 79128
rect 257580 79076 257632 79128
rect 339000 79076 339052 79128
rect 342680 79076 342732 79128
rect 344612 79076 344664 79128
rect 346820 79076 346872 79128
rect 347280 79144 347332 79196
rect 349948 79144 350000 79196
rect 369268 79144 369320 79196
rect 369820 79144 369872 79196
rect 347924 79076 347976 79128
rect 337528 79008 337580 79060
rect 338264 79008 338316 79060
rect 341852 79008 341904 79060
rect 345808 79008 345860 79060
rect 64380 78872 64432 78924
rect 68520 78872 68572 78924
rect 63644 78804 63696 78856
rect 74776 78804 74828 78856
rect 62264 78736 62316 78788
rect 65484 78736 65536 78788
rect 69348 78736 69400 78788
rect 151964 78940 152016 78992
rect 156104 78940 156156 78992
rect 164476 78940 164528 78992
rect 341760 78940 341812 78992
rect 344796 78940 344848 78992
rect 154724 78872 154776 78924
rect 163188 78872 163240 78924
rect 247644 78872 247696 78924
rect 256200 78872 256252 78924
rect 151964 78804 152016 78856
rect 160980 78804 161032 78856
rect 244884 78804 244936 78856
rect 254820 78804 254872 78856
rect 163096 78736 163148 78788
rect 245804 78736 245856 78788
rect 256936 78736 256988 78788
rect 339092 78736 339144 78788
rect 341668 78736 341720 78788
rect 63368 78668 63420 78720
rect 67140 78668 67192 78720
rect 153252 78668 153304 78720
rect 164568 78668 164620 78720
rect 247092 78668 247144 78720
rect 258408 78668 258460 78720
rect 60884 78600 60936 78652
rect 72660 78600 72712 78652
rect 154632 78600 154684 78652
rect 167328 78600 167380 78652
rect 248564 78600 248616 78652
rect 261076 78600 261128 78652
rect 58124 78532 58176 78584
rect 69624 78532 69676 78584
rect 153068 78532 153120 78584
rect 165948 78532 166000 78584
rect 247184 78532 247236 78584
rect 259696 78532 259748 78584
rect 344520 78532 344572 78584
rect 348936 78532 348988 78584
rect 55364 78464 55416 78516
rect 66496 78464 66548 78516
rect 154540 78464 154592 78516
rect 168708 78464 168760 78516
rect 248472 78464 248524 78516
rect 262456 78464 262508 78516
rect 338540 78464 338592 78516
rect 349488 78464 349540 78516
rect 59504 78396 59556 78448
rect 70636 78396 70688 78448
rect 73764 78328 73816 78380
rect 65852 78192 65904 78244
rect 67508 78192 67560 78244
rect 246264 78124 246316 78176
rect 250680 78124 250732 78176
rect 57204 78056 57256 78108
rect 61620 78056 61672 78108
rect 61344 77988 61396 78040
rect 65760 77988 65812 78040
rect 249024 77920 249076 77972
rect 253440 77920 253492 77972
rect 75788 77852 75840 77904
rect 76892 77852 76944 77904
rect 369912 76467 369964 76476
rect 369912 76433 369921 76467
rect 369921 76433 369955 76467
rect 369955 76433 369964 76467
rect 369912 76424 369964 76433
rect 78916 76356 78968 76408
rect 123996 76356 124048 76408
rect 139636 76356 139688 76408
rect 173860 76356 173912 76408
rect 218020 76356 218072 76408
rect 233476 76356 233528 76408
rect 266596 76356 266648 76408
rect 312044 76356 312096 76408
rect 328420 76356 328472 76408
rect 427412 76356 427464 76408
rect 429436 76356 429488 76408
rect 155368 75515 155420 75524
rect 155368 75481 155377 75515
rect 155377 75481 155411 75515
rect 155411 75481 155420 75515
rect 155368 75472 155420 75481
rect 249208 75447 249260 75456
rect 249208 75413 249217 75447
rect 249217 75413 249251 75447
rect 249251 75413 249260 75447
rect 249208 75404 249260 75413
rect 78916 73704 78968 73756
rect 87380 73704 87432 73756
rect 170640 73704 170692 73756
rect 264480 73704 264532 73756
rect 304868 73704 304920 73756
rect 305052 73704 305104 73756
rect 110196 73432 110248 73484
rect 116820 73432 116872 73484
rect 204128 72956 204180 73008
rect 210936 72956 210988 73008
rect 217560 72956 217612 73008
rect 223080 72956 223132 73008
rect 311216 72480 311268 72532
rect 316920 72480 316972 72532
rect 78916 72344 78968 72396
rect 87196 72344 87248 72396
rect 123536 72344 123588 72396
rect 129240 72344 129292 72396
rect 173492 72344 173544 72396
rect 178276 72344 178328 72396
rect 230164 72344 230216 72396
rect 233476 72344 233528 72396
rect 266596 72344 266648 72396
rect 274968 72344 275020 72396
rect 284536 72344 284588 72396
rect 285824 72344 285876 72396
rect 297876 72344 297928 72396
rect 304868 72344 304920 72396
rect 173492 71732 173544 71784
rect 178368 71732 178420 71784
rect 78916 70984 78968 71036
rect 85724 70984 85776 71036
rect 173308 70984 173360 71036
rect 180852 70984 180904 71036
rect 266688 70984 266740 71036
rect 274784 70984 274836 71036
rect 266596 70916 266648 70968
rect 274692 70916 274744 70968
rect 173308 70032 173360 70084
rect 178460 70032 178512 70084
rect 78916 69556 78968 69608
rect 84896 69556 84948 69608
rect 229888 69556 229940 69608
rect 233568 69556 233620 69608
rect 266596 69556 266648 69608
rect 270552 69556 270604 69608
rect 131448 69488 131500 69540
rect 139636 69488 139688 69540
rect 172940 69488 172992 69540
rect 182324 69488 182376 69540
rect 226300 69488 226352 69540
rect 233936 69488 233988 69540
rect 267424 69488 267476 69540
rect 274876 69488 274928 69540
rect 369728 69488 369780 69540
rect 369912 69488 369964 69540
rect 131356 69420 131408 69472
rect 139820 69420 139872 69472
rect 178276 69420 178328 69472
rect 181680 69420 181732 69472
rect 226392 69420 226444 69472
rect 230164 69420 230216 69472
rect 321612 68536 321664 68588
rect 327040 68536 327092 68588
rect 321612 68332 321664 68384
rect 327868 68332 327920 68384
rect 78916 68196 78968 68248
rect 85632 68196 85684 68248
rect 136692 68196 136744 68248
rect 139636 68196 139688 68248
rect 173124 68196 173176 68248
rect 178276 68196 178328 68248
rect 266596 68196 266648 68248
rect 272668 68196 272720 68248
rect 85724 68128 85776 68180
rect 87196 68128 87248 68180
rect 132368 68128 132420 68180
rect 139728 68128 139780 68180
rect 178368 68128 178420 68180
rect 181404 68128 181456 68180
rect 226300 68128 226352 68180
rect 233476 68128 233528 68180
rect 79560 67516 79612 67568
rect 129424 67516 129476 67568
rect 173400 67516 173452 67568
rect 223448 67516 223500 67568
rect 267240 67516 267292 67568
rect 317564 67516 317616 67568
rect 320508 67176 320560 67228
rect 327132 67176 327184 67228
rect 78916 67040 78968 67092
rect 81676 67040 81728 67092
rect 78916 66904 78968 66956
rect 85172 66904 85224 66956
rect 174044 66904 174096 66956
rect 179104 66904 179156 66956
rect 136784 66836 136836 66888
rect 139728 66836 139780 66888
rect 266688 66836 266740 66888
rect 272484 66836 272536 66888
rect 321060 66836 321112 66888
rect 328420 66836 328472 66888
rect 136140 66768 136192 66820
rect 139636 66768 139688 66820
rect 173676 66768 173728 66820
rect 175608 66768 175660 66820
rect 230072 66768 230124 66820
rect 233476 66768 233528 66820
rect 266596 66768 266648 66820
rect 272760 66768 272812 66820
rect 369268 66768 369320 66820
rect 369820 66768 369872 66820
rect 80296 66700 80348 66752
rect 87196 66700 87248 66752
rect 129424 66743 129476 66752
rect 129424 66709 129433 66743
rect 129433 66709 129467 66743
rect 129467 66709 129476 66743
rect 129424 66700 129476 66709
rect 132368 66700 132420 66752
rect 139912 66700 139964 66752
rect 226300 66700 226352 66752
rect 233752 66700 233804 66752
rect 270552 66700 270604 66752
rect 274876 66700 274928 66752
rect 84896 66632 84948 66684
rect 87288 66632 87340 66684
rect 131356 66632 131408 66684
rect 140004 66632 140056 66684
rect 226300 66360 226352 66412
rect 229888 66360 229940 66412
rect 178460 66156 178512 66208
rect 181772 66156 181824 66208
rect 321612 65816 321664 65868
rect 326948 65816 327000 65868
rect 174044 65680 174096 65732
rect 178736 65680 178788 65732
rect 321428 65680 321480 65732
rect 326856 65680 326908 65732
rect 78916 65408 78968 65460
rect 84436 65408 84488 65460
rect 229428 65408 229480 65460
rect 233476 65408 233528 65460
rect 266596 65408 266648 65460
rect 274968 65408 275020 65460
rect 321704 65408 321756 65460
rect 328420 65408 328472 65460
rect 81676 65340 81728 65392
rect 87196 65340 87248 65392
rect 131448 65340 131500 65392
rect 136784 65340 136836 65392
rect 178276 65340 178328 65392
rect 182324 65340 182376 65392
rect 225932 65340 225984 65392
rect 233568 65340 233620 65392
rect 272484 65340 272536 65392
rect 274876 65340 274928 65392
rect 85632 65272 85684 65324
rect 87288 65272 87340 65324
rect 131356 65272 131408 65324
rect 136692 65272 136744 65324
rect 175608 65272 175660 65324
rect 181588 65272 181640 65324
rect 226208 65272 226260 65324
rect 233660 65272 233712 65324
rect 272668 65272 272720 65324
rect 275060 65272 275112 65324
rect 321428 65068 321480 65120
rect 327684 65068 327736 65120
rect 321612 64728 321664 64780
rect 327040 64728 327092 64780
rect 173124 64524 173176 64576
rect 176068 64524 176120 64576
rect 78916 64456 78968 64508
rect 81676 64456 81728 64508
rect 266596 64048 266648 64100
rect 273036 64048 273088 64100
rect 132368 63980 132420 64032
rect 136140 63980 136192 64032
rect 179104 63980 179156 64032
rect 182324 63980 182376 64032
rect 225748 63980 225800 64032
rect 230072 63980 230124 64032
rect 85172 63572 85224 63624
rect 87196 63572 87248 63624
rect 272760 63572 272812 63624
rect 274876 63572 274928 63624
rect 78916 62960 78968 63012
rect 81768 62960 81820 63012
rect 174044 62688 174096 62740
rect 178276 62688 178328 62740
rect 266688 62688 266740 62740
rect 272760 62688 272812 62740
rect 78916 62620 78968 62672
rect 87380 62620 87432 62672
rect 173492 62620 173544 62672
rect 175608 62620 175660 62672
rect 230164 62620 230216 62672
rect 233476 62620 233528 62672
rect 266596 62620 266648 62672
rect 275060 62620 275112 62672
rect 81676 62552 81728 62604
rect 87196 62552 87248 62604
rect 131724 62552 131776 62604
rect 139636 62552 139688 62604
rect 176068 62552 176120 62604
rect 181588 62552 181640 62604
rect 225932 62552 225984 62604
rect 234580 62552 234632 62604
rect 273036 62552 273088 62604
rect 274876 62552 274928 62604
rect 84436 62484 84488 62536
rect 87288 62484 87340 62536
rect 131356 62484 131408 62536
rect 139912 62484 139964 62536
rect 178736 62484 178788 62536
rect 182324 62484 182376 62536
rect 226300 62348 226352 62400
rect 229428 62348 229480 62400
rect 321244 62348 321296 62400
rect 327316 62348 327368 62400
rect 173124 61600 173176 61652
rect 175516 61600 175568 61652
rect 78916 61328 78968 61380
rect 81676 61328 81728 61380
rect 266596 61260 266648 61312
rect 272668 61260 272720 61312
rect 321060 61260 321112 61312
rect 328512 61260 328564 61312
rect 81768 61192 81820 61244
rect 87196 61192 87248 61244
rect 131356 61192 131408 61244
rect 139728 61192 139780 61244
rect 175608 61192 175660 61244
rect 181220 61192 181272 61244
rect 272760 61192 272812 61244
rect 274876 61192 274928 61244
rect 226300 61056 226352 61108
rect 230164 61056 230216 61108
rect 320876 60988 320928 61040
rect 328052 60988 328104 61040
rect 78916 59900 78968 59952
rect 85724 59900 85776 59952
rect 136784 59900 136836 59952
rect 139728 59900 139780 59952
rect 173492 59900 173544 59952
rect 175608 59900 175660 59952
rect 266596 59900 266648 59952
rect 274968 59900 275020 59952
rect 369728 59900 369780 59952
rect 370004 59900 370056 59952
rect 81676 59832 81728 59884
rect 87196 59832 87248 59884
rect 132644 59832 132696 59884
rect 139820 59832 139872 59884
rect 175516 59832 175568 59884
rect 181588 59832 181640 59884
rect 226116 59832 226168 59884
rect 233568 59832 233620 59884
rect 272668 59832 272720 59884
rect 274876 59832 274928 59884
rect 369268 59832 369320 59884
rect 369820 59832 369872 59884
rect 132552 59764 132604 59816
rect 139636 59764 139688 59816
rect 178276 59764 178328 59816
rect 182324 59764 182376 59816
rect 226300 59764 226352 59816
rect 233476 59764 233528 59816
rect 321612 58744 321664 58796
rect 328328 58744 328380 58796
rect 135496 58608 135548 58660
rect 139728 58608 139780 58660
rect 230348 58608 230400 58660
rect 233568 58608 233620 58660
rect 266596 58608 266648 58660
rect 272576 58608 272628 58660
rect 136416 58540 136468 58592
rect 139636 58540 139688 58592
rect 230624 58540 230676 58592
rect 233476 58540 233528 58592
rect 266688 58540 266740 58592
rect 272760 58540 272812 58592
rect 85724 58472 85776 58524
rect 87196 58472 87248 58524
rect 132644 58472 132696 58524
rect 136784 58472 136836 58524
rect 175608 58472 175660 58524
rect 182324 58472 182376 58524
rect 226300 58472 226352 58524
rect 233660 58472 233712 58524
rect 173492 57384 173544 57436
rect 176252 57384 176304 57436
rect 320876 57180 320928 57232
rect 328420 57180 328472 57232
rect 78916 57112 78968 57164
rect 87380 57112 87432 57164
rect 129516 57112 129568 57164
rect 266596 57112 266648 57164
rect 274968 57112 275020 57164
rect 80388 57044 80440 57096
rect 87196 57044 87248 57096
rect 132644 57044 132696 57096
rect 135496 57044 135548 57096
rect 272760 57044 272812 57096
rect 274876 57044 274928 57096
rect 80296 56976 80348 57028
rect 87288 56976 87340 57028
rect 132552 56976 132604 57028
rect 136416 56976 136468 57028
rect 272576 56976 272628 57028
rect 275060 56976 275112 57028
rect 226300 56908 226352 56960
rect 230348 56908 230400 56960
rect 225380 56636 225432 56688
rect 230624 56636 230676 56688
rect 174136 56568 174188 56620
rect 181772 56568 181824 56620
rect 174228 56432 174280 56484
rect 182324 56432 182376 56484
rect 321612 56296 321664 56348
rect 327684 56296 327736 56348
rect 321060 56024 321112 56076
rect 328512 56024 328564 56076
rect 78916 55752 78968 55804
rect 81676 55752 81728 55804
rect 172756 55752 172808 55804
rect 176804 55752 176856 55804
rect 266596 55752 266648 55804
rect 273404 55752 273456 55804
rect 324556 55752 324608 55804
rect 327500 55752 327552 55804
rect 132644 55684 132696 55736
rect 139636 55684 139688 55736
rect 176252 55684 176304 55736
rect 181680 55684 181732 55736
rect 225380 55684 225432 55736
rect 233476 55684 233528 55736
rect 134208 55072 134260 55124
rect 369728 55072 369780 55124
rect 370004 55072 370056 55124
rect 223448 55004 223500 55056
rect 233476 55004 233528 55056
rect 317472 55004 317524 55056
rect 328512 55004 328564 55056
rect 358504 55004 358556 55056
rect 389416 55004 389468 55056
rect 321612 54936 321664 54988
rect 328328 54936 328380 54988
rect 129516 54868 129568 54920
rect 78916 54392 78968 54444
rect 87288 54392 87340 54444
rect 134116 54392 134168 54444
rect 139636 54392 139688 54444
rect 174044 54392 174096 54444
rect 81676 54324 81728 54376
rect 87196 54324 87248 54376
rect 132644 54324 132696 54376
rect 139544 54324 139596 54376
rect 223540 54324 223592 54376
rect 233476 54392 233528 54444
rect 266596 54392 266648 54444
rect 226300 54324 226352 54376
rect 234396 54324 234448 54376
rect 273404 54324 273456 54376
rect 274876 54324 274928 54376
rect 317472 54392 317524 54444
rect 328420 54392 328472 54444
rect 320968 54324 321020 54376
rect 324556 54324 324608 54376
rect 176804 54188 176856 54240
rect 182324 54188 182376 54240
rect 78916 53712 78968 53764
rect 118200 53712 118252 53764
rect 139636 53712 139688 53764
rect 87288 53644 87340 53696
rect 128688 53644 128740 53696
rect 134116 53644 134168 53696
rect 174044 53644 174096 53696
rect 212040 53644 212092 53696
rect 233476 53644 233528 53696
rect 266596 53644 266648 53696
rect 306984 53644 307036 53696
rect 328420 53644 328472 53696
rect 129056 52284 129108 52336
rect 129516 52284 129568 52336
rect 91244 51536 91296 51588
rect 134760 51536 134812 51588
rect 184992 51536 185044 51588
rect 228600 51536 228652 51588
rect 279016 51536 279068 51588
rect 323820 51536 323872 51588
rect 427596 51536 427648 51588
rect 429804 51536 429856 51588
rect 78180 51468 78232 51520
rect 93636 51468 93688 51520
rect 170180 51468 170232 51520
rect 170640 51468 170692 51520
rect 189684 51468 189736 51520
rect 111944 51128 111996 51180
rect 121236 51128 121288 51180
rect 205784 51128 205836 51180
rect 215536 51128 215588 51180
rect 299624 51128 299676 51180
rect 309560 51128 309612 51180
rect 106424 51060 106476 51112
rect 118936 51060 118988 51112
rect 200264 51060 200316 51112
rect 213236 51060 213288 51112
rect 294104 51060 294156 51112
rect 307260 51060 307312 51112
rect 102284 50992 102336 51044
rect 116544 50992 116596 51044
rect 196124 50992 196176 51044
rect 210844 50992 210896 51044
rect 289964 50992 290016 51044
rect 304868 50992 304920 51044
rect 114152 50924 114204 50976
rect 122340 50924 122392 50976
rect 125928 50924 125980 50976
rect 190604 50924 190656 50976
rect 208452 50924 208504 50976
rect 284444 50924 284496 50976
rect 302476 50924 302528 50976
rect 91244 50856 91296 50908
rect 112036 50856 112088 50908
rect 116084 50856 116136 50908
rect 123628 50856 123680 50908
rect 185084 50856 185136 50908
rect 206152 50856 206204 50908
rect 280304 50856 280356 50908
rect 300176 50856 300228 50908
rect 305144 50856 305196 50908
rect 311952 50856 312004 50908
rect 216180 50652 216232 50704
rect 220228 50652 220280 50704
rect 211304 50380 211356 50432
rect 217928 50380 217980 50432
rect 310020 50380 310072 50432
rect 314252 50380 314304 50432
rect 79008 50312 79060 50364
rect 108632 50312 108684 50364
rect 139728 50312 139780 50364
rect 173952 50312 174004 50364
rect 202564 50312 202616 50364
rect 233568 50312 233620 50364
rect 266688 50312 266740 50364
rect 296588 50312 296640 50364
rect 327684 50312 327736 50364
rect 78916 50244 78968 50296
rect 103572 50244 103624 50296
rect 139636 50244 139688 50296
rect 174044 50244 174096 50296
rect 197504 50244 197556 50296
rect 233476 50244 233528 50296
rect 266596 50244 266648 50296
rect 291528 50244 291580 50296
rect 328420 50244 328472 50296
rect 288308 50176 288360 50228
rect 327224 50176 327276 50228
rect 274968 49564 275020 49616
rect 275612 49564 275664 49616
rect 288308 49564 288360 49616
rect 87472 49496 87524 49548
rect 88392 49496 88444 49548
rect 102376 49496 102428 49548
rect 181864 49496 181916 49548
rect 194376 49496 194428 49548
rect 275060 49496 275112 49548
rect 275888 49496 275940 49548
rect 297784 49496 297836 49548
rect 78916 48884 78968 48936
rect 98604 48884 98656 48936
rect 140556 48884 140608 48936
rect 173308 48884 173360 48936
rect 192536 48884 192588 48936
rect 233476 48884 233528 48936
rect 266596 48884 266648 48936
rect 286560 48884 286612 48936
rect 328512 48884 328564 48936
rect 359700 48884 359752 48936
rect 96764 48519 96816 48528
rect 96764 48485 96773 48519
rect 96773 48485 96807 48519
rect 96807 48485 96816 48519
rect 96764 48476 96816 48485
rect 182232 48136 182284 48188
rect 196676 48136 196728 48188
rect 275796 48136 275848 48188
rect 276072 48136 276124 48188
rect 290700 48136 290752 48188
rect 357308 48179 357360 48188
rect 357308 48145 357317 48179
rect 357317 48145 357351 48179
rect 357351 48145 357360 48179
rect 357308 48136 357360 48145
rect 140004 47660 140056 47712
rect 142856 47524 142908 47576
rect 159508 47524 159560 47576
rect 100444 47456 100496 47508
rect 100904 47456 100956 47508
rect 156840 47456 156892 47508
rect 167604 47456 167656 47508
rect 174044 47456 174096 47508
rect 187568 47456 187620 47508
rect 233476 47456 233528 47508
rect 266596 47456 266648 47508
rect 281592 47456 281644 47508
rect 328052 47456 328104 47508
rect 369268 47456 369320 47508
rect 369820 47456 369872 47508
rect 13044 47388 13096 47440
rect 16540 47388 16592 47440
rect 60700 47388 60752 47440
rect 72568 47388 72620 47440
rect 73304 47388 73356 47440
rect 294196 47388 294248 47440
rect 295484 47388 295536 47440
rect 353628 47388 353680 47440
rect 419776 47388 419828 47440
rect 285916 47320 285968 47372
rect 339644 47320 339696 47372
rect 87104 47184 87156 47236
rect 93636 47184 93688 47236
rect 88024 46776 88076 46828
rect 100904 46776 100956 46828
rect 74684 46708 74736 46760
rect 87196 46708 87248 46760
rect 275888 46708 275940 46760
rect 294196 46708 294248 46760
rect 71188 46164 71240 46216
rect 74316 46164 74368 46216
rect 88208 46164 88260 46216
rect 106608 46164 106660 46216
rect 73304 46096 73356 46148
rect 87196 46096 87248 46148
rect 88116 46096 88168 46148
rect 109460 46096 109512 46148
rect 50212 46028 50264 46080
rect 369544 46028 369596 46080
rect 53708 45960 53760 46012
rect 95476 45960 95528 46012
rect 144696 45960 144748 46012
rect 369728 45960 369780 46012
rect 57204 45892 57256 45944
rect 98052 45892 98104 45944
rect 153436 45892 153488 45944
rect 238628 45892 238680 45944
rect 322624 45892 322676 45944
rect 338356 45892 338408 45944
rect 343140 45892 343192 45944
rect 350132 45892 350184 45944
rect 417016 45892 417068 45944
rect 95476 45824 95528 45876
rect 95752 45824 95804 45876
rect 150584 45824 150636 45876
rect 170180 45824 170232 45876
rect 256936 45824 256988 45876
rect 263192 45824 263244 45876
rect 283708 45824 283760 45876
rect 336148 45824 336200 45876
rect 332652 45756 332704 45808
rect 369820 45756 369872 45808
rect 182048 45416 182100 45468
rect 201460 45416 201512 45468
rect 339644 45416 339696 45468
rect 350776 45416 350828 45468
rect 168892 45348 168944 45400
rect 181956 45348 182008 45400
rect 203760 45348 203812 45400
rect 275980 45348 276032 45400
rect 293092 45348 293144 45400
rect 324556 45348 324608 45400
rect 350132 45348 350184 45400
rect 169720 44736 169772 44788
rect 182048 44736 182100 44788
rect 263192 44736 263244 44788
rect 275980 44736 276032 44788
rect 101364 37732 101416 37784
rect 102284 37732 102336 37784
rect 210016 37732 210068 37784
rect 211304 37732 211356 37784
rect 289044 37732 289096 37784
rect 289964 37732 290016 37784
rect 304040 37732 304092 37784
rect 305144 37732 305196 37784
rect 309100 37732 309152 37784
rect 310020 37732 310072 37784
rect 126388 37596 126440 37648
rect 128596 37596 128648 37648
rect 96396 37460 96448 37512
rect 96764 37460 96816 37512
rect 195020 37392 195072 37444
rect 196124 37392 196176 37444
rect 215076 37392 215128 37444
rect 216180 37392 216232 37444
rect 220044 37392 220096 37444
rect 222436 37392 222488 37444
rect 279108 37324 279160 37376
rect 280304 37324 280356 37376
rect 121420 37256 121472 37308
rect 122340 37256 122392 37308
rect 217560 37052 217612 37104
rect 223540 37052 223592 37104
rect 123904 36712 123956 36764
rect 128688 36712 128740 36764
rect 111392 36644 111444 36696
rect 111944 36644 111996 36696
rect 311584 36508 311636 36560
rect 317472 36508 317524 36560
rect 314068 36440 314120 36492
rect 316276 36440 316328 36492
rect 12860 36304 12912 36356
rect 16448 36304 16500 36356
rect 276164 33040 276216 33092
rect 369636 33040 369688 33092
rect 182324 32972 182376 33024
rect 369452 32972 369504 33024
rect 88484 32904 88536 32956
rect 369176 32904 369228 32956
rect 427504 28076 427556 28128
rect 429436 28076 429488 28128
rect 12676 24948 12728 25000
rect 16264 24948 16316 25000
rect 185176 17060 185228 17112
rect 186372 17060 186424 17112
rect 191340 17060 191392 17112
rect 192076 17060 192128 17112
rect 288676 17060 288728 17112
rect 290332 17060 290384 17112
rect 194560 16992 194612 17044
rect 196308 16992 196360 17044
rect 92624 16788 92676 16840
rect 105136 16788 105188 16840
rect 80756 16720 80808 16772
rect 102376 16720 102428 16772
rect 285364 16720 285416 16772
rect 299716 16720 299768 16772
rect 67876 16652 67928 16704
rect 107068 16652 107120 16704
rect 170916 16652 170968 16704
rect 201368 16652 201420 16704
rect 273956 16652 274008 16704
rect 295392 16652 295444 16704
rect 54996 16584 55048 16636
rect 112036 16584 112088 16636
rect 158036 16584 158088 16636
rect 206336 16584 206388 16636
rect 261076 16584 261128 16636
rect 300360 16584 300412 16636
rect 29236 16516 29288 16568
rect 122064 16516 122116 16568
rect 145156 16516 145208 16568
rect 211304 16516 211356 16568
rect 248196 16516 248248 16568
rect 305328 16516 305380 16568
rect 42116 16448 42168 16500
rect 117004 16448 117056 16500
rect 119396 16448 119448 16500
rect 221332 16448 221384 16500
rect 235316 16448 235368 16500
rect 310388 16448 310440 16500
rect 16356 16380 16408 16432
rect 127216 16380 127268 16432
rect 132276 16380 132328 16432
rect 216364 16380 216416 16432
rect 222436 16380 222488 16432
rect 315356 16380 315408 16432
rect 95476 16040 95528 16092
rect 97040 16040 97092 16092
rect 427320 15292 427372 15344
rect 429436 15292 429488 15344
rect 12676 14204 12728 14256
rect 16080 14204 16132 14256
rect 93636 12572 93688 12624
rect 95476 12572 95528 12624
rect 286836 12368 286888 12420
rect 288676 12368 288728 12420
rect 325292 12368 325344 12420
rect 364116 12368 364168 12420
rect 376996 12368 377048 12420
rect 378284 12368 378336 12420
rect 105136 12300 105188 12352
rect 106516 12300 106568 12352
rect 183796 12300 183848 12352
rect 194560 12300 194612 12352
rect 362460 12300 362512 12352
rect 402756 12300 402808 12352
rect 185176 12232 185228 12284
rect 209556 12232 209608 12284
rect 280396 12232 280448 12284
rect 312596 12232 312648 12284
rect 322532 12232 322584 12284
rect 415636 12232 415688 12284
rect 192076 12096 192128 12148
rect 196676 12096 196728 12148
rect 350776 9376 350828 9428
rect 351236 9376 351288 9428
rect 389416 9376 389468 9428
rect 389876 9376 389928 9428
rect 428056 9376 428108 9428
rect 428516 9376 428568 9428
<< metal2 >>
rect 23162 396344 23218 396824
rect 49658 396344 49714 396824
rect 76246 396344 76302 396824
rect 102834 396344 102890 396824
rect 129422 396344 129478 396824
rect 155918 396344 155974 396824
rect 182506 396344 182562 396824
rect 209094 396344 209150 396824
rect 235682 396344 235738 396824
rect 262178 396344 262234 396824
rect 288766 396344 288822 396824
rect 315354 396344 315410 396824
rect 341942 396344 341998 396824
rect 368438 396344 368494 396824
rect 395026 396344 395082 396824
rect 421614 396344 421670 396824
rect 23176 393838 23204 396344
rect 49672 393838 49700 396344
rect 76260 396234 76288 396344
rect 76168 396206 76288 396234
rect 22336 393832 22388 393838
rect 22336 393774 22388 393780
rect 23164 393832 23216 393838
rect 23164 393774 23216 393780
rect 48556 393832 48608 393838
rect 48556 393774 48608 393780
rect 49660 393832 49712 393838
rect 49660 393774 49712 393780
rect 13134 391352 13190 391361
rect 13134 391287 13190 391296
rect 13148 391118 13176 391287
rect 13136 391112 13188 391118
rect 13136 391054 13188 391060
rect 22348 389010 22376 393774
rect 48568 389078 48596 393774
rect 76168 389146 76196 396206
rect 102848 393158 102876 396344
rect 129436 393838 129464 396344
rect 155932 393838 155960 396344
rect 182520 396234 182548 396344
rect 209108 396234 209136 396344
rect 182428 396206 182548 396234
rect 208648 396206 209136 396234
rect 128596 393832 128648 393838
rect 128596 393774 128648 393780
rect 129424 393832 129476 393838
rect 129424 393774 129476 393780
rect 154816 393832 154868 393838
rect 154816 393774 154868 393780
rect 155920 393832 155972 393838
rect 155920 393774 155972 393780
rect 102836 393152 102888 393158
rect 102836 393094 102888 393100
rect 108908 393152 108960 393158
rect 108908 393094 108960 393100
rect 87196 391112 87248 391118
rect 87196 391054 87248 391060
rect 76156 389140 76208 389146
rect 76156 389082 76208 389088
rect 48556 389072 48608 389078
rect 48556 389014 48608 389020
rect 22336 389004 22388 389010
rect 22336 388946 22388 388952
rect 13504 388664 13556 388670
rect 13504 388606 13556 388612
rect 13320 388596 13372 388602
rect 13320 388538 13372 388544
rect 13332 337505 13360 388538
rect 13412 388392 13464 388398
rect 13412 388334 13464 388340
rect 13424 348249 13452 388334
rect 13516 359129 13544 388606
rect 13688 388528 13740 388534
rect 13688 388470 13740 388476
rect 13596 388460 13648 388466
rect 13596 388402 13648 388408
rect 13608 369873 13636 388402
rect 13700 380617 13728 388470
rect 13686 380608 13742 380617
rect 13686 380543 13742 380552
rect 13594 369864 13650 369873
rect 13594 369799 13650 369808
rect 53708 359832 53760 359838
rect 53708 359774 53760 359780
rect 76984 359832 77036 359838
rect 76984 359774 77036 359780
rect 50212 359764 50264 359770
rect 50212 359706 50264 359712
rect 13502 359120 13558 359129
rect 13502 359055 13558 359064
rect 50224 357732 50252 359706
rect 53720 357732 53748 359774
rect 76800 359764 76852 359770
rect 76800 359706 76852 359712
rect 64196 359696 64248 359702
rect 64196 359638 64248 359644
rect 76064 359696 76116 359702
rect 76064 359638 76116 359644
rect 60700 359628 60752 359634
rect 60700 359570 60752 359576
rect 57204 359560 57256 359566
rect 57204 359502 57256 359508
rect 57216 357732 57244 359502
rect 60712 357732 60740 359570
rect 64208 357732 64236 359638
rect 75880 359628 75932 359634
rect 75880 359570 75932 359576
rect 75788 359560 75840 359566
rect 75788 359502 75840 359508
rect 67692 359424 67744 359430
rect 67692 359366 67744 359372
rect 67704 357732 67732 359366
rect 75800 357594 75828 359502
rect 75892 357662 75920 359570
rect 75972 359424 76024 359430
rect 75972 359366 76024 359372
rect 75880 357656 75932 357662
rect 75880 357598 75932 357604
rect 75788 357588 75840 357594
rect 75788 357530 75840 357536
rect 71464 357520 71516 357526
rect 71214 357468 71464 357474
rect 75880 357520 75932 357526
rect 71214 357462 71516 357468
rect 71214 357446 71504 357462
rect 74710 357458 74816 357474
rect 75880 357462 75932 357468
rect 74710 357452 74828 357458
rect 74710 357446 74776 357452
rect 74776 357394 74828 357400
rect 13410 348240 13466 348249
rect 13410 348175 13466 348184
rect 13318 337496 13374 337505
rect 13318 337431 13374 337440
rect 75892 334746 75920 357462
rect 75984 334814 76012 359366
rect 76076 349706 76104 359638
rect 76156 357656 76208 357662
rect 76156 357598 76208 357604
rect 76064 349700 76116 349706
rect 76064 349642 76116 349648
rect 76168 349586 76196 357598
rect 76248 353916 76300 353922
rect 76248 353858 76300 353864
rect 76076 349558 76196 349586
rect 76076 340202 76104 349558
rect 76076 340174 76196 340202
rect 76064 340112 76116 340118
rect 76064 340054 76116 340060
rect 75972 334808 76024 334814
rect 75972 334750 76024 334756
rect 76076 334746 76104 340054
rect 75880 334740 75932 334746
rect 75880 334682 75932 334688
rect 76064 334740 76116 334746
rect 76064 334682 76116 334688
rect 76168 334626 76196 340174
rect 76260 340118 76288 353858
rect 76248 340112 76300 340118
rect 76248 340054 76300 340060
rect 75892 334598 76196 334626
rect 75892 334406 75920 334598
rect 75972 334536 76024 334542
rect 75972 334478 76024 334484
rect 76064 334536 76116 334542
rect 76064 334478 76116 334484
rect 75880 334400 75932 334406
rect 75880 334342 75932 334348
rect 75512 330184 75564 330190
rect 75512 330126 75564 330132
rect 75420 330116 75472 330122
rect 75420 330058 75472 330064
rect 48568 329838 48950 329866
rect 14698 326752 14754 326761
rect 14698 326687 14754 326696
rect 14712 326450 14740 326687
rect 14700 326444 14752 326450
rect 14700 326386 14752 326392
rect 13318 316008 13374 316017
rect 13318 315943 13374 315952
rect 13044 273744 13096 273750
rect 13044 273686 13096 273692
rect 13056 272905 13084 273686
rect 13042 272896 13098 272905
rect 13042 272831 13098 272840
rect 13332 262734 13360 315943
rect 38804 315904 38856 315910
rect 38804 315846 38856 315852
rect 38816 315609 38844 315846
rect 38802 315600 38858 315609
rect 38802 315535 38858 315544
rect 16078 313832 16134 313841
rect 16078 313767 16134 313776
rect 38436 313796 38488 313802
rect 13410 305128 13466 305137
rect 13410 305063 13466 305072
rect 13320 262728 13372 262734
rect 13320 262670 13372 262676
rect 13424 262666 13452 305063
rect 13502 294384 13558 294393
rect 13502 294319 13558 294328
rect 13412 262660 13464 262666
rect 13412 262602 13464 262608
rect 13516 262598 13544 294319
rect 13596 279388 13648 279394
rect 13596 279330 13648 279336
rect 13504 262592 13556 262598
rect 13504 262534 13556 262540
rect 13608 262025 13636 279330
rect 13594 262016 13650 262025
rect 13594 261951 13650 261960
rect 13136 251508 13188 251514
rect 13136 251450 13188 251456
rect 13148 251281 13176 251450
rect 13134 251272 13190 251281
rect 13134 251207 13190 251216
rect 13320 240560 13372 240566
rect 13318 240528 13320 240537
rect 13372 240528 13374 240537
rect 13318 240463 13374 240472
rect 12860 230972 12912 230978
rect 12860 230914 12912 230920
rect 12872 229793 12900 230914
rect 12858 229784 12914 229793
rect 12858 229719 12914 229728
rect 13044 219412 13096 219418
rect 13044 219354 13096 219360
rect 13056 218913 13084 219354
rect 13042 218904 13098 218913
rect 13042 218839 13098 218848
rect 13044 208192 13096 208198
rect 13042 208160 13044 208169
rect 13096 208160 13098 208169
rect 13042 208095 13098 208104
rect 13320 199352 13372 199358
rect 13320 199294 13372 199300
rect 13044 197788 13096 197794
rect 13044 197730 13096 197736
rect 13056 197425 13084 197730
rect 13042 197416 13098 197425
rect 13042 197351 13098 197360
rect 13044 186704 13096 186710
rect 13042 186672 13044 186681
rect 13096 186672 13098 186681
rect 13042 186607 13098 186616
rect 13044 175824 13096 175830
rect 13042 175792 13044 175801
rect 13096 175792 13098 175801
rect 13042 175727 13098 175736
rect 12676 154812 12728 154818
rect 12676 154754 12728 154760
rect 12688 154313 12716 154754
rect 12674 154304 12730 154313
rect 12674 154239 12730 154248
rect 13332 143569 13360 199294
rect 13412 189696 13464 189702
rect 13412 189638 13464 189644
rect 13424 165057 13452 189638
rect 16092 186710 16120 313767
rect 38436 313738 38488 313744
rect 38448 313161 38476 313738
rect 38434 313152 38490 313161
rect 38434 313087 38490 313096
rect 38802 310432 38858 310441
rect 38802 310367 38858 310376
rect 38816 310334 38844 310367
rect 38804 310328 38856 310334
rect 38804 310270 38856 310276
rect 16262 308392 16318 308401
rect 16262 308327 16318 308336
rect 16170 293160 16226 293169
rect 16170 293095 16226 293104
rect 16184 230978 16212 293095
rect 16172 230972 16224 230978
rect 16172 230914 16224 230920
rect 16170 219992 16226 220001
rect 16170 219927 16226 219936
rect 16080 186704 16132 186710
rect 16080 186646 16132 186652
rect 16078 184224 16134 184233
rect 16078 184159 16134 184168
rect 16092 175830 16120 184159
rect 16080 175824 16132 175830
rect 16080 175766 16132 175772
rect 13410 165048 13466 165057
rect 13410 164983 13466 164992
rect 13318 143560 13374 143569
rect 13318 143495 13374 143504
rect 13044 132984 13096 132990
rect 13044 132926 13096 132932
rect 13056 132689 13084 132926
rect 13042 132680 13098 132689
rect 13042 132615 13098 132624
rect 16078 126152 16134 126161
rect 16078 126087 16134 126096
rect 13228 121968 13280 121974
rect 13226 121936 13228 121945
rect 13280 121936 13282 121945
rect 13226 121871 13282 121880
rect 12860 111564 12912 111570
rect 12860 111506 12912 111512
rect 12872 111201 12900 111506
rect 12858 111192 12914 111201
rect 12858 111127 12914 111136
rect 13320 105512 13372 105518
rect 13320 105454 13372 105460
rect 12860 100820 12912 100826
rect 12860 100762 12912 100768
rect 12872 100457 12900 100762
rect 12858 100448 12914 100457
rect 12858 100383 12914 100392
rect 13228 90212 13280 90218
rect 13228 90154 13280 90160
rect 13240 89577 13268 90154
rect 13226 89568 13282 89577
rect 13226 89503 13282 89512
rect 13332 57345 13360 105454
rect 13412 99936 13464 99942
rect 13412 99878 13464 99884
rect 13424 68089 13452 99878
rect 13504 95856 13556 95862
rect 13504 95798 13556 95804
rect 13516 78833 13544 95798
rect 13502 78824 13558 78833
rect 13502 78759 13558 78768
rect 13410 68080 13466 68089
rect 13410 68015 13466 68024
rect 13318 57336 13374 57345
rect 13318 57271 13374 57280
rect 13044 47440 13096 47446
rect 13044 47382 13096 47388
rect 13056 46465 13084 47382
rect 13042 46456 13098 46465
rect 13042 46391 13098 46400
rect 12860 36356 12912 36362
rect 12860 36298 12912 36304
rect 12872 35721 12900 36298
rect 12858 35712 12914 35721
rect 12858 35647 12914 35656
rect 12676 25000 12728 25006
rect 12674 24968 12676 24977
rect 12728 24968 12730 24977
rect 12674 24903 12730 24912
rect 16092 14262 16120 126087
rect 16184 100826 16212 219927
rect 16276 197794 16304 308327
rect 38804 308288 38856 308294
rect 38804 308230 38856 308236
rect 38816 308129 38844 308230
rect 38802 308120 38858 308129
rect 38802 308055 38858 308064
rect 38804 306248 38856 306254
rect 38804 306190 38856 306196
rect 38816 305681 38844 306190
rect 38802 305672 38858 305681
rect 38802 305607 38858 305616
rect 16446 304176 16502 304185
rect 16446 304111 16502 304120
rect 38620 304140 38672 304146
rect 16354 298736 16410 298745
rect 16354 298671 16410 298680
rect 16368 219418 16396 298671
rect 16356 219412 16408 219418
rect 16356 219354 16408 219360
rect 16354 214552 16410 214561
rect 16354 214487 16410 214496
rect 16264 197788 16316 197794
rect 16264 197730 16316 197736
rect 16262 195376 16318 195385
rect 16262 195311 16318 195320
rect 16276 154818 16304 195311
rect 16264 154812 16316 154818
rect 16264 154754 16316 154760
rect 16262 120712 16318 120721
rect 16262 120647 16318 120656
rect 16172 100820 16224 100826
rect 16172 100762 16224 100768
rect 16276 25006 16304 120647
rect 16368 111570 16396 214487
rect 16460 208198 16488 304111
rect 38620 304082 38672 304088
rect 38632 303097 38660 304082
rect 38618 303088 38674 303097
rect 38618 303023 38674 303032
rect 38804 300672 38856 300678
rect 38802 300640 38804 300649
rect 38856 300640 38858 300649
rect 38802 300575 38858 300584
rect 38252 298632 38304 298638
rect 38252 298574 38304 298580
rect 38264 298201 38292 298574
rect 38250 298192 38306 298201
rect 38250 298127 38306 298136
rect 38802 295472 38858 295481
rect 38802 295407 38858 295416
rect 38816 295170 38844 295407
rect 38804 295164 38856 295170
rect 38804 295106 38856 295112
rect 18010 293840 18066 293849
rect 18010 293775 18066 293784
rect 38436 293804 38488 293810
rect 18024 293169 18052 293775
rect 38436 293746 38488 293752
rect 38448 293169 38476 293746
rect 18010 293160 18066 293169
rect 18010 293095 18066 293104
rect 38434 293160 38490 293169
rect 38434 293095 38490 293104
rect 38528 291696 38580 291702
rect 38528 291638 38580 291644
rect 38540 290585 38568 291638
rect 38526 290576 38582 290585
rect 38526 290511 38582 290520
rect 17458 289080 17514 289089
rect 17458 289015 17514 289024
rect 17472 240566 17500 289015
rect 38528 288976 38580 288982
rect 38528 288918 38580 288924
rect 38540 288137 38568 288918
rect 38526 288128 38582 288137
rect 38526 288063 38582 288072
rect 38526 285544 38582 285553
rect 38526 285479 38528 285488
rect 38580 285479 38582 285488
rect 38528 285450 38580 285456
rect 17550 283776 17606 283785
rect 17550 283711 17606 283720
rect 17564 251514 17592 283711
rect 38528 283468 38580 283474
rect 38528 283410 38580 283416
rect 38540 283105 38568 283410
rect 38526 283096 38582 283105
rect 38526 283031 38582 283040
rect 38066 280376 38122 280385
rect 38066 280311 38122 280320
rect 38080 280006 38108 280311
rect 48568 280006 48596 329838
rect 49948 285514 49976 329852
rect 50040 329838 50974 329866
rect 51328 329838 51986 329866
rect 50040 291702 50068 329838
rect 51222 308664 51278 308673
rect 51222 308599 51278 308608
rect 51236 308294 51264 308599
rect 51224 308288 51276 308294
rect 51224 308230 51276 308236
rect 50304 300672 50356 300678
rect 50302 300640 50304 300649
rect 50356 300640 50358 300649
rect 50302 300575 50358 300584
rect 51328 295170 51356 329838
rect 53076 326353 53104 329852
rect 54088 326353 54116 329852
rect 55100 326353 55128 329852
rect 56112 326353 56140 329852
rect 57216 326790 57244 329852
rect 57204 326784 57256 326790
rect 57204 326726 57256 326732
rect 58228 326586 58256 329852
rect 59240 327402 59268 329852
rect 59228 327396 59280 327402
rect 59228 327338 59280 327344
rect 60252 327334 60280 329852
rect 60240 327328 60292 327334
rect 60240 327270 60292 327276
rect 58216 326580 58268 326586
rect 58216 326522 58268 326528
rect 61356 326450 61384 329852
rect 62368 327198 62396 329852
rect 62356 327192 62408 327198
rect 62356 327134 62408 327140
rect 62264 326784 62316 326790
rect 62264 326726 62316 326732
rect 61344 326444 61396 326450
rect 61344 326386 61396 326392
rect 53062 326344 53118 326353
rect 53062 326279 53118 326288
rect 54074 326344 54130 326353
rect 54074 326279 54130 326288
rect 55086 326344 55142 326353
rect 55086 326279 55142 326288
rect 56098 326344 56154 326353
rect 56098 326279 56154 326288
rect 62276 320670 62304 326726
rect 63380 326654 63408 329852
rect 63644 327396 63696 327402
rect 63644 327338 63696 327344
rect 63368 326648 63420 326654
rect 63368 326590 63420 326596
rect 62448 326580 62500 326586
rect 62448 326522 62500 326528
rect 62264 320664 62316 320670
rect 62264 320606 62316 320612
rect 58768 320528 58820 320534
rect 58768 320470 58820 320476
rect 57020 320324 57072 320330
rect 57020 320266 57072 320272
rect 56100 320256 56152 320262
rect 56100 320198 56152 320204
rect 55272 320052 55324 320058
rect 55272 319994 55324 320000
rect 55284 316796 55312 319994
rect 56112 316796 56140 320198
rect 57032 316796 57060 320266
rect 57940 319984 57992 319990
rect 57940 319926 57992 319932
rect 57952 316796 57980 319926
rect 58780 316796 58808 320470
rect 60608 320460 60660 320466
rect 60608 320402 60660 320408
rect 59688 320392 59740 320398
rect 59688 320334 59740 320340
rect 59700 316796 59728 320334
rect 60620 316796 60648 320402
rect 62356 320188 62408 320194
rect 62356 320130 62408 320136
rect 61436 320120 61488 320126
rect 61436 320062 61488 320068
rect 61448 316796 61476 320062
rect 62368 316796 62396 320130
rect 62460 319922 62488 326522
rect 63276 320664 63328 320670
rect 63276 320606 63328 320612
rect 62448 319916 62500 319922
rect 62448 319858 62500 319864
rect 63288 316796 63316 320606
rect 63656 320534 63684 327338
rect 64392 327062 64420 329852
rect 65496 327538 65524 329852
rect 66522 329838 66720 329866
rect 65484 327532 65536 327538
rect 65484 327474 65536 327480
rect 66312 327396 66364 327402
rect 66312 327338 66364 327344
rect 65024 327328 65076 327334
rect 65024 327270 65076 327276
rect 64380 327056 64432 327062
rect 64380 326998 64432 327004
rect 65036 320618 65064 327270
rect 65036 320590 65156 320618
rect 63644 320528 63696 320534
rect 63644 320470 63696 320476
rect 65024 320528 65076 320534
rect 65024 320470 65076 320476
rect 64104 319916 64156 319922
rect 64104 319858 64156 319864
rect 64116 316796 64144 319858
rect 65036 316796 65064 320470
rect 65128 319378 65156 320590
rect 66324 320262 66352 327338
rect 66496 327328 66548 327334
rect 66496 327270 66548 327276
rect 66404 326444 66456 326450
rect 66404 326386 66456 326392
rect 66312 320256 66364 320262
rect 66312 320198 66364 320204
rect 66416 319394 66444 326386
rect 66508 320330 66536 327270
rect 66588 327192 66640 327198
rect 66588 327134 66640 327140
rect 66496 320324 66548 320330
rect 66496 320266 66548 320272
rect 65116 319372 65168 319378
rect 65116 319314 65168 319320
rect 65944 319372 65996 319378
rect 66416 319366 66536 319394
rect 65944 319314 65996 319320
rect 65956 316796 65984 319314
rect 66508 316810 66536 319366
rect 66600 316946 66628 327134
rect 66692 320058 66720 329838
rect 66864 327464 66916 327470
rect 66864 327406 66916 327412
rect 66772 326648 66824 326654
rect 66772 326590 66824 326596
rect 66680 320052 66732 320058
rect 66680 319994 66732 320000
rect 66784 319854 66812 326590
rect 66876 320602 66904 327406
rect 67520 327402 67548 329852
rect 67508 327396 67560 327402
rect 67508 327338 67560 327344
rect 68532 327334 68560 329852
rect 69360 329838 69650 329866
rect 69072 327396 69124 327402
rect 69072 327338 69124 327344
rect 68520 327328 68572 327334
rect 68520 327270 68572 327276
rect 68428 327260 68480 327266
rect 68428 327202 68480 327208
rect 66864 320596 66916 320602
rect 66864 320538 66916 320544
rect 68440 320398 68468 327202
rect 69084 320466 69112 327338
rect 69164 327056 69216 327062
rect 69164 326998 69216 327004
rect 69072 320460 69124 320466
rect 69072 320402 69124 320408
rect 68428 320392 68480 320398
rect 68428 320334 68480 320340
rect 66772 319848 66824 319854
rect 66772 319790 66824 319796
rect 68612 319848 68664 319854
rect 68612 319790 68664 319796
rect 66600 316918 67272 316946
rect 67244 316810 67272 316918
rect 66508 316782 66798 316810
rect 67244 316782 67718 316810
rect 68624 316796 68652 319790
rect 69176 319394 69204 326998
rect 69360 319990 69388 329838
rect 69440 327532 69492 327538
rect 69440 327474 69492 327480
rect 69348 319984 69400 319990
rect 69348 319926 69400 319932
rect 69452 319530 69480 327474
rect 70648 327470 70676 329852
rect 70636 327464 70688 327470
rect 70636 327406 70688 327412
rect 71660 327266 71688 329852
rect 72672 327402 72700 329852
rect 73408 329838 73790 329866
rect 72660 327396 72712 327402
rect 72660 327338 72712 327344
rect 71648 327260 71700 327266
rect 71648 327202 71700 327208
rect 73408 320126 73436 329838
rect 74316 326716 74368 326722
rect 74316 326658 74368 326664
rect 74040 326376 74092 326382
rect 74040 326318 74092 326324
rect 73396 320120 73448 320126
rect 73396 320062 73448 320068
rect 69452 319502 69940 319530
rect 69176 319366 69296 319394
rect 69268 316810 69296 319366
rect 69268 316782 69466 316810
rect 69912 316674 69940 319502
rect 69912 316646 70386 316674
rect 55088 315904 55140 315910
rect 55086 315872 55088 315881
rect 55140 315872 55142 315881
rect 55086 315807 55142 315816
rect 51590 313832 51646 313841
rect 51590 313767 51592 313776
rect 51644 313767 51646 313776
rect 51592 313738 51644 313744
rect 54074 310976 54130 310985
rect 54074 310911 54130 310920
rect 54088 310334 54116 310911
rect 54076 310328 54128 310334
rect 54076 310270 54128 310276
rect 55086 308120 55142 308129
rect 55086 308055 55142 308064
rect 54076 306248 54128 306254
rect 54074 306216 54076 306225
rect 54128 306216 54130 306225
rect 54074 306151 54130 306160
rect 51866 304312 51922 304321
rect 51866 304247 51922 304256
rect 51880 304214 51908 304247
rect 51868 304208 51920 304214
rect 51868 304150 51920 304156
rect 55100 300921 55128 308055
rect 73396 305432 73448 305438
rect 73396 305374 73448 305380
rect 73408 304729 73436 305374
rect 73394 304720 73450 304729
rect 73394 304655 73450 304664
rect 55086 300912 55142 300921
rect 55086 300847 55142 300856
rect 51682 299008 51738 299017
rect 51682 298943 51738 298952
rect 51696 298638 51724 298943
rect 51684 298632 51736 298638
rect 51684 298574 51736 298580
rect 51316 295164 51368 295170
rect 51316 295106 51368 295112
rect 51328 293962 51356 295106
rect 51236 293934 51356 293962
rect 51236 293690 51264 293934
rect 52602 293840 52658 293849
rect 52602 293775 52604 293784
rect 52656 293775 52658 293784
rect 52604 293746 52656 293752
rect 51236 293662 51356 293690
rect 50028 291696 50080 291702
rect 50028 291638 50080 291644
rect 50040 291294 50068 291638
rect 50028 291288 50080 291294
rect 50028 291230 50080 291236
rect 51328 289202 51356 293662
rect 54902 292072 54958 292081
rect 54902 292007 54958 292016
rect 51500 291288 51552 291294
rect 51500 291230 51552 291236
rect 51236 289174 51356 289202
rect 51236 288930 51264 289174
rect 51236 288902 51356 288930
rect 49936 285508 49988 285514
rect 49936 285450 49988 285456
rect 38068 280000 38120 280006
rect 38068 279942 38120 279948
rect 48556 280000 48608 280006
rect 48556 279942 48608 279948
rect 18102 279560 18158 279569
rect 18102 279495 18158 279504
rect 18116 279394 18144 279495
rect 18104 279388 18156 279394
rect 18104 279330 18156 279336
rect 38620 279320 38672 279326
rect 38620 279262 38672 279268
rect 38632 278209 38660 279262
rect 38618 278200 38674 278209
rect 38618 278135 38674 278144
rect 21244 273818 21272 276948
rect 23912 274498 23940 276948
rect 26580 274566 26608 276948
rect 29248 274634 29276 276948
rect 29236 274628 29288 274634
rect 29236 274570 29288 274576
rect 26568 274560 26620 274566
rect 26568 274502 26620 274508
rect 23900 274492 23952 274498
rect 23900 274434 23952 274440
rect 21232 273812 21284 273818
rect 21232 273754 21284 273760
rect 22244 273812 22296 273818
rect 22244 273754 22296 273760
rect 17552 251508 17604 251514
rect 17552 251450 17604 251456
rect 17460 240560 17512 240566
rect 17460 240502 17512 240508
rect 22256 229618 22284 273754
rect 31916 273750 31944 276948
rect 34584 274702 34612 276948
rect 34572 274696 34624 274702
rect 34572 274638 34624 274644
rect 47084 274696 47136 274702
rect 47084 274638 47136 274644
rect 46624 274628 46676 274634
rect 46624 274570 46676 274576
rect 46532 274560 46584 274566
rect 46532 274502 46584 274508
rect 46440 274492 46492 274498
rect 46440 274434 46492 274440
rect 31904 273744 31956 273750
rect 31904 273686 31956 273692
rect 31916 273070 31944 273686
rect 31904 273064 31956 273070
rect 31904 273006 31956 273012
rect 46452 249785 46480 274434
rect 46544 252913 46572 274502
rect 46636 256041 46664 274570
rect 46716 273064 46768 273070
rect 46716 273006 46768 273012
rect 46728 259169 46756 273006
rect 47096 262530 47124 274638
rect 48568 263634 48596 279942
rect 49948 263770 49976 285450
rect 51328 267902 51356 288902
rect 51512 287593 51540 291230
rect 54534 289284 54590 289293
rect 54534 289219 54590 289228
rect 54548 289050 54576 289219
rect 54916 289089 54944 292007
rect 74052 290177 74080 326318
rect 74222 314512 74278 314521
rect 74222 314447 74278 314456
rect 74130 311112 74186 311121
rect 74130 311047 74186 311056
rect 74038 290168 74094 290177
rect 74038 290103 74094 290112
rect 54902 289080 54958 289089
rect 54536 289044 54588 289050
rect 54902 289015 54958 289024
rect 54536 288986 54588 288992
rect 74038 288944 74094 288953
rect 74038 288879 74094 288888
rect 51498 287584 51554 287593
rect 51498 287519 51554 287528
rect 51682 287584 51738 287593
rect 51682 287519 51738 287528
rect 51696 277966 51724 287519
rect 52050 283912 52106 283921
rect 52050 283847 52106 283856
rect 52064 283474 52092 283847
rect 52052 283468 52104 283474
rect 52052 283410 52104 283416
rect 74052 279569 74080 288879
rect 74144 280686 74172 311047
rect 74236 297210 74264 314447
rect 74328 308265 74356 326658
rect 74788 320194 74816 329852
rect 74776 320188 74828 320194
rect 74776 320130 74828 320136
rect 74314 308256 74370 308265
rect 74314 308191 74370 308200
rect 75432 299969 75460 330058
rect 75524 305438 75552 330126
rect 75800 326314 75828 329852
rect 75788 326308 75840 326314
rect 75788 326250 75840 326256
rect 75512 305432 75564 305438
rect 75512 305374 75564 305380
rect 75418 299960 75474 299969
rect 75418 299895 75474 299904
rect 75432 298745 75460 299895
rect 75418 298736 75474 298745
rect 75418 298671 75474 298680
rect 74224 297204 74276 297210
rect 74224 297146 74276 297152
rect 74406 296288 74462 296297
rect 74406 296223 74462 296232
rect 74222 293568 74278 293577
rect 74222 293503 74278 293512
rect 74236 291673 74264 293503
rect 74222 291664 74278 291673
rect 74222 291599 74278 291608
rect 74420 289089 74448 296223
rect 75892 293577 75920 334342
rect 75984 334338 76012 334478
rect 75972 334332 76024 334338
rect 75972 334274 76024 334280
rect 75984 296297 76012 334274
rect 76076 327606 76104 334478
rect 76064 327600 76116 327606
rect 76064 327542 76116 327548
rect 76076 326382 76104 327542
rect 76064 326376 76116 326382
rect 76064 326318 76116 326324
rect 76156 312504 76208 312510
rect 76156 312446 76208 312452
rect 75970 296288 76026 296297
rect 75970 296223 76026 296232
rect 75878 293568 75934 293577
rect 75878 293503 75934 293512
rect 74406 289080 74462 289089
rect 74406 289015 74462 289024
rect 74314 288808 74370 288817
rect 74314 288743 74370 288752
rect 74132 280680 74184 280686
rect 74132 280622 74184 280628
rect 74328 279569 74356 288743
rect 74038 279560 74094 279569
rect 74038 279495 74094 279504
rect 74314 279560 74370 279569
rect 74314 279495 74370 279504
rect 52602 279424 52658 279433
rect 52602 279359 52658 279368
rect 52616 279326 52644 279359
rect 52604 279320 52656 279326
rect 52604 279262 52656 279268
rect 74038 278200 74094 278209
rect 74038 278135 74094 278144
rect 51500 277960 51552 277966
rect 51500 277902 51552 277908
rect 51684 277960 51736 277966
rect 51684 277902 51736 277908
rect 51512 272526 51540 277902
rect 55298 276934 55404 276962
rect 56126 276934 56784 276962
rect 51500 272520 51552 272526
rect 51500 272462 51552 272468
rect 51408 269732 51460 269738
rect 51408 269674 51460 269680
rect 51316 267896 51368 267902
rect 51316 267838 51368 267844
rect 49948 263742 50422 263770
rect 51420 263756 51448 269674
rect 52052 267896 52104 267902
rect 52052 267838 52104 267844
rect 52064 263770 52092 267838
rect 53522 266776 53578 266785
rect 53522 266711 53578 266720
rect 54534 266776 54590 266785
rect 54534 266711 54590 266720
rect 52064 263742 52446 263770
rect 53536 263756 53564 266711
rect 54548 263756 54576 266711
rect 55376 266406 55404 276934
rect 55546 266776 55602 266785
rect 55546 266711 55602 266720
rect 56558 266776 56614 266785
rect 56558 266711 56614 266720
rect 55364 266400 55416 266406
rect 55364 266342 55416 266348
rect 55560 263756 55588 266711
rect 56572 263756 56600 266711
rect 56756 266474 56784 276934
rect 57032 274498 57060 276948
rect 57966 276934 58164 276962
rect 58794 276934 59544 276962
rect 57020 274492 57072 274498
rect 57020 274434 57072 274440
rect 57664 266536 57716 266542
rect 57664 266478 57716 266484
rect 56744 266468 56796 266474
rect 56744 266410 56796 266416
rect 57676 263756 57704 266478
rect 58136 266338 58164 276934
rect 59516 266746 59544 276934
rect 59700 274702 59728 276948
rect 60634 276934 60832 276962
rect 59688 274696 59740 274702
rect 59688 274638 59740 274644
rect 60240 274016 60292 274022
rect 60240 273958 60292 273964
rect 59504 266740 59556 266746
rect 59504 266682 59556 266688
rect 60252 266542 60280 273958
rect 60240 266536 60292 266542
rect 60240 266478 60292 266484
rect 58124 266332 58176 266338
rect 58124 266274 58176 266280
rect 60804 266270 60832 276934
rect 60884 274696 60936 274702
rect 60884 274638 60936 274644
rect 60896 266678 60924 274638
rect 61448 273818 61476 276948
rect 62368 274634 62396 276948
rect 63092 274764 63144 274770
rect 63092 274706 63144 274712
rect 62356 274628 62408 274634
rect 62356 274570 62408 274576
rect 63000 273948 63052 273954
rect 63000 273890 63052 273896
rect 61620 273880 61672 273886
rect 61620 273822 61672 273828
rect 61436 273812 61488 273818
rect 61436 273754 61488 273760
rect 60884 266672 60936 266678
rect 60884 266614 60936 266620
rect 60792 266264 60844 266270
rect 60792 266206 60844 266212
rect 59688 265788 59740 265794
rect 59688 265730 59740 265736
rect 58676 265720 58728 265726
rect 58676 265662 58728 265668
rect 58688 263756 58716 265662
rect 59700 263756 59728 265730
rect 61632 265726 61660 273822
rect 62264 273812 62316 273818
rect 62264 273754 62316 273760
rect 62276 266610 62304 273754
rect 62264 266604 62316 266610
rect 62264 266546 62316 266552
rect 61804 265924 61856 265930
rect 61804 265866 61856 265872
rect 61620 265720 61672 265726
rect 61620 265662 61672 265668
rect 60700 265652 60752 265658
rect 60700 265594 60752 265600
rect 60712 263756 60740 265594
rect 61816 263756 61844 265866
rect 63012 265658 63040 273890
rect 63104 265794 63132 274706
rect 63288 274022 63316 276948
rect 63552 274628 63604 274634
rect 63552 274570 63604 274576
rect 63276 274016 63328 274022
rect 63276 273958 63328 273964
rect 63564 266202 63592 274570
rect 64116 273886 64144 276948
rect 65036 274770 65064 276948
rect 65024 274764 65076 274770
rect 65024 274706 65076 274712
rect 65024 274628 65076 274634
rect 65024 274570 65076 274576
rect 64104 273880 64156 273886
rect 64104 273822 64156 273828
rect 63644 273812 63696 273818
rect 63644 273754 63696 273760
rect 63552 266196 63604 266202
rect 63552 266138 63604 266144
rect 63092 265788 63144 265794
rect 63092 265730 63144 265736
rect 63000 265652 63052 265658
rect 63000 265594 63052 265600
rect 63656 265590 63684 273754
rect 64840 266808 64892 266814
rect 64840 266750 64892 266756
rect 62816 265584 62868 265590
rect 62816 265526 62868 265532
rect 63644 265584 63696 265590
rect 63644 265526 63696 265532
rect 63828 265584 63880 265590
rect 63828 265526 63880 265532
rect 62828 263756 62856 265526
rect 63840 263756 63868 265526
rect 64852 263756 64880 266750
rect 65036 265590 65064 274570
rect 65956 273954 65984 276948
rect 66600 276934 66798 276962
rect 65944 273948 65996 273954
rect 65944 273890 65996 273896
rect 66404 273880 66456 273886
rect 66404 273822 66456 273828
rect 65024 265584 65076 265590
rect 65024 265526 65076 265532
rect 66416 263770 66444 273822
rect 66600 265930 66628 276934
rect 67140 274492 67192 274498
rect 67140 274434 67192 274440
rect 66956 266400 67008 266406
rect 66956 266342 67008 266348
rect 66588 265924 66640 265930
rect 66588 265866 66640 265872
rect 65970 263742 66444 263770
rect 66968 263756 66996 266342
rect 67152 265590 67180 274434
rect 67704 273818 67732 276948
rect 68624 274634 68652 276948
rect 69360 276934 69466 276962
rect 68612 274628 68664 274634
rect 68612 274570 68664 274576
rect 67692 273812 67744 273818
rect 67692 273754 67744 273760
rect 69360 266814 69388 276934
rect 70372 273886 70400 276948
rect 70360 273880 70412 273886
rect 70360 273822 70412 273828
rect 69348 266808 69400 266814
rect 69348 266750 69400 266756
rect 71096 266740 71148 266746
rect 71096 266682 71148 266688
rect 67968 266468 68020 266474
rect 67968 266410 68020 266416
rect 67140 265584 67192 265590
rect 67140 265526 67192 265532
rect 67980 263756 68008 266410
rect 70084 266332 70136 266338
rect 70084 266274 70136 266280
rect 68980 265584 69032 265590
rect 68980 265526 69032 265532
rect 68992 263756 69020 265526
rect 70096 263756 70124 266274
rect 71108 263756 71136 266682
rect 72108 266672 72160 266678
rect 72108 266614 72160 266620
rect 72120 263756 72148 266614
rect 73120 266264 73172 266270
rect 73120 266206 73172 266212
rect 73132 263756 73160 266206
rect 48568 263606 49410 263634
rect 73854 263512 73910 263521
rect 74052 263482 74080 278135
rect 74224 266604 74276 266610
rect 74224 266546 74276 266552
rect 74236 263756 74264 266546
rect 75236 266196 75288 266202
rect 75236 266138 75288 266144
rect 75248 263756 75276 266138
rect 76168 263770 76196 312446
rect 76168 263742 76274 263770
rect 73854 263447 73856 263456
rect 73908 263447 73910 263456
rect 74040 263476 74092 263482
rect 73856 263418 73908 263424
rect 74040 263418 74092 263424
rect 49198 262560 49254 262569
rect 47084 262524 47136 262530
rect 49198 262495 49200 262504
rect 47084 262466 47136 262472
rect 49252 262495 49254 262504
rect 49200 262466 49252 262472
rect 46714 259160 46770 259169
rect 46714 259095 46770 259104
rect 46622 256032 46678 256041
rect 46622 255967 46678 255976
rect 46728 253026 46756 259095
rect 46728 252998 46848 253026
rect 46530 252904 46586 252913
rect 46530 252839 46586 252848
rect 46438 249776 46494 249785
rect 46438 249711 46494 249720
rect 46820 243506 46848 252998
rect 46820 243478 46940 243506
rect 46912 234446 46940 243478
rect 47082 237400 47138 237409
rect 47082 237335 47138 237344
rect 46900 234440 46952 234446
rect 46900 234382 46952 234388
rect 47096 230978 47124 237335
rect 48568 235862 49410 235890
rect 49948 235862 50422 235890
rect 51328 235862 51434 235890
rect 51512 235862 52446 235890
rect 47084 230972 47136 230978
rect 47084 230914 47136 230920
rect 22244 229612 22296 229618
rect 22244 229554 22296 229560
rect 47084 228388 47136 228394
rect 47084 228330 47136 228336
rect 34020 228320 34072 228326
rect 34020 228262 34072 228268
rect 34032 221730 34060 228262
rect 34572 226892 34624 226898
rect 34572 226834 34624 226840
rect 34584 221798 34612 226834
rect 34572 221792 34624 221798
rect 34572 221734 34624 221740
rect 34940 221792 34992 221798
rect 34940 221734 34992 221740
rect 34020 221724 34072 221730
rect 34020 221666 34072 221672
rect 34756 221724 34808 221730
rect 34756 221666 34808 221672
rect 34664 220568 34716 220574
rect 34664 220510 34716 220516
rect 17550 209656 17606 209665
rect 17550 209591 17606 209600
rect 17564 208985 17592 209591
rect 16538 208976 16594 208985
rect 16538 208911 16594 208920
rect 17550 208976 17606 208985
rect 17550 208911 17606 208920
rect 16448 208192 16500 208198
rect 16448 208134 16500 208140
rect 16446 204896 16502 204905
rect 16446 204831 16502 204840
rect 16460 132990 16488 204831
rect 16448 132984 16500 132990
rect 16448 132926 16500 132932
rect 16552 121974 16580 208911
rect 34676 206922 34704 220510
rect 34768 220506 34796 221666
rect 34952 220574 34980 221734
rect 34940 220568 34992 220574
rect 34940 220510 34992 220516
rect 34756 220500 34808 220506
rect 34756 220442 34808 220448
rect 38068 219956 38120 219962
rect 38068 219898 38120 219904
rect 38080 219457 38108 219898
rect 38066 219448 38122 219457
rect 38066 219383 38122 219392
rect 38528 217168 38580 217174
rect 38528 217110 38580 217116
rect 38540 216873 38568 217110
rect 38526 216864 38582 216873
rect 38526 216799 38582 216808
rect 38528 214448 38580 214454
rect 38528 214390 38580 214396
rect 38540 214289 38568 214390
rect 38526 214280 38582 214289
rect 38526 214215 38582 214224
rect 34848 213904 34900 213910
rect 34768 213852 34848 213858
rect 34768 213846 34900 213852
rect 34768 213830 34888 213846
rect 34768 211682 34796 213830
rect 34768 211654 34980 211682
rect 34676 206906 34888 206922
rect 34676 206900 34900 206906
rect 34676 206894 34848 206900
rect 34848 206842 34900 206848
rect 34848 204724 34900 204730
rect 34768 204684 34848 204712
rect 17642 199728 17698 199737
rect 17642 199663 17698 199672
rect 17656 199358 17684 199663
rect 17644 199352 17696 199358
rect 17644 199294 17696 199300
rect 34768 195226 34796 204684
rect 34848 204666 34900 204672
rect 34768 195198 34888 195226
rect 17090 189800 17146 189809
rect 17090 189735 17146 189744
rect 17104 189702 17132 189735
rect 17092 189696 17144 189702
rect 34860 189650 34888 195198
rect 17092 189638 17144 189644
rect 34768 189622 34888 189650
rect 34768 189242 34796 189622
rect 34676 189214 34796 189242
rect 34388 183236 34440 183242
rect 34388 183178 34440 183184
rect 21258 182958 21640 182986
rect 23926 182958 24216 182986
rect 26594 182958 26976 182986
rect 29262 182958 29552 182986
rect 21612 181338 21640 182958
rect 21600 181332 21652 181338
rect 21600 181274 21652 181280
rect 24188 180658 24216 182958
rect 26948 180726 26976 182958
rect 29524 180794 29552 182958
rect 31824 182822 31930 182850
rect 31824 180862 31852 182822
rect 34400 181338 34428 183178
rect 34676 183122 34704 189214
rect 34952 183242 34980 211654
rect 38710 211560 38766 211569
rect 38710 211495 38766 211504
rect 38724 210986 38752 211495
rect 38712 210980 38764 210986
rect 38712 210922 38764 210928
rect 38528 209620 38580 209626
rect 38528 209562 38580 209568
rect 38540 209257 38568 209562
rect 38526 209248 38582 209257
rect 38526 209183 38582 209192
rect 38528 206832 38580 206838
rect 38528 206774 38580 206780
rect 38540 206673 38568 206774
rect 38526 206664 38582 206673
rect 38526 206599 38582 206608
rect 38528 204792 38580 204798
rect 38528 204734 38580 204740
rect 38540 204497 38568 204734
rect 38526 204488 38582 204497
rect 38526 204423 38582 204432
rect 38526 201496 38582 201505
rect 38526 201431 38582 201440
rect 38540 201330 38568 201431
rect 38528 201324 38580 201330
rect 38528 201266 38580 201272
rect 38528 199284 38580 199290
rect 38528 199226 38580 199232
rect 38540 199193 38568 199226
rect 38526 199184 38582 199193
rect 38526 199119 38582 199128
rect 38526 196464 38582 196473
rect 38526 196399 38582 196408
rect 38540 195822 38568 196399
rect 38528 195816 38580 195822
rect 38528 195758 38580 195764
rect 38804 195136 38856 195142
rect 38804 195078 38856 195084
rect 38816 194569 38844 195078
rect 38802 194560 38858 194569
rect 38802 194495 38858 194504
rect 38804 191668 38856 191674
rect 38804 191610 38856 191616
rect 38816 191577 38844 191610
rect 38802 191568 38858 191577
rect 38802 191503 38858 191512
rect 38068 189628 38120 189634
rect 38068 189570 38120 189576
rect 38080 189265 38108 189570
rect 38066 189256 38122 189265
rect 38066 189191 38122 189200
rect 38066 186536 38122 186545
rect 38066 186471 38122 186480
rect 38080 186166 38108 186471
rect 38068 186160 38120 186166
rect 38068 186102 38120 186108
rect 38802 184088 38858 184097
rect 38802 184023 38804 184032
rect 38856 184023 38858 184032
rect 38804 183994 38856 184000
rect 34940 183236 34992 183242
rect 34940 183178 34992 183184
rect 34676 183094 34796 183122
rect 34598 182958 34704 182986
rect 34572 182692 34624 182698
rect 34572 182634 34624 182640
rect 34388 181332 34440 181338
rect 34388 181274 34440 181280
rect 31812 180856 31864 180862
rect 31812 180798 31864 180804
rect 34584 180810 34612 182634
rect 34676 180930 34704 182958
rect 34768 182698 34796 183094
rect 34756 182692 34808 182698
rect 34756 182634 34808 182640
rect 34664 180924 34716 180930
rect 34664 180866 34716 180872
rect 46992 180924 47044 180930
rect 46992 180866 47044 180872
rect 46716 180856 46768 180862
rect 29512 180788 29564 180794
rect 34584 180782 34704 180810
rect 46716 180798 46768 180804
rect 29512 180730 29564 180736
rect 26936 180720 26988 180726
rect 26936 180662 26988 180668
rect 24176 180652 24228 180658
rect 24176 180594 24228 180600
rect 16540 121968 16592 121974
rect 16540 121910 16592 121916
rect 16446 115136 16502 115145
rect 16446 115071 16502 115080
rect 16356 111564 16408 111570
rect 16356 111506 16408 111512
rect 16460 36362 16488 115071
rect 16538 111056 16594 111065
rect 16538 110991 16594 111000
rect 16552 47446 16580 110991
rect 18102 106296 18158 106305
rect 18102 106231 18158 106240
rect 18116 105518 18144 106231
rect 18104 105512 18156 105518
rect 18104 105454 18156 105460
rect 17458 101264 17514 101273
rect 17458 101199 17514 101208
rect 17472 99942 17500 101199
rect 17460 99936 17512 99942
rect 17460 99878 17512 99884
rect 18102 96232 18158 96241
rect 18102 96167 18158 96176
rect 18116 95862 18144 96167
rect 18104 95856 18156 95862
rect 18104 95798 18156 95804
rect 17274 91336 17330 91345
rect 17274 91271 17330 91280
rect 17288 90286 17316 91271
rect 17276 90280 17328 90286
rect 17276 90222 17328 90228
rect 21244 87158 21272 88860
rect 23912 87498 23940 88860
rect 23900 87492 23952 87498
rect 23900 87434 23952 87440
rect 26580 87430 26608 88860
rect 26568 87424 26620 87430
rect 26568 87366 26620 87372
rect 29248 87362 29276 88860
rect 29236 87356 29288 87362
rect 29236 87298 29288 87304
rect 31916 87294 31944 88860
rect 31904 87288 31956 87294
rect 31904 87230 31956 87236
rect 34584 87226 34612 88860
rect 34572 87220 34624 87226
rect 34572 87162 34624 87168
rect 34676 87158 34704 180782
rect 46624 180788 46676 180794
rect 46624 180730 46676 180736
rect 46532 180720 46584 180726
rect 46532 180662 46584 180668
rect 46440 180652 46492 180658
rect 46440 180594 46492 180600
rect 46452 155809 46480 180594
rect 46544 158937 46572 180662
rect 46636 162609 46664 180730
rect 46728 171682 46756 180798
rect 46716 171676 46768 171682
rect 46716 171618 46768 171624
rect 46900 171676 46952 171682
rect 46900 171618 46952 171624
rect 46912 165193 46940 171618
rect 47004 168894 47032 180866
rect 46992 168888 47044 168894
rect 46992 168830 47044 168836
rect 46898 165184 46954 165193
rect 46898 165119 46954 165128
rect 46622 162600 46678 162609
rect 46622 162535 46678 162544
rect 46530 158928 46586 158937
rect 46530 158863 46586 158872
rect 46438 155800 46494 155809
rect 46438 155735 46494 155744
rect 47096 143433 47124 228330
rect 48568 186166 48596 235862
rect 49948 191674 49976 235862
rect 51328 195822 51356 235862
rect 51406 210200 51462 210209
rect 51406 210135 51462 210144
rect 51420 209626 51448 210135
rect 51408 209620 51460 209626
rect 51408 209562 51460 209568
rect 51408 206832 51460 206838
rect 51406 206800 51408 206809
rect 51460 206800 51462 206809
rect 51406 206735 51462 206744
rect 51406 205304 51462 205313
rect 51406 205239 51462 205248
rect 51420 204798 51448 205239
rect 51408 204792 51460 204798
rect 51408 204734 51460 204740
rect 51512 201330 51540 235862
rect 53536 232513 53564 235876
rect 54548 232513 54576 235876
rect 55364 233216 55416 233222
rect 55364 233158 55416 233164
rect 53522 232504 53578 232513
rect 53522 232439 53578 232448
rect 54534 232504 54590 232513
rect 54534 232439 54590 232448
rect 55376 222834 55404 233158
rect 55560 229657 55588 235876
rect 56572 231017 56600 235876
rect 56744 233284 56796 233290
rect 56744 233226 56796 233232
rect 56558 231008 56614 231017
rect 56558 230943 56614 230952
rect 55546 229648 55602 229657
rect 55546 229583 55602 229592
rect 56756 225334 56784 233226
rect 57676 232610 57704 235876
rect 58124 233148 58176 233154
rect 58124 233090 58176 233096
rect 57664 232604 57716 232610
rect 57664 232546 57716 232552
rect 56100 225328 56152 225334
rect 56100 225270 56152 225276
rect 56744 225328 56796 225334
rect 56744 225270 56796 225276
rect 55298 222806 55404 222834
rect 56112 222820 56140 225270
rect 57020 224784 57072 224790
rect 57020 224726 57072 224732
rect 57032 222820 57060 224726
rect 58136 222834 58164 233090
rect 58688 232678 58716 235876
rect 59504 232876 59556 232882
rect 59504 232818 59556 232824
rect 58676 232672 58728 232678
rect 58676 232614 58728 232620
rect 59516 225062 59544 232818
rect 59700 232542 59728 235876
rect 59688 232536 59740 232542
rect 59688 232478 59740 232484
rect 60712 232474 60740 235876
rect 61816 233358 61844 235876
rect 62264 233692 62316 233698
rect 62264 233634 62316 233640
rect 61804 233352 61856 233358
rect 61804 233294 61856 233300
rect 60792 233080 60844 233086
rect 60792 233022 60844 233028
rect 60700 232468 60752 232474
rect 60700 232410 60752 232416
rect 60804 225334 60832 233022
rect 60884 232944 60936 232950
rect 60884 232886 60936 232892
rect 59688 225328 59740 225334
rect 59688 225270 59740 225276
rect 60792 225328 60844 225334
rect 60792 225270 60844 225276
rect 58768 225056 58820 225062
rect 58768 224998 58820 225004
rect 59504 225056 59556 225062
rect 59504 224998 59556 225004
rect 57966 222806 58164 222834
rect 58780 222820 58808 224998
rect 59700 222820 59728 225270
rect 60896 222834 60924 232886
rect 61620 232604 61672 232610
rect 61620 232546 61672 232552
rect 61436 225328 61488 225334
rect 61436 225270 61488 225276
rect 60634 222806 60924 222834
rect 61448 222820 61476 225270
rect 61632 225266 61660 232546
rect 62276 225334 62304 233634
rect 62828 233562 62856 235876
rect 62816 233556 62868 233562
rect 62816 233498 62868 233504
rect 63840 233426 63868 235876
rect 64852 233494 64880 235876
rect 65852 233556 65904 233562
rect 65852 233498 65904 233504
rect 64840 233488 64892 233494
rect 64840 233430 64892 233436
rect 63828 233420 63880 233426
rect 63828 233362 63880 233368
rect 65760 233352 65812 233358
rect 65760 233294 65812 233300
rect 63644 233216 63696 233222
rect 63644 233158 63696 233164
rect 63184 232672 63236 232678
rect 63184 232614 63236 232620
rect 63000 232536 63052 232542
rect 63000 232478 63052 232484
rect 62356 225396 62408 225402
rect 62356 225338 62408 225344
rect 62264 225328 62316 225334
rect 62264 225270 62316 225276
rect 61620 225260 61672 225266
rect 61620 225202 61672 225208
rect 62368 222820 62396 225338
rect 63012 224994 63040 232478
rect 63092 232468 63144 232474
rect 63092 232410 63144 232416
rect 63104 225130 63132 232410
rect 63196 225334 63224 232614
rect 63656 225402 63684 233158
rect 63644 225396 63696 225402
rect 63644 225338 63696 225344
rect 65772 225334 65800 233294
rect 63184 225328 63236 225334
rect 63184 225270 63236 225276
rect 64104 225328 64156 225334
rect 64104 225270 64156 225276
rect 65760 225328 65812 225334
rect 65760 225270 65812 225276
rect 63276 225260 63328 225266
rect 63276 225202 63328 225208
rect 63092 225124 63144 225130
rect 63092 225066 63144 225072
rect 63000 224988 63052 224994
rect 63000 224930 63052 224936
rect 63288 222820 63316 225202
rect 64116 222820 64144 225270
rect 65864 225266 65892 233498
rect 65956 232542 65984 235876
rect 66968 233630 66996 235876
rect 66956 233624 67008 233630
rect 66956 233566 67008 233572
rect 67232 233488 67284 233494
rect 67232 233430 67284 233436
rect 67140 233420 67192 233426
rect 67140 233362 67192 233368
rect 65944 232536 65996 232542
rect 65944 232478 65996 232484
rect 66772 225328 66824 225334
rect 66772 225270 66824 225276
rect 65852 225260 65904 225266
rect 65852 225202 65904 225208
rect 65944 225124 65996 225130
rect 65944 225066 65996 225072
rect 65024 224988 65076 224994
rect 65024 224930 65076 224936
rect 65036 222820 65064 224930
rect 65956 222820 65984 225066
rect 66784 222820 66812 225270
rect 67152 224314 67180 233362
rect 67244 224586 67272 233430
rect 67980 233290 68008 235876
rect 67968 233284 68020 233290
rect 67968 233226 68020 233232
rect 68520 232536 68572 232542
rect 68520 232478 68572 232484
rect 67324 232468 67376 232474
rect 67324 232410 67376 232416
rect 67336 224790 67364 232410
rect 68532 225334 68560 232478
rect 68992 232474 69020 235876
rect 70096 233154 70124 235876
rect 70084 233148 70136 233154
rect 70084 233090 70136 233096
rect 71108 232882 71136 235876
rect 72120 233086 72148 235876
rect 72108 233080 72160 233086
rect 72108 233022 72160 233028
rect 73132 232950 73160 235876
rect 73488 234440 73540 234446
rect 73488 234382 73540 234388
rect 73120 232944 73172 232950
rect 73120 232886 73172 232892
rect 71096 232876 71148 232882
rect 71096 232818 71148 232824
rect 68980 232468 69032 232474
rect 68980 232410 69032 232416
rect 68520 225328 68572 225334
rect 68520 225270 68572 225276
rect 70360 225328 70412 225334
rect 70360 225270 70412 225276
rect 67692 225260 67744 225266
rect 67692 225202 67744 225208
rect 67324 224784 67376 224790
rect 67324 224726 67376 224732
rect 67232 224580 67284 224586
rect 67232 224522 67284 224528
rect 67140 224308 67192 224314
rect 67140 224250 67192 224256
rect 67704 222820 67732 225202
rect 69440 224580 69492 224586
rect 69440 224522 69492 224528
rect 68612 224308 68664 224314
rect 68612 224250 68664 224256
rect 68624 222820 68652 224250
rect 69452 222820 69480 224522
rect 70372 222820 70400 225270
rect 53246 221352 53302 221361
rect 53246 221287 53302 221296
rect 51866 220264 51922 220273
rect 51866 220199 51922 220208
rect 51880 220030 51908 220199
rect 51868 220024 51920 220030
rect 51868 219966 51920 219972
rect 53260 217174 53288 221287
rect 53248 217168 53300 217174
rect 53248 217110 53300 217116
rect 51682 215232 51738 215241
rect 51682 215167 51738 215176
rect 51696 214522 51724 215167
rect 51684 214516 51736 214522
rect 51684 214458 51736 214464
rect 54074 211016 54130 211025
rect 54074 210951 54076 210960
rect 54128 210951 54130 210960
rect 54076 210922 54128 210928
rect 73500 210209 73528 234382
rect 74236 233698 74264 235876
rect 74682 235632 74738 235641
rect 74682 235567 74738 235576
rect 74406 235088 74462 235097
rect 74406 235023 74462 235032
rect 74420 234446 74448 235023
rect 74696 234961 74724 235567
rect 74682 234952 74738 234961
rect 74682 234887 74738 234896
rect 74408 234440 74460 234446
rect 74408 234382 74460 234388
rect 74224 233692 74276 233698
rect 74224 233634 74276 233640
rect 74132 233080 74184 233086
rect 74132 233022 74184 233028
rect 74040 228456 74092 228462
rect 74040 228398 74092 228404
rect 72658 210200 72714 210209
rect 72658 210135 72714 210144
rect 73486 210200 73542 210209
rect 73486 210135 73542 210144
rect 51500 201324 51552 201330
rect 51500 201266 51552 201272
rect 51316 195816 51368 195822
rect 51316 195758 51368 195764
rect 51328 195362 51356 195758
rect 51236 195334 51356 195362
rect 51236 194954 51264 195334
rect 51314 195240 51370 195249
rect 51314 195175 51370 195184
rect 51328 195142 51356 195175
rect 51316 195136 51368 195142
rect 51316 195078 51368 195084
rect 51236 194926 51356 194954
rect 49936 191668 49988 191674
rect 49936 191610 49988 191616
rect 48556 186160 48608 186166
rect 48556 186102 48608 186108
rect 48568 171834 48596 186102
rect 48568 171806 49240 171834
rect 49212 169794 49240 171806
rect 49948 169794 49976 191610
rect 51328 169794 51356 194926
rect 51406 185312 51462 185321
rect 51406 185247 51462 185256
rect 51420 184058 51448 185247
rect 51408 184052 51460 184058
rect 51408 183994 51460 184000
rect 51512 171018 51540 201266
rect 51774 200272 51830 200281
rect 51774 200207 51830 200216
rect 51788 199290 51816 200207
rect 51776 199284 51828 199290
rect 51776 199226 51828 199232
rect 51774 190208 51830 190217
rect 51774 190143 51830 190152
rect 51788 189634 51816 190143
rect 51776 189628 51828 189634
rect 51776 189570 51828 189576
rect 55298 182822 55404 182850
rect 56126 182822 56784 182850
rect 55376 172634 55404 182822
rect 55546 172936 55602 172945
rect 55546 172871 55602 172880
rect 55364 172628 55416 172634
rect 55364 172570 55416 172576
rect 53522 171712 53578 171721
rect 53522 171647 53578 171656
rect 54534 171712 54590 171721
rect 54534 171647 54590 171656
rect 51512 170990 52000 171018
rect 51972 169794 52000 170990
rect 49212 169766 49410 169794
rect 49948 169766 50422 169794
rect 51328 169766 51434 169794
rect 51972 169766 52446 169794
rect 53536 169780 53564 171647
rect 54548 169780 54576 171647
rect 55560 169780 55588 172871
rect 56558 172800 56614 172809
rect 56558 172735 56614 172744
rect 56572 169780 56600 172735
rect 56756 172566 56784 182822
rect 57032 180658 57060 182836
rect 57020 180652 57072 180658
rect 57020 180594 57072 180600
rect 57848 180040 57900 180046
rect 57848 179982 57900 179988
rect 57860 173042 57888 179982
rect 57848 173036 57900 173042
rect 57848 172978 57900 172984
rect 57952 172702 57980 182836
rect 58794 182822 59544 182850
rect 59412 181196 59464 181202
rect 59412 181138 59464 181144
rect 59424 173042 59452 181138
rect 58124 173036 58176 173042
rect 58124 172978 58176 172984
rect 58676 173036 58728 173042
rect 58676 172978 58728 172984
rect 59412 173036 59464 173042
rect 59412 172978 59464 172984
rect 57940 172696 57992 172702
rect 57940 172638 57992 172644
rect 56744 172560 56796 172566
rect 56744 172502 56796 172508
rect 58136 169658 58164 172978
rect 58688 169780 58716 172978
rect 59516 172838 59544 182822
rect 59700 181338 59728 182836
rect 60634 182822 60740 182850
rect 59688 181332 59740 181338
rect 59688 181274 59740 181280
rect 60608 180176 60660 180182
rect 60608 180118 60660 180124
rect 59688 173036 59740 173042
rect 59688 172978 59740 172984
rect 59504 172832 59556 172838
rect 59504 172774 59556 172780
rect 59700 169780 59728 172978
rect 60620 169794 60648 180118
rect 60712 172362 60740 182822
rect 61448 181338 61476 182836
rect 60884 181332 60936 181338
rect 60884 181274 60936 181280
rect 61436 181332 61488 181338
rect 61436 181274 61488 181280
rect 62172 181332 62224 181338
rect 62172 181274 62224 181280
rect 60792 181264 60844 181270
rect 60792 181206 60844 181212
rect 60804 173042 60832 181206
rect 60792 173036 60844 173042
rect 60792 172978 60844 172984
rect 60896 172770 60924 181274
rect 60884 172764 60936 172770
rect 60884 172706 60936 172712
rect 62184 172430 62212 181274
rect 62368 180930 62396 182836
rect 62356 180924 62408 180930
rect 62356 180866 62408 180872
rect 63288 180114 63316 182836
rect 64116 181202 64144 182836
rect 65036 181270 65064 182836
rect 65024 181264 65076 181270
rect 65024 181206 65076 181212
rect 64104 181196 64156 181202
rect 64104 181138 64156 181144
rect 63552 180924 63604 180930
rect 63552 180866 63604 180872
rect 63276 180108 63328 180114
rect 63276 180050 63328 180056
rect 62264 180040 62316 180046
rect 62264 179982 62316 179988
rect 62172 172424 62224 172430
rect 62172 172366 62224 172372
rect 60700 172356 60752 172362
rect 60700 172298 60752 172304
rect 60620 169766 60726 169794
rect 62276 169658 62304 179982
rect 62816 173036 62868 173042
rect 62816 172978 62868 172984
rect 62828 169780 62856 172978
rect 63564 172498 63592 180866
rect 64932 180856 64984 180862
rect 64932 180798 64984 180804
rect 63644 179972 63696 179978
rect 63644 179914 63696 179920
rect 63656 173042 63684 179914
rect 64944 173042 64972 180798
rect 65024 180788 65076 180794
rect 65024 180730 65076 180736
rect 63644 173036 63696 173042
rect 63644 172978 63696 172984
rect 63828 173036 63880 173042
rect 63828 172978 63880 172984
rect 64932 173036 64984 173042
rect 64932 172978 64984 172984
rect 63552 172492 63604 172498
rect 63552 172434 63604 172440
rect 63840 169780 63868 172978
rect 65036 169794 65064 180730
rect 65956 180182 65984 182836
rect 66404 180992 66456 180998
rect 66404 180934 66456 180940
rect 65944 180176 65996 180182
rect 65944 180118 65996 180124
rect 66416 169794 66444 180934
rect 66784 180046 66812 182836
rect 67140 180652 67192 180658
rect 67140 180594 67192 180600
rect 66772 180040 66824 180046
rect 66772 179982 66824 179988
rect 67152 173042 67180 180594
rect 67704 179978 67732 182836
rect 68624 180862 68652 182836
rect 68612 180856 68664 180862
rect 68612 180798 68664 180804
rect 69452 180794 69480 182836
rect 70372 180998 70400 182836
rect 70360 180992 70412 180998
rect 70360 180934 70412 180940
rect 69440 180788 69492 180794
rect 69440 180730 69492 180736
rect 67692 179972 67744 179978
rect 67692 179914 67744 179920
rect 67140 173036 67192 173042
rect 67140 172978 67192 172984
rect 68980 173036 69032 173042
rect 68980 172978 69032 172984
rect 66956 172628 67008 172634
rect 66956 172570 67008 172576
rect 64866 169766 65064 169794
rect 65970 169766 66444 169794
rect 66968 169780 66996 172570
rect 67968 172560 68020 172566
rect 67968 172502 68020 172508
rect 67980 169780 68008 172502
rect 68992 169780 69020 172978
rect 71096 172832 71148 172838
rect 71096 172774 71148 172780
rect 70084 172696 70136 172702
rect 70084 172638 70136 172644
rect 70096 169780 70124 172638
rect 71108 169780 71136 172774
rect 72108 172764 72160 172770
rect 72108 172706 72160 172712
rect 72120 169780 72148 172706
rect 72672 171682 72700 210135
rect 73762 206664 73818 206673
rect 73762 206599 73818 206608
rect 73776 199329 73804 206599
rect 73946 205032 74002 205041
rect 73946 204967 74002 204976
rect 73960 199329 73988 204967
rect 73762 199320 73818 199329
rect 73762 199255 73818 199264
rect 73946 199320 74002 199329
rect 73946 199255 74002 199264
rect 73762 189528 73818 189537
rect 73762 189463 73818 189472
rect 73776 180017 73804 189463
rect 74052 185185 74080 228398
rect 74144 203273 74172 233022
rect 74222 231008 74278 231017
rect 74222 230943 74278 230952
rect 74236 221497 74264 230943
rect 74222 221488 74278 221497
rect 74222 221423 74278 221432
rect 74314 220400 74370 220409
rect 74314 220335 74370 220344
rect 74224 214516 74276 214522
rect 74224 214458 74276 214464
rect 74236 213201 74264 214458
rect 74222 213192 74278 213201
rect 74222 213127 74278 213136
rect 74222 204488 74278 204497
rect 74222 204423 74278 204432
rect 74130 203264 74186 203273
rect 74130 203199 74186 203208
rect 74236 188041 74264 204423
rect 74328 203370 74356 220335
rect 74420 214522 74448 234382
rect 75142 234000 75198 234009
rect 75142 233935 75198 233944
rect 75156 233086 75184 233935
rect 75248 233358 75276 235876
rect 76168 235862 76274 235890
rect 75236 233352 75288 233358
rect 75236 233294 75288 233300
rect 75144 233080 75196 233086
rect 75144 233022 75196 233028
rect 76168 219554 76196 235862
rect 76812 230910 76840 359706
rect 76892 357452 76944 357458
rect 76892 357394 76944 357400
rect 76904 331754 76932 357394
rect 76996 334338 77024 359774
rect 80204 357928 80256 357934
rect 80204 357870 80256 357876
rect 80216 357633 80244 357870
rect 80202 357624 80258 357633
rect 80202 357559 80258 357568
rect 80204 356568 80256 356574
rect 80204 356510 80256 356516
rect 80216 356409 80244 356510
rect 80202 356400 80258 356409
rect 80202 356335 80258 356344
rect 80204 355208 80256 355214
rect 80204 355150 80256 355156
rect 79284 355140 79336 355146
rect 79284 355082 79336 355088
rect 79296 354641 79324 355082
rect 80216 355049 80244 355150
rect 80202 355040 80258 355049
rect 80202 354975 80258 354984
rect 79282 354632 79338 354641
rect 79282 354567 79338 354576
rect 80204 353848 80256 353854
rect 80204 353790 80256 353796
rect 80216 353417 80244 353790
rect 80202 353408 80258 353417
rect 80202 353343 80258 353352
rect 80204 352420 80256 352426
rect 80204 352362 80256 352368
rect 80216 352193 80244 352362
rect 80202 352184 80258 352193
rect 80202 352119 80258 352128
rect 87102 351368 87158 351377
rect 87102 351303 87158 351312
rect 79836 351060 79888 351066
rect 79836 351002 79888 351008
rect 79848 350425 79876 351002
rect 80202 350688 80258 350697
rect 80202 350623 80258 350632
rect 79834 350416 79890 350425
rect 80216 350386 80244 350623
rect 87010 350416 87066 350425
rect 79834 350351 79890 350360
rect 80204 350380 80256 350386
rect 87010 350351 87066 350360
rect 80204 350322 80256 350328
rect 86918 349600 86974 349609
rect 86918 349535 86974 349544
rect 78914 349056 78970 349065
rect 78914 348991 78970 349000
rect 78928 348958 78956 348991
rect 78916 348952 78968 348958
rect 78916 348894 78968 348900
rect 78914 347560 78970 347569
rect 78914 347495 78970 347504
rect 78928 347394 78956 347495
rect 78916 347388 78968 347394
rect 78916 347330 78968 347336
rect 79006 346472 79062 346481
rect 79006 346407 79062 346416
rect 78916 346232 78968 346238
rect 78916 346174 78968 346180
rect 78928 346073 78956 346174
rect 78914 346064 78970 346073
rect 79020 346034 79048 346407
rect 86932 346034 86960 349535
rect 87024 347394 87052 350351
rect 87116 348958 87144 351303
rect 87104 348952 87156 348958
rect 87104 348894 87156 348900
rect 87102 348648 87158 348657
rect 87102 348583 87158 348592
rect 87012 347388 87064 347394
rect 87012 347330 87064 347336
rect 87010 347288 87066 347297
rect 87010 347223 87066 347232
rect 78914 345999 78970 346008
rect 79008 346028 79060 346034
rect 79008 345970 79060 345976
rect 86920 346028 86972 346034
rect 86920 345970 86972 345976
rect 85816 345620 85868 345626
rect 85816 345562 85868 345568
rect 78914 344568 78970 344577
rect 78914 344503 78970 344512
rect 78928 344470 78956 344503
rect 78916 344464 78968 344470
rect 78916 344406 78968 344412
rect 78914 343344 78970 343353
rect 78914 343279 78970 343288
rect 78928 342974 78956 343279
rect 85828 342974 85856 345562
rect 85908 344668 85960 344674
rect 85908 344610 85960 344616
rect 78916 342968 78968 342974
rect 78916 342910 78968 342916
rect 85816 342968 85868 342974
rect 85816 342910 85868 342916
rect 78914 342800 78970 342809
rect 78914 342735 78916 342744
rect 78968 342735 78970 342744
rect 78916 342706 78968 342712
rect 78914 341712 78970 341721
rect 78914 341647 78970 341656
rect 78928 341546 78956 341647
rect 85920 341546 85948 344610
rect 87024 344470 87052 347223
rect 87116 346238 87144 348583
rect 87104 346232 87156 346238
rect 87104 346174 87156 346180
rect 87012 344464 87064 344470
rect 87012 344406 87064 344412
rect 78916 341540 78968 341546
rect 78916 341482 78968 341488
rect 85908 341540 85960 341546
rect 85908 341482 85960 341488
rect 78916 341404 78968 341410
rect 78916 341346 78968 341352
rect 78928 341041 78956 341346
rect 78914 341032 78970 341041
rect 78914 340967 78970 340976
rect 85724 340112 85776 340118
rect 85724 340054 85776 340060
rect 78916 340044 78968 340050
rect 78916 339986 78968 339992
rect 78928 339817 78956 339986
rect 78914 339808 78970 339817
rect 78914 339743 78970 339752
rect 84988 338684 85040 338690
rect 84988 338626 85040 338632
rect 80204 338616 80256 338622
rect 80204 338558 80256 338564
rect 78916 338548 78968 338554
rect 78916 338490 78968 338496
rect 78928 338049 78956 338490
rect 80216 338457 80244 338558
rect 80202 338448 80258 338457
rect 80202 338383 80258 338392
rect 78914 338040 78970 338049
rect 78914 337975 78970 337984
rect 80202 336272 80258 336281
rect 80202 336207 80258 336216
rect 80216 336106 80244 336207
rect 80204 336100 80256 336106
rect 80204 336042 80256 336048
rect 80202 335320 80258 335329
rect 80202 335255 80258 335264
rect 80216 335154 80244 335255
rect 85000 335154 85028 338626
rect 85736 336106 85764 340054
rect 85724 336100 85776 336106
rect 85724 336042 85776 336048
rect 85816 335964 85868 335970
rect 85816 335906 85868 335912
rect 80204 335148 80256 335154
rect 80204 335090 80256 335096
rect 84988 335148 85040 335154
rect 84988 335090 85040 335096
rect 76984 334332 77036 334338
rect 76984 334274 77036 334280
rect 80204 334264 80256 334270
rect 80202 334232 80204 334241
rect 80256 334232 80258 334241
rect 78916 334196 78968 334202
rect 80202 334167 80258 334176
rect 78916 334138 78968 334144
rect 78928 333697 78956 334138
rect 78914 333688 78970 333697
rect 78914 333623 78970 333632
rect 80204 333108 80256 333114
rect 80204 333050 80256 333056
rect 80216 332745 80244 333050
rect 80202 332736 80258 332745
rect 80202 332671 80258 332680
rect 76892 331748 76944 331754
rect 76892 331690 76944 331696
rect 76904 326722 76932 331690
rect 80202 330968 80258 330977
rect 80202 330903 80258 330912
rect 80216 330666 80244 330903
rect 85828 330666 85856 335906
rect 80204 330660 80256 330666
rect 80204 330602 80256 330608
rect 85816 330660 85868 330666
rect 85816 330602 85868 330608
rect 78914 329744 78970 329753
rect 78914 329679 78970 329688
rect 78928 329034 78956 329679
rect 78916 329028 78968 329034
rect 78916 328970 78968 328976
rect 76892 326716 76944 326722
rect 76892 326658 76944 326664
rect 76984 326308 77036 326314
rect 76984 326250 77036 326256
rect 76996 313598 77024 326250
rect 76984 313592 77036 313598
rect 81676 313592 81728 313598
rect 76984 313534 77036 313540
rect 81674 313560 81676 313569
rect 81728 313560 81730 313569
rect 76996 312510 77024 313534
rect 81674 313495 81730 313504
rect 76984 312504 77036 312510
rect 76984 312446 77036 312452
rect 81676 297204 81728 297210
rect 81676 297146 81728 297152
rect 81688 296841 81716 297146
rect 81674 296832 81730 296841
rect 81674 296767 81730 296776
rect 84618 285000 84674 285009
rect 84618 284935 84674 284944
rect 84526 284592 84582 284601
rect 84526 284527 84582 284536
rect 84540 281201 84568 284527
rect 84632 281881 84660 284935
rect 84618 281872 84674 281881
rect 84618 281807 84674 281816
rect 84526 281192 84582 281201
rect 84526 281127 84582 281136
rect 81676 280680 81728 280686
rect 81676 280622 81728 280628
rect 81688 280249 81716 280622
rect 81674 280240 81730 280249
rect 81674 280175 81730 280184
rect 87208 271930 87236 391054
rect 108920 389486 108948 393094
rect 108908 389480 108960 389486
rect 108908 389422 108960 389428
rect 111300 389480 111352 389486
rect 111300 389422 111352 389428
rect 91336 388732 91388 388738
rect 91336 388674 91388 388680
rect 91348 386700 91376 388674
rect 96304 388664 96356 388670
rect 96304 388606 96356 388612
rect 96316 386700 96344 388606
rect 106332 388596 106384 388602
rect 106332 388538 106384 388544
rect 101272 388392 101324 388398
rect 101272 388334 101324 388340
rect 101284 386700 101312 388334
rect 106344 386700 106372 388538
rect 111312 386700 111340 389422
rect 116268 389140 116320 389146
rect 116268 389082 116320 389088
rect 116280 386700 116308 389082
rect 121328 389072 121380 389078
rect 121328 389014 121380 389020
rect 121340 386700 121368 389014
rect 128608 389010 128636 393774
rect 154828 389078 154856 393774
rect 182428 389146 182456 396206
rect 208648 389214 208676 396206
rect 235696 393838 235724 396344
rect 262192 393838 262220 396344
rect 234856 393832 234908 393838
rect 234856 393774 234908 393780
rect 235684 393832 235736 393838
rect 235684 393774 235736 393780
rect 261076 393832 261128 393838
rect 261076 393774 261128 393780
rect 262180 393832 262232 393838
rect 262180 393774 262232 393780
rect 195296 389208 195348 389214
rect 195296 389150 195348 389156
rect 208636 389208 208688 389214
rect 208636 389150 208688 389156
rect 182416 389140 182468 389146
rect 182416 389082 182468 389088
rect 154816 389072 154868 389078
rect 154816 389014 154868 389020
rect 126296 389004 126348 389010
rect 126296 388946 126348 388952
rect 128596 389004 128648 389010
rect 128596 388946 128648 388952
rect 126308 386700 126336 388946
rect 185360 388528 185412 388534
rect 185360 388470 185412 388476
rect 190328 388528 190380 388534
rect 190328 388470 190380 388476
rect 185372 386700 185400 388470
rect 190340 386700 190368 388470
rect 195308 386700 195336 389150
rect 200356 389140 200408 389146
rect 200356 389082 200408 389088
rect 200368 386700 200396 389082
rect 205324 389072 205376 389078
rect 205324 389014 205376 389020
rect 205336 386700 205364 389014
rect 234868 389010 234896 393774
rect 261088 389078 261116 393774
rect 279660 393220 279712 393226
rect 279660 393162 279712 393168
rect 261076 389072 261128 389078
rect 261076 389014 261128 389020
rect 210292 389004 210344 389010
rect 210292 388946 210344 388952
rect 234856 389004 234908 389010
rect 234856 388946 234908 388952
rect 210304 386700 210332 388946
rect 223080 388528 223132 388534
rect 223080 388470 223132 388476
rect 215352 388460 215404 388466
rect 215352 388402 215404 388408
rect 220320 388460 220372 388466
rect 220320 388402 220372 388408
rect 215364 386700 215392 388402
rect 220332 386700 220360 388402
rect 131354 384824 131410 384833
rect 131354 384759 131410 384768
rect 89864 367720 89916 367726
rect 89864 367662 89916 367668
rect 89876 351066 89904 367662
rect 90060 367658 90088 370924
rect 92544 367726 92572 370924
rect 95042 370910 95424 370938
rect 92532 367720 92584 367726
rect 92532 367662 92584 367668
rect 90048 367652 90100 367658
rect 90048 367594 90100 367600
rect 91336 367652 91388 367658
rect 91336 367594 91388 367600
rect 91348 363510 91376 367594
rect 91336 363504 91388 363510
rect 91336 363446 91388 363452
rect 92072 363504 92124 363510
rect 92072 363446 92124 363452
rect 92084 351762 92112 363446
rect 95396 355078 95424 370910
rect 96868 370910 97526 370938
rect 96868 355321 96896 370910
rect 99996 367658 100024 370924
rect 102388 370910 102494 370938
rect 99984 367652 100036 367658
rect 99984 367594 100036 367600
rect 100904 367652 100956 367658
rect 100904 367594 100956 367600
rect 96854 355312 96910 355321
rect 96854 355247 96910 355256
rect 100916 355078 100944 367594
rect 102388 358834 102416 370910
rect 102388 358806 102692 358834
rect 95384 355072 95436 355078
rect 95384 355014 95436 355020
rect 97040 355072 97092 355078
rect 97040 355014 97092 355020
rect 100904 355072 100956 355078
rect 100904 355014 100956 355020
rect 102376 355072 102428 355078
rect 102376 355014 102428 355020
rect 97052 351762 97080 355014
rect 102388 351762 102416 355014
rect 102664 352426 102692 358806
rect 105056 355146 105084 370924
rect 106528 370910 107554 370938
rect 105044 355140 105096 355146
rect 105044 355082 105096 355088
rect 106528 353854 106556 370910
rect 110024 367658 110052 370924
rect 112140 370910 112522 370938
rect 110012 367652 110064 367658
rect 110012 367594 110064 367600
rect 112036 367652 112088 367658
rect 112036 367594 112088 367600
rect 107068 355140 107120 355146
rect 107068 355082 107120 355088
rect 106516 353848 106568 353854
rect 106516 353790 106568 353796
rect 102652 352420 102704 352426
rect 102652 352362 102704 352368
rect 92084 351734 92420 351762
rect 97052 351734 97388 351762
rect 102356 351734 102416 351762
rect 107080 351762 107108 355082
rect 112048 351762 112076 367594
rect 112140 354942 112168 370910
rect 114992 367658 115020 370924
rect 114980 367652 115032 367658
rect 114980 367594 115032 367600
rect 116176 367652 116228 367658
rect 116176 367594 116228 367600
rect 116188 363510 116216 367594
rect 116176 363504 116228 363510
rect 116176 363446 116228 363452
rect 116820 363504 116872 363510
rect 116820 363446 116872 363452
rect 116832 363322 116860 363446
rect 116832 363294 116952 363322
rect 112128 354936 112180 354942
rect 112128 354878 112180 354884
rect 116924 351762 116952 363294
rect 117568 355214 117596 370924
rect 120066 370910 120264 370938
rect 120236 355214 120264 370910
rect 121708 370910 122550 370938
rect 121708 356574 121736 370910
rect 125020 367658 125048 370924
rect 127228 370910 127518 370938
rect 125008 367652 125060 367658
rect 125008 367594 125060 367600
rect 126480 367652 126532 367658
rect 126480 367594 126532 367600
rect 121696 356568 121748 356574
rect 121696 356510 121748 356516
rect 117556 355208 117608 355214
rect 117556 355150 117608 355156
rect 118016 355208 118068 355214
rect 118016 355150 118068 355156
rect 120224 355208 120276 355214
rect 120224 355150 120276 355156
rect 122064 355208 122116 355214
rect 122064 355150 122116 355156
rect 118028 355010 118056 355150
rect 118016 355004 118068 355010
rect 118016 354946 118068 354952
rect 122076 351762 122104 355150
rect 126492 355078 126520 367594
rect 127228 357934 127256 370910
rect 127216 357928 127268 357934
rect 127216 357870 127268 357876
rect 126480 355072 126532 355078
rect 126480 355014 126532 355020
rect 127216 355072 127268 355078
rect 127216 355014 127268 355020
rect 127228 351762 127256 355014
rect 107080 351734 107416 351762
rect 112048 351734 112384 351762
rect 116924 351734 117352 351762
rect 122076 351734 122412 351762
rect 127228 351734 127380 351762
rect 96762 351640 96818 351649
rect 96762 351575 96818 351584
rect 96776 351542 96804 351575
rect 96764 351536 96816 351542
rect 96764 351478 96816 351484
rect 89864 351060 89916 351066
rect 89864 351002 89916 351008
rect 87930 346880 87986 346889
rect 87930 346815 87986 346824
rect 87944 345626 87972 346815
rect 88114 346064 88170 346073
rect 88114 345999 88170 346008
rect 87932 345620 87984 345626
rect 87932 345562 87984 345568
rect 87470 345112 87526 345121
rect 87470 345047 87526 345056
rect 87484 344674 87512 345047
rect 87472 344668 87524 344674
rect 87472 344610 87524 344616
rect 87378 343344 87434 343353
rect 87378 343279 87434 343288
rect 87286 341576 87342 341585
rect 87286 341511 87342 341520
rect 87300 338554 87328 341511
rect 87392 340050 87420 343279
rect 88128 342770 88156 345999
rect 88482 344296 88538 344305
rect 88482 344231 88538 344240
rect 88116 342764 88168 342770
rect 88116 342706 88168 342712
rect 87470 342392 87526 342401
rect 87470 342327 87526 342336
rect 87380 340044 87432 340050
rect 87380 339986 87432 339992
rect 87378 339808 87434 339817
rect 87378 339743 87434 339752
rect 87392 338690 87420 339743
rect 87380 338684 87432 338690
rect 87380 338626 87432 338632
rect 87484 338622 87512 342327
rect 88496 341410 88524 344231
rect 88484 341404 88536 341410
rect 88484 341346 88536 341352
rect 87562 340624 87618 340633
rect 87562 340559 87618 340568
rect 87576 340118 87604 340559
rect 87564 340112 87616 340118
rect 87564 340054 87616 340060
rect 87930 338856 87986 338865
rect 87930 338791 87986 338800
rect 87472 338616 87524 338622
rect 87472 338558 87524 338564
rect 87288 338548 87340 338554
rect 87288 338490 87340 338496
rect 87378 337088 87434 337097
rect 87378 337023 87434 337032
rect 87392 333114 87420 337023
rect 87838 336272 87894 336281
rect 87838 336207 87894 336216
rect 87852 335970 87880 336207
rect 87840 335964 87892 335970
rect 87840 335906 87892 335912
rect 87944 335850 87972 338791
rect 88022 338040 88078 338049
rect 88022 337975 88078 337984
rect 87852 335822 87972 335850
rect 87852 334270 87880 335822
rect 87840 334264 87892 334270
rect 87840 334206 87892 334212
rect 88036 334202 88064 337975
rect 91592 335822 91928 335850
rect 94904 335822 95240 335850
rect 98216 335822 98276 335850
rect 88024 334196 88076 334202
rect 88024 334138 88076 334144
rect 91244 333924 91296 333930
rect 91244 333866 91296 333872
rect 87380 333108 87432 333114
rect 87380 333050 87432 333056
rect 91256 321706 91284 333866
rect 91900 333794 91928 335822
rect 95212 333833 95240 335822
rect 98248 334338 98276 335822
rect 101008 335822 101528 335850
rect 104872 335822 104932 335850
rect 108244 335822 108304 335850
rect 98236 334332 98288 334338
rect 98236 334274 98288 334280
rect 98248 333862 98276 334274
rect 98236 333856 98288 333862
rect 95198 333824 95254 333833
rect 91888 333788 91940 333794
rect 98236 333798 98288 333804
rect 95198 333759 95254 333768
rect 91888 333730 91940 333736
rect 101008 327606 101036 335822
rect 104872 334406 104900 335822
rect 108276 334474 108304 335822
rect 111404 335822 111556 335850
rect 114808 335822 114868 335850
rect 118212 335822 118272 335850
rect 121248 335822 121584 335850
rect 124560 335822 124896 335850
rect 127872 335822 128208 335850
rect 108264 334468 108316 334474
rect 108264 334410 108316 334416
rect 104860 334400 104912 334406
rect 104860 334342 104912 334348
rect 111404 334338 111432 335822
rect 111392 334332 111444 334338
rect 111392 334274 111444 334280
rect 103664 333992 103716 333998
rect 103664 333934 103716 333940
rect 100996 327600 101048 327606
rect 100996 327542 101048 327548
rect 101008 326926 101036 327542
rect 100996 326920 101048 326926
rect 100996 326862 101048 326868
rect 103676 321706 103704 333934
rect 111404 331618 111432 334274
rect 114808 334270 114836 335822
rect 114796 334264 114848 334270
rect 114796 334206 114848 334212
rect 114808 331686 114836 334206
rect 118212 334202 118240 335822
rect 118200 334196 118252 334202
rect 118200 334138 118252 334144
rect 116084 334060 116136 334066
rect 116084 334002 116136 334008
rect 114796 331680 114848 331686
rect 114796 331622 114848 331628
rect 111392 331612 111444 331618
rect 111392 331554 111444 331560
rect 116096 321706 116124 334002
rect 118212 331754 118240 334138
rect 121248 333930 121276 335822
rect 124560 333998 124588 335822
rect 127872 334066 127900 335822
rect 131368 334202 131396 384759
rect 131446 382104 131502 382113
rect 131446 382039 131502 382048
rect 131460 334270 131488 382039
rect 131538 380200 131594 380209
rect 131538 380135 131594 380144
rect 131552 334338 131580 380135
rect 131630 377480 131686 377489
rect 131630 377415 131686 377424
rect 131644 334474 131672 377415
rect 131722 374760 131778 374769
rect 131722 374695 131778 374704
rect 131632 334468 131684 334474
rect 131632 334410 131684 334416
rect 131540 334332 131592 334338
rect 131540 334274 131592 334280
rect 131448 334264 131500 334270
rect 131448 334206 131500 334212
rect 131356 334196 131408 334202
rect 131356 334138 131408 334144
rect 127860 334060 127912 334066
rect 127860 334002 127912 334008
rect 131460 333998 131488 334206
rect 131552 334134 131580 334274
rect 131644 334202 131672 334410
rect 131736 334406 131764 374695
rect 131814 372176 131870 372185
rect 131814 372111 131870 372120
rect 131828 371806 131856 372111
rect 131816 371800 131868 371806
rect 131816 371742 131868 371748
rect 134760 371800 134812 371806
rect 134760 371742 134812 371748
rect 131814 351368 131870 351377
rect 131814 351303 131870 351312
rect 131828 351134 131856 351303
rect 131816 351128 131868 351134
rect 131816 351070 131868 351076
rect 131814 350416 131870 350425
rect 131814 350351 131870 350360
rect 131828 349774 131856 350351
rect 131816 349768 131868 349774
rect 131816 349710 131868 349716
rect 131906 349600 131962 349609
rect 131906 349535 131962 349544
rect 131814 348648 131870 348657
rect 131814 348583 131870 348592
rect 131828 348414 131856 348583
rect 131816 348408 131868 348414
rect 131816 348350 131868 348356
rect 131920 348346 131948 349535
rect 131908 348340 131960 348346
rect 131908 348282 131960 348288
rect 132182 347832 132238 347841
rect 132182 347767 132238 347776
rect 132196 346986 132224 347767
rect 132184 346980 132236 346986
rect 132184 346922 132236 346928
rect 131906 346880 131962 346889
rect 131906 346815 131962 346824
rect 131814 346064 131870 346073
rect 131814 345999 131870 346008
rect 131828 345694 131856 345999
rect 131816 345688 131868 345694
rect 131816 345630 131868 345636
rect 131920 345626 131948 346815
rect 134116 345688 134168 345694
rect 134116 345630 134168 345636
rect 131908 345620 131960 345626
rect 131908 345562 131960 345568
rect 132366 345112 132422 345121
rect 132366 345047 132422 345056
rect 131814 344296 131870 344305
rect 131814 344231 131816 344240
rect 131868 344231 131870 344240
rect 131816 344202 131868 344208
rect 132380 344198 132408 345047
rect 132368 344192 132420 344198
rect 132368 344134 132420 344140
rect 131814 343344 131870 343353
rect 131814 343279 131870 343288
rect 131828 342838 131856 343279
rect 131816 342832 131868 342838
rect 131816 342774 131868 342780
rect 134128 342770 134156 345630
rect 134116 342764 134168 342770
rect 134116 342706 134168 342712
rect 131906 342392 131962 342401
rect 131906 342327 131962 342336
rect 131814 341576 131870 341585
rect 131920 341546 131948 342327
rect 131814 341511 131870 341520
rect 131908 341540 131960 341546
rect 131828 341478 131856 341511
rect 131908 341482 131960 341488
rect 131816 341472 131868 341478
rect 131816 341414 131868 341420
rect 131814 340624 131870 340633
rect 131814 340559 131870 340568
rect 131828 340118 131856 340559
rect 131816 340112 131868 340118
rect 131816 340054 131868 340060
rect 131906 339808 131962 339817
rect 131906 339743 131962 339752
rect 131814 338856 131870 338865
rect 131814 338791 131870 338800
rect 131828 338758 131856 338791
rect 131816 338752 131868 338758
rect 131816 338694 131868 338700
rect 131920 338690 131948 339743
rect 131908 338684 131960 338690
rect 131908 338626 131960 338632
rect 131814 338040 131870 338049
rect 131814 337975 131870 337984
rect 131828 337330 131856 337975
rect 131816 337324 131868 337330
rect 131816 337266 131868 337272
rect 131906 337088 131962 337097
rect 131906 337023 131962 337032
rect 131814 336272 131870 336281
rect 131814 336207 131870 336216
rect 131828 335970 131856 336207
rect 131920 336038 131948 337023
rect 131908 336032 131960 336038
rect 131908 335974 131960 335980
rect 131816 335964 131868 335970
rect 131816 335906 131868 335912
rect 131724 334400 131776 334406
rect 131724 334342 131776 334348
rect 131632 334196 131684 334202
rect 131632 334138 131684 334144
rect 131540 334128 131592 334134
rect 131540 334070 131592 334076
rect 124548 333992 124600 333998
rect 124548 333934 124600 333940
rect 131448 333992 131500 333998
rect 131448 333934 131500 333940
rect 131736 333930 131764 334342
rect 121236 333924 121288 333930
rect 121236 333866 121288 333872
rect 131724 333924 131776 333930
rect 131724 333866 131776 333872
rect 118200 331748 118252 331754
rect 118200 331690 118252 331696
rect 128504 329028 128556 329034
rect 128504 328970 128556 328976
rect 91086 321678 91284 321706
rect 103506 321678 103704 321706
rect 116018 321678 116124 321706
rect 128516 321692 128544 328970
rect 87208 271916 88418 271930
rect 87208 271902 88432 271916
rect 88404 269670 88432 271902
rect 88392 269664 88444 269670
rect 88392 269606 88444 269612
rect 95488 268990 95516 271916
rect 102664 269602 102692 271916
rect 102652 269596 102704 269602
rect 102652 269538 102704 269544
rect 109748 269058 109776 271916
rect 95568 269052 95620 269058
rect 95568 268994 95620 269000
rect 109736 269052 109788 269058
rect 109736 268994 109788 269000
rect 95476 268984 95528 268990
rect 95476 268926 95528 268932
rect 77260 264088 77312 264094
rect 77260 264030 77312 264036
rect 77272 263181 77300 264030
rect 77258 263172 77314 263181
rect 77258 263107 77314 263116
rect 79742 261744 79798 261753
rect 79742 261679 79798 261688
rect 79756 261442 79784 261679
rect 79744 261436 79796 261442
rect 79744 261378 79796 261384
rect 87196 261436 87248 261442
rect 87196 261378 87248 261384
rect 79742 260384 79798 260393
rect 79742 260319 79798 260328
rect 79756 260082 79784 260319
rect 79744 260076 79796 260082
rect 79744 260018 79796 260024
rect 85080 260076 85132 260082
rect 85080 260018 85132 260024
rect 79742 258888 79798 258897
rect 79742 258823 79798 258832
rect 79756 258722 79784 258823
rect 79744 258716 79796 258722
rect 79744 258658 79796 258664
rect 84436 258716 84488 258722
rect 84436 258658 84488 258664
rect 80294 257528 80350 257537
rect 80294 257463 80350 257472
rect 79742 256168 79798 256177
rect 79742 256103 79798 256112
rect 79756 255934 79784 256103
rect 79744 255928 79796 255934
rect 79744 255870 79796 255876
rect 80308 255866 80336 257463
rect 80296 255860 80348 255866
rect 80296 255802 80348 255808
rect 84448 255798 84476 258658
rect 85092 256886 85120 260018
rect 87208 258081 87236 261378
rect 95580 261374 95608 268994
rect 116924 268582 116952 271916
rect 124008 271794 124036 271916
rect 123272 271766 124036 271794
rect 114796 268576 114848 268582
rect 114796 268518 114848 268524
rect 116912 268576 116964 268582
rect 116912 268518 116964 268524
rect 95568 261368 95620 261374
rect 95568 261310 95620 261316
rect 96212 261368 96264 261374
rect 96212 261310 96264 261316
rect 87194 258072 87250 258081
rect 87194 258007 87250 258016
rect 96224 257786 96252 261310
rect 114808 260490 114836 268518
rect 123272 264094 123300 271766
rect 131184 269398 131212 271916
rect 127768 269392 127820 269398
rect 127768 269334 127820 269340
rect 131172 269392 131224 269398
rect 131172 269334 131224 269340
rect 123260 264088 123312 264094
rect 123260 264030 123312 264036
rect 124364 264088 124416 264094
rect 124364 264030 124416 264036
rect 124376 263482 124404 264030
rect 124364 263476 124416 263482
rect 124364 263418 124416 263424
rect 127780 260626 127808 269334
rect 132092 262796 132144 262802
rect 132092 262738 132144 262744
rect 132000 261436 132052 261442
rect 132000 261378 132052 261384
rect 123536 260620 123588 260626
rect 123536 260562 123588 260568
rect 127768 260620 127820 260626
rect 127768 260562 127820 260568
rect 110196 260484 110248 260490
rect 110196 260426 110248 260432
rect 114796 260484 114848 260490
rect 114796 260426 114848 260432
rect 110208 257786 110236 260426
rect 123548 257786 123576 260562
rect 96224 257758 96560 257786
rect 109900 257758 110236 257786
rect 123240 257758 123576 257786
rect 131354 257392 131410 257401
rect 131354 257327 131356 257336
rect 131408 257327 131410 257336
rect 131356 257298 131408 257304
rect 85080 256880 85132 256886
rect 87196 256880 87248 256886
rect 85080 256822 85132 256828
rect 87194 256848 87196 256857
rect 87248 256848 87250 256857
rect 87194 256783 87250 256792
rect 131724 256540 131776 256546
rect 131724 256482 131776 256488
rect 87380 255928 87432 255934
rect 87380 255870 87432 255876
rect 87196 255860 87248 255866
rect 87196 255802 87248 255808
rect 84436 255792 84488 255798
rect 84436 255734 84488 255740
rect 87208 255361 87236 255802
rect 87288 255792 87340 255798
rect 87288 255734 87340 255740
rect 87300 255633 87328 255734
rect 87286 255624 87342 255633
rect 87286 255559 87342 255568
rect 87194 255352 87250 255361
rect 87194 255287 87250 255296
rect 79834 254672 79890 254681
rect 79834 254607 79890 254616
rect 79742 253312 79798 253321
rect 79742 253247 79798 253256
rect 79756 253146 79784 253247
rect 79744 253140 79796 253146
rect 79744 253082 79796 253088
rect 79848 252942 79876 254607
rect 87392 254409 87420 255870
rect 131446 255624 131502 255633
rect 131446 255559 131502 255568
rect 131354 254672 131410 254681
rect 131354 254607 131410 254616
rect 131368 254506 131396 254607
rect 131460 254574 131488 255559
rect 131448 254568 131500 254574
rect 131448 254510 131500 254516
rect 131356 254500 131408 254506
rect 131356 254442 131408 254448
rect 87378 254400 87434 254409
rect 87378 254335 87434 254344
rect 131354 253856 131410 253865
rect 131354 253791 131410 253800
rect 131368 253146 131396 253791
rect 131356 253140 131408 253146
rect 131356 253082 131408 253088
rect 87288 253004 87340 253010
rect 87288 252946 87340 252952
rect 79836 252936 79888 252942
rect 87196 252936 87248 252942
rect 79836 252878 79888 252884
rect 87194 252904 87196 252913
rect 87248 252904 87250 252913
rect 87194 252839 87250 252848
rect 87300 252777 87328 252946
rect 131354 252904 131410 252913
rect 131354 252839 131410 252848
rect 87286 252768 87342 252777
rect 87286 252703 87342 252712
rect 79742 251952 79798 251961
rect 79742 251887 79798 251896
rect 79756 251786 79784 251887
rect 131368 251854 131396 252839
rect 131356 251848 131408 251854
rect 131356 251790 131408 251796
rect 79744 251780 79796 251786
rect 79744 251722 79796 251728
rect 87196 251712 87248 251718
rect 87194 251680 87196 251689
rect 87248 251680 87250 251689
rect 87194 251615 87250 251624
rect 79742 250592 79798 250601
rect 79742 250527 79798 250536
rect 79756 250426 79784 250527
rect 79744 250420 79796 250426
rect 79744 250362 79796 250368
rect 87194 250320 87250 250329
rect 87194 250255 87196 250264
rect 87248 250255 87250 250264
rect 87196 250226 87248 250232
rect 77260 249604 77312 249610
rect 77260 249546 77312 249552
rect 87196 249604 87248 249610
rect 87196 249546 87248 249552
rect 77272 249173 77300 249546
rect 87208 249377 87236 249546
rect 87194 249368 87250 249377
rect 87194 249303 87250 249312
rect 77258 249164 77314 249173
rect 77258 249099 77314 249108
rect 87194 248416 87250 248425
rect 87194 248351 87250 248360
rect 87208 248250 87236 248351
rect 131736 248289 131764 256482
rect 132012 250442 132040 261378
rect 131828 250414 132040 250442
rect 131828 248969 131856 250414
rect 131998 250320 132054 250329
rect 131998 250255 132054 250264
rect 132012 248998 132040 250255
rect 132104 250057 132132 262738
rect 132368 260076 132420 260082
rect 132368 260018 132420 260024
rect 132276 257288 132328 257294
rect 132276 257230 132328 257236
rect 132182 251136 132238 251145
rect 132182 251071 132238 251080
rect 132090 250048 132146 250057
rect 132090 249983 132146 249992
rect 132000 248992 132052 248998
rect 131814 248960 131870 248969
rect 132000 248934 132052 248940
rect 131814 248895 131870 248904
rect 131722 248280 131778 248289
rect 77260 248244 77312 248250
rect 77260 248186 77312 248192
rect 87196 248244 87248 248250
rect 131722 248215 131778 248224
rect 87196 248186 87248 248192
rect 77272 247813 77300 248186
rect 77258 247804 77314 247813
rect 77258 247739 77314 247748
rect 88482 247600 88538 247609
rect 77260 247564 77312 247570
rect 88482 247535 88484 247544
rect 77260 247506 77312 247512
rect 88536 247535 88538 247544
rect 88484 247506 88536 247512
rect 77272 246453 77300 247506
rect 87194 246648 87250 246657
rect 87194 246583 87250 246592
rect 77258 246444 77314 246453
rect 77258 246379 77314 246388
rect 87208 246210 87236 246583
rect 78916 246204 78968 246210
rect 78916 246146 78968 246152
rect 87196 246204 87248 246210
rect 87196 246146 87248 246152
rect 78928 245569 78956 246146
rect 131356 246136 131408 246142
rect 131356 246078 131408 246084
rect 87286 245832 87342 245841
rect 87286 245767 87342 245776
rect 78914 245560 78970 245569
rect 78914 245495 78970 245504
rect 87194 244880 87250 244889
rect 80204 244844 80256 244850
rect 87194 244815 87196 244824
rect 80204 244786 80256 244792
rect 87248 244815 87250 244824
rect 87196 244786 87248 244792
rect 78916 244776 78968 244782
rect 78916 244718 78968 244724
rect 78928 244209 78956 244718
rect 78914 244200 78970 244209
rect 78914 244135 78970 244144
rect 80216 242849 80244 244786
rect 87300 244782 87328 245767
rect 131368 245569 131396 246078
rect 131354 245560 131410 245569
rect 131354 245495 131410 245504
rect 87288 244776 87340 244782
rect 87288 244718 87340 244724
rect 131356 244776 131408 244782
rect 131356 244718 131408 244724
rect 131368 244481 131396 244718
rect 131354 244472 131410 244481
rect 131354 244407 131410 244416
rect 87378 244064 87434 244073
rect 87378 243999 87434 244008
rect 87286 243112 87342 243121
rect 87286 243047 87342 243056
rect 80202 242840 80258 242849
rect 80202 242775 80258 242784
rect 87194 242296 87250 242305
rect 87194 242231 87250 242240
rect 79008 242192 79060 242198
rect 79008 242134 79060 242140
rect 78914 240664 78970 240673
rect 78914 240599 78916 240608
rect 78968 240599 78970 240608
rect 78916 240570 78968 240576
rect 79020 239313 79048 242134
rect 87208 242130 87236 242231
rect 87300 242198 87328 243047
rect 87288 242192 87340 242198
rect 87288 242134 87340 242140
rect 79100 242124 79152 242130
rect 79100 242066 79152 242072
rect 87196 242124 87248 242130
rect 87196 242066 87248 242072
rect 79006 239304 79062 239313
rect 79006 239239 79062 239248
rect 79112 238633 79140 242066
rect 87392 240634 87420 243999
rect 131908 243212 131960 243218
rect 131908 243154 131960 243160
rect 131920 242713 131948 243154
rect 131906 242704 131962 242713
rect 131906 242639 131962 242648
rect 91670 241602 91698 241860
rect 95258 241738 95286 241860
rect 98938 241761 98966 241860
rect 95212 241710 95286 241738
rect 98924 241752 98980 241761
rect 91670 241574 91744 241602
rect 87380 240628 87432 240634
rect 87380 240570 87432 240576
rect 91716 239449 91744 241574
rect 95212 239721 95240 241710
rect 102526 241738 102554 241860
rect 102526 241710 102600 241738
rect 98924 241687 98980 241696
rect 95198 239712 95254 239721
rect 95198 239647 95254 239656
rect 91702 239440 91758 239449
rect 91702 239375 91758 239384
rect 102572 238633 102600 241710
rect 106206 241602 106234 241860
rect 109794 241738 109822 241860
rect 113474 241738 113502 241860
rect 117062 241738 117090 241860
rect 109794 241710 109868 241738
rect 113474 241710 113548 241738
rect 117062 241710 117136 241738
rect 105148 241574 106234 241602
rect 79098 238624 79154 238633
rect 79098 238559 79154 238568
rect 102558 238624 102614 238633
rect 102558 238559 102614 238568
rect 78916 236616 78968 236622
rect 78914 236584 78916 236593
rect 78968 236584 78970 236593
rect 78914 236519 78970 236528
rect 105148 233086 105176 241574
rect 109840 235777 109868 241710
rect 109826 235768 109882 235777
rect 109826 235703 109882 235712
rect 113520 234514 113548 241710
rect 113508 234508 113560 234514
rect 113508 234450 113560 234456
rect 117108 234446 117136 241710
rect 120742 241602 120770 241860
rect 124330 241654 124358 241860
rect 120328 241574 120770 241602
rect 123076 241648 123128 241654
rect 123076 241590 123128 241596
rect 124318 241648 124370 241654
rect 128010 241602 128038 241860
rect 124318 241590 124370 241596
rect 117096 234440 117148 234446
rect 117096 234382 117148 234388
rect 105136 233080 105188 233086
rect 105136 233022 105188 233028
rect 76800 230904 76852 230910
rect 76800 230846 76852 230852
rect 115992 230428 116044 230434
rect 115992 230370 116044 230376
rect 103480 230360 103532 230366
rect 103480 230302 103532 230308
rect 91060 230292 91112 230298
rect 91060 230234 91112 230240
rect 91072 227716 91100 230234
rect 103492 227716 103520 230302
rect 116004 227716 116032 230370
rect 120328 230298 120356 241574
rect 123088 230366 123116 241590
rect 127228 241574 128038 241602
rect 127228 230434 127256 241574
rect 132196 239274 132224 251071
rect 132288 246113 132316 257230
rect 132380 256546 132408 260018
rect 132644 258648 132696 258654
rect 132644 258590 132696 258596
rect 132368 256540 132420 256546
rect 132368 256482 132420 256488
rect 132366 256440 132422 256449
rect 132366 256375 132422 256384
rect 132380 255934 132408 256375
rect 132368 255928 132420 255934
rect 132368 255870 132420 255876
rect 132656 248130 132684 258590
rect 133378 252088 133434 252097
rect 133378 252023 133434 252032
rect 132472 248102 132684 248130
rect 132472 247065 132500 248102
rect 132458 247056 132514 247065
rect 132458 246991 132514 247000
rect 132274 246104 132330 246113
rect 132274 246039 132330 246048
rect 132644 243348 132696 243354
rect 132644 243290 132696 243296
rect 132656 243121 132684 243290
rect 132642 243112 132698 243121
rect 132642 243047 132698 243056
rect 133392 240634 133420 252023
rect 133380 240628 133432 240634
rect 133380 240570 133432 240576
rect 132184 239268 132236 239274
rect 132184 239210 132236 239216
rect 127860 237228 127912 237234
rect 127860 237170 127912 237176
rect 127872 236622 127900 237170
rect 127860 236616 127912 236622
rect 127860 236558 127912 236564
rect 128136 236616 128188 236622
rect 128136 236558 128188 236564
rect 127216 230428 127268 230434
rect 127216 230370 127268 230376
rect 123076 230360 123128 230366
rect 123076 230302 123128 230308
rect 120316 230292 120368 230298
rect 120316 230234 120368 230240
rect 128148 227730 128176 236558
rect 134772 230842 134800 371742
rect 184084 367658 184112 370924
rect 186568 367658 186596 370924
rect 189052 368610 189080 370924
rect 190800 370910 191550 370938
rect 194034 370910 194784 370938
rect 189040 368604 189092 368610
rect 189040 368546 189092 368552
rect 190696 368604 190748 368610
rect 190696 368546 190748 368552
rect 184072 367652 184124 367658
rect 184072 367594 184124 367600
rect 185084 367652 185136 367658
rect 185084 367594 185136 367600
rect 185268 367652 185320 367658
rect 185268 367594 185320 367600
rect 186556 367652 186608 367658
rect 186556 367594 186608 367600
rect 139636 357928 139688 357934
rect 139636 357870 139688 357876
rect 174044 357928 174096 357934
rect 174044 357870 174096 357876
rect 139648 357769 139676 357870
rect 139634 357760 139690 357769
rect 139634 357695 139690 357704
rect 174056 357225 174084 357870
rect 174042 357216 174098 357225
rect 174042 357151 174098 357160
rect 139636 356568 139688 356574
rect 139634 356536 139636 356545
rect 173492 356568 173544 356574
rect 139688 356536 139690 356545
rect 173492 356510 173544 356516
rect 139634 356471 139690 356480
rect 173504 356137 173532 356510
rect 173490 356128 173546 356137
rect 173490 356063 173546 356072
rect 139636 355208 139688 355214
rect 139634 355176 139636 355185
rect 174044 355208 174096 355214
rect 139688 355176 139690 355185
rect 174042 355176 174044 355185
rect 174096 355176 174098 355185
rect 139634 355111 139690 355120
rect 139728 355140 139780 355146
rect 139728 355082 139780 355088
rect 173768 355140 173820 355146
rect 174042 355111 174098 355120
rect 173768 355082 173820 355088
rect 139740 354641 139768 355082
rect 139726 354632 139782 354641
rect 139726 354567 139782 354576
rect 173780 354097 173808 355082
rect 185096 355078 185124 367594
rect 185084 355072 185136 355078
rect 185084 355014 185136 355020
rect 173766 354088 173822 354097
rect 173766 354023 173822 354032
rect 139636 353848 139688 353854
rect 139636 353790 139688 353796
rect 174044 353848 174096 353854
rect 174044 353790 174096 353796
rect 139648 353553 139676 353790
rect 139634 353544 139690 353553
rect 139634 353479 139690 353488
rect 174056 353009 174084 353790
rect 174042 353000 174098 353009
rect 174042 352935 174098 352944
rect 139636 352420 139688 352426
rect 139636 352362 139688 352368
rect 174044 352420 174096 352426
rect 174044 352362 174096 352368
rect 139648 352329 139676 352362
rect 139634 352320 139690 352329
rect 139634 352255 139690 352264
rect 174056 352057 174084 352362
rect 174042 352048 174098 352057
rect 174042 351983 174098 351992
rect 182322 351368 182378 351377
rect 182322 351303 182378 351312
rect 139452 351128 139504 351134
rect 139452 351070 139504 351076
rect 139464 349609 139492 351070
rect 139636 351060 139688 351066
rect 139636 351002 139688 351008
rect 173860 351060 173912 351066
rect 173860 351002 173912 351008
rect 139648 350561 139676 351002
rect 139726 350960 139782 350969
rect 139726 350895 139782 350904
rect 173674 350960 173730 350969
rect 173674 350895 173730 350904
rect 139634 350552 139690 350561
rect 139634 350487 139690 350496
rect 139740 350386 139768 350895
rect 173688 350386 173716 350895
rect 139728 350380 139780 350386
rect 139728 350322 139780 350328
rect 173676 350380 173728 350386
rect 173676 350322 173728 350328
rect 173872 349881 173900 351002
rect 180758 350008 180814 350017
rect 180758 349943 180814 349952
rect 173858 349872 173914 349881
rect 173858 349807 173914 349816
rect 139544 349768 139596 349774
rect 139544 349710 139596 349716
rect 139450 349600 139506 349609
rect 139450 349535 139506 349544
rect 137244 348408 137296 348414
rect 137244 348350 137296 348356
rect 137256 346850 137284 348350
rect 137520 348340 137572 348346
rect 137520 348282 137572 348288
rect 137532 346918 137560 348282
rect 139556 348249 139584 349710
rect 172848 349700 172900 349706
rect 172848 349642 172900 349648
rect 172860 348929 172888 349642
rect 172846 348920 172902 348929
rect 172846 348855 172902 348864
rect 139542 348240 139598 348249
rect 139542 348175 139598 348184
rect 180772 348006 180800 349943
rect 182336 349706 182364 351303
rect 185280 351066 185308 367594
rect 186372 355072 186424 355078
rect 186372 355014 186424 355020
rect 186384 351748 186412 355014
rect 190708 351626 190736 368546
rect 190800 359401 190828 370910
rect 190786 359392 190842 359401
rect 190786 359327 190842 359336
rect 194756 355078 194784 370910
rect 196320 370910 196518 370938
rect 196320 355162 196348 370910
rect 199080 367658 199108 370924
rect 200368 370910 201578 370938
rect 199068 367652 199120 367658
rect 199068 367594 199120 367600
rect 200264 367652 200316 367658
rect 200264 367594 200316 367600
rect 196320 355134 196532 355162
rect 194744 355072 194796 355078
rect 194744 355014 194796 355020
rect 196308 355072 196360 355078
rect 196308 355014 196360 355020
rect 196216 353916 196268 353922
rect 196216 353858 196268 353864
rect 196228 352426 196256 353858
rect 196216 352420 196268 352426
rect 196216 352362 196268 352368
rect 191246 351912 191302 351921
rect 191246 351847 191248 351856
rect 191300 351847 191302 351856
rect 191248 351818 191300 351824
rect 196320 351748 196348 355014
rect 196504 353922 196532 355134
rect 200276 354058 200304 367594
rect 200264 354052 200316 354058
rect 200264 353994 200316 354000
rect 196492 353916 196544 353922
rect 196492 353858 196544 353864
rect 200368 353854 200396 370910
rect 204048 367658 204076 370924
rect 205980 370910 206546 370938
rect 204036 367652 204088 367658
rect 204036 367594 204088 367600
rect 205876 367652 205928 367658
rect 205876 367594 205928 367600
rect 201368 354052 201420 354058
rect 201368 353994 201420 354000
rect 200356 353848 200408 353854
rect 200356 353790 200408 353796
rect 201380 351748 201408 353994
rect 205888 351626 205916 367594
rect 205980 355146 206008 370910
rect 209016 368610 209044 370924
rect 211408 370910 211606 370938
rect 209004 368604 209056 368610
rect 209004 368546 209056 368552
rect 210016 368604 210068 368610
rect 210016 368546 210068 368552
rect 210028 363510 210056 368546
rect 210016 363504 210068 363510
rect 210016 363446 210068 363452
rect 210844 363504 210896 363510
rect 210844 363446 210896 363452
rect 210856 363322 210884 363446
rect 210856 363294 210976 363322
rect 205968 355140 206020 355146
rect 205968 355082 206020 355088
rect 210948 351762 210976 363294
rect 211408 355214 211436 370910
rect 214076 355214 214104 370924
rect 215548 370910 216574 370938
rect 215548 356574 215576 370910
rect 219044 368610 219072 370924
rect 221068 370910 221542 370938
rect 219032 368604 219084 368610
rect 219032 368546 219084 368552
rect 220320 368604 220372 368610
rect 220320 368546 220372 368552
rect 215536 356568 215588 356574
rect 215536 356510 215588 356516
rect 211396 355208 211448 355214
rect 211396 355150 211448 355156
rect 212684 355208 212736 355214
rect 212684 355150 212736 355156
rect 214064 355208 214116 355214
rect 214064 355150 214116 355156
rect 216364 355208 216416 355214
rect 216364 355150 216416 355156
rect 212696 355010 212724 355150
rect 212684 355004 212736 355010
rect 212684 354946 212736 354952
rect 210948 351734 211330 351762
rect 216376 351748 216404 355150
rect 220332 355078 220360 368546
rect 221068 357934 221096 370910
rect 223092 367590 223120 388470
rect 279672 386714 279700 393162
rect 288780 392546 288808 396344
rect 315368 393226 315396 396344
rect 341956 393809 341984 396344
rect 368452 396234 368480 396344
rect 395040 396234 395068 396344
rect 368452 396206 368664 396234
rect 395040 396206 395160 396234
rect 341942 393800 341998 393809
rect 341942 393735 341998 393744
rect 315356 393220 315408 393226
rect 315356 393162 315408 393168
rect 314620 393152 314672 393158
rect 314620 393094 314672 393100
rect 284444 392540 284496 392546
rect 284444 392482 284496 392488
rect 288768 392540 288820 392546
rect 288768 392482 288820 392488
rect 284456 386714 284484 392482
rect 299624 389752 299676 389758
rect 299624 389694 299676 389700
rect 288952 389072 289004 389078
rect 288952 389014 289004 389020
rect 279364 386686 279700 386714
rect 284332 386686 284484 386714
rect 288964 386714 288992 389014
rect 294196 389004 294248 389010
rect 294196 388946 294248 388952
rect 294208 386714 294236 388946
rect 299636 386714 299664 389694
rect 304592 388528 304644 388534
rect 304592 388470 304644 388476
rect 304604 386714 304632 388470
rect 309284 388392 309336 388398
rect 309284 388334 309336 388340
rect 288964 386686 289300 386714
rect 294208 386686 294360 386714
rect 299328 386686 299664 386714
rect 304296 386686 304632 386714
rect 309296 386714 309324 388334
rect 314632 386714 314660 393094
rect 358504 388732 358556 388738
rect 358504 388674 358556 388680
rect 322532 388528 322584 388534
rect 322532 388470 322584 388476
rect 315632 388392 315684 388398
rect 315632 388334 315684 388340
rect 309296 386686 309356 386714
rect 314324 386686 314660 386714
rect 225286 384824 225342 384833
rect 225286 384759 225342 384768
rect 225194 382104 225250 382113
rect 225194 382039 225250 382048
rect 223080 367584 223132 367590
rect 223080 367526 223132 367532
rect 221056 357928 221108 357934
rect 221056 357870 221108 357876
rect 220320 355072 220372 355078
rect 220320 355014 220372 355020
rect 221332 355072 221384 355078
rect 221332 355014 221384 355020
rect 221344 351748 221372 355014
rect 190708 351598 191366 351626
rect 205888 351598 206362 351626
rect 185268 351060 185320 351066
rect 185268 351002 185320 351008
rect 182324 349700 182376 349706
rect 182324 349642 182376 349648
rect 180942 349056 180998 349065
rect 180942 348991 180998 349000
rect 180850 348376 180906 348385
rect 180850 348311 180906 348320
rect 174044 348000 174096 348006
rect 174044 347942 174096 347948
rect 180760 348000 180812 348006
rect 180760 347942 180812 347948
rect 174056 347841 174084 347942
rect 174042 347832 174098 347841
rect 174042 347767 174098 347776
rect 180758 347288 180814 347297
rect 180758 347223 180814 347232
rect 139728 346980 139780 346986
rect 139728 346922 139780 346928
rect 137520 346912 137572 346918
rect 139636 346912 139688 346918
rect 137520 346854 137572 346860
rect 139634 346880 139636 346889
rect 139688 346880 139690 346889
rect 137244 346844 137296 346850
rect 139634 346815 139690 346824
rect 137244 346786 137296 346792
rect 139636 345620 139688 345626
rect 139636 345562 139688 345568
rect 138164 344260 138216 344266
rect 138164 344202 138216 344208
rect 138176 341410 138204 344202
rect 139648 344169 139676 345562
rect 139740 345393 139768 346922
rect 174044 346912 174096 346918
rect 174042 346880 174044 346889
rect 174096 346880 174098 346889
rect 139820 346844 139872 346850
rect 174042 346815 174098 346824
rect 139820 346786 139872 346792
rect 139832 346345 139860 346786
rect 139818 346336 139874 346345
rect 139818 346271 139874 346280
rect 173124 346300 173176 346306
rect 173124 346242 173176 346248
rect 173136 345801 173164 346242
rect 173122 345792 173178 345801
rect 173122 345727 173178 345736
rect 173032 345620 173084 345626
rect 173032 345562 173084 345568
rect 139726 345384 139782 345393
rect 139726 345319 139782 345328
rect 139728 344192 139780 344198
rect 139634 344160 139690 344169
rect 139728 344134 139780 344140
rect 172940 344192 172992 344198
rect 172940 344134 172992 344140
rect 139634 344095 139690 344104
rect 139636 342764 139688 342770
rect 139636 342706 139688 342712
rect 139648 342673 139676 342706
rect 139634 342664 139690 342673
rect 139634 342599 139690 342608
rect 139740 342265 139768 344134
rect 139820 342832 139872 342838
rect 139820 342774 139872 342780
rect 139726 342256 139782 342265
rect 139726 342191 139782 342200
rect 139728 341540 139780 341546
rect 139728 341482 139780 341488
rect 138164 341404 138216 341410
rect 138164 341346 138216 341352
rect 139636 341404 139688 341410
rect 139636 341346 139688 341352
rect 139648 341313 139676 341346
rect 139634 341304 139690 341313
rect 139634 341239 139690 341248
rect 137336 340112 137388 340118
rect 137336 340054 137388 340060
rect 136140 338752 136192 338758
rect 136140 338694 136192 338700
rect 136152 334474 136180 338694
rect 136232 337324 136284 337330
rect 136232 337266 136284 337272
rect 136140 334468 136192 334474
rect 136140 334410 136192 334416
rect 136244 334270 136272 337266
rect 137348 337262 137376 340054
rect 139636 338684 139688 338690
rect 139636 338626 139688 338632
rect 137336 337256 137388 337262
rect 137336 337198 137388 337204
rect 138072 336032 138124 336038
rect 138072 335974 138124 335980
rect 136232 334264 136284 334270
rect 136232 334206 136284 334212
rect 136968 334196 137020 334202
rect 136968 334138 137020 334144
rect 134852 333788 134904 333794
rect 134852 333730 134904 333736
rect 134864 232406 134892 333730
rect 136980 332201 137008 334138
rect 137060 334128 137112 334134
rect 137060 334070 137112 334076
rect 136966 332192 137022 332201
rect 136966 332127 137022 332136
rect 136876 326920 136928 326926
rect 136876 326862 136928 326868
rect 136888 326314 136916 326862
rect 136876 326308 136928 326314
rect 136876 326250 136928 326256
rect 136416 308288 136468 308294
rect 136416 308230 136468 308236
rect 136428 301601 136456 308230
rect 136888 304729 136916 326250
rect 136980 310985 137008 332127
rect 137072 330841 137100 334070
rect 137244 334060 137296 334066
rect 137244 334002 137296 334008
rect 137152 333992 137204 333998
rect 137152 333934 137204 333940
rect 137058 330832 137114 330841
rect 137058 330767 137114 330776
rect 137072 314113 137100 330767
rect 137164 328121 137192 333934
rect 137256 328801 137284 334002
rect 137520 333924 137572 333930
rect 137520 333866 137572 333872
rect 137532 329102 137560 333866
rect 137980 333856 138032 333862
rect 137980 333798 138032 333804
rect 137520 329096 137572 329102
rect 137520 329038 137572 329044
rect 137242 328792 137298 328801
rect 137242 328727 137298 328736
rect 137150 328112 137206 328121
rect 137150 328047 137206 328056
rect 137164 317241 137192 328047
rect 137256 320369 137284 328727
rect 137242 320360 137298 320369
rect 137242 320295 137298 320304
rect 137150 317232 137206 317241
rect 137150 317167 137206 317176
rect 137058 314104 137114 314113
rect 137058 314039 137114 314048
rect 136966 310976 137022 310985
rect 136966 310911 137022 310920
rect 136968 310872 137020 310878
rect 136968 310814 137020 310820
rect 136980 308294 137008 310814
rect 136968 308288 137020 308294
rect 136968 308230 137020 308236
rect 137532 307857 137560 329038
rect 137992 327538 138020 333798
rect 138084 333114 138112 335974
rect 138164 335964 138216 335970
rect 138164 335906 138216 335912
rect 138072 333108 138124 333114
rect 138072 333050 138124 333056
rect 138176 331754 138204 335906
rect 139648 335873 139676 338626
rect 139740 338593 139768 341482
rect 139832 339953 139860 342774
rect 172756 342288 172808 342294
rect 172756 342230 172808 342236
rect 172768 341585 172796 342230
rect 172754 341576 172810 341585
rect 172754 341511 172810 341520
rect 139912 341472 139964 341478
rect 139912 341414 139964 341420
rect 139818 339944 139874 339953
rect 139818 339879 139874 339888
rect 139726 338584 139782 338593
rect 139726 338519 139782 338528
rect 139924 338185 139952 341414
rect 172952 340633 172980 344134
rect 173044 342673 173072 345562
rect 180772 345218 180800 347223
rect 180864 346306 180892 348311
rect 180956 346918 180984 348991
rect 180944 346912 180996 346918
rect 180944 346854 180996 346860
rect 181034 346880 181090 346889
rect 181034 346815 181090 346824
rect 180852 346300 180904 346306
rect 180852 346242 180904 346248
rect 181048 345801 181076 346815
rect 182322 346064 182378 346073
rect 182322 345999 182378 346008
rect 180850 345792 180906 345801
rect 180850 345727 180906 345736
rect 181034 345792 181090 345801
rect 181034 345727 181090 345736
rect 173308 345212 173360 345218
rect 173308 345154 173360 345160
rect 180760 345212 180812 345218
rect 180760 345154 180812 345160
rect 173320 344713 173348 345154
rect 173306 344704 173362 344713
rect 173306 344639 173362 344648
rect 180864 343790 180892 345727
rect 182336 345626 182364 345999
rect 182324 345620 182376 345626
rect 182324 345562 182376 345568
rect 180942 344704 180998 344713
rect 180942 344639 180998 344648
rect 173676 343784 173728 343790
rect 173674 343752 173676 343761
rect 180852 343784 180904 343790
rect 173728 343752 173730 343761
rect 180852 343726 180904 343732
rect 173674 343687 173730 343696
rect 173676 342832 173728 342838
rect 173676 342774 173728 342780
rect 173030 342664 173086 342673
rect 173030 342599 173086 342608
rect 172938 340624 172994 340633
rect 172938 340559 172994 340568
rect 173492 340112 173544 340118
rect 173492 340054 173544 340060
rect 173308 338752 173360 338758
rect 173308 338694 173360 338700
rect 139910 338176 139966 338185
rect 139910 338111 139966 338120
rect 139728 337256 139780 337262
rect 139728 337198 139780 337204
rect 139740 336825 139768 337198
rect 139726 336816 139782 336825
rect 139726 336751 139782 336760
rect 172848 335964 172900 335970
rect 172848 335906 172900 335912
rect 139634 335864 139690 335873
rect 139634 335799 139690 335808
rect 139636 334468 139688 334474
rect 139636 334410 139688 334416
rect 139648 334377 139676 334410
rect 139634 334368 139690 334377
rect 139634 334303 139690 334312
rect 139636 334264 139688 334270
rect 139636 334206 139688 334212
rect 139648 333969 139676 334206
rect 139634 333960 139690 333969
rect 139634 333895 139690 333904
rect 139636 333108 139688 333114
rect 139636 333050 139688 333056
rect 139648 333017 139676 333050
rect 139634 333008 139690 333017
rect 139634 332943 139690 332952
rect 172860 332337 172888 335906
rect 173320 335465 173348 338694
rect 173400 338684 173452 338690
rect 173400 338626 173452 338632
rect 173306 335456 173362 335465
rect 173306 335391 173362 335400
rect 173412 334377 173440 338626
rect 173504 336417 173532 340054
rect 173688 339545 173716 342774
rect 180956 342294 180984 344639
rect 182322 344296 182378 344305
rect 182322 344231 182378 344240
rect 182336 344198 182364 344231
rect 182324 344192 182376 344198
rect 182324 344134 182376 344140
rect 181402 343344 181458 343353
rect 181402 343279 181458 343288
rect 181416 342838 181444 343279
rect 181404 342832 181456 342838
rect 181404 342774 181456 342780
rect 182138 342392 182194 342401
rect 182138 342327 182194 342336
rect 180944 342288 180996 342294
rect 180944 342230 180996 342236
rect 181770 341576 181826 341585
rect 181770 341511 181826 341520
rect 181402 340624 181458 340633
rect 181402 340559 181458 340568
rect 181416 340118 181444 340559
rect 181404 340112 181456 340118
rect 181404 340054 181456 340060
rect 181586 339808 181642 339817
rect 181586 339743 181642 339752
rect 173674 339536 173730 339545
rect 173674 339471 173730 339480
rect 181600 338758 181628 339743
rect 181588 338752 181640 338758
rect 181588 338694 181640 338700
rect 181784 338622 181812 341511
rect 173952 338616 174004 338622
rect 181772 338616 181824 338622
rect 173952 338558 174004 338564
rect 174042 338584 174098 338593
rect 173964 337505 173992 338558
rect 181772 338558 181824 338564
rect 182152 338554 182180 342327
rect 182322 338856 182378 338865
rect 182322 338791 182378 338800
rect 182336 338690 182364 338791
rect 182324 338684 182376 338690
rect 182324 338626 182376 338632
rect 174042 338519 174044 338528
rect 174096 338519 174098 338528
rect 182140 338548 182192 338554
rect 174044 338490 174096 338496
rect 182140 338490 182192 338496
rect 173950 337496 174006 337505
rect 173950 337431 174006 337440
rect 180390 337496 180446 337505
rect 180390 337431 180446 337440
rect 173490 336408 173546 336417
rect 173490 336343 173546 336352
rect 173398 334368 173454 334377
rect 173398 334303 173454 334312
rect 180404 333522 180432 337431
rect 181586 337088 181642 337097
rect 181586 337023 181642 337032
rect 180942 336136 180998 336145
rect 180942 336071 180998 336080
rect 173308 333516 173360 333522
rect 173308 333458 173360 333464
rect 180392 333516 180444 333522
rect 180392 333458 180444 333464
rect 173320 333289 173348 333458
rect 173306 333280 173362 333289
rect 173306 333215 173362 333224
rect 172846 332328 172902 332337
rect 172846 332263 172902 332272
rect 180956 331754 180984 336071
rect 181600 335970 181628 337023
rect 198712 336094 198910 336122
rect 181588 335964 181640 335970
rect 181588 335906 181640 335912
rect 187948 335958 188882 335986
rect 192088 335958 192194 335986
rect 194848 335958 195506 335986
rect 185570 335822 185952 335850
rect 185084 333856 185136 333862
rect 185084 333798 185136 333804
rect 138164 331748 138216 331754
rect 138164 331690 138216 331696
rect 139636 331748 139688 331754
rect 139636 331690 139688 331696
rect 173676 331748 173728 331754
rect 173676 331690 173728 331696
rect 180944 331748 180996 331754
rect 180944 331690 180996 331696
rect 139648 331657 139676 331690
rect 139634 331648 139690 331657
rect 139634 331583 139690 331592
rect 173688 331249 173716 331690
rect 173674 331240 173730 331249
rect 173674 331175 173730 331184
rect 140370 330288 140426 330297
rect 140370 330223 140426 330232
rect 172110 330288 172166 330297
rect 172110 330223 172166 330232
rect 140384 329034 140412 330223
rect 158586 330152 158642 330161
rect 159598 330152 159654 330161
rect 158642 330110 158752 330138
rect 158586 330087 158642 330096
rect 159654 330110 159764 330138
rect 159598 330087 159654 330096
rect 155900 329974 155960 330002
rect 156820 329974 156880 330002
rect 142408 329838 143388 329866
rect 144308 329838 144644 329866
rect 145228 329838 145564 329866
rect 140372 329028 140424 329034
rect 140372 328970 140424 328976
rect 137704 327532 137756 327538
rect 137704 327474 137756 327480
rect 137980 327532 138032 327538
rect 137980 327474 138032 327480
rect 137612 326988 137664 326994
rect 137612 326930 137664 326936
rect 137518 307848 137574 307857
rect 137518 307783 137574 307792
rect 136874 304720 136930 304729
rect 136874 304655 136930 304664
rect 137518 304720 137574 304729
rect 137518 304655 137574 304664
rect 136414 301592 136470 301601
rect 136414 301527 136470 301536
rect 136428 298706 136456 301527
rect 136416 298700 136468 298706
rect 136416 298642 136468 298648
rect 136876 298700 136928 298706
rect 136876 298642 136928 298648
rect 136888 284873 136916 298642
rect 136874 284864 136930 284873
rect 136874 284799 136930 284808
rect 136874 282552 136930 282561
rect 136874 282487 136930 282496
rect 136888 282386 136916 282487
rect 136876 282380 136928 282386
rect 136876 282322 136928 282328
rect 136874 282280 136930 282289
rect 136874 282215 136930 282224
rect 135128 257356 135180 257362
rect 135128 257298 135180 257304
rect 135036 254568 135088 254574
rect 135036 254510 135088 254516
rect 134944 254500 134996 254506
rect 134944 254442 134996 254448
rect 134956 246210 134984 254442
rect 135048 247366 135076 254510
rect 135140 250290 135168 257298
rect 136232 255996 136284 256002
rect 136232 255938 136284 255944
rect 135128 250284 135180 250290
rect 135128 250226 135180 250232
rect 136140 248992 136192 248998
rect 136140 248934 136192 248940
rect 135036 247360 135088 247366
rect 135036 247302 135088 247308
rect 134944 246204 134996 246210
rect 134944 246146 134996 246152
rect 136152 239206 136180 248934
rect 136244 246142 136272 255938
rect 136324 251848 136376 251854
rect 136324 251790 136376 251796
rect 136232 246136 136284 246142
rect 136232 246078 136284 246084
rect 136336 243422 136364 251790
rect 136324 243416 136376 243422
rect 136324 243358 136376 243364
rect 136140 239200 136192 239206
rect 136140 239142 136192 239148
rect 134852 232400 134904 232406
rect 134852 232342 134904 232348
rect 134760 230836 134812 230842
rect 134760 230778 134812 230784
rect 128148 227702 128530 227730
rect 76800 226960 76852 226966
rect 76800 226902 76852 226908
rect 76156 219548 76208 219554
rect 76156 219490 76208 219496
rect 75418 217408 75474 217417
rect 75418 217343 75474 217352
rect 74408 214516 74460 214522
rect 74408 214458 74460 214464
rect 74406 211696 74462 211705
rect 74406 211631 74462 211640
rect 74420 205449 74448 211631
rect 74406 205440 74462 205449
rect 74406 205375 74462 205384
rect 74316 203364 74368 203370
rect 74316 203306 74368 203312
rect 74314 200544 74370 200553
rect 74314 200479 74370 200488
rect 74328 191985 74356 200479
rect 74314 191976 74370 191985
rect 74314 191911 74370 191920
rect 74328 191033 74356 191911
rect 74314 191024 74370 191033
rect 74314 190959 74370 190968
rect 74222 188032 74278 188041
rect 74222 187967 74278 187976
rect 74236 186953 74264 187967
rect 74498 187080 74554 187089
rect 74498 187015 74554 187024
rect 74222 186944 74278 186953
rect 74222 186879 74278 186888
rect 74038 185176 74094 185185
rect 74038 185111 74094 185120
rect 74406 181232 74462 181241
rect 74406 181167 74462 181176
rect 73762 180008 73818 180017
rect 73762 179943 73818 179952
rect 74224 172424 74276 172430
rect 74224 172366 74276 172372
rect 73120 172356 73172 172362
rect 73120 172298 73172 172304
rect 72660 171676 72712 171682
rect 72660 171618 72712 171624
rect 72672 169817 72700 171618
rect 72658 169808 72714 169817
rect 73132 169780 73160 172298
rect 74236 169780 74264 172366
rect 74420 171721 74448 181167
rect 74512 180017 74540 187015
rect 75432 186846 75460 217343
rect 75420 186840 75472 186846
rect 75420 186782 75472 186788
rect 74498 180008 74554 180017
rect 74498 179943 74554 179952
rect 75236 172492 75288 172498
rect 75236 172434 75288 172440
rect 74406 171712 74462 171721
rect 74406 171647 74462 171656
rect 75248 169780 75276 172434
rect 76168 169794 76196 219490
rect 76168 169766 76274 169794
rect 72658 169743 72714 169752
rect 57690 169630 58164 169658
rect 61830 169630 62304 169658
rect 73486 169536 73542 169545
rect 73486 169471 73542 169480
rect 73500 169438 73528 169471
rect 73488 169432 73540 169438
rect 73488 169374 73540 169380
rect 49200 168888 49252 168894
rect 49198 168856 49200 168865
rect 49252 168856 49254 168865
rect 49198 168791 49254 168800
rect 47082 143424 47138 143433
rect 47082 143359 47138 143368
rect 48568 141886 49410 141914
rect 49948 141886 50422 141914
rect 51328 141886 51434 141914
rect 51604 141886 52446 141914
rect 38802 127512 38858 127521
rect 38802 127447 38858 127456
rect 38816 126802 38844 127447
rect 38804 126796 38856 126802
rect 38804 126738 38856 126744
rect 38252 126116 38304 126122
rect 38252 126058 38304 126064
rect 38264 125617 38292 126058
rect 38250 125608 38306 125617
rect 38250 125543 38306 125552
rect 38802 122752 38858 122761
rect 38802 122687 38858 122696
rect 38816 122654 38844 122687
rect 38804 122648 38856 122654
rect 38804 122590 38856 122596
rect 38804 120608 38856 120614
rect 38804 120550 38856 120556
rect 38816 120313 38844 120550
rect 38802 120304 38858 120313
rect 38802 120239 38858 120248
rect 38250 117584 38306 117593
rect 38250 117519 38306 117528
rect 38264 117146 38292 117519
rect 38252 117140 38304 117146
rect 38252 117082 38304 117088
rect 38804 115100 38856 115106
rect 38804 115042 38856 115048
rect 38816 115009 38844 115042
rect 38802 115000 38858 115009
rect 38802 114935 38858 114944
rect 38804 112992 38856 112998
rect 38804 112934 38856 112940
rect 38816 112833 38844 112934
rect 38802 112824 38858 112833
rect 38802 112759 38858 112768
rect 38252 110952 38304 110958
rect 38252 110894 38304 110900
rect 38264 110521 38292 110894
rect 38250 110512 38306 110521
rect 38250 110447 38306 110456
rect 38802 107520 38858 107529
rect 38802 107455 38804 107464
rect 38856 107455 38858 107464
rect 38804 107426 38856 107432
rect 38804 105444 38856 105450
rect 38804 105386 38856 105392
rect 38816 105353 38844 105386
rect 38802 105344 38858 105353
rect 38802 105279 38858 105288
rect 38618 102488 38674 102497
rect 38618 102423 38674 102432
rect 38632 101370 38660 102423
rect 38620 101364 38672 101370
rect 38620 101306 38672 101312
rect 38804 100616 38856 100622
rect 38804 100558 38856 100564
rect 38816 100321 38844 100558
rect 38802 100312 38858 100321
rect 38802 100247 38858 100256
rect 38802 97864 38858 97873
rect 38802 97799 38804 97808
rect 38856 97799 38858 97808
rect 38804 97770 38856 97776
rect 38068 95788 38120 95794
rect 38068 95730 38120 95736
rect 38080 95425 38108 95730
rect 38066 95416 38122 95425
rect 38066 95351 38122 95360
rect 37606 92560 37662 92569
rect 37606 92495 37662 92504
rect 37620 92326 37648 92495
rect 48568 92326 48596 141886
rect 49948 97834 49976 141886
rect 51222 126288 51278 126297
rect 51222 126223 51278 126232
rect 51236 126122 51264 126223
rect 51224 126116 51276 126122
rect 51224 126058 51276 126064
rect 51222 116224 51278 116233
rect 51222 116159 51278 116168
rect 51236 115106 51264 116159
rect 51224 115100 51276 115106
rect 51224 115042 51276 115048
rect 51328 101574 51356 141886
rect 51604 134418 51632 141886
rect 53536 139625 53564 141900
rect 54548 139625 54576 141900
rect 55468 141886 55574 141914
rect 55652 141886 56586 141914
rect 53522 139616 53578 139625
rect 53522 139551 53578 139560
rect 54534 139616 54590 139625
rect 54534 139551 54590 139560
rect 55364 139308 55416 139314
rect 55364 139250 55416 139256
rect 51592 134412 51644 134418
rect 51592 134354 51644 134360
rect 51868 134412 51920 134418
rect 51868 134354 51920 134360
rect 51880 124778 51908 134354
rect 55376 128722 55404 139250
rect 55468 131601 55496 141886
rect 55652 132417 55680 141886
rect 57676 139586 57704 141900
rect 57664 139580 57716 139586
rect 57664 139522 57716 139528
rect 58124 139444 58176 139450
rect 58124 139386 58176 139392
rect 56744 139376 56796 139382
rect 56744 139318 56796 139324
rect 55638 132408 55694 132417
rect 55638 132343 55694 132352
rect 55454 131592 55510 131601
rect 55454 131527 55510 131536
rect 56756 128858 56784 139318
rect 57020 130944 57072 130950
rect 57020 130886 57072 130892
rect 56388 128830 56784 128858
rect 56388 128722 56416 128830
rect 55298 128694 55404 128722
rect 56126 128694 56416 128722
rect 57032 128708 57060 130886
rect 58136 128722 58164 139386
rect 58688 138702 58716 141900
rect 59504 139648 59556 139654
rect 59504 139590 59556 139596
rect 58676 138696 58728 138702
rect 58676 138638 58728 138644
rect 59516 128858 59544 139590
rect 59700 138838 59728 141900
rect 60240 139580 60292 139586
rect 60240 139522 60292 139528
rect 59688 138832 59740 138838
rect 59688 138774 59740 138780
rect 59688 131624 59740 131630
rect 59688 131566 59740 131572
rect 59148 128830 59544 128858
rect 59148 128722 59176 128830
rect 57966 128694 58164 128722
rect 58794 128694 59176 128722
rect 59700 128708 59728 131566
rect 60252 130542 60280 139522
rect 60712 138634 60740 141900
rect 60884 139648 60936 139654
rect 60884 139590 60936 139596
rect 60792 139240 60844 139246
rect 60792 139182 60844 139188
rect 60700 138628 60752 138634
rect 60700 138570 60752 138576
rect 60804 131630 60832 139182
rect 60792 131624 60844 131630
rect 60792 131566 60844 131572
rect 60240 130536 60292 130542
rect 60240 130478 60292 130484
rect 60896 128722 60924 139590
rect 61816 138770 61844 141900
rect 62264 139716 62316 139722
rect 62264 139658 62316 139664
rect 61804 138764 61856 138770
rect 61804 138706 61856 138712
rect 62276 130338 62304 139658
rect 62828 138906 62856 141900
rect 63644 139512 63696 139518
rect 63644 139454 63696 139460
rect 62816 138900 62868 138906
rect 62816 138842 62868 138848
rect 63000 138832 63052 138838
rect 63000 138774 63052 138780
rect 63012 130474 63040 138774
rect 63092 138696 63144 138702
rect 63092 138638 63144 138644
rect 63000 130468 63052 130474
rect 63000 130410 63052 130416
rect 62356 130400 62408 130406
rect 62356 130342 62408 130348
rect 61436 130332 61488 130338
rect 61436 130274 61488 130280
rect 62264 130332 62316 130338
rect 62264 130274 62316 130280
rect 60634 128694 60924 128722
rect 61448 128708 61476 130274
rect 62368 128708 62396 130342
rect 63104 130338 63132 138638
rect 63184 138628 63236 138634
rect 63184 138570 63236 138576
rect 63196 131562 63224 138570
rect 63184 131556 63236 131562
rect 63184 131498 63236 131504
rect 63276 130536 63328 130542
rect 63276 130478 63328 130484
rect 63092 130332 63144 130338
rect 63092 130274 63144 130280
rect 63288 128708 63316 130478
rect 63656 130406 63684 139454
rect 63840 139178 63868 141900
rect 64852 139790 64880 141900
rect 64840 139784 64892 139790
rect 64840 139726 64892 139732
rect 65956 139654 65984 141900
rect 65944 139648 65996 139654
rect 65944 139590 65996 139596
rect 66968 139314 66996 141900
rect 67980 139382 68008 141900
rect 68072 141886 69006 141914
rect 67968 139376 68020 139382
rect 67968 139318 68020 139324
rect 66956 139308 67008 139314
rect 66956 139250 67008 139256
rect 63828 139172 63880 139178
rect 63828 139114 63880 139120
rect 67692 138832 67744 138838
rect 67692 138774 67744 138780
rect 65760 138764 65812 138770
rect 65760 138706 65812 138712
rect 65024 130468 65076 130474
rect 65024 130410 65076 130416
rect 63644 130400 63696 130406
rect 63644 130342 63696 130348
rect 64104 130332 64156 130338
rect 64104 130274 64156 130280
rect 64116 128708 64144 130274
rect 65036 128708 65064 130410
rect 65772 130338 65800 138706
rect 65944 131556 65996 131562
rect 65944 131498 65996 131504
rect 65760 130332 65812 130338
rect 65760 130274 65812 130280
rect 65956 128708 65984 131498
rect 66772 130332 66824 130338
rect 66772 130274 66824 130280
rect 66784 128708 66812 130274
rect 67704 128708 67732 138774
rect 68072 130950 68100 141886
rect 70096 139450 70124 141900
rect 70452 139852 70504 139858
rect 70452 139794 70504 139800
rect 70084 139444 70136 139450
rect 70084 139386 70136 139392
rect 68612 139172 68664 139178
rect 68612 139114 68664 139120
rect 68060 130944 68112 130950
rect 68060 130886 68112 130892
rect 68624 128708 68652 139114
rect 70464 129674 70492 139794
rect 70544 139648 70596 139654
rect 70544 139590 70596 139596
rect 69820 129646 70492 129674
rect 69820 128722 69848 129646
rect 70556 128722 70584 139590
rect 71108 139586 71136 141900
rect 71096 139580 71148 139586
rect 71096 139522 71148 139528
rect 72120 139246 72148 141900
rect 73132 139722 73160 141900
rect 74038 141656 74094 141665
rect 74038 141591 74094 141600
rect 73120 139716 73172 139722
rect 73120 139658 73172 139664
rect 72108 139240 72160 139246
rect 72108 139182 72160 139188
rect 74052 137154 74080 141591
rect 74130 141520 74186 141529
rect 74130 141455 74186 141464
rect 69466 128694 69848 128722
rect 70386 128694 70584 128722
rect 73868 137126 74080 137154
rect 74144 137138 74172 141455
rect 74236 139790 74264 141900
rect 74314 141792 74370 141801
rect 74314 141727 74370 141736
rect 74224 139784 74276 139790
rect 74224 139726 74276 139732
rect 74328 139246 74356 141727
rect 75248 139518 75276 141900
rect 76168 141886 76274 141914
rect 75236 139512 75288 139518
rect 75236 139454 75288 139460
rect 74316 139240 74368 139246
rect 74316 139182 74368 139188
rect 74132 137132 74184 137138
rect 73868 127550 73896 137126
rect 74132 137074 74184 137080
rect 73856 127544 73908 127550
rect 73856 127486 73908 127492
rect 74224 127544 74276 127550
rect 74224 127486 74276 127492
rect 74040 127408 74092 127414
rect 74040 127350 74092 127356
rect 54074 127240 54130 127249
rect 54074 127175 54130 127184
rect 54088 126802 54116 127175
rect 54076 126796 54128 126802
rect 54076 126738 54128 126744
rect 51880 124750 52000 124778
rect 74052 124762 74080 127350
rect 51972 117842 52000 124750
rect 74040 124756 74092 124762
rect 74040 124698 74092 124704
rect 53154 122752 53210 122761
rect 53154 122687 53210 122696
rect 74130 122752 74186 122761
rect 74130 122687 74186 122696
rect 53168 122654 53196 122687
rect 53156 122648 53208 122654
rect 53156 122590 53208 122596
rect 52602 121256 52658 121265
rect 52602 121191 52658 121200
rect 52616 120614 52644 121191
rect 52604 120608 52656 120614
rect 52604 120550 52656 120556
rect 73394 120576 73450 120585
rect 73394 120511 73450 120520
rect 73408 119769 73436 120511
rect 73394 119760 73450 119769
rect 73394 119695 73450 119704
rect 51880 117814 52000 117842
rect 51880 115106 51908 117814
rect 54074 117176 54130 117185
rect 54074 117111 54076 117120
rect 54128 117111 54130 117120
rect 54076 117082 54128 117088
rect 51868 115100 51920 115106
rect 51868 115042 51920 115048
rect 52142 113096 52198 113105
rect 52142 113031 52198 113040
rect 52156 112998 52184 113031
rect 52144 112992 52196 112998
rect 52144 112934 52196 112940
rect 52602 111328 52658 111337
rect 52602 111263 52658 111272
rect 52616 110958 52644 111263
rect 52604 110952 52656 110958
rect 52604 110894 52656 110900
rect 51684 108028 51736 108034
rect 51684 107970 51736 107976
rect 51696 107490 51724 107970
rect 51684 107484 51736 107490
rect 51684 107426 51736 107432
rect 50028 101568 50080 101574
rect 50028 101510 50080 101516
rect 51316 101568 51368 101574
rect 51316 101510 51368 101516
rect 50040 101370 50068 101510
rect 50028 101364 50080 101370
rect 50028 101306 50080 101312
rect 49936 97828 49988 97834
rect 49936 97770 49988 97776
rect 37608 92320 37660 92326
rect 37608 92262 37660 92268
rect 48556 92320 48608 92326
rect 48556 92262 48608 92268
rect 38804 90212 38856 90218
rect 38804 90154 38856 90160
rect 38816 90121 38844 90154
rect 38802 90112 38858 90121
rect 38802 90047 38858 90056
rect 21232 87152 21284 87158
rect 21232 87094 21284 87100
rect 34664 87152 34716 87158
rect 34664 87094 34716 87100
rect 48568 75818 48596 92262
rect 48568 75790 48950 75818
rect 49948 75804 49976 97770
rect 50040 75682 50068 101306
rect 51696 91458 51724 107426
rect 52602 106296 52658 106305
rect 52602 106231 52658 106240
rect 52616 105450 52644 106231
rect 52604 105444 52656 105450
rect 52604 105386 52656 105392
rect 52602 101264 52658 101273
rect 52602 101199 52658 101208
rect 52616 100622 52644 101199
rect 52604 100616 52656 100622
rect 52604 100558 52656 100564
rect 52602 96232 52658 96241
rect 52602 96167 52658 96176
rect 52616 95794 52644 96167
rect 52604 95788 52656 95794
rect 52604 95730 52656 95736
rect 72568 94360 72620 94366
rect 72568 94302 72620 94308
rect 51236 91430 51724 91458
rect 51236 90098 51264 91430
rect 52602 91336 52658 91345
rect 52602 91271 52658 91280
rect 52616 90286 52644 91271
rect 52604 90280 52656 90286
rect 52604 90222 52656 90228
rect 51236 90070 51356 90098
rect 51328 75682 51356 90070
rect 69544 88982 70386 89010
rect 55298 88846 55404 88874
rect 53062 79096 53118 79105
rect 53062 79031 53118 79040
rect 54074 79096 54130 79105
rect 54074 79031 54130 79040
rect 53076 75804 53104 79031
rect 54088 75804 54116 79031
rect 55086 78960 55142 78969
rect 55086 78895 55142 78904
rect 55100 75804 55128 78895
rect 55376 78522 55404 88846
rect 56112 86954 56140 88860
rect 56100 86948 56152 86954
rect 56100 86890 56152 86896
rect 57032 86818 57060 88860
rect 57966 88846 58164 88874
rect 58794 88846 59544 88874
rect 57020 86812 57072 86818
rect 57020 86754 57072 86760
rect 56098 79096 56154 79105
rect 56098 79031 56154 79040
rect 55364 78516 55416 78522
rect 55364 78458 55416 78464
rect 56112 75804 56140 79031
rect 58136 78590 58164 88846
rect 59228 79128 59280 79134
rect 59228 79070 59280 79076
rect 58216 78992 58268 78998
rect 58216 78934 58268 78940
rect 58124 78584 58176 78590
rect 58124 78526 58176 78532
rect 57204 78108 57256 78114
rect 57204 78050 57256 78056
rect 57216 75804 57244 78050
rect 58228 75804 58256 78934
rect 59240 75804 59268 79070
rect 59516 78454 59544 88846
rect 59700 86886 59728 88860
rect 60634 88846 60924 88874
rect 59688 86880 59740 86886
rect 59688 86822 59740 86828
rect 60240 79196 60292 79202
rect 60240 79138 60292 79144
rect 59504 78448 59556 78454
rect 59504 78390 59556 78396
rect 60252 75804 60280 79138
rect 60896 78658 60924 88846
rect 61448 86138 61476 88860
rect 61620 86200 61672 86206
rect 61620 86142 61672 86148
rect 61436 86132 61488 86138
rect 61436 86074 61488 86080
rect 60884 78652 60936 78658
rect 60884 78594 60936 78600
rect 61632 78114 61660 86142
rect 62368 86138 62396 88860
rect 63288 86206 63316 88860
rect 63748 88846 64130 88874
rect 64300 88846 65050 88874
rect 63276 86200 63328 86206
rect 63276 86142 63328 86148
rect 62264 86132 62316 86138
rect 62264 86074 62316 86080
rect 62356 86132 62408 86138
rect 62356 86074 62408 86080
rect 63644 86132 63696 86138
rect 63644 86074 63696 86080
rect 62276 78794 62304 86074
rect 62356 78924 62408 78930
rect 62356 78866 62408 78872
rect 62264 78788 62316 78794
rect 62264 78730 62316 78736
rect 61620 78108 61672 78114
rect 61620 78050 61672 78056
rect 61344 78040 61396 78046
rect 61344 77982 61396 77988
rect 61356 75804 61384 77982
rect 62368 75804 62396 78866
rect 63656 78862 63684 86074
rect 63748 78998 63776 88846
rect 64300 86154 64328 88846
rect 65956 87158 65984 88860
rect 64380 87152 64432 87158
rect 64380 87094 64432 87100
rect 65944 87152 65996 87158
rect 65944 87094 65996 87100
rect 63840 86126 64328 86154
rect 63840 79134 63868 86126
rect 64392 79202 64420 87094
rect 65852 86948 65904 86954
rect 65852 86890 65904 86896
rect 65760 86132 65812 86138
rect 65760 86074 65812 86080
rect 64380 79196 64432 79202
rect 64380 79138 64432 79144
rect 63828 79128 63880 79134
rect 63828 79070 63880 79076
rect 63736 78992 63788 78998
rect 63736 78934 63788 78940
rect 64380 78924 64432 78930
rect 64380 78866 64432 78872
rect 63644 78856 63696 78862
rect 63644 78798 63696 78804
rect 63368 78720 63420 78726
rect 63368 78662 63420 78668
rect 63380 75804 63408 78662
rect 64392 75804 64420 78866
rect 65484 78788 65536 78794
rect 65484 78730 65536 78736
rect 65496 75804 65524 78730
rect 65772 78046 65800 86074
rect 65864 78250 65892 86890
rect 66784 86138 66812 88860
rect 67336 88846 67718 88874
rect 67140 86200 67192 86206
rect 67140 86142 67192 86148
rect 66772 86132 66824 86138
rect 66772 86074 66824 86080
rect 66680 86064 66732 86070
rect 66680 86006 66732 86012
rect 66692 79134 66720 86006
rect 66680 79128 66732 79134
rect 66680 79070 66732 79076
rect 67152 78726 67180 86142
rect 67336 86070 67364 88846
rect 67876 86812 67928 86818
rect 67876 86754 67928 86760
rect 67324 86064 67376 86070
rect 67324 86006 67376 86012
rect 67140 78720 67192 78726
rect 67140 78662 67192 78668
rect 66496 78516 66548 78522
rect 66496 78458 66548 78464
rect 65852 78244 65904 78250
rect 65852 78186 65904 78192
rect 65760 78040 65812 78046
rect 65760 77982 65812 77988
rect 66508 75804 66536 78458
rect 67508 78244 67560 78250
rect 67508 78186 67560 78192
rect 67520 75804 67548 78186
rect 67888 75682 67916 86754
rect 68624 86206 68652 88860
rect 68612 86200 68664 86206
rect 68612 86142 68664 86148
rect 69452 86138 69480 88860
rect 68520 86132 68572 86138
rect 68520 86074 68572 86080
rect 69440 86132 69492 86138
rect 69440 86074 69492 86080
rect 68532 78930 68560 86074
rect 69544 86018 69572 88982
rect 72580 88353 72608 94302
rect 73408 93754 73436 119695
rect 73488 117820 73540 117826
rect 73488 117762 73540 117768
rect 73500 116233 73528 117762
rect 74040 117752 74092 117758
rect 74040 117694 74092 117700
rect 73486 116224 73542 116233
rect 73486 116159 73542 116168
rect 73396 93748 73448 93754
rect 73396 93690 73448 93696
rect 72566 88344 72622 88353
rect 72566 88279 72622 88288
rect 72580 87498 72608 88279
rect 72568 87492 72620 87498
rect 72568 87434 72620 87440
rect 73500 87294 73528 116159
rect 74052 115106 74080 117694
rect 74040 115100 74092 115106
rect 74040 115042 74092 115048
rect 73578 112824 73634 112833
rect 73578 112759 73634 112768
rect 73592 93890 73620 112759
rect 73670 109560 73726 109569
rect 73670 109495 73726 109504
rect 73684 108889 73712 109495
rect 73670 108880 73726 108889
rect 73670 108815 73726 108824
rect 73580 93884 73632 93890
rect 73580 93826 73632 93832
rect 73580 93748 73632 93754
rect 73580 93690 73632 93696
rect 73488 87288 73540 87294
rect 73488 87230 73540 87236
rect 70728 86880 70780 86886
rect 70728 86822 70780 86828
rect 69360 85990 69572 86018
rect 68520 78924 68572 78930
rect 68520 78866 68572 78872
rect 69360 78794 69388 85990
rect 69348 78788 69400 78794
rect 69348 78730 69400 78736
rect 69624 78584 69676 78590
rect 69624 78526 69676 78532
rect 69636 75804 69664 78526
rect 70636 78448 70688 78454
rect 70636 78390 70688 78396
rect 70648 75804 70676 78390
rect 70740 75954 70768 86822
rect 73500 86177 73528 87230
rect 73592 87226 73620 93690
rect 73684 87430 73712 108815
rect 73948 98440 74000 98446
rect 73948 98382 74000 98388
rect 73960 94366 73988 98382
rect 73948 94360 74000 94366
rect 73948 94302 74000 94308
rect 73764 93884 73816 93890
rect 73764 93826 73816 93832
rect 73672 87424 73724 87430
rect 73672 87366 73724 87372
rect 73580 87220 73632 87226
rect 73580 87162 73632 87168
rect 73592 86449 73620 87162
rect 73578 86440 73634 86449
rect 73578 86375 73634 86384
rect 73684 86313 73712 87366
rect 73776 87362 73804 93826
rect 74144 93006 74172 122687
rect 74236 117826 74264 127486
rect 74328 120585 74356 139182
rect 74408 137132 74460 137138
rect 74408 137074 74460 137080
rect 74420 127550 74448 137074
rect 74408 127544 74460 127550
rect 74408 127486 74460 127492
rect 74406 126424 74462 126433
rect 74406 126359 74462 126368
rect 74314 120576 74370 120585
rect 74314 120511 74370 120520
rect 74224 117820 74276 117826
rect 74224 117762 74276 117768
rect 74224 115100 74276 115106
rect 74224 115042 74276 115048
rect 74236 105489 74264 115042
rect 74420 109530 74448 126359
rect 76168 125102 76196 141886
rect 76156 125096 76208 125102
rect 76156 125038 76208 125044
rect 74408 109524 74460 109530
rect 74408 109466 74460 109472
rect 74222 105480 74278 105489
rect 74222 105415 74278 105424
rect 74222 105344 74278 105353
rect 74222 105279 74278 105288
rect 74236 98446 74264 105279
rect 74224 98440 74276 98446
rect 74224 98382 74276 98388
rect 74684 94360 74736 94366
rect 74682 94328 74684 94337
rect 74736 94328 74738 94337
rect 74682 94263 74738 94272
rect 74132 93000 74184 93006
rect 74132 92942 74184 92948
rect 76812 91306 76840 226902
rect 134760 225532 134812 225538
rect 134760 225474 134812 225480
rect 81674 219584 81730 219593
rect 81674 219519 81676 219528
rect 81728 219519 81730 219528
rect 81676 219490 81728 219496
rect 81676 203364 81728 203370
rect 81676 203306 81728 203312
rect 81688 202865 81716 203306
rect 81674 202856 81730 202865
rect 81674 202791 81730 202800
rect 81676 186840 81728 186846
rect 81676 186782 81728 186788
rect 81688 186273 81716 186782
rect 81674 186264 81730 186273
rect 81674 186199 81730 186208
rect 88404 175830 88432 177940
rect 88392 175824 88444 175830
rect 88392 175766 88444 175772
rect 95488 175762 95516 177940
rect 95476 175756 95528 175762
rect 95476 175698 95528 175704
rect 96764 175212 96816 175218
rect 96764 175154 96816 175160
rect 79192 170248 79244 170254
rect 79192 170190 79244 170196
rect 79204 169137 79232 170190
rect 79190 169128 79246 169137
rect 79190 169063 79246 169072
rect 77258 167700 77314 167709
rect 77258 167635 77314 167644
rect 77272 167602 77300 167635
rect 77260 167596 77312 167602
rect 77260 167538 77312 167544
rect 87196 167596 87248 167602
rect 87196 167538 87248 167544
rect 77258 166340 77314 166349
rect 77258 166275 77314 166284
rect 77272 166242 77300 166275
rect 77260 166236 77312 166242
rect 77260 166178 77312 166184
rect 87104 166236 87156 166242
rect 87104 166178 87156 166184
rect 77258 164844 77314 164853
rect 77258 164779 77260 164788
rect 77312 164779 77314 164788
rect 77260 164750 77312 164756
rect 77258 163484 77314 163493
rect 77258 163419 77260 163428
rect 77312 163419 77314 163428
rect 77260 163390 77312 163396
rect 87116 163153 87144 166178
rect 87208 164105 87236 167538
rect 87288 164808 87340 164814
rect 87288 164750 87340 164756
rect 87194 164096 87250 164105
rect 87194 164031 87250 164040
rect 87196 163448 87248 163454
rect 87196 163390 87248 163396
rect 87102 163144 87158 163153
rect 87102 163079 87158 163088
rect 77258 162124 77314 162133
rect 77258 162059 77314 162068
rect 77272 160598 77300 162059
rect 87208 161385 87236 163390
rect 87300 161929 87328 164750
rect 96776 163810 96804 175154
rect 102664 175150 102692 177940
rect 109748 175218 109776 177940
rect 116924 175218 116952 177940
rect 109736 175212 109788 175218
rect 109736 175154 109788 175160
rect 112680 175212 112732 175218
rect 112680 175154 112732 175160
rect 116912 175212 116964 175218
rect 116912 175154 116964 175160
rect 102652 175144 102704 175150
rect 102652 175086 102704 175092
rect 112692 166854 112720 175154
rect 124008 170254 124036 177940
rect 131184 174470 131212 177940
rect 129240 174464 129292 174470
rect 129240 174406 129292 174412
rect 131172 174464 131224 174470
rect 131172 174406 131224 174412
rect 123996 170248 124048 170254
rect 123996 170190 124048 170196
rect 124008 169574 124036 170190
rect 123996 169568 124048 169574
rect 123996 169510 124048 169516
rect 128136 168548 128188 168554
rect 128136 168490 128188 168496
rect 110196 166848 110248 166854
rect 110196 166790 110248 166796
rect 112680 166848 112732 166854
rect 112680 166790 112732 166796
rect 110208 163810 110236 166790
rect 123536 166576 123588 166582
rect 123536 166518 123588 166524
rect 123548 163810 123576 166518
rect 96560 163782 96804 163810
rect 109900 163782 110236 163810
rect 123240 163782 123576 163810
rect 87286 161920 87342 161929
rect 87286 161855 87342 161864
rect 87194 161376 87250 161385
rect 87194 161311 87250 161320
rect 77260 160592 77312 160598
rect 77260 160534 77312 160540
rect 87196 160592 87248 160598
rect 87196 160534 87248 160540
rect 87208 160433 87236 160534
rect 87194 160424 87250 160433
rect 87194 160359 87250 160368
rect 81766 160016 81822 160025
rect 81766 159951 81822 159960
rect 79282 159336 79338 159345
rect 79282 159271 79284 159280
rect 79336 159271 79338 159280
rect 79284 159242 79336 159248
rect 81780 159102 81808 159951
rect 87288 159164 87340 159170
rect 87288 159106 87340 159112
rect 81768 159096 81820 159102
rect 81768 159038 81820 159044
rect 87196 159096 87248 159102
rect 87196 159038 87248 159044
rect 87208 158937 87236 159038
rect 87194 158928 87250 158937
rect 87194 158863 87250 158872
rect 87300 158665 87328 159106
rect 87286 158656 87342 158665
rect 87286 158591 87342 158600
rect 79742 157976 79798 157985
rect 79742 157911 79744 157920
rect 79796 157911 79798 157920
rect 79744 157882 79796 157888
rect 87196 157804 87248 157810
rect 87196 157746 87248 157752
rect 87208 157713 87236 157746
rect 87194 157704 87250 157713
rect 87194 157639 87250 157648
rect 77258 156548 77314 156557
rect 77258 156483 77260 156492
rect 77312 156483 77314 156492
rect 77260 156454 77312 156460
rect 87196 156444 87248 156450
rect 87196 156386 87248 156392
rect 87208 156353 87236 156386
rect 87194 156344 87250 156353
rect 87194 156279 87250 156288
rect 87194 155392 87250 155401
rect 87194 155327 87250 155336
rect 79742 155120 79798 155129
rect 87208 155090 87236 155327
rect 79742 155055 79744 155064
rect 79796 155055 79798 155064
rect 87196 155084 87248 155090
rect 79744 155026 79796 155032
rect 87196 155026 87248 155032
rect 87194 154440 87250 154449
rect 81768 154404 81820 154410
rect 87194 154375 87196 154384
rect 81768 154346 81820 154352
rect 87248 154375 87250 154384
rect 87196 154346 87248 154352
rect 81780 153769 81808 154346
rect 81766 153760 81822 153769
rect 81766 153695 81822 153704
rect 87194 153624 87250 153633
rect 87194 153559 87250 153568
rect 87208 153050 87236 153559
rect 81768 153044 81820 153050
rect 81768 152986 81820 152992
rect 87196 153044 87248 153050
rect 87196 152986 87248 152992
rect 79744 152432 79796 152438
rect 81780 152409 81808 152986
rect 87194 152672 87250 152681
rect 87194 152607 87250 152616
rect 87208 152438 87236 152607
rect 87196 152432 87248 152438
rect 79744 152374 79796 152380
rect 81766 152400 81822 152409
rect 79756 150913 79784 152374
rect 87196 152374 87248 152380
rect 81766 152335 81822 152344
rect 88114 151856 88170 151865
rect 88114 151791 88170 151800
rect 79742 150904 79798 150913
rect 79742 150839 79798 150848
rect 87102 150904 87158 150913
rect 87102 150839 87158 150848
rect 80112 149644 80164 149650
rect 80112 149586 80164 149592
rect 79742 148184 79798 148193
rect 79742 148119 79744 148128
rect 79796 148119 79798 148128
rect 79744 148090 79796 148096
rect 80124 146697 80152 149586
rect 81768 149576 81820 149582
rect 81766 149544 81768 149553
rect 81820 149544 81822 149553
rect 81766 149479 81822 149488
rect 87116 148154 87144 150839
rect 87194 150088 87250 150097
rect 87194 150023 87250 150032
rect 87208 149650 87236 150023
rect 87196 149644 87248 149650
rect 87196 149586 87248 149592
rect 88128 149582 88156 151791
rect 88116 149576 88168 149582
rect 88116 149518 88168 149524
rect 87194 149136 87250 149145
rect 87194 149071 87250 149080
rect 87104 148148 87156 148154
rect 87104 148090 87156 148096
rect 80110 146688 80166 146697
rect 80110 146623 80166 146632
rect 87208 145434 87236 149071
rect 87286 148320 87342 148329
rect 87286 148255 87342 148264
rect 79744 145428 79796 145434
rect 79744 145370 79796 145376
rect 87196 145428 87248 145434
rect 87196 145370 87248 145376
rect 79756 145337 79784 145370
rect 79742 145328 79798 145337
rect 79742 145263 79798 145272
rect 87300 144074 87328 148255
rect 91670 147626 91698 147884
rect 95258 147762 95286 147884
rect 98938 147762 98966 147884
rect 95212 147734 95286 147762
rect 98892 147734 98966 147762
rect 91670 147598 91744 147626
rect 91716 145434 91744 147598
rect 91704 145428 91756 145434
rect 91704 145370 91756 145376
rect 91244 144748 91296 144754
rect 91244 144690 91296 144696
rect 79744 144068 79796 144074
rect 79744 144010 79796 144016
rect 87288 144068 87340 144074
rect 87288 144010 87340 144016
rect 79756 143977 79784 144010
rect 79742 143968 79798 143977
rect 79742 143903 79798 143912
rect 77258 142540 77314 142549
rect 77258 142475 77314 142484
rect 77272 141354 77300 142475
rect 82318 141656 82374 141665
rect 82318 141591 82374 141600
rect 77718 141520 77774 141529
rect 77718 141455 77774 141464
rect 77260 141348 77312 141354
rect 77260 141290 77312 141296
rect 77732 141286 77760 141455
rect 77720 141280 77772 141286
rect 77720 141222 77772 141228
rect 82332 140810 82360 141591
rect 82320 140804 82372 140810
rect 82320 140746 82372 140752
rect 91256 133754 91284 144690
rect 95212 144521 95240 147734
rect 98892 145201 98920 147734
rect 102526 147626 102554 147884
rect 106206 147762 106234 147884
rect 109794 147762 109822 147884
rect 102388 147598 102554 147626
rect 106160 147734 106234 147762
rect 109748 147734 109822 147762
rect 98878 145192 98934 145201
rect 98878 145127 98934 145136
rect 95198 144512 95254 144521
rect 95198 144447 95254 144456
rect 102388 140606 102416 147598
rect 103664 144816 103716 144822
rect 103664 144758 103716 144764
rect 102284 140600 102336 140606
rect 102376 140600 102428 140606
rect 102336 140560 102376 140588
rect 102284 140542 102336 140548
rect 102376 140542 102428 140548
rect 102388 140477 102416 140542
rect 103676 133754 103704 144758
rect 106160 142617 106188 147734
rect 109748 143161 109776 147734
rect 113474 147626 113502 147884
rect 117062 147626 117090 147884
rect 120742 147626 120770 147884
rect 124330 147626 124358 147884
rect 128024 147870 128084 147898
rect 113428 147598 113502 147626
rect 116188 147598 117090 147626
rect 120696 147598 120770 147626
rect 124284 147598 124358 147626
rect 109734 143152 109790 143161
rect 109734 143087 109790 143096
rect 106146 142608 106202 142617
rect 106146 142543 106202 142552
rect 113428 141286 113456 147598
rect 116084 144884 116136 144890
rect 116084 144826 116136 144832
rect 113416 141280 113468 141286
rect 113416 141222 113468 141228
rect 114704 141280 114756 141286
rect 114704 141222 114756 141228
rect 114716 140674 114744 141222
rect 114704 140668 114756 140674
rect 114704 140610 114756 140616
rect 116096 133754 116124 144826
rect 116188 139246 116216 147598
rect 120696 144754 120724 147598
rect 124284 144822 124312 147598
rect 128056 144890 128084 147870
rect 128148 145434 128176 168490
rect 129252 166582 129280 174406
rect 132184 168956 132236 168962
rect 132184 168898 132236 168904
rect 129240 166576 129292 166582
rect 129240 166518 129292 166524
rect 132092 166236 132144 166242
rect 132092 166178 132144 166184
rect 131356 163516 131408 163522
rect 131356 163458 131408 163464
rect 131368 163425 131396 163458
rect 131908 163448 131960 163454
rect 131354 163416 131410 163425
rect 131908 163390 131960 163396
rect 131354 163351 131410 163360
rect 131446 161648 131502 161657
rect 131446 161583 131502 161592
rect 131356 160728 131408 160734
rect 131354 160696 131356 160705
rect 131408 160696 131410 160705
rect 131460 160666 131488 161583
rect 131354 160631 131410 160640
rect 131448 160660 131500 160666
rect 131448 160602 131500 160608
rect 131354 159880 131410 159889
rect 131354 159815 131410 159824
rect 131368 159374 131396 159815
rect 131920 159458 131948 163390
rect 131998 162464 132054 162473
rect 131998 162399 132054 162408
rect 132012 162162 132040 162399
rect 132000 162156 132052 162162
rect 132000 162098 132052 162104
rect 132000 162020 132052 162026
rect 132000 161962 132052 161968
rect 131644 159430 131948 159458
rect 131356 159368 131408 159374
rect 131356 159310 131408 159316
rect 131644 152273 131672 159430
rect 131816 159300 131868 159306
rect 131816 159242 131868 159248
rect 131630 152264 131686 152273
rect 131630 152199 131686 152208
rect 131356 150936 131408 150942
rect 131356 150878 131408 150884
rect 131368 150505 131396 150878
rect 131354 150496 131410 150505
rect 131354 150431 131410 150440
rect 131356 149576 131408 149582
rect 131828 149553 131856 159242
rect 131908 159164 131960 159170
rect 131908 159106 131960 159112
rect 131920 153633 131948 159106
rect 132012 155129 132040 161962
rect 132104 159170 132132 166178
rect 132092 159164 132144 159170
rect 132092 159106 132144 159112
rect 132196 159050 132224 168898
rect 132276 167596 132328 167602
rect 132276 167538 132328 167544
rect 132288 162026 132316 167538
rect 132644 164808 132696 164814
rect 132644 164750 132696 164756
rect 132368 162088 132420 162094
rect 132368 162030 132420 162036
rect 132276 162020 132328 162026
rect 132276 161962 132328 161968
rect 132104 159022 132224 159050
rect 132104 156081 132132 159022
rect 132182 158928 132238 158937
rect 132182 158863 132238 158872
rect 132196 157946 132224 158863
rect 132184 157940 132236 157946
rect 132184 157882 132236 157888
rect 132274 157160 132330 157169
rect 132274 157095 132330 157104
rect 132090 156072 132146 156081
rect 132090 156007 132146 156016
rect 131998 155120 132054 155129
rect 131998 155055 132054 155064
rect 131906 153624 131962 153633
rect 131906 153559 131962 153568
rect 131356 149518 131408 149524
rect 131814 149544 131870 149553
rect 131368 148873 131396 149518
rect 131814 149479 131870 149488
rect 131354 148864 131410 148873
rect 131354 148799 131410 148808
rect 132288 145434 132316 157095
rect 132380 156466 132408 162030
rect 132550 158112 132606 158121
rect 132550 158047 132606 158056
rect 132380 156438 132500 156466
rect 132366 156344 132422 156353
rect 132366 156279 132422 156288
rect 128136 145428 128188 145434
rect 128136 145370 128188 145376
rect 132276 145428 132328 145434
rect 132276 145370 132328 145376
rect 128044 144884 128096 144890
rect 128044 144826 128096 144832
rect 124272 144816 124324 144822
rect 124272 144758 124324 144764
rect 120684 144748 120736 144754
rect 120684 144690 120736 144696
rect 132380 144074 132408 156279
rect 132472 150913 132500 156438
rect 132458 150904 132514 150913
rect 132458 150839 132514 150848
rect 132564 146794 132592 158047
rect 132656 153361 132684 164750
rect 132642 153352 132698 153361
rect 132642 153287 132698 153296
rect 132552 146788 132604 146794
rect 132552 146730 132604 146736
rect 132368 144068 132420 144074
rect 132368 144010 132420 144016
rect 127216 142028 127268 142034
rect 127216 141970 127268 141976
rect 127228 141354 127256 141970
rect 127216 141348 127268 141354
rect 127216 141290 127268 141296
rect 116176 139240 116228 139246
rect 116176 139182 116228 139188
rect 127228 134434 127256 141290
rect 127228 134406 128084 134434
rect 91086 133726 91284 133754
rect 103506 133726 103704 133754
rect 116018 133726 116124 133754
rect 128056 133618 128084 134406
rect 128056 133590 128530 133618
rect 76892 125504 76944 125510
rect 81676 125504 81728 125510
rect 76892 125446 76944 125452
rect 81674 125472 81676 125481
rect 81728 125472 81730 125481
rect 76904 125102 76932 125446
rect 81674 125407 81730 125416
rect 76892 125096 76944 125102
rect 76892 125038 76944 125044
rect 73856 91300 73908 91306
rect 73856 91242 73908 91248
rect 76800 91300 76852 91306
rect 76800 91242 76852 91248
rect 73868 91209 73896 91242
rect 73854 91200 73910 91209
rect 73854 91135 73910 91144
rect 73764 87356 73816 87362
rect 73764 87298 73816 87304
rect 73670 86304 73726 86313
rect 73670 86239 73726 86248
rect 73776 86177 73804 87298
rect 73486 86168 73542 86177
rect 73486 86103 73542 86112
rect 73762 86168 73818 86177
rect 73762 86103 73818 86112
rect 72842 85896 72898 85905
rect 72842 85831 72898 85840
rect 72660 78652 72712 78658
rect 72660 78594 72712 78600
rect 70740 75926 71136 75954
rect 71108 75818 71136 75926
rect 71108 75790 71674 75818
rect 72672 75804 72700 78594
rect 72856 76521 72884 85831
rect 74776 78856 74828 78862
rect 74776 78798 74828 78804
rect 73764 78380 73816 78386
rect 73764 78322 73816 78328
rect 72842 76512 72898 76521
rect 72842 76447 72898 76456
rect 73776 75804 73804 78322
rect 74788 75804 74816 78798
rect 76904 77910 76932 125038
rect 78178 110920 78234 110929
rect 78178 110855 78234 110864
rect 78192 109705 78220 110855
rect 78178 109696 78234 109705
rect 78178 109631 78234 109640
rect 78192 94366 78220 109631
rect 81676 109524 81728 109530
rect 81676 109466 81728 109472
rect 81688 108889 81716 109466
rect 81674 108880 81730 108889
rect 81674 108815 81730 108824
rect 78180 94360 78232 94366
rect 78180 94302 78232 94308
rect 75788 77904 75840 77910
rect 75788 77846 75840 77852
rect 76892 77904 76944 77910
rect 76892 77846 76944 77852
rect 75800 75804 75828 77846
rect 50040 75654 50974 75682
rect 51328 75654 51986 75682
rect 67888 75654 68546 75682
rect 78192 51526 78220 94302
rect 81676 93000 81728 93006
rect 81676 92942 81728 92948
rect 81688 92297 81716 92942
rect 81674 92288 81730 92297
rect 81674 92223 81730 92232
rect 88418 83814 88524 83842
rect 95502 83814 95792 83842
rect 102678 83814 102968 83842
rect 109762 83814 109868 83842
rect 116938 83814 117136 83842
rect 124022 83814 124128 83842
rect 131198 83814 131304 83842
rect 88496 81990 88524 83814
rect 88484 81984 88536 81990
rect 88484 81926 88536 81932
rect 95764 81922 95792 83814
rect 95752 81916 95804 81922
rect 95752 81858 95804 81864
rect 102940 81854 102968 83814
rect 102928 81848 102980 81854
rect 102928 81790 102980 81796
rect 109840 81310 109868 83814
rect 96764 81304 96816 81310
rect 96764 81246 96816 81252
rect 109828 81304 109880 81310
rect 109828 81246 109880 81252
rect 78916 76408 78968 76414
rect 78916 76350 78968 76356
rect 78928 75841 78956 76350
rect 78914 75832 78970 75841
rect 78914 75767 78970 75776
rect 78914 73928 78970 73937
rect 78914 73863 78970 73872
rect 78928 73762 78956 73863
rect 78916 73756 78968 73762
rect 78916 73698 78968 73704
rect 87380 73756 87432 73762
rect 87380 73698 87432 73704
rect 78914 72840 78970 72849
rect 78914 72775 78970 72784
rect 78928 72402 78956 72775
rect 78916 72396 78968 72402
rect 78916 72338 78968 72344
rect 87196 72396 87248 72402
rect 87196 72338 87248 72344
rect 78914 71616 78970 71625
rect 78914 71551 78970 71560
rect 78928 71042 78956 71551
rect 80202 71208 80258 71217
rect 80258 71166 80336 71194
rect 80202 71143 80258 71152
rect 78916 71036 78968 71042
rect 78916 70978 78968 70984
rect 78914 69848 78970 69857
rect 78914 69783 78970 69792
rect 78928 69614 78956 69783
rect 78916 69608 78968 69614
rect 78916 69550 78968 69556
rect 78914 68624 78970 68633
rect 78914 68559 78970 68568
rect 78928 68254 78956 68559
rect 78916 68248 78968 68254
rect 78916 68190 78968 68196
rect 79560 67568 79612 67574
rect 78914 67536 78970 67545
rect 79560 67510 79612 67516
rect 78914 67471 78970 67480
rect 78928 67098 78956 67471
rect 78916 67092 78968 67098
rect 78916 67034 78968 67040
rect 78916 66956 78968 66962
rect 78916 66898 78968 66904
rect 78928 66865 78956 66898
rect 78914 66856 78970 66865
rect 78914 66791 78970 66800
rect 78914 65632 78970 65641
rect 78914 65567 78970 65576
rect 78928 65466 78956 65567
rect 78916 65460 78968 65466
rect 78916 65402 78968 65408
rect 78914 64680 78970 64689
rect 78914 64615 78970 64624
rect 78928 64514 78956 64615
rect 78916 64508 78968 64514
rect 78916 64450 78968 64456
rect 78914 63456 78970 63465
rect 78914 63391 78970 63400
rect 78928 63018 78956 63391
rect 78916 63012 78968 63018
rect 78916 62954 78968 62960
rect 78914 62912 78970 62921
rect 78914 62847 78970 62856
rect 78928 62678 78956 62847
rect 78916 62672 78968 62678
rect 78916 62614 78968 62620
rect 78914 61552 78970 61561
rect 78914 61487 78970 61496
rect 78928 61386 78956 61487
rect 78916 61380 78968 61386
rect 78916 61322 78968 61328
rect 78914 60328 78970 60337
rect 78914 60263 78970 60272
rect 78928 59958 78956 60263
rect 78916 59952 78968 59958
rect 78916 59894 78968 59900
rect 78914 57336 78970 57345
rect 78914 57271 78970 57280
rect 78928 57170 78956 57271
rect 78916 57164 78968 57170
rect 78916 57106 78968 57112
rect 78914 56248 78970 56257
rect 78914 56183 78970 56192
rect 78928 55810 78956 56183
rect 78916 55804 78968 55810
rect 78916 55746 78968 55752
rect 79572 55713 79600 67510
rect 80308 66758 80336 71166
rect 85724 71036 85776 71042
rect 85724 70978 85776 70984
rect 84896 69608 84948 69614
rect 84896 69550 84948 69556
rect 81676 67092 81728 67098
rect 81676 67034 81728 67040
rect 80296 66752 80348 66758
rect 80296 66694 80348 66700
rect 81688 65398 81716 67034
rect 84908 66690 84936 69550
rect 85632 68248 85684 68254
rect 85632 68190 85684 68196
rect 85172 66956 85224 66962
rect 85172 66898 85224 66904
rect 84896 66684 84948 66690
rect 84896 66626 84948 66632
rect 84436 65460 84488 65466
rect 84436 65402 84488 65408
rect 81676 65392 81728 65398
rect 81676 65334 81728 65340
rect 81676 64508 81728 64514
rect 81676 64450 81728 64456
rect 81688 62610 81716 64450
rect 81768 63012 81820 63018
rect 81768 62954 81820 62960
rect 81676 62604 81728 62610
rect 81676 62546 81728 62552
rect 81676 61380 81728 61386
rect 81676 61322 81728 61328
rect 81688 59890 81716 61322
rect 81780 61250 81808 62954
rect 84448 62542 84476 65402
rect 85184 63630 85212 66898
rect 85644 65330 85672 68190
rect 85736 68186 85764 70978
rect 87208 68497 87236 72338
rect 87392 69449 87420 73698
rect 96776 69834 96804 81246
rect 117108 79354 117136 83814
rect 124100 83706 124128 83814
rect 116924 79326 117136 79354
rect 124008 83678 124128 83706
rect 116924 79218 116952 79326
rect 116832 79190 116952 79218
rect 116832 73490 116860 79190
rect 124008 76414 124036 83678
rect 131276 80630 131304 83814
rect 129240 80624 129292 80630
rect 129240 80566 129292 80572
rect 131264 80624 131316 80630
rect 131264 80566 131316 80572
rect 123996 76408 124048 76414
rect 123996 76350 124048 76356
rect 110196 73484 110248 73490
rect 110196 73426 110248 73432
rect 116820 73484 116872 73490
rect 116820 73426 116872 73432
rect 110208 69834 110236 73426
rect 129252 72402 129280 80566
rect 123536 72396 123588 72402
rect 123536 72338 123588 72344
rect 129240 72396 129292 72402
rect 129240 72338 129292 72344
rect 123548 69834 123576 72338
rect 96560 69806 96804 69834
rect 109900 69806 110236 69834
rect 123240 69806 123576 69834
rect 131448 69540 131500 69546
rect 131448 69482 131500 69488
rect 131356 69472 131408 69478
rect 87378 69440 87434 69449
rect 87378 69375 87434 69384
rect 131354 69440 131356 69449
rect 131408 69440 131410 69449
rect 131354 69375 131410 69384
rect 131460 68497 131488 69482
rect 87194 68488 87250 68497
rect 87194 68423 87250 68432
rect 131446 68488 131502 68497
rect 131446 68423 131502 68432
rect 85724 68180 85776 68186
rect 85724 68122 85776 68128
rect 87196 68180 87248 68186
rect 87196 68122 87248 68128
rect 132368 68180 132420 68186
rect 132368 68122 132420 68128
rect 87208 67681 87236 68122
rect 132380 67681 132408 68122
rect 87194 67672 87250 67681
rect 87194 67607 87250 67616
rect 132366 67672 132422 67681
rect 132366 67607 132422 67616
rect 129424 67568 129476 67574
rect 129424 67510 129476 67516
rect 129436 66758 129464 67510
rect 87196 66752 87248 66758
rect 87194 66720 87196 66729
rect 129424 66752 129476 66758
rect 87248 66720 87250 66729
rect 132368 66752 132420 66758
rect 129424 66694 129476 66700
rect 131354 66720 131410 66729
rect 87194 66655 87250 66664
rect 87288 66684 87340 66690
rect 132368 66694 132420 66700
rect 131354 66655 131356 66664
rect 87288 66626 87340 66632
rect 131408 66655 131410 66664
rect 131356 66626 131408 66632
rect 87300 65913 87328 66626
rect 132380 65913 132408 66694
rect 87286 65904 87342 65913
rect 87286 65839 87342 65848
rect 132366 65904 132422 65913
rect 132366 65839 132422 65848
rect 87196 65392 87248 65398
rect 87196 65334 87248 65340
rect 131448 65392 131500 65398
rect 131448 65334 131500 65340
rect 85632 65324 85684 65330
rect 85632 65266 85684 65272
rect 87208 64145 87236 65334
rect 87288 65324 87340 65330
rect 87288 65266 87340 65272
rect 131356 65324 131408 65330
rect 131356 65266 131408 65272
rect 87300 64961 87328 65266
rect 131368 64961 131396 65266
rect 87286 64952 87342 64961
rect 87286 64887 87342 64896
rect 131354 64952 131410 64961
rect 131354 64887 131410 64896
rect 131460 64145 131488 65334
rect 87194 64136 87250 64145
rect 87194 64071 87250 64080
rect 131446 64136 131502 64145
rect 131446 64071 131502 64080
rect 132368 64032 132420 64038
rect 132368 63974 132420 63980
rect 85172 63624 85224 63630
rect 85172 63566 85224 63572
rect 87196 63624 87248 63630
rect 87196 63566 87248 63572
rect 87208 63193 87236 63566
rect 132380 63193 132408 63974
rect 87194 63184 87250 63193
rect 87194 63119 87250 63128
rect 132366 63184 132422 63193
rect 132366 63119 132422 63128
rect 87380 62672 87432 62678
rect 87380 62614 87432 62620
rect 87196 62604 87248 62610
rect 87196 62546 87248 62552
rect 84436 62536 84488 62542
rect 84436 62478 84488 62484
rect 87208 61425 87236 62546
rect 87288 62536 87340 62542
rect 87288 62478 87340 62484
rect 87300 62377 87328 62478
rect 87286 62368 87342 62377
rect 87286 62303 87342 62312
rect 87194 61416 87250 61425
rect 87194 61351 87250 61360
rect 81768 61244 81820 61250
rect 81768 61186 81820 61192
rect 87196 61244 87248 61250
rect 87196 61186 87248 61192
rect 87208 60473 87236 61186
rect 87194 60464 87250 60473
rect 87194 60399 87250 60408
rect 85724 59952 85776 59958
rect 85724 59894 85776 59900
rect 81676 59884 81728 59890
rect 81676 59826 81728 59832
rect 80202 59104 80258 59113
rect 80258 59062 80428 59090
rect 80202 59039 80258 59048
rect 80202 58560 80258 58569
rect 80258 58518 80336 58546
rect 80202 58495 80258 58504
rect 80308 57034 80336 58518
rect 80400 57102 80428 59062
rect 85736 58530 85764 59894
rect 87196 59884 87248 59890
rect 87196 59826 87248 59832
rect 87208 58705 87236 59826
rect 87392 59657 87420 62614
rect 131724 62604 131776 62610
rect 131724 62546 131776 62552
rect 131356 62536 131408 62542
rect 131356 62478 131408 62484
rect 131368 62377 131396 62478
rect 131354 62368 131410 62377
rect 131354 62303 131410 62312
rect 131736 61425 131764 62546
rect 131722 61416 131778 61425
rect 131722 61351 131778 61360
rect 131356 61244 131408 61250
rect 131356 61186 131408 61192
rect 131368 60473 131396 61186
rect 131354 60464 131410 60473
rect 131354 60399 131410 60408
rect 132644 59884 132696 59890
rect 132644 59826 132696 59832
rect 132552 59816 132604 59822
rect 132552 59758 132604 59764
rect 87378 59648 87434 59657
rect 87378 59583 87434 59592
rect 132564 58705 132592 59758
rect 132656 59657 132684 59826
rect 132642 59648 132698 59657
rect 132642 59583 132698 59592
rect 87194 58696 87250 58705
rect 87194 58631 87250 58640
rect 132550 58696 132606 58705
rect 132550 58631 132606 58640
rect 85724 58524 85776 58530
rect 85724 58466 85776 58472
rect 87196 58524 87248 58530
rect 87196 58466 87248 58472
rect 132644 58524 132696 58530
rect 132644 58466 132696 58472
rect 87208 57889 87236 58466
rect 132656 57889 132684 58466
rect 87194 57880 87250 57889
rect 87194 57815 87250 57824
rect 132642 57880 132698 57889
rect 132642 57815 132698 57824
rect 87380 57164 87432 57170
rect 87380 57106 87432 57112
rect 129516 57164 129568 57170
rect 129516 57106 129568 57112
rect 80388 57096 80440 57102
rect 80388 57038 80440 57044
rect 87196 57096 87248 57102
rect 87196 57038 87248 57044
rect 80296 57028 80348 57034
rect 80296 56970 80348 56976
rect 87208 56937 87236 57038
rect 87288 57028 87340 57034
rect 87288 56970 87340 56976
rect 87194 56928 87250 56937
rect 87194 56863 87250 56872
rect 87300 56121 87328 56970
rect 87286 56112 87342 56121
rect 87286 56047 87342 56056
rect 81676 55804 81728 55810
rect 81676 55746 81728 55752
rect 79558 55704 79614 55713
rect 79558 55639 79614 55648
rect 78914 54616 78970 54625
rect 78914 54551 78970 54560
rect 78928 54450 78956 54551
rect 78916 54444 78968 54450
rect 78916 54386 78968 54392
rect 81688 54382 81716 55746
rect 87392 55169 87420 57106
rect 87378 55160 87434 55169
rect 87378 55095 87434 55104
rect 129528 54926 129556 57106
rect 132644 57096 132696 57102
rect 132644 57038 132696 57044
rect 132552 57028 132604 57034
rect 132552 56970 132604 56976
rect 132564 56121 132592 56970
rect 132656 56937 132684 57038
rect 132642 56928 132698 56937
rect 132642 56863 132698 56872
rect 132550 56112 132606 56121
rect 132550 56047 132606 56056
rect 132644 55736 132696 55742
rect 132644 55678 132696 55684
rect 132656 55169 132684 55678
rect 132642 55160 132698 55169
rect 132642 55095 132698 55104
rect 134206 55160 134262 55169
rect 134206 55095 134208 55104
rect 134260 55095 134262 55104
rect 134208 55066 134260 55072
rect 129516 54920 129568 54926
rect 129516 54862 129568 54868
rect 87288 54444 87340 54450
rect 87288 54386 87340 54392
rect 81676 54376 81728 54382
rect 87196 54376 87248 54382
rect 81676 54318 81728 54324
rect 87194 54344 87196 54353
rect 87248 54344 87250 54353
rect 87194 54279 87250 54288
rect 78916 53764 78968 53770
rect 78916 53706 78968 53712
rect 78928 53673 78956 53706
rect 87300 53702 87328 54386
rect 100424 54030 100484 54058
rect 91040 53894 91284 53922
rect 93340 53894 93676 53922
rect 95732 53894 95792 53922
rect 98032 53894 98092 53922
rect 87288 53696 87340 53702
rect 78914 53664 78970 53673
rect 87288 53638 87340 53644
rect 78914 53599 78970 53608
rect 91256 51594 91284 53894
rect 91244 51588 91296 51594
rect 91244 51530 91296 51536
rect 93648 51526 93676 53894
rect 78180 51520 78232 51526
rect 78180 51462 78232 51468
rect 93636 51520 93688 51526
rect 93636 51462 93688 51468
rect 91244 50908 91296 50914
rect 91244 50850 91296 50856
rect 79006 50808 79062 50817
rect 79006 50743 79062 50752
rect 79020 50370 79048 50743
rect 79008 50364 79060 50370
rect 79008 50306 79060 50312
rect 78916 50296 78968 50302
rect 78914 50264 78916 50273
rect 78968 50264 78970 50273
rect 78914 50199 78970 50208
rect 87472 49548 87524 49554
rect 87472 49490 87524 49496
rect 88392 49548 88444 49554
rect 88392 49490 88444 49496
rect 87484 49321 87512 49490
rect 87470 49312 87526 49321
rect 87470 49247 87526 49256
rect 78914 49176 78970 49185
rect 78914 49111 78970 49120
rect 78928 48942 78956 49111
rect 78916 48936 78968 48942
rect 78916 48878 78968 48884
rect 67874 48088 67930 48097
rect 67718 48046 67874 48074
rect 67874 48023 67930 48032
rect 74314 48088 74370 48097
rect 74314 48023 74370 48032
rect 87102 48088 87158 48097
rect 87102 48023 87158 48032
rect 88298 48088 88354 48097
rect 88298 48023 88354 48032
rect 16540 47440 16592 47446
rect 16540 47382 16592 47388
rect 50224 46086 50252 47924
rect 50212 46080 50264 46086
rect 50212 46022 50264 46028
rect 53720 46018 53748 47924
rect 53708 46012 53760 46018
rect 53708 45954 53760 45960
rect 57216 45950 57244 47924
rect 60712 47446 60740 47924
rect 60700 47440 60752 47446
rect 60700 47382 60752 47388
rect 57204 45944 57256 45950
rect 64208 45921 64236 47924
rect 71200 46222 71228 47924
rect 72568 47440 72620 47446
rect 72566 47408 72568 47417
rect 73304 47440 73356 47446
rect 72620 47408 72622 47417
rect 73304 47382 73356 47388
rect 72566 47343 72622 47352
rect 71188 46216 71240 46222
rect 71188 46158 71240 46164
rect 73316 46154 73344 47382
rect 74328 46222 74356 48023
rect 74696 47417 74724 47924
rect 74682 47408 74738 47417
rect 74682 47343 74738 47352
rect 74696 46766 74724 47343
rect 87116 47242 87144 48023
rect 87104 47236 87156 47242
rect 87104 47178 87156 47184
rect 88024 46828 88076 46834
rect 88024 46770 88076 46776
rect 74684 46760 74736 46766
rect 74684 46702 74736 46708
rect 87196 46760 87248 46766
rect 87196 46702 87248 46708
rect 74316 46216 74368 46222
rect 74316 46158 74368 46164
rect 87208 46154 87236 46702
rect 73304 46148 73356 46154
rect 73304 46090 73356 46096
rect 87196 46148 87248 46154
rect 87196 46090 87248 46096
rect 57204 45886 57256 45892
rect 64194 45912 64250 45921
rect 64194 45847 64250 45856
rect 16448 36356 16500 36362
rect 16448 36298 16500 36304
rect 16264 25000 16316 25006
rect 16264 24942 16316 24948
rect 88036 23345 88064 46770
rect 88208 46216 88260 46222
rect 88208 46158 88260 46164
rect 88116 46148 88168 46154
rect 88116 46090 88168 46096
rect 88128 33681 88156 46090
rect 88114 33672 88170 33681
rect 88114 33607 88170 33616
rect 88220 30825 88248 46158
rect 88206 30816 88262 30825
rect 88206 30751 88262 30760
rect 88312 28105 88340 48023
rect 88298 28096 88354 28105
rect 88298 28031 88354 28040
rect 88404 26065 88432 49490
rect 91256 34746 91284 50850
rect 93648 50681 93676 51462
rect 93634 50672 93690 50681
rect 93634 50607 93690 50616
rect 93636 47236 93688 47242
rect 93636 47178 93688 47184
rect 93648 34746 93676 47178
rect 95476 46012 95528 46018
rect 95476 45954 95528 45960
rect 95488 45882 95516 45954
rect 95764 45882 95792 53894
rect 96764 48528 96816 48534
rect 96764 48470 96816 48476
rect 95476 45876 95528 45882
rect 95476 45818 95528 45824
rect 95752 45876 95804 45882
rect 95752 45818 95804 45824
rect 96776 37518 96804 48470
rect 98064 45950 98092 53894
rect 98604 48936 98656 48942
rect 98604 48878 98656 48884
rect 98052 45944 98104 45950
rect 98052 45886 98104 45892
rect 96396 37512 96448 37518
rect 96396 37454 96448 37460
rect 96764 37512 96816 37518
rect 96764 37454 96816 37460
rect 96408 34746 96436 37454
rect 98616 34746 98644 48878
rect 100456 47514 100484 54030
rect 102388 53894 102724 53922
rect 105116 53894 105176 53922
rect 107508 53894 107568 53922
rect 102388 51361 102416 53894
rect 102374 51352 102430 51361
rect 102374 51287 102430 51296
rect 102284 51044 102336 51050
rect 102284 50986 102336 50992
rect 100444 47508 100496 47514
rect 100444 47450 100496 47456
rect 100904 47508 100956 47514
rect 100904 47450 100956 47456
rect 100916 46834 100944 47450
rect 100904 46828 100956 46834
rect 100904 46770 100956 46776
rect 102296 37790 102324 50986
rect 102388 49554 102416 51287
rect 103572 50296 103624 50302
rect 103572 50238 103624 50244
rect 102376 49548 102428 49554
rect 102376 49490 102428 49496
rect 101364 37784 101416 37790
rect 101364 37726 101416 37732
rect 102284 37784 102336 37790
rect 102284 37726 102336 37732
rect 101376 34746 101404 37726
rect 103584 34746 103612 50238
rect 105148 49321 105176 53894
rect 106424 51112 106476 51118
rect 106424 51054 106476 51060
rect 105134 49312 105190 49321
rect 105134 49247 105190 49256
rect 105148 48097 105176 49247
rect 105134 48088 105190 48097
rect 105134 48023 105190 48032
rect 106436 34746 106464 51054
rect 107540 50273 107568 53894
rect 109472 53894 109808 53922
rect 112048 53894 112200 53922
rect 114164 53894 114500 53922
rect 116556 53894 116892 53922
rect 118948 53894 119284 53922
rect 121248 53894 121584 53922
rect 123640 53894 123976 53922
rect 125940 53894 126276 53922
rect 108632 50364 108684 50370
rect 108632 50306 108684 50312
rect 107526 50264 107582 50273
rect 107526 50199 107582 50208
rect 106606 47408 106662 47417
rect 106606 47343 106662 47352
rect 106620 46222 106648 47343
rect 106608 46216 106660 46222
rect 106608 46158 106660 46164
rect 108644 34746 108672 50306
rect 109472 50273 109500 53894
rect 111944 51180 111996 51186
rect 111944 51122 111996 51128
rect 109458 50264 109514 50273
rect 109458 50199 109514 50208
rect 109458 47272 109514 47281
rect 109458 47207 109514 47216
rect 109472 46154 109500 47207
rect 109460 46148 109512 46154
rect 109460 46090 109512 46096
rect 111956 36702 111984 51122
rect 112048 50914 112076 53894
rect 114164 50982 114192 53894
rect 116556 51050 116584 53894
rect 118200 53764 118252 53770
rect 118200 53706 118252 53712
rect 118212 53129 118240 53706
rect 118198 53120 118254 53129
rect 118198 53055 118254 53064
rect 118948 51118 118976 53894
rect 121248 51186 121276 53894
rect 121236 51180 121288 51186
rect 121236 51122 121288 51128
rect 118936 51112 118988 51118
rect 118936 51054 118988 51060
rect 116544 51044 116596 51050
rect 116544 50986 116596 50992
rect 114152 50976 114204 50982
rect 114152 50918 114204 50924
rect 122340 50976 122392 50982
rect 122340 50918 122392 50924
rect 112036 50908 112088 50914
rect 112036 50850 112088 50856
rect 116084 50908 116136 50914
rect 116084 50850 116136 50856
rect 113598 47544 113654 47553
rect 113598 47479 113654 47488
rect 111392 36696 111444 36702
rect 111392 36638 111444 36644
rect 111944 36696 111996 36702
rect 111944 36638 111996 36644
rect 111404 34746 111432 36638
rect 113612 34746 113640 47479
rect 116096 34746 116124 50850
rect 118658 44688 118714 44697
rect 118658 44623 118714 44632
rect 118672 34746 118700 44623
rect 122352 37314 122380 50918
rect 123640 50914 123668 53894
rect 125940 50982 125968 53894
rect 128654 53786 128682 53908
rect 128608 53758 128682 53786
rect 125928 50976 125980 50982
rect 125928 50918 125980 50924
rect 123628 50908 123680 50914
rect 123628 50850 123680 50856
rect 128608 37654 128636 53758
rect 128688 53696 128740 53702
rect 128688 53638 128740 53644
rect 126388 37648 126440 37654
rect 126388 37590 126440 37596
rect 128596 37648 128648 37654
rect 128596 37590 128648 37596
rect 121420 37308 121472 37314
rect 121420 37250 121472 37256
rect 122340 37308 122392 37314
rect 122340 37250 122392 37256
rect 121432 34746 121460 37250
rect 123904 36764 123956 36770
rect 123904 36706 123956 36712
rect 123916 34746 123944 36706
rect 126400 34746 126428 37590
rect 128700 36770 128728 53638
rect 129528 52342 129556 54862
rect 134116 54444 134168 54450
rect 134116 54386 134168 54392
rect 132644 54376 132696 54382
rect 132642 54344 132644 54353
rect 132696 54344 132698 54353
rect 132642 54279 132698 54288
rect 134128 53702 134156 54386
rect 134116 53696 134168 53702
rect 134116 53638 134168 53644
rect 129056 52336 129108 52342
rect 129056 52278 129108 52284
rect 129516 52336 129568 52342
rect 129516 52278 129568 52284
rect 128688 36764 128740 36770
rect 128688 36706 128740 36712
rect 91132 34718 91284 34746
rect 93616 34718 93676 34746
rect 96100 34718 96436 34746
rect 98584 34718 98644 34746
rect 101068 34718 101404 34746
rect 103552 34718 103612 34746
rect 106128 34718 106464 34746
rect 108612 34718 108672 34746
rect 111096 34718 111432 34746
rect 113580 34718 113640 34746
rect 116064 34718 116124 34746
rect 118640 34718 118700 34746
rect 121124 34718 121460 34746
rect 123608 34718 123944 34746
rect 126092 34718 126428 34746
rect 129068 34610 129096 52278
rect 134772 51594 134800 225474
rect 136888 204882 136916 282215
rect 137532 275178 137560 304655
rect 137624 298609 137652 326930
rect 137716 326246 137744 327474
rect 137704 326240 137756 326246
rect 137704 326182 137756 326188
rect 137796 316652 137848 316658
rect 137796 316594 137848 316600
rect 137808 311150 137836 316594
rect 137796 311144 137848 311150
rect 137796 311086 137848 311092
rect 137704 309716 137756 309722
rect 137704 309658 137756 309664
rect 137610 298600 137666 298609
rect 137610 298535 137666 298544
rect 137610 285272 137666 285281
rect 137610 285207 137666 285216
rect 137520 275172 137572 275178
rect 137520 275114 137572 275120
rect 137532 273857 137560 275114
rect 137518 273848 137574 273857
rect 137518 273783 137574 273792
rect 137520 254500 137572 254506
rect 137520 254442 137572 254448
rect 137532 244782 137560 254442
rect 137520 244776 137572 244782
rect 137520 244718 137572 244724
rect 136968 238656 137020 238662
rect 136966 238624 136968 238633
rect 137020 238624 137022 238633
rect 137022 238582 137100 238610
rect 136966 238559 137022 238568
rect 136966 235768 137022 235777
rect 136966 235703 137022 235712
rect 136980 235262 137008 235703
rect 136968 235256 137020 235262
rect 136968 235198 137020 235204
rect 136966 235088 137022 235097
rect 136966 235023 137022 235032
rect 136980 210753 137008 235023
rect 137072 213881 137100 238582
rect 137152 235256 137204 235262
rect 137152 235198 137204 235204
rect 137164 233306 137192 235198
rect 137336 234508 137388 234514
rect 137336 234450 137388 234456
rect 137164 233278 137284 233306
rect 137164 233086 137192 233117
rect 137152 233080 137204 233086
rect 137150 233048 137152 233057
rect 137204 233048 137206 233057
rect 137150 232983 137206 232992
rect 137164 217009 137192 232983
rect 137256 220137 137284 233278
rect 137348 223265 137376 234450
rect 137624 226150 137652 285207
rect 137716 279705 137744 309658
rect 137796 295912 137848 295918
rect 137796 295854 137848 295860
rect 137702 279696 137758 279705
rect 137702 279631 137758 279640
rect 137808 276577 137836 295854
rect 141660 283536 141712 283542
rect 141660 283478 141712 283484
rect 138622 278200 138678 278209
rect 138622 278135 138678 278144
rect 137794 276568 137850 276577
rect 137794 276503 137850 276512
rect 138636 275110 138664 278135
rect 138624 275104 138676 275110
rect 138624 275046 138676 275052
rect 138072 273744 138124 273750
rect 138072 273686 138124 273692
rect 138084 273449 138112 273686
rect 138070 273440 138126 273449
rect 138070 273375 138126 273384
rect 138636 269777 138664 275046
rect 141672 273750 141700 283478
rect 142408 282386 142436 329838
rect 144616 326722 144644 329838
rect 144604 326716 144656 326722
rect 144604 326658 144656 326664
rect 145536 326654 145564 329838
rect 145904 329838 146240 329866
rect 147160 329838 147496 329866
rect 148172 329838 148508 329866
rect 145524 326648 145576 326654
rect 145524 326590 145576 326596
rect 145904 326382 145932 329838
rect 147468 326382 147496 329838
rect 148480 326518 148508 329838
rect 148756 329838 149092 329866
rect 150104 329838 150440 329866
rect 151024 329838 151360 329866
rect 152036 329838 152372 329866
rect 152956 329838 153292 329866
rect 153968 329838 154304 329866
rect 148468 326512 148520 326518
rect 148468 326454 148520 326460
rect 148756 326450 148784 329838
rect 149388 327260 149440 327266
rect 149388 327202 149440 327208
rect 147916 326444 147968 326450
rect 147916 326386 147968 326392
rect 148744 326444 148796 326450
rect 148744 326386 148796 326392
rect 145156 326376 145208 326382
rect 145156 326318 145208 326324
rect 145892 326376 145944 326382
rect 145892 326318 145944 326324
rect 147456 326376 147508 326382
rect 147456 326318 147508 326324
rect 145168 319922 145196 326318
rect 147928 320058 147956 326386
rect 149296 320120 149348 320126
rect 149296 320062 149348 320068
rect 147916 320052 147968 320058
rect 147916 319994 147968 320000
rect 145156 319916 145208 319922
rect 145156 319858 145208 319864
rect 149308 316796 149336 320062
rect 149400 318578 149428 327202
rect 150412 326586 150440 329838
rect 151332 327334 151360 329838
rect 151964 327396 152016 327402
rect 151964 327338 152016 327344
rect 151320 327328 151372 327334
rect 151320 327270 151372 327276
rect 150768 327124 150820 327130
rect 150768 327066 150820 327072
rect 150400 326580 150452 326586
rect 150400 326522 150452 326528
rect 149400 318550 149796 318578
rect 149768 316810 149796 318550
rect 150780 316810 150808 327066
rect 149768 316782 150150 316810
rect 150780 316782 151070 316810
rect 151976 316796 152004 327338
rect 152056 326784 152108 326790
rect 152056 326726 152108 326732
rect 152068 319378 152096 326726
rect 152344 326450 152372 329838
rect 153264 327062 153292 329838
rect 154172 327192 154224 327198
rect 154172 327134 154224 327140
rect 153252 327056 153304 327062
rect 153252 326998 153304 327004
rect 153528 326852 153580 326858
rect 153528 326794 153580 326800
rect 152332 326444 152384 326450
rect 152332 326386 152384 326392
rect 152056 319372 152108 319378
rect 152056 319314 152108 319320
rect 152792 319372 152844 319378
rect 152792 319314 152844 319320
rect 152804 316796 152832 319314
rect 153540 316810 153568 326794
rect 154184 316946 154212 327134
rect 154276 326926 154304 329838
rect 154874 329594 154902 329852
rect 154828 329566 154902 329594
rect 154828 327470 154856 329566
rect 155932 327538 155960 329974
rect 156852 327606 156880 329974
rect 157832 329838 158260 329866
rect 160684 329838 160744 329866
rect 161696 329838 161756 329866
rect 158232 329238 158260 329838
rect 158220 329232 158272 329238
rect 158220 329174 158272 329180
rect 158232 329102 158260 329174
rect 158220 329096 158272 329102
rect 158220 329038 158272 329044
rect 160716 328121 160744 329838
rect 161728 328801 161756 329838
rect 162280 329838 162616 329866
rect 163292 329838 163628 329866
rect 164548 329838 164608 329866
rect 161714 328792 161770 328801
rect 161714 328727 161770 328736
rect 160702 328112 160758 328121
rect 160702 328047 160758 328056
rect 156288 327600 156340 327606
rect 156288 327542 156340 327548
rect 156840 327600 156892 327606
rect 156840 327542 156892 327548
rect 155920 327532 155972 327538
rect 155920 327474 155972 327480
rect 154816 327464 154868 327470
rect 154816 327406 154868 327412
rect 154828 326994 154856 327406
rect 154816 326988 154868 326994
rect 154816 326930 154868 326936
rect 154908 326988 154960 326994
rect 154908 326930 154960 326936
rect 154264 326920 154316 326926
rect 154264 326862 154316 326868
rect 154920 316946 154948 326930
rect 155552 326716 155604 326722
rect 155552 326658 155604 326664
rect 156196 326716 156248 326722
rect 156196 326658 156248 326664
rect 155564 319378 155592 326658
rect 155552 319372 155604 319378
rect 155552 319314 155604 319320
rect 154184 316918 154396 316946
rect 154920 316918 155132 316946
rect 154368 316810 154396 316918
rect 155104 316810 155132 316918
rect 156208 316810 156236 326658
rect 156300 326314 156328 327542
rect 157576 326648 157628 326654
rect 157576 326590 157628 326596
rect 156932 326376 156984 326382
rect 156932 326318 156984 326324
rect 156288 326308 156340 326314
rect 156288 326250 156340 326256
rect 156944 320262 156972 326318
rect 156932 320256 156984 320262
rect 156932 320198 156984 320204
rect 157300 319372 157352 319378
rect 157300 319314 157352 319320
rect 153540 316782 153738 316810
rect 154368 316782 154658 316810
rect 155104 316782 155486 316810
rect 156208 316782 156406 316810
rect 157312 316796 157340 319314
rect 157588 316946 157616 326590
rect 161624 326580 161676 326586
rect 161624 326522 161676 326528
rect 160244 326512 160296 326518
rect 160244 326454 160296 326460
rect 159968 320256 160020 320262
rect 159968 320198 160020 320204
rect 159048 319780 159100 319786
rect 159048 319722 159100 319728
rect 157588 316918 157892 316946
rect 157864 316810 157892 316918
rect 157864 316782 158154 316810
rect 159060 316796 159088 319722
rect 159980 316796 160008 320198
rect 160256 319394 160284 326454
rect 161532 326308 161584 326314
rect 161532 326250 161584 326256
rect 161544 320126 161572 326250
rect 161532 320120 161584 320126
rect 161532 320062 161584 320068
rect 160256 319366 160468 319394
rect 161636 319378 161664 326522
rect 162280 326314 162308 329838
rect 163188 327328 163240 327334
rect 163188 327270 163240 327276
rect 163096 326444 163148 326450
rect 163096 326386 163148 326392
rect 162268 326308 162320 326314
rect 162268 326250 162320 326256
rect 161716 319916 161768 319922
rect 161716 319858 161768 319864
rect 160440 316810 160468 319366
rect 161624 319372 161676 319378
rect 161624 319314 161676 319320
rect 160440 316782 160822 316810
rect 161728 316796 161756 319858
rect 162636 319372 162688 319378
rect 162636 319314 162688 319320
rect 162648 316796 162676 319314
rect 163108 318562 163136 326386
rect 163096 318556 163148 318562
rect 163096 318498 163148 318504
rect 163200 316810 163228 327270
rect 163292 327266 163320 329838
rect 163280 327260 163332 327266
rect 163280 327202 163332 327208
rect 164580 327130 164608 329838
rect 165224 329838 165560 329866
rect 166144 329838 166480 329866
rect 167340 329838 167492 329866
rect 168076 329838 168412 329866
rect 169088 329838 169424 329866
rect 170008 329838 170344 329866
rect 165224 327402 165252 329838
rect 165212 327396 165264 327402
rect 165212 327338 165264 327344
rect 164568 327124 164620 327130
rect 164568 327066 164620 327072
rect 165120 327056 165172 327062
rect 165120 326998 165172 327004
rect 164108 318556 164160 318562
rect 164108 318498 164160 318504
rect 164120 316810 164148 318498
rect 163200 316782 163490 316810
rect 164120 316782 164410 316810
rect 165132 313122 165160 326998
rect 166144 326790 166172 329838
rect 167340 326858 167368 329838
rect 168076 327198 168104 329838
rect 168064 327192 168116 327198
rect 168064 327134 168116 327140
rect 167328 326852 167380 326858
rect 167328 326794 167380 326800
rect 166132 326784 166184 326790
rect 166132 326726 166184 326732
rect 169088 326654 169116 329838
rect 170008 326722 170036 329838
rect 172124 329102 172152 330223
rect 172112 329096 172164 329102
rect 172112 329038 172164 329044
rect 169996 326716 170048 326722
rect 169996 326658 170048 326664
rect 169076 326648 169128 326654
rect 169076 326590 169128 326596
rect 185096 321692 185124 333798
rect 185924 333794 185952 335822
rect 185912 333788 185964 333794
rect 185912 333730 185964 333736
rect 187948 326994 187976 335958
rect 192088 327470 192116 335958
rect 194848 327606 194876 335958
rect 197504 333924 197556 333930
rect 197504 333866 197556 333872
rect 194836 327600 194888 327606
rect 194836 327542 194888 327548
rect 192076 327464 192128 327470
rect 192076 327406 192128 327412
rect 194848 327130 194876 327542
rect 194836 327124 194888 327130
rect 194836 327066 194888 327072
rect 187936 326988 187988 326994
rect 187936 326930 187988 326936
rect 197516 321692 197544 333866
rect 198712 331754 198740 336094
rect 201840 335958 202222 335986
rect 208740 335958 208846 335986
rect 218584 335958 218874 335986
rect 221896 335958 222186 335986
rect 201840 333153 201868 335958
rect 205534 335822 205640 335850
rect 201826 333144 201882 333153
rect 201826 333079 201882 333088
rect 201840 332201 201868 333079
rect 201826 332192 201882 332201
rect 201826 332127 201882 332136
rect 198700 331748 198752 331754
rect 198700 331690 198752 331696
rect 198712 330410 198740 331690
rect 205612 331657 205640 335822
rect 205598 331648 205654 331657
rect 205598 331583 205654 331592
rect 198712 330382 198924 330410
rect 198896 329170 198924 330382
rect 198884 329164 198936 329170
rect 198884 329106 198936 329112
rect 208740 328966 208768 335958
rect 212250 335822 212356 335850
rect 215562 335822 215668 335850
rect 212328 334474 212356 335822
rect 212316 334468 212368 334474
rect 212316 334410 212368 334416
rect 211304 333992 211356 333998
rect 211304 333934 211356 333940
rect 208728 328960 208780 328966
rect 208728 328902 208780 328908
rect 208740 328121 208768 328902
rect 208726 328112 208782 328121
rect 208726 328047 208782 328056
rect 211316 323526 211344 333934
rect 212328 333561 212356 334410
rect 215640 333862 215668 335822
rect 218584 333930 218612 335958
rect 221896 333998 221924 335958
rect 221884 333992 221936 333998
rect 221884 333934 221936 333940
rect 218572 333924 218624 333930
rect 218572 333866 218624 333872
rect 215628 333856 215680 333862
rect 215628 333798 215680 333804
rect 212314 333552 212370 333561
rect 212314 333487 212370 333496
rect 222528 329096 222580 329102
rect 222528 329038 222580 329044
rect 210016 323520 210068 323526
rect 210016 323462 210068 323468
rect 211304 323520 211356 323526
rect 211304 323462 211356 323468
rect 210028 321692 210056 323462
rect 222540 321692 222568 329038
rect 225208 328966 225236 382039
rect 225300 334270 225328 384759
rect 225378 380200 225434 380209
rect 225378 380135 225434 380144
rect 225288 334264 225340 334270
rect 225288 334206 225340 334212
rect 225392 331657 225420 380135
rect 315644 378554 315672 388334
rect 319034 384824 319090 384833
rect 319034 384759 319090 384768
rect 315816 378668 315868 378674
rect 315816 378610 315868 378616
rect 315828 378554 315856 378610
rect 315644 378526 315856 378554
rect 225470 377480 225526 377489
rect 225470 377415 225526 377424
rect 225484 333153 225512 377415
rect 225562 374760 225618 374769
rect 225562 374695 225618 374704
rect 225470 333144 225526 333153
rect 225470 333079 225526 333088
rect 225378 331648 225434 331657
rect 225576 331618 225604 374695
rect 225838 372176 225894 372185
rect 225838 372111 225894 372120
rect 225852 371806 225880 372111
rect 225840 371800 225892 371806
rect 225840 371742 225892 371748
rect 265860 371800 265912 371806
rect 265860 371742 265912 371748
rect 233476 357928 233528 357934
rect 233476 357870 233528 357876
rect 233488 357769 233516 357870
rect 233474 357760 233530 357769
rect 233474 357695 233530 357704
rect 233476 356568 233528 356574
rect 233474 356536 233476 356545
rect 233528 356536 233530 356545
rect 233474 356471 233530 356480
rect 233476 355208 233528 355214
rect 233474 355176 233476 355185
rect 233528 355176 233530 355185
rect 233474 355111 233530 355120
rect 233568 355140 233620 355146
rect 233568 355082 233620 355088
rect 233580 354641 233608 355082
rect 233566 354632 233622 354641
rect 233566 354567 233622 354576
rect 233476 353848 233528 353854
rect 233476 353790 233528 353796
rect 233488 353553 233516 353790
rect 233474 353544 233530 353553
rect 233474 353479 233530 353488
rect 233476 352420 233528 352426
rect 233476 352362 233528 352368
rect 233488 352329 233516 352362
rect 233474 352320 233530 352329
rect 233474 352255 233530 352264
rect 226298 351368 226354 351377
rect 226298 351303 226300 351312
rect 226352 351303 226354 351312
rect 231636 351332 231688 351338
rect 226300 351274 226352 351280
rect 231636 351274 231688 351280
rect 226574 350416 226630 350425
rect 226574 350351 226630 350360
rect 226482 349600 226538 349609
rect 226482 349535 226538 349544
rect 226390 348648 226446 348657
rect 226390 348583 226446 348592
rect 226404 348346 226432 348583
rect 226496 348414 226524 349535
rect 226484 348408 226536 348414
rect 226484 348350 226536 348356
rect 226392 348340 226444 348346
rect 226392 348282 226444 348288
rect 226588 348278 226616 350351
rect 231648 349706 231676 351274
rect 233568 351060 233620 351066
rect 233568 351002 233620 351008
rect 233474 350960 233530 350969
rect 233474 350895 233530 350904
rect 233488 350386 233516 350895
rect 233580 350561 233608 351002
rect 233566 350552 233622 350561
rect 233566 350487 233622 350496
rect 233476 350380 233528 350386
rect 233476 350322 233528 350328
rect 231636 349700 231688 349706
rect 231636 349642 231688 349648
rect 233476 349700 233528 349706
rect 233476 349642 233528 349648
rect 233488 349609 233516 349642
rect 233474 349600 233530 349609
rect 233474 349535 233530 349544
rect 232004 348408 232056 348414
rect 232004 348350 232056 348356
rect 231636 348340 231688 348346
rect 231636 348282 231688 348288
rect 226576 348272 226628 348278
rect 226576 348214 226628 348220
rect 226390 347832 226446 347841
rect 226390 347767 226446 347776
rect 226404 346986 226432 347767
rect 226392 346980 226444 346986
rect 226392 346922 226444 346928
rect 228600 346980 228652 346986
rect 228600 346922 228652 346928
rect 226482 346880 226538 346889
rect 226482 346815 226538 346824
rect 226390 346064 226446 346073
rect 226390 345999 226446 346008
rect 226404 345626 226432 345999
rect 226496 345694 226524 346815
rect 226484 345688 226536 345694
rect 226484 345630 226536 345636
rect 228048 345688 228100 345694
rect 228048 345630 228100 345636
rect 226392 345620 226444 345626
rect 226392 345562 226444 345568
rect 226022 345112 226078 345121
rect 226022 345047 226078 345056
rect 226036 344674 226064 345047
rect 226024 344668 226076 344674
rect 226024 344610 226076 344616
rect 226390 344296 226446 344305
rect 226390 344231 226392 344240
rect 226444 344231 226446 344240
rect 227956 344260 228008 344266
rect 226392 344202 226444 344208
rect 227956 344202 228008 344208
rect 226390 343344 226446 343353
rect 226390 343279 226446 343288
rect 226404 342838 226432 343279
rect 226392 342832 226444 342838
rect 226392 342774 226444 342780
rect 226482 342392 226538 342401
rect 226482 342327 226538 342336
rect 226390 341576 226446 341585
rect 226496 341546 226524 342327
rect 226390 341511 226446 341520
rect 226484 341540 226536 341546
rect 226404 341478 226432 341511
rect 226484 341482 226536 341488
rect 226392 341472 226444 341478
rect 226392 341414 226444 341420
rect 227968 341410 227996 344202
rect 228060 344130 228088 345630
rect 228612 345558 228640 346922
rect 231648 346850 231676 348282
rect 232016 346918 232044 348350
rect 233476 348272 233528 348278
rect 233474 348240 233476 348249
rect 233528 348240 233530 348249
rect 233474 348175 233530 348184
rect 232004 346912 232056 346918
rect 233476 346912 233528 346918
rect 232004 346854 232056 346860
rect 233474 346880 233476 346889
rect 233528 346880 233530 346889
rect 231636 346844 231688 346850
rect 233474 346815 233530 346824
rect 233568 346844 233620 346850
rect 231636 346786 231688 346792
rect 233568 346786 233620 346792
rect 233580 346481 233608 346786
rect 233566 346472 233622 346481
rect 233566 346407 233622 346416
rect 234580 345620 234632 345626
rect 234580 345562 234632 345568
rect 228600 345552 228652 345558
rect 228600 345494 228652 345500
rect 233476 345552 233528 345558
rect 233476 345494 233528 345500
rect 233488 345257 233516 345494
rect 233474 345248 233530 345257
rect 233474 345183 233530 345192
rect 228508 344668 228560 344674
rect 228508 344610 228560 344616
rect 228048 344124 228100 344130
rect 228048 344066 228100 344072
rect 228520 342770 228548 344610
rect 233476 344124 233528 344130
rect 233476 344066 233528 344072
rect 233488 344033 233516 344066
rect 233474 344024 233530 344033
rect 233474 343959 233530 343968
rect 233660 342832 233712 342838
rect 233660 342774 233712 342780
rect 228508 342764 228560 342770
rect 228508 342706 228560 342712
rect 233476 342764 233528 342770
rect 233476 342706 233528 342712
rect 233488 342265 233516 342706
rect 233474 342256 233530 342265
rect 233474 342191 233530 342200
rect 233568 341540 233620 341546
rect 233568 341482 233620 341488
rect 227956 341404 228008 341410
rect 227956 341346 228008 341352
rect 233476 341404 233528 341410
rect 233476 341346 233528 341352
rect 233488 341177 233516 341346
rect 233474 341168 233530 341177
rect 233474 341103 233530 341112
rect 226390 340624 226446 340633
rect 226390 340559 226446 340568
rect 226404 340118 226432 340559
rect 226392 340112 226444 340118
rect 226392 340054 226444 340060
rect 231912 340112 231964 340118
rect 231912 340054 231964 340060
rect 225930 339808 225986 339817
rect 225930 339743 225986 339752
rect 225944 338690 225972 339743
rect 226482 338856 226538 338865
rect 226482 338791 226484 338800
rect 226536 338791 226538 338800
rect 226484 338762 226536 338768
rect 225932 338684 225984 338690
rect 225932 338626 225984 338632
rect 230808 338684 230860 338690
rect 230808 338626 230860 338632
rect 225930 338040 225986 338049
rect 225930 337975 225986 337984
rect 225944 337330 225972 337975
rect 225932 337324 225984 337330
rect 225932 337266 225984 337272
rect 230716 337324 230768 337330
rect 230716 337266 230768 337272
rect 225930 337088 225986 337097
rect 225930 337023 225986 337032
rect 225944 335970 225972 337023
rect 226482 336272 226538 336281
rect 226538 336230 226616 336258
rect 226482 336207 226538 336216
rect 225932 335964 225984 335970
rect 225932 335906 225984 335912
rect 226588 331754 226616 336230
rect 230728 334474 230756 337266
rect 230820 335902 230848 338626
rect 231924 337262 231952 340054
rect 233580 338593 233608 341482
rect 233672 339953 233700 342774
rect 234592 342673 234620 345562
rect 234578 342664 234634 342673
rect 234578 342599 234634 342608
rect 233752 341472 233804 341478
rect 233752 341414 233804 341420
rect 233658 339944 233714 339953
rect 233658 339879 233714 339888
rect 233660 338820 233712 338826
rect 233660 338762 233712 338768
rect 233566 338584 233622 338593
rect 233566 338519 233622 338528
rect 231912 337256 231964 337262
rect 231912 337198 231964 337204
rect 233476 337256 233528 337262
rect 233476 337198 233528 337204
rect 233488 337097 233516 337198
rect 233474 337088 233530 337097
rect 233474 337023 233530 337032
rect 230900 335964 230952 335970
rect 230900 335906 230952 335912
rect 230808 335896 230860 335902
rect 230808 335838 230860 335844
rect 230716 334468 230768 334474
rect 230716 334410 230768 334416
rect 228600 333788 228652 333794
rect 228600 333730 228652 333736
rect 226576 331748 226628 331754
rect 226576 331690 226628 331696
rect 225378 331583 225434 331592
rect 225564 331612 225616 331618
rect 225564 331554 225616 331560
rect 225196 328960 225248 328966
rect 225196 328902 225248 328908
rect 175514 313560 175570 313569
rect 175514 313495 175570 313504
rect 175528 313122 175556 313495
rect 165120 313116 165172 313122
rect 165120 313058 165172 313064
rect 175516 313116 175568 313122
rect 175516 313058 175568 313064
rect 145522 310160 145578 310169
rect 145522 310095 145578 310104
rect 145536 309722 145564 310095
rect 145524 309716 145576 309722
rect 145524 309658 145576 309664
rect 145430 296832 145486 296841
rect 145430 296767 145486 296776
rect 145444 295918 145472 296767
rect 145432 295912 145484 295918
rect 145432 295854 145484 295860
rect 145616 283536 145668 283542
rect 145614 283504 145616 283513
rect 145668 283504 145670 283513
rect 145614 283439 145670 283448
rect 142396 282380 142448 282386
rect 142396 282322 142448 282328
rect 143040 282380 143092 282386
rect 143040 282322 143092 282328
rect 141660 273744 141712 273750
rect 141660 273686 141712 273692
rect 138622 269768 138678 269777
rect 138622 269703 138678 269712
rect 143052 266542 143080 282322
rect 149124 276934 149230 276962
rect 147824 274696 147876 274702
rect 147824 274638 147876 274644
rect 145064 274628 145116 274634
rect 145064 274570 145116 274576
rect 143684 274492 143736 274498
rect 143684 274434 143736 274440
rect 143040 266536 143092 266542
rect 143040 266478 143092 266484
rect 143696 263770 143724 274434
rect 145076 263770 145104 274570
rect 146444 274560 146496 274566
rect 146444 274502 146496 274508
rect 146456 263770 146484 274502
rect 147836 263770 147864 274638
rect 149124 274362 149152 276934
rect 149768 274974 149796 276948
rect 150426 276934 150624 276962
rect 149756 274968 149808 274974
rect 149756 274910 149808 274916
rect 149204 274424 149256 274430
rect 149204 274366 149256 274372
rect 149112 274356 149164 274362
rect 149112 274298 149164 274304
rect 149216 263770 149244 274366
rect 150492 274288 150544 274294
rect 150492 274230 150544 274236
rect 150504 264042 150532 274230
rect 150596 266678 150624 276934
rect 151056 274770 151084 276948
rect 151622 276934 151912 276962
rect 151044 274764 151096 274770
rect 151044 274706 151096 274712
rect 151780 274764 151832 274770
rect 151780 274706 151832 274712
rect 150584 266672 150636 266678
rect 150584 266614 150636 266620
rect 151792 266134 151820 274706
rect 151884 266406 151912 276934
rect 151964 274900 152016 274906
rect 151964 274842 152016 274848
rect 151872 266400 151924 266406
rect 151872 266342 151924 266348
rect 151780 266128 151832 266134
rect 151780 266070 151832 266076
rect 150504 264014 150578 264042
rect 143572 263742 143724 263770
rect 144952 263742 145104 263770
rect 146332 263742 146484 263770
rect 147712 263742 147864 263770
rect 149092 263742 149244 263770
rect 150550 263756 150578 264014
rect 151976 263770 152004 274842
rect 152252 274770 152280 276948
rect 152910 276934 153200 276962
rect 152240 274764 152292 274770
rect 152240 274706 152292 274712
rect 153172 266338 153200 276934
rect 153448 274838 153476 276948
rect 153436 274832 153488 274838
rect 153436 274774 153488 274780
rect 154092 274770 154120 276948
rect 154460 276934 154750 276962
rect 153344 274764 153396 274770
rect 153344 274706 153396 274712
rect 154080 274764 154132 274770
rect 154080 274706 154132 274712
rect 153252 266740 153304 266746
rect 153252 266682 153304 266688
rect 153160 266332 153212 266338
rect 153160 266274 153212 266280
rect 153264 264314 153292 266682
rect 153356 266474 153384 274706
rect 153344 266468 153396 266474
rect 153344 266410 153396 266416
rect 153264 264286 153384 264314
rect 151944 263742 152004 263770
rect 142394 263648 142450 263657
rect 153356 263634 153384 264286
rect 153324 263606 153384 263634
rect 154460 263618 154488 276934
rect 155288 275110 155316 276948
rect 155932 275178 155960 276948
rect 156208 276934 156590 276962
rect 155920 275172 155972 275178
rect 155920 275114 155972 275120
rect 155276 275104 155328 275110
rect 155276 275046 155328 275052
rect 154540 274832 154592 274838
rect 154540 274774 154592 274780
rect 154552 266270 154580 274774
rect 154632 274764 154684 274770
rect 154632 274706 154684 274712
rect 154540 266264 154592 266270
rect 154540 266206 154592 266212
rect 154644 266202 154672 274706
rect 155736 266536 155788 266542
rect 155736 266478 155788 266484
rect 154632 266196 154684 266202
rect 154632 266138 154684 266144
rect 154724 265652 154776 265658
rect 154724 265594 154776 265600
rect 154736 263770 154764 265594
rect 154704 263742 154764 263770
rect 155748 263770 155776 266478
rect 156208 263929 156236 276934
rect 157220 274401 157248 276948
rect 157772 274537 157800 276948
rect 158416 274537 158444 276948
rect 159060 274673 159088 276948
rect 159336 276934 159626 276962
rect 159046 274664 159102 274673
rect 159046 274599 159102 274608
rect 157758 274528 157814 274537
rect 157758 274463 157814 274472
rect 158402 274528 158458 274537
rect 159336 274498 159364 276934
rect 160256 274634 160284 276948
rect 160520 274968 160572 274974
rect 160520 274910 160572 274916
rect 160244 274628 160296 274634
rect 160244 274570 160296 274576
rect 158402 274463 158458 274472
rect 159324 274492 159376 274498
rect 159324 274434 159376 274440
rect 159600 274492 159652 274498
rect 159600 274434 159652 274440
rect 157206 274392 157262 274401
rect 156840 274356 156892 274362
rect 157206 274327 157262 274336
rect 156840 274298 156892 274304
rect 156852 265590 156880 274298
rect 157852 265720 157904 265726
rect 157852 265662 157904 265668
rect 156840 265584 156892 265590
rect 156840 265526 156892 265532
rect 156194 263920 156250 263929
rect 156194 263855 156250 263864
rect 157864 263770 157892 265662
rect 159612 265658 159640 274434
rect 159600 265652 159652 265658
rect 159600 265594 159652 265600
rect 158956 265584 159008 265590
rect 158956 265526 159008 265532
rect 158968 263770 158996 265526
rect 160532 263770 160560 274910
rect 160900 274566 160928 276948
rect 161452 274702 161480 276948
rect 162096 274770 162124 276948
rect 162740 274906 162768 276948
rect 162728 274900 162780 274906
rect 162728 274842 162780 274848
rect 163292 274838 163320 276948
rect 163280 274832 163332 274838
rect 163280 274774 163332 274780
rect 162084 274764 162136 274770
rect 162084 274706 162136 274712
rect 161440 274696 161492 274702
rect 161440 274638 161492 274644
rect 160888 274560 160940 274566
rect 160888 274502 160940 274508
rect 163936 273818 163964 276948
rect 164580 274498 164608 276948
rect 164568 274492 164620 274498
rect 164568 274434 164620 274440
rect 162360 273812 162412 273818
rect 162360 273754 162412 273760
rect 163924 273812 163976 273818
rect 163924 273754 163976 273760
rect 162372 266746 162400 273754
rect 162360 266740 162412 266746
rect 162360 266682 162412 266688
rect 161716 266672 161768 266678
rect 161716 266614 161768 266620
rect 161728 263770 161756 266614
rect 164568 266400 164620 266406
rect 164568 266342 164620 266348
rect 163096 266128 163148 266134
rect 163096 266070 163148 266076
rect 163108 263770 163136 266070
rect 164580 263770 164608 266342
rect 165132 265726 165160 313058
rect 167878 306216 167934 306225
rect 167878 306151 167934 306160
rect 167892 297210 167920 306151
rect 167880 297204 167932 297210
rect 167880 297146 167932 297152
rect 175516 297204 175568 297210
rect 175516 297146 175568 297152
rect 175528 296841 175556 297146
rect 175514 296832 175570 296841
rect 175514 296767 175570 296776
rect 168062 286360 168118 286369
rect 168062 286295 168118 286304
rect 168076 286262 168104 286295
rect 168064 286256 168116 286262
rect 168064 286198 168116 286204
rect 172756 286256 172808 286262
rect 172756 286198 172808 286204
rect 172768 280686 172796 286198
rect 172756 280680 172808 280686
rect 172756 280622 172808 280628
rect 175792 280680 175844 280686
rect 175792 280622 175844 280628
rect 175804 280249 175832 280622
rect 175790 280240 175846 280249
rect 175790 280175 175846 280184
rect 182428 269670 182456 271916
rect 182416 269664 182468 269670
rect 182416 269606 182468 269612
rect 189512 269534 189540 271916
rect 196688 269602 196716 271916
rect 196676 269596 196728 269602
rect 196676 269538 196728 269544
rect 197504 269596 197556 269602
rect 197504 269538 197556 269544
rect 189500 269528 189552 269534
rect 189500 269470 189552 269476
rect 189316 269052 189368 269058
rect 189316 268994 189368 269000
rect 174872 268984 174924 268990
rect 174872 268926 174924 268932
rect 165948 266468 166000 266474
rect 165948 266410 166000 266416
rect 165120 265720 165172 265726
rect 165120 265662 165172 265668
rect 165960 263770 165988 266410
rect 167328 266332 167380 266338
rect 167328 266274 167380 266280
rect 167340 263770 167368 266274
rect 168708 266264 168760 266270
rect 168708 266206 168760 266212
rect 168720 263770 168748 266206
rect 170088 266196 170140 266202
rect 170088 266138 170140 266144
rect 170100 263770 170128 266138
rect 155748 263742 156084 263770
rect 157556 263742 157892 263770
rect 158936 263742 158996 263770
rect 160316 263742 160560 263770
rect 161696 263742 161756 263770
rect 163076 263742 163136 263770
rect 164548 263742 164608 263770
rect 165928 263742 165988 263770
rect 167308 263742 167368 263770
rect 168688 263742 168748 263770
rect 170068 263742 170128 263770
rect 154448 263612 154500 263618
rect 142394 263583 142450 263592
rect 140280 263476 140332 263482
rect 140280 263418 140332 263424
rect 139818 263104 139874 263113
rect 139818 263039 139874 263048
rect 139832 262802 139860 263039
rect 139820 262796 139872 262802
rect 139820 262738 139872 262744
rect 138806 259976 138862 259985
rect 138806 259911 138862 259920
rect 138820 250465 138848 259911
rect 139544 255928 139596 255934
rect 139544 255870 139596 255876
rect 138900 253140 138952 253146
rect 138900 253082 138952 253088
rect 138806 250456 138862 250465
rect 138806 250391 138862 250400
rect 138912 244209 138940 253082
rect 139556 248425 139584 255870
rect 139542 248416 139598 248425
rect 139542 248351 139598 248360
rect 138898 244200 138954 244209
rect 138898 244135 138954 244144
rect 140188 239200 140240 239206
rect 140188 239142 140240 239148
rect 140200 238497 140228 239142
rect 140186 238488 140242 238497
rect 140186 238423 140242 238432
rect 140292 237273 140320 263418
rect 140370 261744 140426 261753
rect 140370 261679 140426 261688
rect 140384 261442 140412 261679
rect 140372 261436 140424 261442
rect 140372 261378 140424 261384
rect 140370 260384 140426 260393
rect 140370 260319 140426 260328
rect 140384 260082 140412 260319
rect 140372 260076 140424 260082
rect 140372 260018 140424 260024
rect 140554 258888 140610 258897
rect 140554 258823 140610 258832
rect 140568 258654 140596 258823
rect 140556 258648 140608 258654
rect 140556 258590 140608 258596
rect 140554 257528 140610 257537
rect 140554 257463 140610 257472
rect 140568 257294 140596 257463
rect 140556 257288 140608 257294
rect 140556 257230 140608 257236
rect 140554 256168 140610 256177
rect 140554 256103 140610 256112
rect 140568 256002 140596 256103
rect 140556 255996 140608 256002
rect 140556 255938 140608 255944
rect 140554 254672 140610 254681
rect 140554 254607 140610 254616
rect 140568 254506 140596 254607
rect 140556 254500 140608 254506
rect 140556 254442 140608 254448
rect 140462 253312 140518 253321
rect 140462 253247 140518 253256
rect 140370 250592 140426 250601
rect 140370 250527 140426 250536
rect 140278 237264 140334 237273
rect 140384 237234 140412 250527
rect 140476 243354 140504 253247
rect 140738 251952 140794 251961
rect 140738 251887 140794 251896
rect 140556 250284 140608 250290
rect 140556 250226 140608 250232
rect 140568 249649 140596 250226
rect 140554 249640 140610 249649
rect 140554 249575 140610 249584
rect 140648 247360 140700 247366
rect 140648 247302 140700 247308
rect 140660 246929 140688 247302
rect 140646 246920 140702 246929
rect 140646 246855 140702 246864
rect 140556 246204 140608 246210
rect 140556 246146 140608 246152
rect 140568 245569 140596 246146
rect 140554 245560 140610 245569
rect 140554 245495 140610 245504
rect 140752 245410 140780 251887
rect 140568 245382 140780 245410
rect 140464 243348 140516 243354
rect 140464 243290 140516 243296
rect 140568 243218 140596 245382
rect 140648 243416 140700 243422
rect 140648 243358 140700 243364
rect 140556 243212 140608 243218
rect 140556 243154 140608 243160
rect 140660 242849 140688 243358
rect 140646 242840 140702 242849
rect 140646 242775 140702 242784
rect 140554 240664 140610 240673
rect 140554 240599 140556 240608
rect 140608 240599 140610 240608
rect 140556 240570 140608 240576
rect 140554 239304 140610 239313
rect 140554 239239 140556 239248
rect 140608 239239 140610 239248
rect 140556 239210 140608 239216
rect 142408 238662 142436 263583
rect 154448 263554 154500 263560
rect 173398 263104 173454 263113
rect 173398 263039 173454 263048
rect 173124 255588 173176 255594
rect 173124 255530 173176 255536
rect 172938 253312 172994 253321
rect 172938 253247 172940 253256
rect 172992 253247 172994 253256
rect 172940 253218 172992 253224
rect 173136 250601 173164 255530
rect 173308 254568 173360 254574
rect 173308 254510 173360 254516
rect 173122 250592 173178 250601
rect 173122 250527 173178 250536
rect 173320 249626 173348 254510
rect 173412 250290 173440 263039
rect 173490 261744 173546 261753
rect 173490 261679 173546 261688
rect 173400 250284 173452 250290
rect 173400 250226 173452 250232
rect 173320 249598 173440 249626
rect 173308 249468 173360 249474
rect 173308 249410 173360 249416
rect 173320 249105 173348 249410
rect 173306 249096 173362 249105
rect 173306 249031 173362 249040
rect 173308 247904 173360 247910
rect 173308 247846 173360 247852
rect 173320 247745 173348 247846
rect 173306 247736 173362 247745
rect 173306 247671 173362 247680
rect 173412 247586 173440 249598
rect 173504 248930 173532 261679
rect 173766 260384 173822 260393
rect 173766 260319 173822 260328
rect 173780 254794 173808 260319
rect 173858 258888 173914 258897
rect 173858 258823 173914 258832
rect 173596 254766 173808 254794
rect 173596 254250 173624 254766
rect 173766 254672 173822 254681
rect 173766 254607 173822 254616
rect 173780 254506 173808 254607
rect 173768 254500 173820 254506
rect 173768 254442 173820 254448
rect 173596 254222 173808 254250
rect 173674 251952 173730 251961
rect 173674 251887 173676 251896
rect 173728 251887 173730 251896
rect 173676 251858 173728 251864
rect 173584 251780 173636 251786
rect 173584 251722 173636 251728
rect 173492 248924 173544 248930
rect 173492 248866 173544 248872
rect 173320 247558 173440 247586
rect 173320 244889 173348 247558
rect 173306 244880 173362 244889
rect 173306 244815 173362 244824
rect 173308 244436 173360 244442
rect 173308 244378 173360 244384
rect 173320 243529 173348 244378
rect 173306 243520 173362 243529
rect 173306 243455 173362 243464
rect 172940 242804 172992 242810
rect 172940 242746 172992 242752
rect 172952 242169 172980 242746
rect 172938 242160 172994 242169
rect 172938 242095 172994 242104
rect 173596 240673 173624 251722
rect 173676 250352 173728 250358
rect 173676 250294 173728 250300
rect 173688 247042 173716 250294
rect 173780 248862 173808 254222
rect 173768 248856 173820 248862
rect 173768 248798 173820 248804
rect 173872 247570 173900 258823
rect 173950 257528 174006 257537
rect 173950 257463 174006 257472
rect 173860 247564 173912 247570
rect 173860 247506 173912 247512
rect 173688 247014 173900 247042
rect 173676 246952 173728 246958
rect 173676 246894 173728 246900
rect 173688 246385 173716 246894
rect 173674 246376 173730 246385
rect 173674 246311 173730 246320
rect 173582 240664 173638 240673
rect 173582 240599 173638 240608
rect 173872 239313 173900 247014
rect 173964 246210 173992 257463
rect 174042 256168 174098 256177
rect 174042 256103 174098 256112
rect 174056 256002 174084 256103
rect 174044 255996 174096 256002
rect 174044 255938 174096 255944
rect 174780 253276 174832 253282
rect 174780 253218 174832 253224
rect 174044 248992 174096 248998
rect 174044 248934 174096 248940
rect 173952 246204 174004 246210
rect 173952 246146 174004 246152
rect 173858 239304 173914 239313
rect 173858 239239 173914 239248
rect 142396 238656 142448 238662
rect 142396 238598 142448 238604
rect 142764 238656 142816 238662
rect 142764 238598 142816 238604
rect 142776 238361 142804 238598
rect 142762 238352 142818 238361
rect 142762 238287 142818 238296
rect 174056 237953 174084 248934
rect 174792 243422 174820 253218
rect 174780 243416 174832 243422
rect 174780 243358 174832 243364
rect 174042 237944 174098 237953
rect 174042 237879 174098 237888
rect 140278 237199 140334 237208
rect 140372 237228 140424 237234
rect 140372 237170 140424 237176
rect 172940 237228 172992 237234
rect 172940 237170 172992 237176
rect 172952 236593 172980 237170
rect 172938 236584 172994 236593
rect 172938 236519 172994 236528
rect 147454 236176 147510 236185
rect 148374 236176 148430 236185
rect 147454 236111 147510 236120
rect 147836 236134 148374 236162
rect 147468 235890 147496 236111
rect 142408 235862 143388 235890
rect 144308 235862 144644 235890
rect 145228 235862 145288 235890
rect 137702 234952 137758 234961
rect 137702 234887 137758 234896
rect 139266 234952 139322 234961
rect 139266 234887 139322 234896
rect 137716 234446 137744 234887
rect 139280 234514 139308 234887
rect 139268 234508 139320 234514
rect 139268 234450 139320 234456
rect 137704 234440 137756 234446
rect 137704 234382 137756 234388
rect 137716 226393 137744 234382
rect 138164 233760 138216 233766
rect 138164 233702 138216 233708
rect 137702 226384 137758 226393
rect 137702 226319 137758 226328
rect 137612 226144 137664 226150
rect 137612 226086 137664 226092
rect 137520 225600 137572 225606
rect 137520 225542 137572 225548
rect 137334 223256 137390 223265
rect 137334 223191 137390 223200
rect 137242 220128 137298 220137
rect 137242 220063 137298 220072
rect 137150 217000 137206 217009
rect 137150 216935 137206 216944
rect 137058 213872 137114 213881
rect 137058 213807 137114 213816
rect 136966 210744 137022 210753
rect 136966 210679 137022 210688
rect 136796 204854 136916 204882
rect 136796 204338 136824 204854
rect 136876 204792 136928 204798
rect 136876 204734 136928 204740
rect 136888 204497 136916 204734
rect 136874 204488 136930 204497
rect 136874 204423 136930 204432
rect 136796 204310 136916 204338
rect 136888 200961 136916 204310
rect 136874 200952 136930 200961
rect 136874 200887 136930 200896
rect 136966 141928 137022 141937
rect 136966 141863 137022 141872
rect 136980 141354 137008 141863
rect 136968 141348 137020 141354
rect 136968 141290 137020 141296
rect 136874 139888 136930 139897
rect 136874 139823 136930 139832
rect 136888 139246 136916 139823
rect 136876 139240 136928 139246
rect 136876 139182 136928 139188
rect 136888 132961 136916 139182
rect 136874 132952 136930 132961
rect 136874 132887 136930 132896
rect 136876 132372 136928 132378
rect 136876 132314 136928 132320
rect 136888 120449 136916 132314
rect 136980 123305 137008 141290
rect 137334 141112 137390 141121
rect 137334 141047 137390 141056
rect 137348 140606 137376 141047
rect 137336 140600 137388 140606
rect 137336 140542 137388 140548
rect 137242 134448 137298 134457
rect 137242 134383 137298 134392
rect 137256 127550 137284 134383
rect 137348 132378 137376 140542
rect 137336 132372 137388 132378
rect 137336 132314 137388 132320
rect 137060 127544 137112 127550
rect 137060 127486 137112 127492
rect 137244 127544 137296 127550
rect 137244 127486 137296 127492
rect 137072 126025 137100 127486
rect 137058 126016 137114 126025
rect 137058 125951 137114 125960
rect 136966 123296 137022 123305
rect 136966 123231 137022 123240
rect 136874 120440 136930 120449
rect 136874 120375 136930 120384
rect 136874 113232 136930 113241
rect 136874 113167 136930 113176
rect 136888 112998 136916 113167
rect 136876 112992 136928 112998
rect 136876 112934 136928 112940
rect 136876 110952 136928 110958
rect 136876 110894 136928 110900
rect 136888 110793 136916 110894
rect 136874 110784 136930 110793
rect 136874 110719 136930 110728
rect 137532 98553 137560 225542
rect 137702 216592 137758 216601
rect 137702 216527 137758 216536
rect 137612 215876 137664 215882
rect 137612 215818 137664 215824
rect 137624 185729 137652 215818
rect 137716 191985 137744 216527
rect 138176 208305 138204 233702
rect 138162 208296 138218 208305
rect 138162 208231 138218 208240
rect 138176 207625 138204 208231
rect 138162 207616 138218 207625
rect 138162 207551 138218 207560
rect 137796 202072 137848 202078
rect 137796 202014 137848 202020
rect 137702 191976 137758 191985
rect 137702 191911 137758 191920
rect 137808 188698 137836 202014
rect 137808 188670 137928 188698
rect 137794 188576 137850 188585
rect 137794 188511 137850 188520
rect 137808 188342 137836 188511
rect 137796 188336 137848 188342
rect 137796 188278 137848 188284
rect 137610 185720 137666 185729
rect 137610 185655 137666 185664
rect 137900 182601 137928 188670
rect 142408 188342 142436 235862
rect 144616 233154 144644 235862
rect 144604 233148 144656 233154
rect 144604 233090 144656 233096
rect 145260 233086 145288 235862
rect 145352 235862 146240 235890
rect 146824 235862 147496 235890
rect 145248 233080 145300 233086
rect 145248 233022 145300 233028
rect 145154 216184 145210 216193
rect 145154 216119 145210 216128
rect 145168 215882 145196 216119
rect 145156 215876 145208 215882
rect 145156 215818 145208 215824
rect 145352 204798 145380 235862
rect 146824 233766 146852 235862
rect 147836 235097 147864 236134
rect 148374 236111 148430 236120
rect 148650 236040 148706 236049
rect 148650 235975 148706 235984
rect 148664 235262 148692 235975
rect 148742 235904 148798 235913
rect 148798 235862 149244 235890
rect 150104 235862 150164 235890
rect 148742 235839 148798 235848
rect 148652 235256 148704 235262
rect 148652 235198 148704 235204
rect 149216 235194 149244 235862
rect 149204 235188 149256 235194
rect 149204 235130 149256 235136
rect 147822 235088 147878 235097
rect 147822 235023 147878 235032
rect 146812 233760 146864 233766
rect 150136 233737 150164 235862
rect 150688 235862 151024 235890
rect 152036 235862 152096 235890
rect 152956 235862 153292 235890
rect 153968 235862 154304 235890
rect 154888 235862 155224 235890
rect 155900 235862 156144 235890
rect 156820 235862 157156 235890
rect 157832 235862 158168 235890
rect 158752 235862 158904 235890
rect 159764 235862 160100 235890
rect 160684 235862 161020 235890
rect 161696 235862 162032 235890
rect 150688 235262 150716 235862
rect 150676 235256 150728 235262
rect 150676 235198 150728 235204
rect 152068 234961 152096 235862
rect 152054 234952 152110 234961
rect 152054 234887 152110 234896
rect 150584 233760 150636 233766
rect 146812 233702 146864 233708
rect 149294 233728 149350 233737
rect 149294 233663 149350 233672
rect 150122 233728 150178 233737
rect 150584 233702 150636 233708
rect 150122 233663 150178 233672
rect 149308 233057 149336 233663
rect 150492 233352 150544 233358
rect 150492 233294 150544 233300
rect 149294 233048 149350 233057
rect 149294 232983 149350 232992
rect 149296 224852 149348 224858
rect 149296 224794 149348 224800
rect 149308 222820 149336 224794
rect 150504 222698 150532 233294
rect 150596 224858 150624 233702
rect 153264 233601 153292 235862
rect 153250 233592 153306 233601
rect 153250 233527 153306 233536
rect 153344 233556 153396 233562
rect 153344 233498 153396 233504
rect 151964 233488 152016 233494
rect 151964 233430 152016 233436
rect 151872 233284 151924 233290
rect 151872 233226 151924 233232
rect 151884 225198 151912 233226
rect 151044 225192 151096 225198
rect 151044 225134 151096 225140
rect 151872 225192 151924 225198
rect 151872 225134 151924 225140
rect 150584 224852 150636 224858
rect 150584 224794 150636 224800
rect 151056 222820 151084 225134
rect 151976 222820 152004 233430
rect 150150 222670 150532 222698
rect 153356 222562 153384 233498
rect 154276 232474 154304 235862
rect 154724 233420 154776 233426
rect 154724 233362 154776 233368
rect 154632 233216 154684 233222
rect 154632 233158 154684 233164
rect 154264 232468 154316 232474
rect 154264 232410 154316 232416
rect 153712 225328 153764 225334
rect 153712 225270 153764 225276
rect 153724 222820 153752 225270
rect 154644 222820 154672 233158
rect 154736 225334 154764 233362
rect 155196 232542 155224 235862
rect 156012 232876 156064 232882
rect 156012 232818 156064 232824
rect 155184 232536 155236 232542
rect 155184 232478 155236 232484
rect 156024 230586 156052 232818
rect 156116 232678 156144 235862
rect 156104 232672 156156 232678
rect 156104 232614 156156 232620
rect 157128 232610 157156 235862
rect 157484 233692 157536 233698
rect 157484 233634 157536 233640
rect 157116 232604 157168 232610
rect 157116 232546 157168 232552
rect 156380 232468 156432 232474
rect 156380 232410 156432 232416
rect 156024 230558 156144 230586
rect 156116 225334 156144 230558
rect 156392 225418 156420 232410
rect 156392 225390 156696 225418
rect 154724 225328 154776 225334
rect 154724 225270 154776 225276
rect 155460 225328 155512 225334
rect 155460 225270 155512 225276
rect 156104 225328 156156 225334
rect 156104 225270 156156 225276
rect 156380 225328 156432 225334
rect 156380 225270 156432 225276
rect 155472 222820 155500 225270
rect 156392 222820 156420 225270
rect 156668 222834 156696 225390
rect 157496 225334 157524 233634
rect 158140 232542 158168 235862
rect 158220 232672 158272 232678
rect 158220 232614 158272 232620
rect 157576 232536 157628 232542
rect 157576 232478 157628 232484
rect 158128 232536 158180 232542
rect 158128 232478 158180 232484
rect 157484 225328 157536 225334
rect 157484 225270 157536 225276
rect 156668 222806 157326 222834
rect 157588 222698 157616 232478
rect 158232 224246 158260 232614
rect 158876 232474 158904 235862
rect 160072 232814 160100 235862
rect 160992 233630 161020 235862
rect 160980 233624 161032 233630
rect 160980 233566 161032 233572
rect 160060 232808 160112 232814
rect 160060 232750 160112 232756
rect 161808 232808 161860 232814
rect 161808 232750 161860 232756
rect 159048 232604 159100 232610
rect 159048 232546 159100 232552
rect 158864 232468 158916 232474
rect 158864 232410 158916 232416
rect 159060 224330 159088 232546
rect 160336 232536 160388 232542
rect 160336 232478 160388 232484
rect 159060 224302 159456 224330
rect 158220 224240 158272 224246
rect 158220 224182 158272 224188
rect 159048 224240 159100 224246
rect 159048 224182 159100 224188
rect 159060 222820 159088 224182
rect 159428 222698 159456 224302
rect 160348 222834 160376 232478
rect 160980 232468 161032 232474
rect 160980 232410 161032 232416
rect 160992 224382 161020 232410
rect 160980 224376 161032 224382
rect 160980 224318 161032 224324
rect 161716 224376 161768 224382
rect 161716 224318 161768 224324
rect 160348 222806 160822 222834
rect 161728 222820 161756 224318
rect 161820 222698 161848 232750
rect 162004 232474 162032 235862
rect 162280 235862 162616 235890
rect 163292 235862 163628 235890
rect 164548 235862 164608 235890
rect 162280 233766 162308 235862
rect 162268 233760 162320 233766
rect 162268 233702 162320 233708
rect 163188 233624 163240 233630
rect 163188 233566 163240 233572
rect 161992 232468 162044 232474
rect 161992 232410 162044 232416
rect 163004 232468 163056 232474
rect 163004 232410 163056 232416
rect 163016 225198 163044 232410
rect 163004 225192 163056 225198
rect 163004 225134 163056 225140
rect 163200 222834 163228 233566
rect 163292 232950 163320 235862
rect 164580 233290 164608 235862
rect 165224 235862 165560 235890
rect 166144 235862 166480 235890
rect 167248 235862 167492 235890
rect 168076 235862 168412 235890
rect 169088 235862 169424 235890
rect 170008 235862 170344 235890
rect 165224 233494 165252 235862
rect 166144 233562 166172 235862
rect 166132 233556 166184 233562
rect 166132 233498 166184 233504
rect 165212 233488 165264 233494
rect 165212 233430 165264 233436
rect 167248 233426 167276 235862
rect 167236 233420 167288 233426
rect 167236 233362 167288 233368
rect 164568 233284 164620 233290
rect 164568 233226 164620 233232
rect 168076 233222 168104 235862
rect 168064 233216 168116 233222
rect 168064 233158 168116 233164
rect 165120 233148 165172 233154
rect 165120 233090 165172 233096
rect 163280 232944 163332 232950
rect 163280 232886 163332 232892
rect 164384 225192 164436 225198
rect 164384 225134 164436 225140
rect 163200 222806 163490 222834
rect 164396 222820 164424 225134
rect 157588 222670 158154 222698
rect 159428 222670 159994 222698
rect 161820 222670 162662 222698
rect 152818 222534 153384 222562
rect 165132 219282 165160 233090
rect 169088 232882 169116 235862
rect 170008 233698 170036 235862
rect 169996 233692 170048 233698
rect 169996 233634 170048 233640
rect 169076 232876 169128 232882
rect 169076 232818 169128 232824
rect 172020 225668 172072 225674
rect 172020 225610 172072 225616
rect 165120 219276 165172 219282
rect 165120 219218 165172 219224
rect 145340 204792 145392 204798
rect 145340 204734 145392 204740
rect 145430 202856 145486 202865
rect 145430 202791 145486 202800
rect 145444 202078 145472 202791
rect 145432 202072 145484 202078
rect 145432 202014 145484 202020
rect 145614 189528 145670 189537
rect 145614 189463 145670 189472
rect 142396 188336 142448 188342
rect 142396 188278 142448 188284
rect 143040 188336 143092 188342
rect 143040 188278 143092 188284
rect 138900 188268 138952 188274
rect 138900 188210 138952 188216
rect 137886 182592 137942 182601
rect 137886 182527 137942 182536
rect 138912 179473 138940 188210
rect 138898 179464 138954 179473
rect 138898 179399 138954 179408
rect 143052 172702 143080 188278
rect 145628 188274 145656 189463
rect 145616 188268 145668 188274
rect 145616 188210 145668 188216
rect 149216 181134 149244 182836
rect 149768 181202 149796 182836
rect 149756 181196 149808 181202
rect 149756 181138 149808 181144
rect 149204 181128 149256 181134
rect 149204 181070 149256 181076
rect 150308 180992 150360 180998
rect 150308 180934 150360 180940
rect 147824 180924 147876 180930
rect 147824 180866 147876 180872
rect 145064 180788 145116 180794
rect 145064 180730 145116 180736
rect 143684 180652 143736 180658
rect 143684 180594 143736 180600
rect 143040 172696 143092 172702
rect 143040 172638 143092 172644
rect 143696 169794 143724 180594
rect 145076 169794 145104 180730
rect 146444 180720 146496 180726
rect 146444 180662 146496 180668
rect 146456 169794 146484 180662
rect 147836 169794 147864 180866
rect 149204 180856 149256 180862
rect 149204 180798 149256 180804
rect 148742 180008 148798 180017
rect 148742 179943 148798 179952
rect 148756 173081 148784 179943
rect 148742 173072 148798 173081
rect 148742 173007 148798 173016
rect 149216 169794 149244 180798
rect 143572 169766 143724 169794
rect 144952 169766 145104 169794
rect 146332 169766 146484 169794
rect 147712 169766 147864 169794
rect 149092 169766 149244 169794
rect 150320 169794 150348 180934
rect 150412 172838 150440 182836
rect 151070 182822 151360 182850
rect 150400 172832 150452 172838
rect 150400 172774 150452 172780
rect 151332 172770 151360 182822
rect 151320 172764 151372 172770
rect 151320 172706 151372 172712
rect 151608 172566 151636 182836
rect 151964 181060 152016 181066
rect 151964 181002 152016 181008
rect 151596 172560 151648 172566
rect 151596 172502 151648 172508
rect 151976 169794 152004 181002
rect 152252 179978 152280 182836
rect 152910 182822 153384 182850
rect 152240 179972 152292 179978
rect 152240 179914 152292 179920
rect 153252 179972 153304 179978
rect 153252 179914 153304 179920
rect 153160 173036 153212 173042
rect 153160 172978 153212 172984
rect 153172 172498 153200 172978
rect 153264 172634 153292 179914
rect 153356 173042 153384 182822
rect 153448 179978 153476 182836
rect 154106 182822 154672 182850
rect 154644 180130 154672 182822
rect 154736 182057 154764 182836
rect 154722 182048 154778 182057
rect 154722 181983 154778 181992
rect 155288 181241 155316 182836
rect 155274 181232 155330 181241
rect 155274 181167 155330 181176
rect 154644 180102 154764 180130
rect 153436 179972 153488 179978
rect 153436 179914 153488 179920
rect 154632 179972 154684 179978
rect 154632 179914 154684 179920
rect 154644 174282 154672 179914
rect 154552 174254 154672 174282
rect 153344 173036 153396 173042
rect 153344 172978 153396 172984
rect 153344 172900 153396 172906
rect 153344 172842 153396 172848
rect 153252 172628 153304 172634
rect 153252 172570 153304 172576
rect 153160 172492 153212 172498
rect 153160 172434 153212 172440
rect 153356 169794 153384 172842
rect 154552 172430 154580 174254
rect 154736 174146 154764 180102
rect 155932 180017 155960 182836
rect 156576 180697 156604 182836
rect 157220 180969 157248 182836
rect 157206 180960 157262 180969
rect 157206 180895 157262 180904
rect 157772 180833 157800 182836
rect 158416 181105 158444 182836
rect 158956 181128 159008 181134
rect 158402 181096 158458 181105
rect 158956 181070 159008 181076
rect 158402 181031 158458 181040
rect 157758 180824 157814 180833
rect 157758 180759 157814 180768
rect 156562 180688 156618 180697
rect 156562 180623 156618 180632
rect 155918 180008 155974 180017
rect 155918 179943 155974 179952
rect 154644 174118 154764 174146
rect 154540 172424 154592 172430
rect 154540 172366 154592 172372
rect 154644 172362 154672 174118
rect 154724 172968 154776 172974
rect 154724 172910 154776 172916
rect 154632 172356 154684 172362
rect 154632 172298 154684 172304
rect 154736 169794 154764 172910
rect 155736 172696 155788 172702
rect 155736 172638 155788 172644
rect 157852 172696 157904 172702
rect 157852 172638 157904 172644
rect 150320 169766 150564 169794
rect 151944 169766 152004 169794
rect 153324 169766 153384 169794
rect 154704 169766 154764 169794
rect 155748 169794 155776 172638
rect 157864 169794 157892 172638
rect 158968 169794 158996 181070
rect 159060 180561 159088 182836
rect 159336 182822 159626 182850
rect 159336 180658 159364 182822
rect 159600 181196 159652 181202
rect 159600 181138 159652 181144
rect 159324 180652 159376 180658
rect 159324 180594 159376 180600
rect 159046 180552 159102 180561
rect 159046 180487 159102 180496
rect 159612 173042 159640 181138
rect 160256 180794 160284 182836
rect 160244 180788 160296 180794
rect 160244 180730 160296 180736
rect 160900 180726 160928 182836
rect 161452 180930 161480 182836
rect 161440 180924 161492 180930
rect 161440 180866 161492 180872
rect 162096 180862 162124 182836
rect 162740 180998 162768 182836
rect 163292 181066 163320 182836
rect 163280 181060 163332 181066
rect 163280 181002 163332 181008
rect 162728 180992 162780 180998
rect 162728 180934 162780 180940
rect 162084 180856 162136 180862
rect 162084 180798 162136 180804
rect 160888 180720 160940 180726
rect 160888 180662 160940 180668
rect 159600 173036 159652 173042
rect 159600 172978 159652 172984
rect 160336 173036 160388 173042
rect 160336 172978 160388 172984
rect 160348 169794 160376 172978
rect 163936 172906 163964 182836
rect 164594 182822 164700 182850
rect 164672 172974 164700 182822
rect 164660 172968 164712 172974
rect 164660 172910 164712 172916
rect 163924 172900 163976 172906
rect 163924 172842 163976 172848
rect 161716 172832 161768 172838
rect 161716 172774 161768 172780
rect 161728 169794 161756 172774
rect 163096 172764 163148 172770
rect 163096 172706 163148 172712
rect 163108 169794 163136 172706
rect 165132 172702 165160 219218
rect 167970 212784 168026 212793
rect 167970 212719 168026 212728
rect 167984 211734 168012 212719
rect 167972 211728 168024 211734
rect 167972 211670 168024 211676
rect 169258 192792 169314 192801
rect 169258 192727 169314 192736
rect 169272 186846 169300 192727
rect 169260 186840 169312 186846
rect 169260 186782 169312 186788
rect 165120 172696 165172 172702
rect 165120 172638 165172 172644
rect 165856 172628 165908 172634
rect 165856 172570 165908 172576
rect 164476 172560 164528 172566
rect 164476 172502 164528 172508
rect 164488 169930 164516 172502
rect 165868 169930 165896 172570
rect 167328 172492 167380 172498
rect 167328 172434 167380 172440
rect 164488 169902 164562 169930
rect 165868 169902 165942 169930
rect 155748 169766 156084 169794
rect 157556 169766 157892 169794
rect 158936 169766 158996 169794
rect 160316 169766 160376 169794
rect 161696 169766 161756 169794
rect 163076 169766 163136 169794
rect 164534 169780 164562 169902
rect 165914 169780 165942 169902
rect 167340 169794 167368 172434
rect 168708 172424 168760 172430
rect 168708 172366 168760 172372
rect 168720 169794 168748 172366
rect 170088 172356 170140 172362
rect 170088 172298 170140 172304
rect 170100 169794 170128 172298
rect 167308 169766 167368 169794
rect 168688 169766 168748 169794
rect 170068 169766 170128 169794
rect 140280 169568 140332 169574
rect 140280 169510 140332 169516
rect 139634 164912 139690 164921
rect 139634 164847 139690 164856
rect 139648 164814 139676 164847
rect 139636 164808 139688 164814
rect 139636 164750 139688 164756
rect 139634 163552 139690 163561
rect 137612 163516 137664 163522
rect 139634 163487 139690 163496
rect 137612 163458 137664 163464
rect 137624 155090 137652 163458
rect 139648 163454 139676 163487
rect 139636 163448 139688 163454
rect 139636 163390 139688 163396
rect 139634 162192 139690 162201
rect 139544 162156 139596 162162
rect 139634 162127 139690 162136
rect 139544 162098 139596 162104
rect 138900 157940 138952 157946
rect 138900 157882 138952 157888
rect 137612 155084 137664 155090
rect 137612 155026 137664 155032
rect 138912 148193 138940 157882
rect 139556 153769 139584 162098
rect 139648 162094 139676 162127
rect 139636 162088 139688 162094
rect 139636 162030 139688 162036
rect 139634 159336 139690 159345
rect 139634 159271 139636 159280
rect 139688 159271 139690 159280
rect 139636 159242 139688 159248
rect 139634 155120 139690 155129
rect 139634 155055 139636 155064
rect 139688 155055 139690 155064
rect 139636 155026 139688 155032
rect 139542 153760 139598 153769
rect 139542 153695 139598 153704
rect 138898 148184 138954 148193
rect 138898 148119 138954 148128
rect 139636 146788 139688 146794
rect 139636 146730 139688 146736
rect 139648 146697 139676 146730
rect 139634 146688 139690 146697
rect 139634 146623 139690 146632
rect 139636 145428 139688 145434
rect 139636 145370 139688 145376
rect 139648 145337 139676 145370
rect 139634 145328 139690 145337
rect 139634 145263 139690 145272
rect 139636 144068 139688 144074
rect 139636 144010 139688 144016
rect 139648 143977 139676 144010
rect 139634 143968 139690 143977
rect 139634 143903 139690 143912
rect 140292 142617 140320 169510
rect 140554 169128 140610 169137
rect 140554 169063 140610 169072
rect 140568 168962 140596 169063
rect 140556 168956 140608 168962
rect 140556 168898 140608 168904
rect 140554 167768 140610 167777
rect 140554 167703 140610 167712
rect 140568 167602 140596 167703
rect 140556 167596 140608 167602
rect 140556 167538 140608 167544
rect 140554 166408 140610 166417
rect 140554 166343 140610 166352
rect 140568 166242 140596 166343
rect 140556 166236 140608 166242
rect 140556 166178 140608 166184
rect 140464 160728 140516 160734
rect 140464 160670 140516 160676
rect 140646 160696 140702 160705
rect 140370 156616 140426 156625
rect 140370 156551 140426 156560
rect 140278 142608 140334 142617
rect 140278 142543 140334 142552
rect 140384 142034 140412 156551
rect 140476 150913 140504 160670
rect 140646 160631 140702 160640
rect 140832 160660 140884 160666
rect 140556 159368 140608 159374
rect 140556 159310 140608 159316
rect 140462 150904 140518 150913
rect 140462 150839 140518 150848
rect 140568 149553 140596 159310
rect 140660 150942 140688 160631
rect 140832 160602 140884 160608
rect 140738 157976 140794 157985
rect 140738 157911 140794 157920
rect 140648 150936 140700 150942
rect 140648 150878 140700 150884
rect 140752 149582 140780 157911
rect 140844 152409 140872 160602
rect 140830 152400 140886 152409
rect 140830 152335 140886 152344
rect 140740 149576 140792 149582
rect 140554 149544 140610 149553
rect 140740 149518 140792 149524
rect 140554 149479 140610 149488
rect 167788 142232 167840 142238
rect 147914 142200 147970 142209
rect 147914 142135 147970 142144
rect 150674 142200 150730 142209
rect 167786 142200 167788 142209
rect 167840 142200 167842 142209
rect 150730 142158 151024 142186
rect 150674 142135 150730 142144
rect 167786 142135 167842 142144
rect 147454 142064 147510 142073
rect 140372 142028 140424 142034
rect 147160 142022 147454 142050
rect 147454 141999 147510 142008
rect 140372 141970 140424 141976
rect 147928 141914 147956 142135
rect 142408 141886 143388 141914
rect 144308 141886 144644 141914
rect 145228 141886 145288 141914
rect 137612 140668 137664 140674
rect 137612 140610 137664 140616
rect 137624 140441 137652 140610
rect 137610 140432 137666 140441
rect 137610 140367 137666 140376
rect 137624 129833 137652 140367
rect 141844 139920 141896 139926
rect 141842 139888 141844 139897
rect 141896 139888 141898 139897
rect 141842 139823 141898 139832
rect 137610 129824 137666 129833
rect 137610 129759 137666 129768
rect 137612 122036 137664 122042
rect 137612 121978 137664 121984
rect 137518 98544 137574 98553
rect 137518 98479 137574 98488
rect 137624 92297 137652 121978
rect 137704 108232 137756 108238
rect 137704 108174 137756 108180
rect 137610 92288 137666 92297
rect 137610 92223 137666 92232
rect 137716 88897 137744 108174
rect 137794 104120 137850 104129
rect 137794 104055 137850 104064
rect 137808 95289 137836 104055
rect 137794 95280 137850 95289
rect 137794 95215 137850 95224
rect 138162 94600 138218 94609
rect 138162 94535 138218 94544
rect 138176 94434 138204 94535
rect 142408 94434 142436 141886
rect 144616 139246 144644 141886
rect 144604 139240 144656 139246
rect 144604 139182 144656 139188
rect 145260 138770 145288 141886
rect 145352 141886 146240 141914
rect 147928 141886 148232 141914
rect 149092 141886 149152 141914
rect 150104 141886 150440 141914
rect 152036 141886 152096 141914
rect 145248 138764 145300 138770
rect 145248 138706 145300 138712
rect 144234 122344 144290 122353
rect 144234 122279 144290 122288
rect 144248 122042 144276 122279
rect 144236 122036 144288 122042
rect 144236 121978 144288 121984
rect 145352 110958 145380 141886
rect 148204 139897 148232 141886
rect 149124 141121 149152 141886
rect 150412 141354 150440 141886
rect 150400 141348 150452 141354
rect 150400 141290 150452 141296
rect 152068 141121 152096 141886
rect 152620 141886 152956 141914
rect 153968 141886 154580 141914
rect 154888 141886 155224 141914
rect 155900 141886 156144 141914
rect 156820 141886 157524 141914
rect 157832 141886 158168 141914
rect 158752 141886 158812 141914
rect 159764 141886 160284 141914
rect 160684 141886 161020 141914
rect 161696 141886 162032 141914
rect 149110 141112 149166 141121
rect 149110 141047 149166 141056
rect 152054 141112 152110 141121
rect 152054 141047 152110 141056
rect 152620 139926 152648 141886
rect 152608 139920 152660 139926
rect 148190 139888 148246 139897
rect 152608 139862 152660 139868
rect 148190 139823 148246 139832
rect 150492 139852 150544 139858
rect 150492 139794 150544 139800
rect 150504 130338 150532 139794
rect 151780 139784 151832 139790
rect 151780 139726 151832 139732
rect 150584 139580 150636 139586
rect 150584 139522 150636 139528
rect 149296 130332 149348 130338
rect 149296 130274 149348 130280
rect 150492 130332 150544 130338
rect 150492 130274 150544 130280
rect 149308 128708 149336 130274
rect 150596 128722 150624 139522
rect 151792 130338 151820 139726
rect 153344 139648 153396 139654
rect 153344 139590 153396 139596
rect 151872 139512 151924 139518
rect 151872 139454 151924 139460
rect 151044 130332 151096 130338
rect 151044 130274 151096 130280
rect 151780 130332 151832 130338
rect 151780 130274 151832 130280
rect 150150 128694 150624 128722
rect 151056 128708 151084 130274
rect 151884 128722 151912 139454
rect 153356 130082 153384 139590
rect 154552 130406 154580 141886
rect 154724 139716 154776 139722
rect 154724 139658 154776 139664
rect 154632 139376 154684 139382
rect 154632 139318 154684 139324
rect 154540 130400 154592 130406
rect 154540 130342 154592 130348
rect 153712 130332 153764 130338
rect 153712 130274 153764 130280
rect 153264 130054 153384 130082
rect 153264 128722 153292 130054
rect 151884 128694 151990 128722
rect 152818 128694 153292 128722
rect 153724 128708 153752 130274
rect 154644 128708 154672 139318
rect 154736 130338 154764 139658
rect 155196 139450 155224 141886
rect 155184 139444 155236 139450
rect 155184 139386 155236 139392
rect 156012 139444 156064 139450
rect 156012 139386 156064 139392
rect 155920 139308 155972 139314
rect 155920 139250 155972 139256
rect 154724 130332 154776 130338
rect 154724 130274 154776 130280
rect 155932 130082 155960 139250
rect 156024 130474 156052 139386
rect 156116 130542 156144 141886
rect 157392 139512 157444 139518
rect 157392 139454 157444 139460
rect 156104 130536 156156 130542
rect 156104 130478 156156 130484
rect 156012 130468 156064 130474
rect 156012 130410 156064 130416
rect 157300 130400 157352 130406
rect 157300 130342 157352 130348
rect 156380 130332 156432 130338
rect 156380 130274 156432 130280
rect 155840 130054 155960 130082
rect 155840 128722 155868 130054
rect 155486 128694 155868 128722
rect 156392 128708 156420 130274
rect 157312 128708 157340 130342
rect 157404 130338 157432 139454
rect 157496 130406 157524 141886
rect 158140 139586 158168 141886
rect 158128 139580 158180 139586
rect 158128 139522 158180 139528
rect 158784 131358 158812 141886
rect 158864 139580 158916 139586
rect 158864 139522 158916 139528
rect 158772 131352 158824 131358
rect 158772 131294 158824 131300
rect 158128 130468 158180 130474
rect 158128 130410 158180 130416
rect 157484 130400 157536 130406
rect 157484 130342 157536 130348
rect 157392 130332 157444 130338
rect 157392 130274 157444 130280
rect 158140 128708 158168 130410
rect 158876 130338 158904 139522
rect 160256 130746 160284 141886
rect 160992 139586 161020 141886
rect 162004 139586 162032 141886
rect 162280 141886 162616 141914
rect 163292 141886 163628 141914
rect 164548 141886 164608 141914
rect 162280 139858 162308 141886
rect 162268 139852 162320 139858
rect 162268 139794 162320 139800
rect 163292 139654 163320 141886
rect 164580 139790 164608 141886
rect 165224 141886 165560 141914
rect 166144 141886 166480 141914
rect 167340 141886 167492 141914
rect 164568 139784 164620 139790
rect 164568 139726 164620 139732
rect 163280 139648 163332 139654
rect 163280 139590 163332 139596
rect 160980 139580 161032 139586
rect 160980 139522 161032 139528
rect 161624 139580 161676 139586
rect 161624 139522 161676 139528
rect 161992 139580 162044 139586
rect 161992 139522 162044 139528
rect 163004 139580 163056 139586
rect 163004 139522 163056 139528
rect 161636 131426 161664 139522
rect 161624 131420 161676 131426
rect 161624 131362 161676 131368
rect 161716 131352 161768 131358
rect 161716 131294 161768 131300
rect 160244 130740 160296 130746
rect 160244 130682 160296 130688
rect 159048 130536 159100 130542
rect 159048 130478 159100 130484
rect 158864 130332 158916 130338
rect 158864 130274 158916 130280
rect 159060 128708 159088 130478
rect 159968 130400 160020 130406
rect 159968 130342 160020 130348
rect 159980 128708 160008 130342
rect 160796 130332 160848 130338
rect 160796 130274 160848 130280
rect 160808 128708 160836 130274
rect 161728 128708 161756 131294
rect 162636 130740 162688 130746
rect 162636 130682 162688 130688
rect 162648 128708 162676 130682
rect 163016 130338 163044 139522
rect 165224 139450 165252 141886
rect 166144 139926 166172 141886
rect 166132 139920 166184 139926
rect 166132 139862 166184 139868
rect 167340 139722 167368 141886
rect 167800 141354 167828 142135
rect 168076 141886 168412 141914
rect 169088 141886 169424 141914
rect 170008 141886 170344 141914
rect 167788 141348 167840 141354
rect 167788 141290 167840 141296
rect 167328 139716 167380 139722
rect 167328 139658 167380 139664
rect 165212 139444 165264 139450
rect 165212 139386 165264 139392
rect 168076 139382 168104 141886
rect 168064 139376 168116 139382
rect 168064 139318 168116 139324
rect 169088 139314 169116 141886
rect 170008 139518 170036 141886
rect 169996 139512 170048 139518
rect 169996 139454 170048 139460
rect 169076 139308 169128 139314
rect 169076 139250 169128 139256
rect 170640 139240 170692 139246
rect 170640 139182 170692 139188
rect 163464 131420 163516 131426
rect 163464 131362 163516 131368
rect 163004 130332 163056 130338
rect 163004 130274 163056 130280
rect 163476 128708 163504 131362
rect 164384 130332 164436 130338
rect 164384 130274 164436 130280
rect 164396 128708 164424 130274
rect 170652 125442 170680 139182
rect 169996 125436 170048 125442
rect 169996 125378 170048 125384
rect 170640 125436 170692 125442
rect 170640 125378 170692 125384
rect 167878 118808 167934 118817
rect 167878 118743 167934 118752
rect 167892 117894 167920 118743
rect 167880 117888 167932 117894
rect 167880 117830 167932 117836
rect 147362 113640 147418 113649
rect 147362 113575 147418 113584
rect 147376 112998 147404 113575
rect 147364 112992 147416 112998
rect 147364 112934 147416 112940
rect 147376 112561 147404 112934
rect 147362 112552 147418 112561
rect 147362 112487 147418 112496
rect 145340 110952 145392 110958
rect 145340 110894 145392 110900
rect 143958 108880 144014 108889
rect 143958 108815 144014 108824
rect 143972 108238 144000 108815
rect 143960 108232 144012 108238
rect 143960 108174 144012 108180
rect 168246 98816 168302 98825
rect 168246 98751 168302 98760
rect 168260 98650 168288 98751
rect 168248 98644 168300 98650
rect 168248 98586 168300 98592
rect 169260 98644 169312 98650
rect 169260 98586 169312 98592
rect 144418 95552 144474 95561
rect 144418 95487 144474 95496
rect 138164 94428 138216 94434
rect 138164 94370 138216 94376
rect 142396 94428 142448 94434
rect 142396 94370 142448 94376
rect 137702 88888 137758 88897
rect 137702 88823 137758 88832
rect 138164 85520 138216 85526
rect 138162 85488 138164 85497
rect 138216 85488 138218 85497
rect 138162 85423 138218 85432
rect 139636 76408 139688 76414
rect 139636 76350 139688 76356
rect 139648 75297 139676 76350
rect 142408 75682 142436 94370
rect 144432 85526 144460 95487
rect 169272 93006 169300 98586
rect 169260 93000 169312 93006
rect 169260 92942 169312 92948
rect 155366 89160 155422 89169
rect 155302 89118 155366 89146
rect 155366 89095 155422 89104
rect 149216 87362 149244 88860
rect 149204 87356 149256 87362
rect 149204 87298 149256 87304
rect 149768 87294 149796 88860
rect 149756 87288 149808 87294
rect 149756 87230 149808 87236
rect 150412 87158 150440 88860
rect 151056 87226 151084 88860
rect 151622 88846 152004 88874
rect 151044 87220 151096 87226
rect 151044 87162 151096 87168
rect 150400 87152 150452 87158
rect 150400 87094 150452 87100
rect 150584 87084 150636 87090
rect 150584 87026 150636 87032
rect 149204 87016 149256 87022
rect 149204 86958 149256 86964
rect 146444 86948 146496 86954
rect 146444 86890 146496 86896
rect 145064 86812 145116 86818
rect 145064 86754 145116 86760
rect 144420 85520 144472 85526
rect 144420 85462 144472 85468
rect 145076 75818 145104 86754
rect 146456 75818 146484 86890
rect 147824 86880 147876 86886
rect 147824 86822 147876 86828
rect 147836 75818 147864 86822
rect 149216 75818 149244 86958
rect 150596 75818 150624 87026
rect 151976 78998 152004 88846
rect 152252 86274 152280 88860
rect 152910 88846 153292 88874
rect 152240 86268 152292 86274
rect 152240 86210 152292 86216
rect 153264 81122 153292 88846
rect 153448 86750 153476 88860
rect 154106 88846 154672 88874
rect 154644 87378 154672 88846
rect 154736 87498 154764 88860
rect 154724 87492 154776 87498
rect 154724 87434 154776 87440
rect 155932 87401 155960 88860
rect 155918 87392 155974 87401
rect 154644 87350 154764 87378
rect 153436 86744 153488 86750
rect 153436 86686 153488 86692
rect 154632 86744 154684 86750
rect 154632 86686 154684 86692
rect 153344 86268 153396 86274
rect 153344 86210 153396 86216
rect 153080 81094 153292 81122
rect 151964 78992 152016 78998
rect 151964 78934 152016 78940
rect 151964 78856 152016 78862
rect 151964 78798 152016 78804
rect 151976 75818 152004 78798
rect 153080 78590 153108 81094
rect 153356 80986 153384 86210
rect 153264 80958 153384 80986
rect 153264 78726 153292 80958
rect 153344 79196 153396 79202
rect 153344 79138 153396 79144
rect 153252 78720 153304 78726
rect 153252 78662 153304 78668
rect 153068 78584 153120 78590
rect 153068 78526 153120 78532
rect 153356 75818 153384 79138
rect 154540 79128 154592 79134
rect 154540 79070 154592 79076
rect 154552 78522 154580 79070
rect 154644 78658 154672 86686
rect 154736 79134 154764 87350
rect 155918 87327 155974 87336
rect 156576 86857 156604 88860
rect 156932 87356 156984 87362
rect 156932 87298 156984 87304
rect 156562 86848 156618 86857
rect 156562 86783 156618 86792
rect 156840 86336 156892 86342
rect 156840 86278 156892 86284
rect 156852 79202 156880 86278
rect 156944 79202 156972 87298
rect 157220 86721 157248 88860
rect 157772 87129 157800 88860
rect 157758 87120 157814 87129
rect 157758 87055 157814 87064
rect 158416 86993 158444 88860
rect 158956 87288 159008 87294
rect 158956 87230 159008 87236
rect 158402 86984 158458 86993
rect 158402 86919 158458 86928
rect 157206 86712 157262 86721
rect 157206 86647 157262 86656
rect 156840 79196 156892 79202
rect 156840 79138 156892 79144
rect 156932 79196 156984 79202
rect 156932 79138 156984 79144
rect 157576 79196 157628 79202
rect 157576 79138 157628 79144
rect 154724 79128 154776 79134
rect 154724 79070 154776 79076
rect 156104 78992 156156 78998
rect 156104 78934 156156 78940
rect 154724 78924 154776 78930
rect 154724 78866 154776 78872
rect 154632 78652 154684 78658
rect 154632 78594 154684 78600
rect 154540 78516 154592 78522
rect 154540 78458 154592 78464
rect 154736 75818 154764 78866
rect 156116 75818 156144 78934
rect 157588 75818 157616 79138
rect 158968 75818 158996 87230
rect 159060 87129 159088 88860
rect 159336 88846 159626 88874
rect 159046 87120 159102 87129
rect 159046 87055 159102 87064
rect 159336 86818 159364 88846
rect 159600 87152 159652 87158
rect 159600 87094 159652 87100
rect 159324 86812 159376 86818
rect 159324 86754 159376 86760
rect 159612 79202 159640 87094
rect 160256 86954 160284 88860
rect 160244 86948 160296 86954
rect 160244 86890 160296 86896
rect 160900 86886 160928 88860
rect 161452 87022 161480 88860
rect 161716 87220 161768 87226
rect 161716 87162 161768 87168
rect 161440 87016 161492 87022
rect 161440 86958 161492 86964
rect 160888 86880 160940 86886
rect 160888 86822 160940 86828
rect 160980 86880 161032 86886
rect 160980 86822 161032 86828
rect 159600 79196 159652 79202
rect 159600 79138 159652 79144
rect 160336 79196 160388 79202
rect 160336 79138 160388 79144
rect 160348 75818 160376 79138
rect 160992 78862 161020 86822
rect 160980 78856 161032 78862
rect 160980 78798 161032 78804
rect 161728 75818 161756 87162
rect 162096 87090 162124 88860
rect 162084 87084 162136 87090
rect 162084 87026 162136 87032
rect 162740 86886 162768 88860
rect 162728 86880 162780 86886
rect 162728 86822 162780 86828
rect 163292 86342 163320 88860
rect 163476 88846 163950 88874
rect 164488 88846 164594 88874
rect 163280 86336 163332 86342
rect 163280 86278 163332 86284
rect 163476 86154 163504 88846
rect 163200 86126 163504 86154
rect 163200 78930 163228 86126
rect 164488 78998 164516 88846
rect 164476 78992 164528 78998
rect 164476 78934 164528 78940
rect 163188 78924 163240 78930
rect 163188 78866 163240 78872
rect 163096 78788 163148 78794
rect 163096 78730 163148 78736
rect 163108 75818 163136 78730
rect 164568 78720 164620 78726
rect 164568 78662 164620 78668
rect 164580 75818 164608 78662
rect 167328 78652 167380 78658
rect 167328 78594 167380 78600
rect 165948 78584 166000 78590
rect 165948 78526 166000 78532
rect 165960 75818 165988 78526
rect 167340 75818 167368 78594
rect 168708 78516 168760 78522
rect 168708 78458 168760 78464
rect 168720 75818 168748 78458
rect 170008 76090 170036 125378
rect 172032 87498 172060 225610
rect 174780 211728 174832 211734
rect 174780 211670 174832 211676
rect 174792 209694 174820 211670
rect 174780 209688 174832 209694
rect 174780 209630 174832 209636
rect 174884 175762 174912 268926
rect 189328 260898 189356 268994
rect 189512 268990 189540 269470
rect 197516 268990 197544 269538
rect 203772 269058 203800 271916
rect 203760 269052 203812 269058
rect 203760 268994 203812 269000
rect 189500 268984 189552 268990
rect 189500 268926 189552 268932
rect 197504 268984 197556 268990
rect 197504 268926 197556 268932
rect 210948 268310 210976 271916
rect 218032 268417 218060 271916
rect 218018 268408 218074 268417
rect 218018 268343 218074 268352
rect 209924 268304 209976 268310
rect 209924 268246 209976 268252
rect 210936 268304 210988 268310
rect 210936 268246 210988 268252
rect 209936 261306 209964 268246
rect 203852 261300 203904 261306
rect 203852 261242 203904 261248
rect 209924 261300 209976 261306
rect 209924 261242 209976 261248
rect 189316 260892 189368 260898
rect 189316 260834 189368 260840
rect 190512 260892 190564 260898
rect 190512 260834 190564 260840
rect 190524 257772 190552 260834
rect 203864 257772 203892 261242
rect 225208 260694 225236 271916
rect 225932 262932 225984 262938
rect 225932 262874 225984 262880
rect 225840 261436 225892 261442
rect 225840 261378 225892 261384
rect 217192 260688 217244 260694
rect 217192 260630 217244 260636
rect 225196 260688 225248 260694
rect 225196 260630 225248 260636
rect 217204 257772 217232 260630
rect 182322 257392 182378 257401
rect 182322 257327 182378 257336
rect 182336 257294 182364 257327
rect 179196 257288 179248 257294
rect 179196 257230 179248 257236
rect 182324 257288 182376 257294
rect 182324 257230 182376 257236
rect 178276 255928 178328 255934
rect 178276 255870 178328 255876
rect 176160 254500 176212 254506
rect 176160 254442 176212 254448
rect 176252 254500 176304 254506
rect 176252 254442 176304 254448
rect 176172 244714 176200 254442
rect 176264 246958 176292 254442
rect 178288 247910 178316 255870
rect 178920 253140 178972 253146
rect 178920 253082 178972 253088
rect 178276 247904 178328 247910
rect 178276 247846 178328 247852
rect 176252 246952 176304 246958
rect 176252 246894 176304 246900
rect 176160 244708 176212 244714
rect 176160 244650 176212 244656
rect 178932 244442 178960 253082
rect 179012 251848 179064 251854
rect 179012 251790 179064 251796
rect 178920 244436 178972 244442
rect 178920 244378 178972 244384
rect 179024 242810 179052 251790
rect 179208 249474 179236 257230
rect 225656 256540 225708 256546
rect 225656 256482 225708 256488
rect 182322 256440 182378 256449
rect 182322 256375 182378 256384
rect 181036 256132 181088 256138
rect 181036 256074 181088 256080
rect 181680 256132 181732 256138
rect 181680 256074 181732 256080
rect 181048 256002 181076 256074
rect 181036 255996 181088 256002
rect 181036 255938 181088 255944
rect 181586 255624 181642 255633
rect 181586 255559 181642 255568
rect 181600 254506 181628 255559
rect 181588 254500 181640 254506
rect 181588 254442 181640 254448
rect 181586 252904 181642 252913
rect 181586 252839 181642 252848
rect 180300 251916 180352 251922
rect 180300 251858 180352 251864
rect 179196 249468 179248 249474
rect 179196 249410 179248 249416
rect 180312 242849 180340 251858
rect 181600 251854 181628 252839
rect 181588 251848 181640 251854
rect 181588 251790 181640 251796
rect 181496 250284 181548 250290
rect 181496 250226 181548 250232
rect 181508 249785 181536 250226
rect 181494 249776 181550 249785
rect 181494 249711 181550 249720
rect 181692 246362 181720 256074
rect 182336 255934 182364 256375
rect 182324 255928 182376 255934
rect 182324 255870 182376 255876
rect 225562 255624 225618 255633
rect 222712 255588 222764 255594
rect 225562 255559 225618 255568
rect 222712 255530 222764 255536
rect 182322 254672 182378 254681
rect 182322 254607 182378 254616
rect 182336 254574 182364 254607
rect 182324 254568 182376 254574
rect 182324 254510 182376 254516
rect 181770 253856 181826 253865
rect 181770 253791 181826 253800
rect 181784 253146 181812 253791
rect 181772 253140 181824 253146
rect 181772 253082 181824 253088
rect 222724 253026 222752 255530
rect 225576 254574 225604 255559
rect 225564 254568 225616 254574
rect 225564 254510 225616 254516
rect 225378 253856 225434 253865
rect 225378 253791 225434 253800
rect 225392 253146 225420 253791
rect 225380 253140 225432 253146
rect 225380 253082 225432 253088
rect 222632 252998 222752 253026
rect 181770 252088 181826 252097
rect 181770 252023 181826 252032
rect 181784 251786 181812 252023
rect 181772 251780 181824 251786
rect 181772 251722 181824 251728
rect 182322 251136 182378 251145
rect 182322 251071 182378 251080
rect 222632 251122 222660 252998
rect 222632 251094 222844 251122
rect 182336 250358 182364 251071
rect 182324 250352 182376 250358
rect 182230 250320 182286 250329
rect 182324 250294 182376 250300
rect 182230 250255 182286 250264
rect 182244 248998 182272 250255
rect 182232 248992 182284 248998
rect 182232 248934 182284 248940
rect 181956 248924 182008 248930
rect 181956 248866 182008 248872
rect 181864 248856 181916 248862
rect 181864 248798 181916 248804
rect 181876 248289 181904 248798
rect 181968 248697 181996 248866
rect 181954 248688 182010 248697
rect 181954 248623 182010 248632
rect 181862 248280 181918 248289
rect 181862 248215 181918 248224
rect 182324 247564 182376 247570
rect 182324 247506 182376 247512
rect 182336 247337 182364 247506
rect 182322 247328 182378 247337
rect 182322 247263 182378 247272
rect 181600 246334 181720 246362
rect 181600 245569 181628 246334
rect 181680 246204 181732 246210
rect 181680 246146 181732 246152
rect 181692 246113 181720 246146
rect 181678 246104 181734 246113
rect 181678 246039 181734 246048
rect 181586 245560 181642 245569
rect 181586 245495 181642 245504
rect 182048 244708 182100 244714
rect 182048 244650 182100 244656
rect 182060 244617 182088 244650
rect 182046 244608 182102 244617
rect 182046 244543 182102 244552
rect 222632 243506 222660 251094
rect 222816 251038 222844 251094
rect 222804 251032 222856 251038
rect 222804 250974 222856 250980
rect 225378 250320 225434 250329
rect 225378 250255 225434 250264
rect 225392 248998 225420 250255
rect 225380 248992 225432 248998
rect 225380 248934 225432 248940
rect 225668 247609 225696 256482
rect 225746 252904 225802 252913
rect 225746 252839 225802 252848
rect 225760 251786 225788 252839
rect 225748 251780 225800 251786
rect 225748 251722 225800 251728
rect 225852 248425 225880 261378
rect 225944 249377 225972 262874
rect 228612 262326 228640 333730
rect 230806 333144 230862 333153
rect 230912 333114 230940 335906
rect 233476 335896 233528 335902
rect 233474 335864 233476 335873
rect 233528 335864 233530 335873
rect 233474 335799 233530 335808
rect 233476 334468 233528 334474
rect 233476 334410 233528 334416
rect 231360 334264 231412 334270
rect 231360 334206 231412 334212
rect 230806 333079 230862 333088
rect 230900 333108 230952 333114
rect 230820 332994 230848 333079
rect 230900 333050 230952 333056
rect 230820 332966 230940 332994
rect 230912 332201 230940 332966
rect 230898 332192 230954 332201
rect 230898 332127 230954 332136
rect 230808 331612 230860 331618
rect 230808 331554 230860 331560
rect 230820 330841 230848 331554
rect 230806 330832 230862 330841
rect 230806 330767 230862 330776
rect 230716 326988 230768 326994
rect 230716 326930 230768 326936
rect 230728 298473 230756 326930
rect 230820 307857 230848 330767
rect 230912 310985 230940 332127
rect 231372 329034 231400 334206
rect 233488 333969 233516 334410
rect 233672 334377 233700 338762
rect 233764 338185 233792 341414
rect 233750 338176 233806 338185
rect 233750 338111 233806 338120
rect 233658 334368 233714 334377
rect 233658 334303 233714 334312
rect 233474 333960 233530 333969
rect 233474 333895 233530 333904
rect 233476 333108 233528 333114
rect 233476 333050 233528 333056
rect 233488 333017 233516 333050
rect 233474 333008 233530 333017
rect 233474 332943 233530 332952
rect 233476 331748 233528 331754
rect 233476 331690 233528 331696
rect 233488 331521 233516 331690
rect 233474 331512 233530 331521
rect 233474 331447 233530 331456
rect 233474 330288 233530 330297
rect 233474 330223 233530 330232
rect 233488 329102 233516 330223
rect 251966 330152 252022 330161
rect 251856 330110 251966 330138
rect 251966 330087 252022 330096
rect 252610 330152 252666 330161
rect 252666 330110 252776 330138
rect 252610 330087 252666 330096
rect 248852 329974 248912 330002
rect 250784 329974 250844 330002
rect 236248 329838 237412 329866
rect 238332 329838 238668 329866
rect 239252 329838 239588 329866
rect 233476 329096 233528 329102
rect 233476 329038 233528 329044
rect 231360 329028 231412 329034
rect 231360 328970 231412 328976
rect 231084 328960 231136 328966
rect 231084 328902 231136 328908
rect 230990 328792 231046 328801
rect 230990 328727 231046 328736
rect 231004 314113 231032 328727
rect 231096 317950 231124 328902
rect 231372 320369 231400 328970
rect 232004 327464 232056 327470
rect 232004 327406 232056 327412
rect 232016 326994 232044 327406
rect 232096 327124 232148 327130
rect 232096 327066 232148 327072
rect 232004 326988 232056 326994
rect 232004 326930 232056 326936
rect 231358 320360 231414 320369
rect 231358 320295 231414 320304
rect 231084 317944 231136 317950
rect 231084 317886 231136 317892
rect 231360 317944 231412 317950
rect 231360 317886 231412 317892
rect 231372 317241 231400 317886
rect 231358 317232 231414 317241
rect 231358 317167 231414 317176
rect 230990 314104 231046 314113
rect 230990 314039 231046 314048
rect 230898 310976 230954 310985
rect 230898 310911 230954 310920
rect 231452 309716 231504 309722
rect 231452 309658 231504 309664
rect 230806 307848 230862 307857
rect 230806 307783 230862 307792
rect 230714 298464 230770 298473
rect 230714 298399 230770 298408
rect 230716 289112 230768 289118
rect 230714 289080 230716 289089
rect 230768 289080 230770 289089
rect 230714 289015 230770 289024
rect 231358 285272 231414 285281
rect 231358 285207 231414 285216
rect 228600 262320 228652 262326
rect 228600 262262 228652 262268
rect 226300 260076 226352 260082
rect 226300 260018 226352 260024
rect 226208 258648 226260 258654
rect 226208 258590 226260 258596
rect 226116 257288 226168 257294
rect 226116 257230 226168 257236
rect 226022 251136 226078 251145
rect 226022 251071 226078 251080
rect 225930 249368 225986 249377
rect 225930 249303 225986 249312
rect 225838 248416 225894 248425
rect 225838 248351 225894 248360
rect 225654 247600 225710 247609
rect 225654 247535 225710 247544
rect 225380 245524 225432 245530
rect 225380 245466 225432 245472
rect 225392 244889 225420 245466
rect 225378 244880 225434 244889
rect 225378 244815 225434 244824
rect 225564 244776 225616 244782
rect 225564 244718 225616 244724
rect 225576 244073 225604 244718
rect 225562 244064 225618 244073
rect 225562 243999 225618 244008
rect 222448 243478 222660 243506
rect 181036 243416 181088 243422
rect 181034 243384 181036 243393
rect 181088 243384 181090 243393
rect 181034 243319 181090 243328
rect 180298 242840 180354 242849
rect 179012 242804 179064 242810
rect 180298 242775 180354 242784
rect 179012 242746 179064 242752
rect 222002 241982 222200 242010
rect 185648 239342 185676 241860
rect 189236 239721 189264 241860
rect 189222 239712 189278 239721
rect 189222 239647 189278 239656
rect 185636 239336 185688 239342
rect 185636 239278 185688 239284
rect 186464 239336 186516 239342
rect 186464 239278 186516 239284
rect 185084 230292 185136 230298
rect 185084 230234 185136 230240
rect 185096 227716 185124 230234
rect 186476 227578 186504 239278
rect 192916 237001 192944 241860
rect 192902 236992 192958 237001
rect 192902 236927 192958 236936
rect 196504 235194 196532 241860
rect 200184 238594 200212 241860
rect 200172 238588 200224 238594
rect 200172 238530 200224 238536
rect 200184 238361 200212 238530
rect 200170 238352 200226 238361
rect 200170 238287 200226 238296
rect 203772 235874 203800 241860
rect 207452 241738 207480 241860
rect 207268 241710 207480 241738
rect 203760 235868 203812 235874
rect 203760 235810 203812 235816
rect 196492 235188 196544 235194
rect 196492 235130 196544 235136
rect 207268 234961 207296 241710
rect 211040 239721 211068 241860
rect 214720 241738 214748 241860
rect 214168 241710 214748 241738
rect 211026 239712 211082 239721
rect 211026 239647 211082 239656
rect 207254 234952 207310 234961
rect 207254 234887 207310 234896
rect 207268 234446 207296 234887
rect 207256 234440 207308 234446
rect 207256 234382 207308 234388
rect 210016 230428 210068 230434
rect 210016 230370 210068 230376
rect 197504 230360 197556 230366
rect 197504 230302 197556 230308
rect 197516 227716 197544 230302
rect 210028 227716 210056 230370
rect 214168 230298 214196 241710
rect 218308 230366 218336 241860
rect 219766 237808 219822 237817
rect 219766 237743 219822 237752
rect 219780 237234 219808 237743
rect 219768 237228 219820 237234
rect 219768 237170 219820 237176
rect 222172 233834 222200 241982
rect 222448 240673 222476 243478
rect 222434 240664 222490 240673
rect 222434 240599 222490 240608
rect 222802 240664 222858 240673
rect 222802 240599 222858 240608
rect 221056 233828 221108 233834
rect 221056 233770 221108 233776
rect 222160 233828 222212 233834
rect 222160 233770 222212 233776
rect 221068 230434 221096 233770
rect 222816 231046 222844 240599
rect 226036 239274 226064 251071
rect 226128 245841 226156 257230
rect 226220 246657 226248 258590
rect 226312 256546 226340 260018
rect 226390 257392 226446 257401
rect 226390 257327 226446 257336
rect 226300 256540 226352 256546
rect 226300 256482 226352 256488
rect 226298 256440 226354 256449
rect 226298 256375 226354 256384
rect 226312 255934 226340 256375
rect 226300 255928 226352 255934
rect 226300 255870 226352 255876
rect 226298 254672 226354 254681
rect 226298 254607 226300 254616
rect 226352 254607 226354 254616
rect 226300 254578 226352 254584
rect 226404 250290 226432 257327
rect 229980 255996 230032 256002
rect 229980 255938 230032 255944
rect 227218 252088 227274 252097
rect 227218 252023 227274 252032
rect 226392 250284 226444 250290
rect 226392 250226 226444 250232
rect 226206 246648 226262 246657
rect 226206 246583 226262 246592
rect 226114 245832 226170 245841
rect 226114 245767 226170 245776
rect 226392 243416 226444 243422
rect 226392 243358 226444 243364
rect 226300 243144 226352 243150
rect 226298 243112 226300 243121
rect 226352 243112 226354 243121
rect 226298 243047 226354 243056
rect 226404 242305 226432 243358
rect 226390 242296 226446 242305
rect 226390 242231 226446 242240
rect 227232 240634 227260 252023
rect 227312 248992 227364 248998
rect 227312 248934 227364 248940
rect 227220 240628 227272 240634
rect 227220 240570 227272 240576
rect 226024 239268 226076 239274
rect 226024 239210 226076 239216
rect 227324 239206 227352 248934
rect 229992 245530 230020 255938
rect 230072 253140 230124 253146
rect 230072 253082 230124 253088
rect 229980 245524 230032 245530
rect 229980 245466 230032 245472
rect 230084 244714 230112 253082
rect 230072 244708 230124 244714
rect 230072 244650 230124 244656
rect 227312 239200 227364 239206
rect 227312 239142 227364 239148
rect 230990 239032 231046 239041
rect 230990 238967 231046 238976
rect 230900 238588 230952 238594
rect 230900 238530 230952 238536
rect 230912 238361 230940 238530
rect 230898 238352 230954 238361
rect 230898 238287 230954 238296
rect 230912 236026 230940 238287
rect 230728 235998 230940 236026
rect 222620 231040 222672 231046
rect 222620 230982 222672 230988
rect 222804 231040 222856 231046
rect 222804 230982 222856 230988
rect 221056 230428 221108 230434
rect 221056 230370 221108 230376
rect 218296 230360 218348 230366
rect 218296 230302 218348 230308
rect 214156 230292 214208 230298
rect 214156 230234 214208 230240
rect 222632 227646 222660 230982
rect 222436 227640 222488 227646
rect 222620 227640 222672 227646
rect 222488 227588 222554 227594
rect 222436 227582 222554 227588
rect 222620 227582 222672 227588
rect 186464 227572 186516 227578
rect 222448 227566 222554 227582
rect 186464 227514 186516 227520
rect 228600 225328 228652 225334
rect 228600 225270 228652 225276
rect 179286 219584 179342 219593
rect 179286 219519 179342 219528
rect 179300 219282 179328 219519
rect 179288 219276 179340 219282
rect 179288 219218 179340 219224
rect 178920 209688 178972 209694
rect 178920 209630 178972 209636
rect 178932 202865 178960 209630
rect 178918 202856 178974 202865
rect 178918 202791 178974 202800
rect 178920 186840 178972 186846
rect 178920 186782 178972 186788
rect 178932 186273 178960 186782
rect 178918 186264 178974 186273
rect 178918 186199 178974 186208
rect 182428 175830 182456 177940
rect 182416 175824 182468 175830
rect 182416 175766 182468 175772
rect 182968 175824 183020 175830
rect 182968 175766 183020 175772
rect 174872 175756 174924 175762
rect 174872 175698 174924 175704
rect 174884 175218 174912 175698
rect 174872 175212 174924 175218
rect 174872 175154 174924 175160
rect 176160 175212 176212 175218
rect 176160 175154 176212 175160
rect 174780 175144 174832 175150
rect 174780 175086 174832 175092
rect 173582 169128 173638 169137
rect 173582 169063 173638 169072
rect 173490 167768 173546 167777
rect 173490 167703 173546 167712
rect 173398 166408 173454 166417
rect 173398 166343 173454 166352
rect 172938 164912 172994 164921
rect 172938 164847 172994 164856
rect 172756 159300 172808 159306
rect 172756 159242 172808 159248
rect 172768 149553 172796 159242
rect 172952 153730 172980 164847
rect 173122 163552 173178 163561
rect 173122 163487 173178 163496
rect 173136 156518 173164 163487
rect 173412 161634 173440 166343
rect 173228 161606 173440 161634
rect 173124 156512 173176 156518
rect 173124 156454 173176 156460
rect 172940 153724 172992 153730
rect 172940 153666 172992 153672
rect 173228 153662 173256 161606
rect 173308 161544 173360 161550
rect 173308 161486 173360 161492
rect 173320 156625 173348 161486
rect 173504 161362 173532 167703
rect 173412 161334 173532 161362
rect 173306 156616 173362 156625
rect 173306 156551 173362 156560
rect 173308 156512 173360 156518
rect 173308 156454 173360 156460
rect 173216 153656 173268 153662
rect 173216 153598 173268 153604
rect 173320 152370 173348 156454
rect 173412 155090 173440 161334
rect 173492 157940 173544 157946
rect 173492 157882 173544 157888
rect 173400 155084 173452 155090
rect 173400 155026 173452 155032
rect 173400 154948 173452 154954
rect 173400 154890 173452 154896
rect 173412 153769 173440 154890
rect 173398 153760 173454 153769
rect 173398 153695 173454 153704
rect 173308 152364 173360 152370
rect 173308 152306 173360 152312
rect 173504 150618 173532 157882
rect 173596 156450 173624 169063
rect 173766 162192 173822 162201
rect 173766 162127 173822 162136
rect 173676 159368 173728 159374
rect 173674 159336 173676 159345
rect 173728 159336 173730 159345
rect 173674 159271 173730 159280
rect 173676 158076 173728 158082
rect 173676 158018 173728 158024
rect 173688 157985 173716 158018
rect 173674 157976 173730 157985
rect 173674 157911 173730 157920
rect 173676 156512 173728 156518
rect 173676 156454 173728 156460
rect 173584 156444 173636 156450
rect 173584 156386 173636 156392
rect 173582 155120 173638 155129
rect 173582 155055 173584 155064
rect 173636 155055 173638 155064
rect 173584 155026 173636 155032
rect 173584 152432 173636 152438
rect 173582 152400 173584 152409
rect 173636 152400 173638 152409
rect 173582 152335 173638 152344
rect 173688 151690 173716 156454
rect 173676 151684 173728 151690
rect 173676 151626 173728 151632
rect 173780 150942 173808 162127
rect 174042 160696 174098 160705
rect 174042 160631 174044 160640
rect 174096 160631 174098 160640
rect 174044 160602 174096 160608
rect 173860 155152 173912 155158
rect 173860 155094 173912 155100
rect 173768 150936 173820 150942
rect 173582 150904 173638 150913
rect 173768 150878 173820 150884
rect 173582 150839 173638 150848
rect 173596 150806 173624 150839
rect 173584 150800 173636 150806
rect 173584 150742 173636 150748
rect 173872 150754 173900 155094
rect 173872 150726 174084 150754
rect 173952 150664 174004 150670
rect 173504 150590 173900 150618
rect 173952 150606 174004 150612
rect 172754 149544 172810 149553
rect 172754 149479 172810 149488
rect 173584 148216 173636 148222
rect 173582 148184 173584 148193
rect 173636 148184 173638 148193
rect 173582 148119 173638 148128
rect 173872 146697 173900 150590
rect 173858 146688 173914 146697
rect 173858 146623 173914 146632
rect 173964 145337 173992 150606
rect 173950 145328 174006 145337
rect 173950 145263 174006 145272
rect 174056 143977 174084 150726
rect 174042 143968 174098 143977
rect 174042 143903 174098 143912
rect 173582 142608 173638 142617
rect 173582 142543 173638 142552
rect 173596 142034 173624 142543
rect 173584 142028 173636 142034
rect 173584 141970 173636 141976
rect 172020 87492 172072 87498
rect 172020 87434 172072 87440
rect 174792 81854 174820 175086
rect 175514 125472 175570 125481
rect 175514 125407 175516 125416
rect 175568 125407 175570 125416
rect 175516 125378 175568 125384
rect 174872 117888 174924 117894
rect 174872 117830 174924 117836
rect 174884 108889 174912 117830
rect 174870 108880 174926 108889
rect 174870 108815 174926 108824
rect 175516 93000 175568 93006
rect 175516 92942 175568 92948
rect 175528 92297 175556 92942
rect 175514 92288 175570 92297
rect 175514 92223 175570 92232
rect 176172 81922 176200 175154
rect 182980 174985 183008 175766
rect 189512 175762 189540 177940
rect 189316 175756 189368 175762
rect 189316 175698 189368 175704
rect 189500 175756 189552 175762
rect 189500 175698 189552 175704
rect 189328 175218 189356 175698
rect 196688 175694 196716 177940
rect 196676 175688 196728 175694
rect 196676 175630 196728 175636
rect 189316 175212 189368 175218
rect 189316 175154 189368 175160
rect 190604 175212 190656 175218
rect 190604 175154 190656 175160
rect 182966 174976 183022 174985
rect 182966 174911 183022 174920
rect 190616 163946 190644 175154
rect 196688 175150 196716 175630
rect 203772 175218 203800 177940
rect 203760 175212 203812 175218
rect 203760 175154 203812 175160
rect 196676 175144 196728 175150
rect 196676 175086 196728 175092
rect 210948 174810 210976 177940
rect 218032 175529 218060 177940
rect 218018 175520 218074 175529
rect 218018 175455 218074 175464
rect 206520 174804 206572 174810
rect 206520 174746 206572 174752
rect 210936 174804 210988 174810
rect 210936 174746 210988 174752
rect 206532 166854 206560 174746
rect 222160 168616 222212 168622
rect 222160 168558 222212 168564
rect 203852 166848 203904 166854
rect 203852 166790 203904 166796
rect 206520 166848 206572 166854
rect 206520 166790 206572 166796
rect 217192 166848 217244 166854
rect 217192 166790 217244 166796
rect 190616 163918 190736 163946
rect 190708 163674 190736 163918
rect 203864 163796 203892 166790
rect 217204 163796 217232 166790
rect 190538 163646 190736 163674
rect 181770 163416 181826 163425
rect 181770 163351 181826 163360
rect 181310 162464 181366 162473
rect 181310 162399 181366 162408
rect 180298 160968 180354 160977
rect 180298 160903 180354 160912
rect 176252 160660 176304 160666
rect 176252 160602 176304 160608
rect 179012 160660 179064 160666
rect 179012 160602 179064 160608
rect 176264 150874 176292 160602
rect 178920 158008 178972 158014
rect 178920 157950 178972 157956
rect 176252 150868 176304 150874
rect 176252 150810 176304 150816
rect 178932 148222 178960 157950
rect 179024 150806 179052 160602
rect 180312 152438 180340 160903
rect 181324 154954 181352 162399
rect 181678 159880 181734 159889
rect 181678 159815 181734 159824
rect 181496 159368 181548 159374
rect 181496 159310 181548 159316
rect 181402 158928 181458 158937
rect 181402 158863 181458 158872
rect 181416 158014 181444 158863
rect 181508 158234 181536 159310
rect 181692 159306 181720 159815
rect 181680 159300 181732 159306
rect 181680 159242 181732 159248
rect 181508 158206 181720 158234
rect 181404 158008 181456 158014
rect 181404 157950 181456 157956
rect 181312 154948 181364 154954
rect 181312 154890 181364 154896
rect 181404 153724 181456 153730
rect 181404 153666 181456 153672
rect 181416 153225 181444 153666
rect 181402 153216 181458 153225
rect 181402 153151 181458 153160
rect 180300 152432 180352 152438
rect 180300 152374 180352 152380
rect 179012 150800 179064 150806
rect 179012 150742 179064 150748
rect 181692 149553 181720 158206
rect 181784 155090 181812 163351
rect 182322 160696 182378 160705
rect 182322 160631 182324 160640
rect 182376 160631 182378 160640
rect 182324 160602 182376 160608
rect 182322 158112 182378 158121
rect 181864 158076 181916 158082
rect 182322 158047 182378 158056
rect 181864 158018 181916 158024
rect 181772 155084 181824 155090
rect 181772 155026 181824 155032
rect 181678 149544 181734 149553
rect 181678 149479 181734 149488
rect 181876 148873 181904 158018
rect 182336 157946 182364 158047
rect 182324 157940 182376 157946
rect 182324 157882 182376 157888
rect 182322 157160 182378 157169
rect 182322 157095 182378 157104
rect 182336 156518 182364 157095
rect 182324 156512 182376 156518
rect 182324 156454 182376 156460
rect 182140 156444 182192 156450
rect 182140 156386 182192 156392
rect 182152 156081 182180 156386
rect 182322 156344 182378 156353
rect 182322 156279 182378 156288
rect 182138 156072 182194 156081
rect 182138 156007 182194 156016
rect 182336 155158 182364 156279
rect 182324 155152 182376 155158
rect 182324 155094 182376 155100
rect 182324 155016 182376 155022
rect 182322 154984 182324 154993
rect 182376 154984 182378 154993
rect 182322 154919 182378 154928
rect 182324 153656 182376 153662
rect 182322 153624 182324 153633
rect 182376 153624 182378 153633
rect 182322 153559 182378 153568
rect 182324 152364 182376 152370
rect 182324 152306 182376 152312
rect 182336 152137 182364 152306
rect 182322 152128 182378 152137
rect 182322 152063 182378 152072
rect 182324 150936 182376 150942
rect 182322 150904 182324 150913
rect 182376 150904 182378 150913
rect 182232 150868 182284 150874
rect 182322 150839 182378 150848
rect 182232 150810 182284 150816
rect 182244 150641 182272 150810
rect 182230 150632 182286 150641
rect 182230 150567 182286 150576
rect 181862 148864 181918 148873
rect 181862 148799 181918 148808
rect 178920 148216 178972 148222
rect 178920 148158 178972 148164
rect 185648 145434 185676 147884
rect 185636 145428 185688 145434
rect 185636 145370 185688 145376
rect 185084 144748 185136 144754
rect 185084 144690 185136 144696
rect 185096 133740 185124 144690
rect 189236 144521 189264 147884
rect 192916 144657 192944 147884
rect 196504 147762 196532 147884
rect 196228 147734 196532 147762
rect 192902 144648 192958 144657
rect 192902 144583 192958 144592
rect 189222 144512 189278 144521
rect 189222 144447 189278 144456
rect 196228 140577 196256 147734
rect 197504 144816 197556 144822
rect 197504 144758 197556 144764
rect 196214 140568 196270 140577
rect 196214 140503 196270 140512
rect 197516 133740 197544 144758
rect 200184 142850 200212 147884
rect 203772 143297 203800 147884
rect 207452 147762 207480 147884
rect 207268 147734 207480 147762
rect 203758 143288 203814 143297
rect 203758 143223 203814 143232
rect 200172 142844 200224 142850
rect 200172 142786 200224 142792
rect 207268 141121 207296 147734
rect 211040 144890 211068 147884
rect 211028 144884 211080 144890
rect 211028 144826 211080 144832
rect 214720 144754 214748 147884
rect 218308 144822 218336 147884
rect 218296 144816 218348 144822
rect 218296 144758 218348 144764
rect 214708 144748 214760 144754
rect 214708 144690 214760 144696
rect 221988 144414 222016 147884
rect 222172 145434 222200 168558
rect 225208 166854 225236 177940
rect 226024 168956 226076 168962
rect 226024 168898 226076 168904
rect 225932 167596 225984 167602
rect 225932 167538 225984 167544
rect 225196 166848 225248 166854
rect 225196 166790 225248 166796
rect 225840 166236 225892 166242
rect 225840 166178 225892 166184
rect 225656 164808 225708 164814
rect 225656 164750 225708 164756
rect 222436 161612 222488 161618
rect 222436 161554 222488 161560
rect 222448 157146 222476 161554
rect 222804 157192 222856 157198
rect 222448 157140 222804 157146
rect 222448 157134 222856 157140
rect 222448 157118 222844 157134
rect 222160 145428 222212 145434
rect 222160 145370 222212 145376
rect 216180 144408 216232 144414
rect 216180 144350 216232 144356
rect 221976 144408 222028 144414
rect 221976 144350 222028 144356
rect 207254 141112 207310 141121
rect 207254 141047 207310 141056
rect 207898 141112 207954 141121
rect 207898 141047 207954 141056
rect 207912 140606 207940 141047
rect 207900 140600 207952 140606
rect 207900 140542 207952 140548
rect 216192 136458 216220 144350
rect 219674 142064 219730 142073
rect 219674 141999 219676 142008
rect 219728 141999 219730 142008
rect 219676 141970 219728 141976
rect 210016 136452 210068 136458
rect 210016 136394 210068 136400
rect 216180 136452 216232 136458
rect 216180 136394 216232 136400
rect 210028 133740 210056 136394
rect 222448 133754 222476 157118
rect 225668 152681 225696 164750
rect 225746 160696 225802 160705
rect 225746 160631 225802 160640
rect 225654 152672 225710 152681
rect 225654 152607 225710 152616
rect 225760 150942 225788 160631
rect 225852 153633 225880 166178
rect 225944 154449 225972 167538
rect 226036 155401 226064 168898
rect 226300 163516 226352 163522
rect 226300 163458 226352 163464
rect 226312 163425 226340 163458
rect 226392 163448 226444 163454
rect 226298 163416 226354 163425
rect 226392 163390 226444 163396
rect 226298 163351 226354 163360
rect 226206 162464 226262 162473
rect 226206 162399 226262 162408
rect 226220 162094 226248 162399
rect 226404 162314 226432 163390
rect 226312 162286 226432 162314
rect 226208 162088 226260 162094
rect 226208 162030 226260 162036
rect 226312 161906 226340 162286
rect 226392 162156 226444 162162
rect 226392 162098 226444 162104
rect 226220 161878 226340 161906
rect 226114 159880 226170 159889
rect 226114 159815 226170 159824
rect 226128 159306 226156 159815
rect 226116 159300 226168 159306
rect 226116 159242 226168 159248
rect 226114 157160 226170 157169
rect 226114 157095 226170 157104
rect 226022 155392 226078 155401
rect 226022 155327 226078 155336
rect 225930 154440 225986 154449
rect 225930 154375 225986 154384
rect 225838 153624 225894 153633
rect 225838 153559 225894 153568
rect 225748 150936 225800 150942
rect 225748 150878 225800 150884
rect 225564 150868 225616 150874
rect 225564 150810 225616 150816
rect 225576 150097 225604 150810
rect 225562 150088 225618 150097
rect 225562 150023 225618 150032
rect 225932 149576 225984 149582
rect 225932 149518 225984 149524
rect 225944 148329 225972 149518
rect 225930 148320 225986 148329
rect 225930 148255 225986 148264
rect 226128 145434 226156 157095
rect 226220 151865 226248 161878
rect 226298 161648 226354 161657
rect 226298 161583 226354 161592
rect 226312 160666 226340 161583
rect 226300 160660 226352 160666
rect 226300 160602 226352 160608
rect 226298 158112 226354 158121
rect 226298 158047 226354 158056
rect 226206 151856 226262 151865
rect 226206 151791 226262 151800
rect 226312 149258 226340 158047
rect 226404 156466 226432 162098
rect 227218 158928 227274 158937
rect 227218 158863 227274 158872
rect 226404 156438 226524 156466
rect 226390 156344 226446 156353
rect 226390 156279 226446 156288
rect 226404 149394 226432 156279
rect 226496 150913 226524 156438
rect 226482 150904 226538 150913
rect 226482 150839 226538 150848
rect 226404 149366 226524 149394
rect 226312 149230 226432 149258
rect 226300 149168 226352 149174
rect 226298 149136 226300 149145
rect 226352 149136 226354 149145
rect 226298 149071 226354 149080
rect 226404 146794 226432 149230
rect 226392 146788 226444 146794
rect 226392 146730 226444 146736
rect 226116 145428 226168 145434
rect 226116 145370 226168 145376
rect 226496 144074 226524 149366
rect 227232 148222 227260 158863
rect 227220 148216 227272 148222
rect 227220 148158 227272 148164
rect 226484 144068 226536 144074
rect 226484 144010 226536 144016
rect 222448 133726 222554 133754
rect 177630 114864 177686 114873
rect 177630 114799 177686 114808
rect 177644 105489 177672 114799
rect 177630 105480 177686 105489
rect 177630 105415 177686 105424
rect 182442 83828 182548 83842
rect 182428 83814 182548 83828
rect 182428 81990 182456 83814
rect 182520 83729 182548 83814
rect 182506 83720 182562 83729
rect 182506 83655 182562 83664
rect 182416 81984 182468 81990
rect 182416 81926 182468 81932
rect 189512 81922 189540 83828
rect 176160 81916 176212 81922
rect 176160 81858 176212 81864
rect 189500 81916 189552 81922
rect 189500 81858 189552 81864
rect 196688 81854 196716 83828
rect 174780 81848 174832 81854
rect 174780 81790 174832 81796
rect 196676 81848 196728 81854
rect 196676 81790 196728 81796
rect 203772 81310 203800 83828
rect 190604 81304 190656 81310
rect 190604 81246 190656 81252
rect 203760 81304 203812 81310
rect 203760 81246 203812 81252
rect 173860 76408 173912 76414
rect 173860 76350 173912 76356
rect 170008 76062 170082 76090
rect 144952 75790 145104 75818
rect 146332 75790 146484 75818
rect 147712 75790 147864 75818
rect 149092 75790 149244 75818
rect 150564 75790 150624 75818
rect 151944 75790 152004 75818
rect 153324 75790 153384 75818
rect 154704 75790 154764 75818
rect 156084 75790 156144 75818
rect 157556 75790 157616 75818
rect 158936 75790 158996 75818
rect 160316 75790 160376 75818
rect 161696 75790 161756 75818
rect 163076 75790 163136 75818
rect 164548 75790 164608 75818
rect 165928 75790 165988 75818
rect 167308 75790 167368 75818
rect 168688 75790 168748 75818
rect 170054 75804 170082 76062
rect 142408 75654 143572 75682
rect 155366 75560 155422 75569
rect 155366 75495 155368 75504
rect 155420 75495 155422 75504
rect 155368 75466 155420 75472
rect 173872 75297 173900 76350
rect 139634 75288 139690 75297
rect 139634 75223 139690 75232
rect 173858 75288 173914 75297
rect 173858 75223 173914 75232
rect 172938 74200 172994 74209
rect 172938 74135 172994 74144
rect 139818 73792 139874 73801
rect 139818 73727 139874 73736
rect 170640 73756 170692 73762
rect 139634 72568 139690 72577
rect 139634 72503 139690 72512
rect 139648 69546 139676 72503
rect 139726 71480 139782 71489
rect 139726 71415 139782 71424
rect 139636 69540 139688 69546
rect 139636 69482 139688 69488
rect 139634 68352 139690 68361
rect 139634 68287 139690 68296
rect 139648 68254 139676 68287
rect 136692 68248 136744 68254
rect 136692 68190 136744 68196
rect 139636 68248 139688 68254
rect 139636 68190 139688 68196
rect 136140 66820 136192 66826
rect 136140 66762 136192 66768
rect 136152 64038 136180 66762
rect 136704 65330 136732 68190
rect 139740 68186 139768 71415
rect 139832 69478 139860 73727
rect 170640 73698 170692 73704
rect 140002 71072 140058 71081
rect 140002 71007 140058 71016
rect 139910 69576 139966 69585
rect 139910 69511 139966 69520
rect 139820 69472 139872 69478
rect 139820 69414 139872 69420
rect 139728 68180 139780 68186
rect 139728 68122 139780 68128
rect 139726 67400 139782 67409
rect 139726 67335 139782 67344
rect 139634 67128 139690 67137
rect 139634 67063 139690 67072
rect 136784 66888 136836 66894
rect 136784 66830 136836 66836
rect 136796 65398 136824 66830
rect 139648 66826 139676 67063
rect 139740 66894 139768 67335
rect 139728 66888 139780 66894
rect 139728 66830 139780 66836
rect 139636 66820 139688 66826
rect 139636 66762 139688 66768
rect 139924 66758 139952 69511
rect 139912 66752 139964 66758
rect 139912 66694 139964 66700
rect 140016 66690 140044 71007
rect 140004 66684 140056 66690
rect 140004 66626 140056 66632
rect 139910 65496 139966 65505
rect 139910 65431 139966 65440
rect 136784 65392 136836 65398
rect 136784 65334 136836 65340
rect 136692 65324 136744 65330
rect 136692 65266 136744 65272
rect 139634 64272 139690 64281
rect 139634 64207 139690 64216
rect 136140 64032 136192 64038
rect 136140 63974 136192 63980
rect 139648 62610 139676 64207
rect 139726 63184 139782 63193
rect 139726 63119 139782 63128
rect 139636 62604 139688 62610
rect 139636 62546 139688 62552
rect 139634 61416 139690 61425
rect 139634 61351 139690 61360
rect 136784 59952 136836 59958
rect 136784 59894 136836 59900
rect 135496 58660 135548 58666
rect 135496 58602 135548 58608
rect 135508 57102 135536 58602
rect 136416 58592 136468 58598
rect 136416 58534 136468 58540
rect 135496 57096 135548 57102
rect 135496 57038 135548 57044
rect 136428 57034 136456 58534
rect 136796 58530 136824 59894
rect 139648 59822 139676 61351
rect 139740 61250 139768 63119
rect 139818 62776 139874 62785
rect 139818 62711 139874 62720
rect 139728 61244 139780 61250
rect 139728 61186 139780 61192
rect 139726 60056 139782 60065
rect 139726 59991 139782 60000
rect 139740 59958 139768 59991
rect 139728 59952 139780 59958
rect 139728 59894 139780 59900
rect 139832 59890 139860 62711
rect 139924 62542 139952 65431
rect 139912 62536 139964 62542
rect 139912 62478 139964 62484
rect 139820 59884 139872 59890
rect 139820 59826 139872 59832
rect 139636 59816 139688 59822
rect 139636 59758 139688 59764
rect 139726 58968 139782 58977
rect 139726 58903 139782 58912
rect 139634 58696 139690 58705
rect 139740 58666 139768 58903
rect 139634 58631 139690 58640
rect 139728 58660 139780 58666
rect 139648 58598 139676 58631
rect 139728 58602 139780 58608
rect 139636 58592 139688 58598
rect 139636 58534 139688 58540
rect 136784 58524 136836 58530
rect 136784 58466 136836 58472
rect 139634 57336 139690 57345
rect 139634 57271 139690 57280
rect 136416 57028 136468 57034
rect 136416 56970 136468 56976
rect 139542 55976 139598 55985
rect 139542 55911 139598 55920
rect 139556 54382 139584 55911
rect 139648 55742 139676 57271
rect 139636 55736 139688 55742
rect 139636 55678 139688 55684
rect 139634 54480 139690 54489
rect 139634 54415 139636 54424
rect 139688 54415 139690 54424
rect 139636 54386 139688 54392
rect 139544 54376 139596 54382
rect 139544 54318 139596 54324
rect 139636 53764 139688 53770
rect 139636 53706 139688 53712
rect 139648 53537 139676 53706
rect 139634 53528 139690 53537
rect 139634 53463 139690 53472
rect 134760 51588 134812 51594
rect 134760 51530 134812 51536
rect 170652 51526 170680 73698
rect 172952 69546 172980 74135
rect 173490 73248 173546 73257
rect 173490 73183 173546 73192
rect 173504 72402 173532 73183
rect 173492 72396 173544 72402
rect 173492 72338 173544 72344
rect 178276 72396 178328 72402
rect 178276 72338 178328 72344
rect 173490 72160 173546 72169
rect 173490 72095 173546 72104
rect 173504 71790 173532 72095
rect 173492 71784 173544 71790
rect 173492 71726 173544 71732
rect 173306 71072 173362 71081
rect 173306 71007 173308 71016
rect 173360 71007 173362 71016
rect 173308 70978 173360 70984
rect 173306 70120 173362 70129
rect 173306 70055 173308 70064
rect 173360 70055 173362 70064
rect 173308 70026 173360 70032
rect 172940 69540 172992 69546
rect 172940 69482 172992 69488
rect 178288 69478 178316 72338
rect 178368 71784 178420 71790
rect 178368 71726 178420 71732
rect 178276 69472 178328 69478
rect 178276 69414 178328 69420
rect 173122 69032 173178 69041
rect 173122 68967 173178 68976
rect 173136 68254 173164 68967
rect 173124 68248 173176 68254
rect 173124 68190 173176 68196
rect 178276 68248 178328 68254
rect 178276 68190 178328 68196
rect 173674 67944 173730 67953
rect 173674 67879 173730 67888
rect 173400 67568 173452 67574
rect 173400 67510 173452 67516
rect 173122 64952 173178 64961
rect 173122 64887 173178 64896
rect 173136 64582 173164 64887
rect 173124 64576 173176 64582
rect 173124 64518 173176 64524
rect 173122 61824 173178 61833
rect 173122 61759 173178 61768
rect 173136 61658 173164 61759
rect 173124 61652 173176 61658
rect 173124 61594 173176 61600
rect 172754 56656 172810 56665
rect 172754 56591 172810 56600
rect 172768 55810 172796 56591
rect 172756 55804 172808 55810
rect 172756 55746 172808 55752
rect 173412 55577 173440 67510
rect 173688 66826 173716 67879
rect 174042 66992 174098 67001
rect 174042 66927 174044 66936
rect 174096 66927 174098 66936
rect 174044 66898 174096 66904
rect 173676 66820 173728 66826
rect 173676 66762 173728 66768
rect 175608 66820 175660 66826
rect 175608 66762 175660 66768
rect 174042 65904 174098 65913
rect 174042 65839 174098 65848
rect 174056 65738 174084 65839
rect 174044 65732 174096 65738
rect 174044 65674 174096 65680
rect 175620 65330 175648 66762
rect 178288 65398 178316 68190
rect 178380 68186 178408 71726
rect 180852 71036 180904 71042
rect 180852 70978 180904 70984
rect 178460 70084 178512 70090
rect 178460 70026 178512 70032
rect 178368 68180 178420 68186
rect 178368 68122 178420 68128
rect 178472 66214 178500 70026
rect 179104 66956 179156 66962
rect 179104 66898 179156 66904
rect 178460 66208 178512 66214
rect 178460 66150 178512 66156
rect 178736 65732 178788 65738
rect 178736 65674 178788 65680
rect 178276 65392 178328 65398
rect 178276 65334 178328 65340
rect 175608 65324 175660 65330
rect 175608 65266 175660 65272
rect 176068 64576 176120 64582
rect 176068 64518 176120 64524
rect 173490 63864 173546 63873
rect 173490 63799 173546 63808
rect 173504 62678 173532 63799
rect 174042 62776 174098 62785
rect 174042 62711 174044 62720
rect 174096 62711 174098 62720
rect 174044 62682 174096 62688
rect 173492 62672 173544 62678
rect 173492 62614 173544 62620
rect 175608 62672 175660 62678
rect 175608 62614 175660 62620
rect 175516 61652 175568 61658
rect 175516 61594 175568 61600
rect 173490 60736 173546 60745
rect 173490 60671 173546 60680
rect 173504 59958 173532 60671
rect 173492 59952 173544 59958
rect 173492 59894 173544 59900
rect 175528 59890 175556 61594
rect 175620 61250 175648 62614
rect 176080 62610 176108 64518
rect 178276 62740 178328 62746
rect 178276 62682 178328 62688
rect 176068 62604 176120 62610
rect 176068 62546 176120 62552
rect 175608 61244 175660 61250
rect 175608 61186 175660 61192
rect 175608 59952 175660 59958
rect 175608 59894 175660 59900
rect 175516 59884 175568 59890
rect 175516 59826 175568 59832
rect 174042 59648 174098 59657
rect 174042 59583 174098 59592
rect 174056 59498 174084 59583
rect 174056 59470 174268 59498
rect 174042 58696 174098 58705
rect 174098 58654 174176 58682
rect 174042 58631 174098 58640
rect 173490 57608 173546 57617
rect 173490 57543 173546 57552
rect 173504 57442 173532 57543
rect 173492 57436 173544 57442
rect 173492 57378 173544 57384
rect 174148 56626 174176 58654
rect 174136 56620 174188 56626
rect 174136 56562 174188 56568
rect 174240 56490 174268 59470
rect 175620 58530 175648 59894
rect 178288 59822 178316 62682
rect 178748 62542 178776 65674
rect 179116 64038 179144 66898
rect 180864 65505 180892 70978
rect 190616 69834 190644 81246
rect 210948 73014 210976 83828
rect 218032 76414 218060 83828
rect 225208 80630 225236 83828
rect 223080 80624 223132 80630
rect 223080 80566 223132 80572
rect 225196 80624 225248 80630
rect 225196 80566 225248 80572
rect 218020 76408 218072 76414
rect 218020 76350 218072 76356
rect 223092 73014 223120 80566
rect 204128 73008 204180 73014
rect 204128 72950 204180 72956
rect 210936 73008 210988 73014
rect 210936 72950 210988 72956
rect 217560 73008 217612 73014
rect 217560 72950 217612 72956
rect 223080 73008 223132 73014
rect 223080 72950 223132 72956
rect 204140 69834 204168 72950
rect 217572 69834 217600 72950
rect 190538 69806 190644 69834
rect 203878 69806 204168 69834
rect 217218 69806 217600 69834
rect 182324 69540 182376 69546
rect 182324 69482 182376 69488
rect 226300 69540 226352 69546
rect 226300 69482 226352 69488
rect 181680 69472 181732 69478
rect 182336 69449 182364 69482
rect 226312 69449 226340 69482
rect 226392 69472 226444 69478
rect 181680 69414 181732 69420
rect 182322 69440 182378 69449
rect 181692 68497 181720 69414
rect 182322 69375 182378 69384
rect 226298 69440 226354 69449
rect 226392 69414 226444 69420
rect 226298 69375 226354 69384
rect 226404 68497 226432 69414
rect 181678 68488 181734 68497
rect 181678 68423 181734 68432
rect 226390 68488 226446 68497
rect 226390 68423 226446 68432
rect 181404 68180 181456 68186
rect 181404 68122 181456 68128
rect 226300 68180 226352 68186
rect 226300 68122 226352 68128
rect 181416 67681 181444 68122
rect 226312 67681 226340 68122
rect 181402 67672 181458 67681
rect 181402 67607 181458 67616
rect 226298 67672 226354 67681
rect 226298 67607 226354 67616
rect 223448 67568 223500 67574
rect 223448 67510 223500 67516
rect 181772 66208 181824 66214
rect 181034 66176 181090 66185
rect 181772 66150 181824 66156
rect 181034 66111 181090 66120
rect 181048 65505 181076 66111
rect 181784 65913 181812 66150
rect 181770 65904 181826 65913
rect 181770 65839 181826 65848
rect 180850 65496 180906 65505
rect 180850 65431 180906 65440
rect 181034 65496 181090 65505
rect 181034 65431 181090 65440
rect 182324 65392 182376 65398
rect 182324 65334 182376 65340
rect 181588 65324 181640 65330
rect 181588 65266 181640 65272
rect 181600 64145 181628 65266
rect 182336 64961 182364 65334
rect 182322 64952 182378 64961
rect 182322 64887 182378 64896
rect 181586 64136 181642 64145
rect 181586 64071 181642 64080
rect 179104 64032 179156 64038
rect 179104 63974 179156 63980
rect 182324 64032 182376 64038
rect 182324 63974 182376 63980
rect 182336 63193 182364 63974
rect 182322 63184 182378 63193
rect 182322 63119 182378 63128
rect 181588 62604 181640 62610
rect 181588 62546 181640 62552
rect 178736 62536 178788 62542
rect 178736 62478 178788 62484
rect 181600 61425 181628 62546
rect 182324 62536 182376 62542
rect 182324 62478 182376 62484
rect 182336 62377 182364 62478
rect 182322 62368 182378 62377
rect 182322 62303 182378 62312
rect 181586 61416 181642 61425
rect 181586 61351 181642 61360
rect 181220 61244 181272 61250
rect 181220 61186 181272 61192
rect 181232 60473 181260 61186
rect 181218 60464 181274 60473
rect 181218 60399 181274 60408
rect 181588 59884 181640 59890
rect 181588 59826 181640 59832
rect 178276 59816 178328 59822
rect 178276 59758 178328 59764
rect 181600 58705 181628 59826
rect 182324 59816 182376 59822
rect 182324 59758 182376 59764
rect 182336 59657 182364 59758
rect 182322 59648 182378 59657
rect 182322 59583 182378 59592
rect 181586 58696 181642 58705
rect 181586 58631 181642 58640
rect 175608 58524 175660 58530
rect 175608 58466 175660 58472
rect 182324 58524 182376 58530
rect 182324 58466 182376 58472
rect 182336 57889 182364 58466
rect 182322 57880 182378 57889
rect 182322 57815 182378 57824
rect 176252 57436 176304 57442
rect 176252 57378 176304 57384
rect 174228 56484 174280 56490
rect 174228 56426 174280 56432
rect 176264 55742 176292 57378
rect 181772 56620 181824 56626
rect 181772 56562 181824 56568
rect 181784 56121 181812 56562
rect 182322 56520 182378 56529
rect 182322 56455 182324 56464
rect 182376 56455 182378 56464
rect 182324 56426 182376 56432
rect 181770 56112 181826 56121
rect 181770 56047 181826 56056
rect 176804 55804 176856 55810
rect 176804 55746 176856 55752
rect 176252 55736 176304 55742
rect 176252 55678 176304 55684
rect 173398 55568 173454 55577
rect 173398 55503 173454 55512
rect 174042 54480 174098 54489
rect 174042 54415 174044 54424
rect 174096 54415 174098 54424
rect 174044 54386 174096 54392
rect 176816 54246 176844 55746
rect 181680 55736 181732 55742
rect 181680 55678 181732 55684
rect 181692 55169 181720 55678
rect 181678 55160 181734 55169
rect 181678 55095 181734 55104
rect 223460 55062 223488 67510
rect 226300 66752 226352 66758
rect 226298 66720 226300 66729
rect 226352 66720 226354 66729
rect 226298 66655 226354 66664
rect 226300 66412 226352 66418
rect 226300 66354 226352 66360
rect 226312 65913 226340 66354
rect 226298 65904 226354 65913
rect 226298 65839 226354 65848
rect 225932 65392 225984 65398
rect 225932 65334 225984 65340
rect 225944 64145 225972 65334
rect 226208 65324 226260 65330
rect 226208 65266 226260 65272
rect 226220 64961 226248 65266
rect 226206 64952 226262 64961
rect 226206 64887 226262 64896
rect 225930 64136 225986 64145
rect 225930 64071 225986 64080
rect 225748 64032 225800 64038
rect 225748 63974 225800 63980
rect 225760 63193 225788 63974
rect 225746 63184 225802 63193
rect 225746 63119 225802 63128
rect 225932 62604 225984 62610
rect 225932 62546 225984 62552
rect 225944 61425 225972 62546
rect 226300 62400 226352 62406
rect 226298 62368 226300 62377
rect 226352 62368 226354 62377
rect 226298 62303 226354 62312
rect 225930 61416 225986 61425
rect 225930 61351 225986 61360
rect 226300 61108 226352 61114
rect 226300 61050 226352 61056
rect 226312 60473 226340 61050
rect 226298 60464 226354 60473
rect 226298 60399 226354 60408
rect 226116 59884 226168 59890
rect 226116 59826 226168 59832
rect 226128 59657 226156 59826
rect 226300 59816 226352 59822
rect 226300 59758 226352 59764
rect 226114 59648 226170 59657
rect 226114 59583 226170 59592
rect 226312 58705 226340 59758
rect 226298 58696 226354 58705
rect 226298 58631 226354 58640
rect 226300 58524 226352 58530
rect 226300 58466 226352 58472
rect 226312 57889 226340 58466
rect 226298 57880 226354 57889
rect 226298 57815 226354 57824
rect 226300 56960 226352 56966
rect 226298 56928 226300 56937
rect 226352 56928 226354 56937
rect 226298 56863 226354 56872
rect 225380 56688 225432 56694
rect 225380 56630 225432 56636
rect 225392 56121 225420 56630
rect 225378 56112 225434 56121
rect 225378 56047 225434 56056
rect 225380 55736 225432 55742
rect 225380 55678 225432 55684
rect 225392 55169 225420 55678
rect 225378 55160 225434 55169
rect 225378 55095 225434 55104
rect 223448 55056 223500 55062
rect 223448 54998 223500 55004
rect 182322 54344 182378 54353
rect 182322 54279 182378 54288
rect 182336 54246 182364 54279
rect 176804 54240 176856 54246
rect 176804 54182 176856 54188
rect 182324 54240 182376 54246
rect 182324 54182 182376 54188
rect 174044 53696 174096 53702
rect 174044 53638 174096 53644
rect 174056 53537 174084 53638
rect 174042 53528 174098 53537
rect 174042 53463 174098 53472
rect 185004 51594 185032 53908
rect 184992 51588 185044 51594
rect 184992 51530 185044 51536
rect 170180 51520 170232 51526
rect 170180 51462 170232 51468
rect 170640 51520 170692 51526
rect 170640 51462 170692 51468
rect 142854 51080 142910 51089
rect 142854 51015 142910 51024
rect 139726 50672 139782 50681
rect 139726 50607 139782 50616
rect 139634 50400 139690 50409
rect 139740 50370 139768 50607
rect 139634 50335 139690 50344
rect 139728 50364 139780 50370
rect 139648 50302 139676 50335
rect 139728 50306 139780 50312
rect 139636 50296 139688 50302
rect 139636 50238 139688 50244
rect 140554 49040 140610 49049
rect 140554 48975 140610 48984
rect 140568 48942 140596 48975
rect 140556 48936 140608 48942
rect 140556 48878 140608 48884
rect 140002 48088 140058 48097
rect 140002 48023 140058 48032
rect 140016 47718 140044 48023
rect 140004 47712 140056 47718
rect 140004 47654 140056 47660
rect 142868 47582 142896 51015
rect 147730 48088 147786 48097
rect 147436 48046 147730 48074
rect 153986 48088 154042 48097
rect 150564 48046 150624 48074
rect 147730 48023 147786 48032
rect 144400 47910 144736 47938
rect 142856 47576 142908 47582
rect 142856 47518 142908 47524
rect 144708 46018 144736 47910
rect 144696 46012 144748 46018
rect 144696 45954 144748 45960
rect 150596 45882 150624 48046
rect 153448 48046 153986 48074
rect 153448 45950 153476 48046
rect 167602 48088 167658 48097
rect 153986 48023 154042 48032
rect 165960 48046 166448 48074
rect 160058 47952 160114 47961
rect 156820 47910 156880 47938
rect 156852 47514 156880 47910
rect 159520 47910 160058 47938
rect 159520 47582 159548 47910
rect 162984 47910 163044 47938
rect 160058 47887 160114 47896
rect 159508 47576 159560 47582
rect 159508 47518 159560 47524
rect 156840 47508 156892 47514
rect 156840 47450 156892 47456
rect 163016 47281 163044 47910
rect 163002 47272 163058 47281
rect 163002 47207 163058 47216
rect 153436 45944 153488 45950
rect 153436 45886 153488 45892
rect 150584 45876 150636 45882
rect 150584 45818 150636 45824
rect 163016 45785 163044 47207
rect 165960 45921 165988 48046
rect 166420 47825 166448 48046
rect 167602 48023 167658 48032
rect 166406 47816 166462 47825
rect 166406 47751 166462 47760
rect 167616 47514 167644 48023
rect 168890 47952 168946 47961
rect 168946 47910 169240 47938
rect 168890 47887 168946 47896
rect 167604 47508 167656 47514
rect 167604 47450 167656 47456
rect 168904 46057 168932 47887
rect 168890 46048 168946 46057
rect 168890 45983 168946 45992
rect 165946 45912 166002 45921
rect 165946 45847 166002 45856
rect 163002 45776 163058 45785
rect 163002 45711 163058 45720
rect 168904 45406 168932 45983
rect 170192 45882 170220 51462
rect 173950 51352 174006 51361
rect 173950 51287 174006 51296
rect 173964 50370 173992 51287
rect 185084 50908 185136 50914
rect 185084 50850 185136 50856
rect 174042 50400 174098 50409
rect 173952 50364 174004 50370
rect 174042 50335 174098 50344
rect 173952 50306 174004 50312
rect 174056 50302 174084 50335
rect 174044 50296 174096 50302
rect 174044 50238 174096 50244
rect 181864 49548 181916 49554
rect 181864 49490 181916 49496
rect 181876 49321 181904 49490
rect 173306 49312 173362 49321
rect 173306 49247 173362 49256
rect 181862 49312 181918 49321
rect 181862 49247 181918 49256
rect 173320 48942 173348 49247
rect 173308 48936 173360 48942
rect 173308 48878 173360 48884
rect 174042 48360 174098 48369
rect 174042 48295 174098 48304
rect 174056 47514 174084 48295
rect 174044 47508 174096 47514
rect 174044 47450 174096 47456
rect 170180 45876 170232 45882
rect 170180 45818 170232 45824
rect 168892 45400 168944 45406
rect 168892 45342 168944 45348
rect 169718 44824 169774 44833
rect 169718 44759 169720 44768
rect 169772 44759 169774 44768
rect 169720 44730 169772 44736
rect 128576 34582 129096 34610
rect 88484 32956 88536 32962
rect 88484 32898 88536 32904
rect 88390 26056 88446 26065
rect 88390 25991 88446 26000
rect 88022 23336 88078 23345
rect 88022 23271 88078 23280
rect 88496 20761 88524 32898
rect 181876 23345 181904 49247
rect 182232 48188 182284 48194
rect 182232 48130 182284 48136
rect 182244 47961 182272 48130
rect 182230 47952 182286 47961
rect 182230 47887 182286 47896
rect 182138 46592 182194 46601
rect 182138 46527 182194 46536
rect 182048 45468 182100 45474
rect 182048 45410 182100 45416
rect 181956 45400 182008 45406
rect 181956 45342 182008 45348
rect 181968 33681 181996 45342
rect 182060 44794 182088 45410
rect 182048 44788 182100 44794
rect 182048 44730 182100 44736
rect 181954 33672 182010 33681
rect 181954 33607 182010 33616
rect 182060 30825 182088 44730
rect 182046 30816 182102 30825
rect 182046 30751 182102 30760
rect 182152 28105 182180 46527
rect 182138 28096 182194 28105
rect 182138 28031 182194 28040
rect 182244 26065 182272 47887
rect 185096 34732 185124 50850
rect 187304 50681 187332 53908
rect 189696 51526 189724 53908
rect 189684 51520 189736 51526
rect 189684 51462 189736 51468
rect 190604 50976 190656 50982
rect 190604 50918 190656 50924
rect 187290 50672 187346 50681
rect 187290 50607 187346 50616
rect 187568 47508 187620 47514
rect 187568 47450 187620 47456
rect 187580 34732 187608 47450
rect 190616 34610 190644 50918
rect 191996 50409 192024 53908
rect 191982 50400 192038 50409
rect 191982 50335 192038 50344
rect 194388 49554 194416 53908
rect 196124 51044 196176 51050
rect 196124 50986 196176 50992
rect 194376 49548 194428 49554
rect 194376 49490 194428 49496
rect 192536 48936 192588 48942
rect 192536 48878 192588 48884
rect 192548 34732 192576 48878
rect 196136 37450 196164 50986
rect 196688 48194 196716 53908
rect 197504 50296 197556 50302
rect 199080 50273 199108 53908
rect 200264 51112 200316 51118
rect 200264 51054 200316 51060
rect 197504 50238 197556 50244
rect 199066 50264 199122 50273
rect 196676 48188 196728 48194
rect 196676 48130 196728 48136
rect 195020 37444 195072 37450
rect 195020 37386 195072 37392
rect 196124 37444 196176 37450
rect 196124 37386 196176 37392
rect 195032 34732 195060 37386
rect 197516 34732 197544 50238
rect 199066 50199 199122 50208
rect 200276 34746 200304 51054
rect 201472 45474 201500 53908
rect 202564 50364 202616 50370
rect 202564 50306 202616 50312
rect 201460 45468 201512 45474
rect 201460 45410 201512 45416
rect 200106 34718 200304 34746
rect 202576 34732 202604 50306
rect 203772 49321 203800 53908
rect 205784 51180 205836 51186
rect 205784 51122 205836 51128
rect 203758 49312 203814 49321
rect 203758 49247 203814 49256
rect 203772 45406 203800 49247
rect 203760 45400 203812 45406
rect 203760 45342 203812 45348
rect 205796 44674 205824 51122
rect 206164 50914 206192 53908
rect 208464 50982 208492 53908
rect 210856 51050 210884 53908
rect 212040 53696 212092 53702
rect 212040 53638 212092 53644
rect 212052 53129 212080 53638
rect 212038 53120 212094 53129
rect 212038 53055 212094 53064
rect 213248 51118 213276 53908
rect 215548 51186 215576 53908
rect 215536 51180 215588 51186
rect 215536 51122 215588 51128
rect 213236 51112 213288 51118
rect 213236 51054 213288 51060
rect 210844 51044 210896 51050
rect 210844 50986 210896 50992
rect 208452 50976 208504 50982
rect 208452 50918 208504 50924
rect 206152 50908 206204 50914
rect 206152 50850 206204 50856
rect 216180 50704 216232 50710
rect 216180 50646 216232 50652
rect 211304 50432 211356 50438
rect 211304 50374 211356 50380
rect 205612 44646 205824 44674
rect 205612 35154 205640 44646
rect 207530 39112 207586 39121
rect 207530 39047 207586 39056
rect 205520 35126 205640 35154
rect 205520 34746 205548 35126
rect 205074 34718 205548 34746
rect 207544 34732 207572 39047
rect 211316 37790 211344 50374
rect 212590 43464 212646 43473
rect 212590 43399 212646 43408
rect 210016 37784 210068 37790
rect 210016 37726 210068 37732
rect 211304 37784 211356 37790
rect 211304 37726 211356 37732
rect 210028 34732 210056 37726
rect 212604 34732 212632 43399
rect 216192 37450 216220 50646
rect 217940 50438 217968 53908
rect 220240 50710 220268 53908
rect 222448 53894 222646 53922
rect 220228 50704 220280 50710
rect 220228 50646 220280 50652
rect 217928 50432 217980 50438
rect 217928 50374 217980 50380
rect 222448 37450 222476 53894
rect 223460 44674 223488 54998
rect 223540 54376 223592 54382
rect 226300 54376 226352 54382
rect 223540 54318 223592 54324
rect 226298 54344 226300 54353
rect 226352 54344 226354 54353
rect 223092 44646 223488 44674
rect 215076 37444 215128 37450
rect 215076 37386 215128 37392
rect 216180 37444 216232 37450
rect 216180 37386 216232 37392
rect 220044 37444 220096 37450
rect 220044 37386 220096 37392
rect 222436 37444 222488 37450
rect 222436 37386 222488 37392
rect 215088 34732 215116 37386
rect 217560 37104 217612 37110
rect 217560 37046 217612 37052
rect 217572 34732 217600 37046
rect 220056 34732 220084 37386
rect 223092 35154 223120 44646
rect 223552 37110 223580 54318
rect 226298 54279 226354 54288
rect 228612 51594 228640 225270
rect 230728 217009 230756 235998
rect 230808 235868 230860 235874
rect 230808 235810 230860 235816
rect 230820 220137 230848 235810
rect 231004 233034 231032 238967
rect 231176 234440 231228 234446
rect 231176 234382 231228 234388
rect 230912 233006 231032 233034
rect 230912 226393 230940 233006
rect 231188 232490 231216 234382
rect 231004 232462 231216 232490
rect 230898 226384 230954 226393
rect 230898 226319 230954 226328
rect 231004 223265 231032 232462
rect 231372 226218 231400 285207
rect 231464 279705 231492 309658
rect 232002 304720 232058 304729
rect 232108 304706 232136 327066
rect 233476 327056 233528 327062
rect 233476 326998 233528 327004
rect 232058 304678 232136 304706
rect 232002 304655 232058 304664
rect 232108 304214 232136 304678
rect 232096 304208 232148 304214
rect 232096 304150 232148 304156
rect 232740 304208 232792 304214
rect 232740 304150 232792 304156
rect 232002 301592 232058 301601
rect 232002 301527 232058 301536
rect 232016 301426 232044 301527
rect 232004 301420 232056 301426
rect 232004 301362 232056 301368
rect 231544 295912 231596 295918
rect 231544 295854 231596 295860
rect 231450 279696 231506 279705
rect 231450 279631 231506 279640
rect 231556 276577 231584 295854
rect 231820 283536 231872 283542
rect 231820 283478 231872 283484
rect 231636 282856 231688 282862
rect 231634 282824 231636 282833
rect 231688 282824 231690 282833
rect 231634 282759 231690 282768
rect 231832 282674 231860 283478
rect 231648 282646 231860 282674
rect 231542 276568 231598 276577
rect 231542 276503 231598 276512
rect 231648 273449 231676 282646
rect 232752 274401 232780 304150
rect 233488 301426 233516 326998
rect 233476 301420 233528 301426
rect 233476 301362 233528 301368
rect 234120 301420 234172 301426
rect 234120 301362 234172 301368
rect 234132 275178 234160 301362
rect 236052 289112 236104 289118
rect 236050 289080 236052 289089
rect 236104 289080 236106 289089
rect 236050 289015 236106 289024
rect 236248 282862 236276 329838
rect 238640 327538 238668 329838
rect 238628 327532 238680 327538
rect 238628 327474 238680 327480
rect 238996 327396 239048 327402
rect 238996 327338 239048 327344
rect 239008 320058 239036 327338
rect 239560 326790 239588 329838
rect 239928 329838 240264 329866
rect 241184 329838 241520 329866
rect 242196 329838 242532 329866
rect 239928 327402 239956 329838
rect 241492 327606 241520 329838
rect 241480 327600 241532 327606
rect 241480 327542 241532 327548
rect 239916 327396 239968 327402
rect 239916 327338 239968 327344
rect 239548 326784 239600 326790
rect 239548 326726 239600 326732
rect 241940 326716 241992 326722
rect 241940 326658 241992 326664
rect 238996 320052 239048 320058
rect 238996 319994 239048 320000
rect 241952 319990 241980 326658
rect 242504 326382 242532 329838
rect 242780 329838 243116 329866
rect 244128 329838 244464 329866
rect 245048 329838 245384 329866
rect 246060 329838 246396 329866
rect 246980 329838 247224 329866
rect 247992 329838 248328 329866
rect 242780 326722 242808 329838
rect 244436 327402 244464 329838
rect 244424 327396 244476 327402
rect 244424 327338 244476 327344
rect 245356 327334 245384 329838
rect 245344 327328 245396 327334
rect 245344 327270 245396 327276
rect 244608 326988 244660 326994
rect 244608 326930 244660 326936
rect 243136 326852 243188 326858
rect 243136 326794 243188 326800
rect 242768 326716 242820 326722
rect 242768 326658 242820 326664
rect 242492 326376 242544 326382
rect 242492 326318 242544 326324
rect 243148 320330 243176 326794
rect 243136 320324 243188 320330
rect 243136 320266 243188 320272
rect 243780 320324 243832 320330
rect 243780 320266 243832 320272
rect 243596 320120 243648 320126
rect 243596 320062 243648 320068
rect 241940 319984 241992 319990
rect 241940 319926 241992 319932
rect 243608 316810 243636 320062
rect 243300 316782 243636 316810
rect 243792 316810 243820 320266
rect 244620 316810 244648 326930
rect 245896 326784 245948 326790
rect 245896 326726 245948 326732
rect 245908 320330 245936 326726
rect 246368 326654 246396 329838
rect 246908 327396 246960 327402
rect 246908 327338 246960 327344
rect 246356 326648 246408 326654
rect 246356 326590 246408 326596
rect 245896 320324 245948 320330
rect 245896 320266 245948 320272
rect 246448 320324 246500 320330
rect 246448 320266 246500 320272
rect 246264 320188 246316 320194
rect 246264 320130 246316 320136
rect 246172 317944 246224 317950
rect 246172 317886 246224 317892
rect 246184 316969 246212 317886
rect 246170 316960 246226 316969
rect 246170 316895 246226 316904
rect 246276 316810 246304 320130
rect 243792 316782 244128 316810
rect 244620 316782 245048 316810
rect 245968 316782 246304 316810
rect 246460 316810 246488 320266
rect 246920 320262 246948 327338
rect 247196 327198 247224 329838
rect 247920 327328 247972 327334
rect 247920 327270 247972 327276
rect 247368 327260 247420 327266
rect 247368 327202 247420 327208
rect 247184 327192 247236 327198
rect 247184 327134 247236 327140
rect 246908 320256 246960 320262
rect 246908 320198 246960 320204
rect 247380 316810 247408 327202
rect 247932 320398 247960 327270
rect 248300 326994 248328 329838
rect 248852 327554 248880 329974
rect 248668 327526 248880 327554
rect 248668 327470 248696 327526
rect 248656 327464 248708 327470
rect 248656 327406 248708 327412
rect 248748 327464 248800 327470
rect 248748 327406 248800 327412
rect 248760 327146 248788 327406
rect 248668 327118 248788 327146
rect 248668 327062 248696 327118
rect 248656 327056 248708 327062
rect 248656 326998 248708 327004
rect 248748 327056 248800 327062
rect 248748 326998 248800 327004
rect 248288 326988 248340 326994
rect 248288 326930 248340 326936
rect 248760 320602 248788 326998
rect 248852 326518 248880 327526
rect 249864 329838 249924 329866
rect 249864 327470 249892 329838
rect 250784 327538 250812 329974
rect 253544 329838 253788 329866
rect 254708 329838 254860 329866
rect 253544 328801 253572 329838
rect 253530 328792 253586 328801
rect 253530 328727 253586 328736
rect 254832 327606 254860 329838
rect 255568 329838 255720 329866
rect 256304 329838 256640 329866
rect 257316 329838 257652 329866
rect 258420 329838 258572 329866
rect 259248 329838 259584 329866
rect 260168 329838 260504 329866
rect 261180 329838 261516 329866
rect 262100 329838 262436 329866
rect 263112 329838 263448 329866
rect 264032 329838 264368 329866
rect 255568 329034 255596 329838
rect 255556 329028 255608 329034
rect 255556 328970 255608 328976
rect 252888 327600 252940 327606
rect 252888 327542 252940 327548
rect 254820 327600 254872 327606
rect 254820 327542 254872 327548
rect 249944 327532 249996 327538
rect 249944 327474 249996 327480
rect 250036 327532 250088 327538
rect 250036 327474 250088 327480
rect 250772 327532 250824 327538
rect 250772 327474 250824 327480
rect 249852 327464 249904 327470
rect 249852 327406 249904 327412
rect 248840 326512 248892 326518
rect 248840 326454 248892 326460
rect 248932 320664 248984 320670
rect 248932 320606 248984 320612
rect 248748 320596 248800 320602
rect 248748 320538 248800 320544
rect 247920 320392 247972 320398
rect 247920 320334 247972 320340
rect 248944 316810 248972 320606
rect 249208 320596 249260 320602
rect 249208 320538 249260 320544
rect 246460 316782 246796 316810
rect 247380 316782 247716 316810
rect 248636 316782 248972 316810
rect 249220 316810 249248 320538
rect 249956 319514 249984 327474
rect 250048 327130 250076 327474
rect 250036 327124 250088 327130
rect 250036 327066 250088 327072
rect 250128 327124 250180 327130
rect 250128 327066 250180 327072
rect 250036 326716 250088 326722
rect 250036 326658 250088 326664
rect 250048 319786 250076 326658
rect 250036 319780 250088 319786
rect 250036 319722 250088 319728
rect 249944 319508 249996 319514
rect 249944 319450 249996 319456
rect 250140 316810 250168 327066
rect 250220 326376 250272 326382
rect 250220 326318 250272 326324
rect 250232 319922 250260 326318
rect 252796 320052 252848 320058
rect 252796 319994 252848 320000
rect 250220 319916 250272 319922
rect 250220 319858 250272 319864
rect 251784 319780 251836 319786
rect 251784 319722 251836 319728
rect 250956 319508 251008 319514
rect 250956 319450 251008 319456
rect 250968 316810 250996 319450
rect 251796 316810 251824 319722
rect 252808 316810 252836 319994
rect 252900 316946 252928 327542
rect 254452 319916 254504 319922
rect 254452 319858 254504 319864
rect 252900 316918 253388 316946
rect 249220 316782 249464 316810
rect 250140 316782 250384 316810
rect 250968 316782 251304 316810
rect 251796 316782 252132 316810
rect 252808 316782 253052 316810
rect 253360 316674 253388 316918
rect 254464 316810 254492 319858
rect 254832 317950 254860 327542
rect 256304 326858 256332 329838
rect 255464 326852 255516 326858
rect 255464 326794 255516 326800
rect 256292 326852 256344 326858
rect 256292 326794 256344 326800
rect 256936 326852 256988 326858
rect 256936 326794 256988 326800
rect 254912 326308 254964 326314
rect 254912 326250 254964 326256
rect 254924 320194 254952 326250
rect 254912 320188 254964 320194
rect 254912 320130 254964 320136
rect 255476 320126 255504 326794
rect 256948 320670 256976 326794
rect 257316 326722 257344 329838
rect 258420 327266 258448 329838
rect 258408 327260 258460 327266
rect 258408 327202 258460 327208
rect 258960 327192 259012 327198
rect 258960 327134 259012 327140
rect 257304 326716 257356 326722
rect 257304 326658 257356 326664
rect 258224 326648 258276 326654
rect 258224 326590 258276 326596
rect 256936 320664 256988 320670
rect 256936 320606 256988 320612
rect 258236 320618 258264 326590
rect 258236 320590 258356 320618
rect 257120 320392 257172 320398
rect 257120 320334 257172 320340
rect 256292 320256 256344 320262
rect 256292 320198 256344 320204
rect 255464 320120 255516 320126
rect 255464 320062 255516 320068
rect 255556 319984 255608 319990
rect 255556 319926 255608 319932
rect 254820 317944 254872 317950
rect 254820 317886 254872 317892
rect 255568 316810 255596 319926
rect 256304 316810 256332 320198
rect 257132 316810 257160 320334
rect 258328 317082 258356 320590
rect 258328 317054 258402 317082
rect 254464 316782 254800 316810
rect 255568 316782 255720 316810
rect 256304 316782 256640 316810
rect 257132 316782 257468 316810
rect 258374 316796 258402 317054
rect 253360 316646 253972 316674
rect 258972 313122 259000 327134
rect 259248 326314 259276 329838
rect 260168 326790 260196 329838
rect 261180 327334 261208 329838
rect 261168 327328 261220 327334
rect 261168 327270 261220 327276
rect 262100 326858 262128 329838
rect 263112 327062 263140 329838
rect 264032 327130 264060 329838
rect 264020 327124 264072 327130
rect 264020 327066 264072 327072
rect 263100 327056 263152 327062
rect 263100 326998 263152 327004
rect 262088 326852 262140 326858
rect 262088 326794 262140 326800
rect 260156 326784 260208 326790
rect 260156 326726 260208 326732
rect 259236 326308 259288 326314
rect 259236 326250 259288 326256
rect 258960 313116 259012 313122
rect 258960 313058 259012 313064
rect 240650 310160 240706 310169
rect 240650 310095 240706 310104
rect 240664 309722 240692 310095
rect 240652 309716 240704 309722
rect 240652 309658 240704 309664
rect 240926 296832 240982 296841
rect 240926 296767 240982 296776
rect 240940 295918 240968 296767
rect 240928 295912 240980 295918
rect 240928 295854 240980 295860
rect 240928 283536 240980 283542
rect 240926 283504 240928 283513
rect 240980 283504 240982 283513
rect 240926 283439 240982 283448
rect 236236 282856 236288 282862
rect 236236 282798 236288 282804
rect 236248 282114 236276 282798
rect 236236 282108 236288 282114
rect 236236 282050 236288 282056
rect 236880 282108 236932 282114
rect 236880 282050 236932 282056
rect 234120 275172 234172 275178
rect 234120 275114 234172 275120
rect 232738 274392 232794 274401
rect 232738 274327 232794 274336
rect 234132 273886 234160 275114
rect 234120 273880 234172 273886
rect 234120 273822 234172 273828
rect 234764 273880 234816 273886
rect 234764 273822 234816 273828
rect 231634 273440 231690 273449
rect 231634 273375 231690 273384
rect 233474 263104 233530 263113
rect 233474 263039 233530 263048
rect 233488 262938 233516 263039
rect 233476 262932 233528 262938
rect 233476 262874 233528 262880
rect 233474 261744 233530 261753
rect 233474 261679 233530 261688
rect 233488 261442 233516 261679
rect 233476 261436 233528 261442
rect 233476 261378 233528 261384
rect 233474 260384 233530 260393
rect 233474 260319 233530 260328
rect 233488 260082 233516 260319
rect 233476 260076 233528 260082
rect 233476 260018 233528 260024
rect 233474 258888 233530 258897
rect 233474 258823 233530 258832
rect 233488 258654 233516 258823
rect 233476 258648 233528 258654
rect 233476 258590 233528 258596
rect 233474 257528 233530 257537
rect 233474 257463 233530 257472
rect 233488 257294 233516 257463
rect 233476 257288 233528 257294
rect 233476 257230 233528 257236
rect 233474 256168 233530 256177
rect 233474 256103 233530 256112
rect 233488 256002 233516 256103
rect 233476 255996 233528 256002
rect 233476 255938 233528 255944
rect 233568 255928 233620 255934
rect 233568 255870 233620 255876
rect 232738 254672 232794 254681
rect 232738 254607 232794 254616
rect 231452 253140 231504 253146
rect 231452 253082 231504 253088
rect 231464 243150 231492 253082
rect 232752 244782 232780 254607
rect 232830 251952 232886 251961
rect 232830 251887 232886 251896
rect 232740 244776 232792 244782
rect 232740 244718 232792 244724
rect 232844 243422 232872 251887
rect 233476 251032 233528 251038
rect 233474 251000 233476 251009
rect 233528 251000 233530 251009
rect 233474 250935 233530 250944
rect 233476 250284 233528 250290
rect 233476 250226 233528 250232
rect 233488 249785 233516 250226
rect 233474 249776 233530 249785
rect 233474 249711 233530 249720
rect 233580 248425 233608 255870
rect 234120 254636 234172 254642
rect 234120 254578 234172 254584
rect 234132 253026 234160 254578
rect 234304 254568 234356 254574
rect 234304 254510 234356 254516
rect 234210 253312 234266 253321
rect 234210 253247 234266 253256
rect 234224 253146 234252 253247
rect 234212 253140 234264 253146
rect 234212 253082 234264 253088
rect 234132 252998 234252 253026
rect 234120 251780 234172 251786
rect 234120 251722 234172 251728
rect 233566 248416 233622 248425
rect 233566 248351 233622 248360
rect 233568 244708 233620 244714
rect 233568 244650 233620 244656
rect 233580 244209 233608 244650
rect 233566 244200 233622 244209
rect 233566 244135 233622 244144
rect 232832 243416 232884 243422
rect 232832 243358 232884 243364
rect 231452 243144 231504 243150
rect 231452 243086 231504 243092
rect 234132 242849 234160 251722
rect 234224 245569 234252 252998
rect 234316 246929 234344 254510
rect 234302 246920 234358 246929
rect 234302 246855 234358 246864
rect 234210 245560 234266 245569
rect 234210 245495 234266 245504
rect 234118 242840 234174 242849
rect 234118 242775 234174 242784
rect 233474 240664 233530 240673
rect 233474 240599 233476 240608
rect 233528 240599 233530 240608
rect 233476 240570 233528 240576
rect 233474 239304 233530 239313
rect 233474 239239 233476 239248
rect 233528 239239 233530 239248
rect 233476 239210 233528 239216
rect 233568 239200 233620 239206
rect 233568 239142 233620 239148
rect 233580 238633 233608 239142
rect 233566 238624 233622 238633
rect 233566 238559 233622 238568
rect 233476 237228 233528 237234
rect 233476 237170 233528 237176
rect 233488 237137 233516 237170
rect 233474 237128 233530 237137
rect 233474 237063 233530 237072
rect 232004 235868 232056 235874
rect 232004 235810 232056 235816
rect 232016 235194 232044 235810
rect 232004 235188 232056 235194
rect 232004 235130 232056 235136
rect 231818 234952 231874 234961
rect 231818 234887 231874 234896
rect 231832 234446 231860 234887
rect 231820 234440 231872 234446
rect 231820 234382 231872 234388
rect 234776 233766 234804 273822
rect 236892 266406 236920 282050
rect 243208 276934 243544 276962
rect 243760 276934 244096 276962
rect 244404 276934 244464 276962
rect 245048 276934 245384 276962
rect 245600 276934 245752 276962
rect 246244 276934 246580 276962
rect 246888 276934 247132 276962
rect 247440 276934 247776 276962
rect 248084 276934 248512 276962
rect 248728 276934 249064 276962
rect 243044 274764 243096 274770
rect 243044 274706 243096 274712
rect 240284 274696 240336 274702
rect 240284 274638 240336 274644
rect 238904 274560 238956 274566
rect 238904 274502 238956 274508
rect 237524 274492 237576 274498
rect 237524 274434 237576 274440
rect 236880 266400 236932 266406
rect 236880 266342 236932 266348
rect 237536 263770 237564 274434
rect 238916 263770 238944 274502
rect 240296 263770 240324 274638
rect 241664 274628 241716 274634
rect 241664 274570 241716 274576
rect 241676 263770 241704 274570
rect 243056 263770 243084 274706
rect 243516 273886 243544 276934
rect 244068 274838 244096 276934
rect 244056 274832 244108 274838
rect 244056 274774 244108 274780
rect 243504 273880 243556 273886
rect 243504 273822 243556 273828
rect 244436 266610 244464 276934
rect 245356 274362 245384 276934
rect 245344 274356 245396 274362
rect 245344 274298 245396 274304
rect 245724 266814 245752 276934
rect 245804 274356 245856 274362
rect 245804 274298 245856 274304
rect 245712 266808 245764 266814
rect 245712 266750 245764 266756
rect 245816 266678 245844 274298
rect 246552 273954 246580 276934
rect 246540 273948 246592 273954
rect 246540 273890 246592 273896
rect 246264 266740 246316 266746
rect 246264 266682 246316 266688
rect 245804 266672 245856 266678
rect 245804 266614 245856 266620
rect 244424 266604 244476 266610
rect 244424 266546 244476 266552
rect 244884 266196 244936 266202
rect 244884 266138 244936 266144
rect 244896 263770 244924 266138
rect 246276 263770 246304 266682
rect 247104 266338 247132 276934
rect 247748 274498 247776 276934
rect 247920 274900 247972 274906
rect 247920 274842 247972 274848
rect 247932 274673 247960 274842
rect 247918 274664 247974 274673
rect 247918 274599 247974 274608
rect 247736 274492 247788 274498
rect 247736 274434 247788 274440
rect 247184 273948 247236 273954
rect 247184 273890 247236 273896
rect 247196 266474 247224 273890
rect 247276 273744 247328 273750
rect 247274 273712 247276 273721
rect 247328 273712 247330 273721
rect 247274 273647 247330 273656
rect 247644 266536 247696 266542
rect 247644 266478 247696 266484
rect 247184 266468 247236 266474
rect 247184 266410 247236 266416
rect 247092 266332 247144 266338
rect 247092 266274 247144 266280
rect 247656 263770 247684 266478
rect 248484 266134 248512 276934
rect 248564 274492 248616 274498
rect 248564 274434 248616 274440
rect 248576 266270 248604 274434
rect 249036 274090 249064 276934
rect 249128 276934 249280 276962
rect 249588 276934 249924 276962
rect 250568 276934 250904 276962
rect 249128 275178 249156 276934
rect 249116 275172 249168 275178
rect 249116 275114 249168 275120
rect 249588 274906 249616 276934
rect 249576 274900 249628 274906
rect 249576 274842 249628 274848
rect 250876 274401 250904 276934
rect 250968 276934 251212 276962
rect 251764 276934 252100 276962
rect 250862 274392 250918 274401
rect 250862 274327 250918 274336
rect 249024 274084 249076 274090
rect 249024 274026 249076 274032
rect 249944 274084 249996 274090
rect 249944 274026 249996 274032
rect 248564 266264 248616 266270
rect 248564 266206 248616 266212
rect 248472 266128 248524 266134
rect 248472 266070 248524 266076
rect 249024 265652 249076 265658
rect 249024 265594 249076 265600
rect 249036 263770 249064 265594
rect 237536 263742 237596 263770
rect 238916 263742 238976 263770
rect 240296 263742 240356 263770
rect 241676 263742 241736 263770
rect 243056 263742 243116 263770
rect 244588 263742 244924 263770
rect 245968 263742 246304 263770
rect 247348 263742 247684 263770
rect 248728 263742 249064 263770
rect 249956 263550 249984 274026
rect 250680 274016 250732 274022
rect 250680 273958 250732 273964
rect 250036 266400 250088 266406
rect 250036 266342 250088 266348
rect 250048 263770 250076 266342
rect 250692 266202 250720 273958
rect 250772 273880 250824 273886
rect 250968 273857 250996 276934
rect 252072 274537 252100 276934
rect 252164 276934 252408 276962
rect 253052 276934 253388 276962
rect 252058 274528 252114 274537
rect 252058 274463 252114 274472
rect 250772 273822 250824 273828
rect 250954 273848 251010 273857
rect 250784 266338 250812 273822
rect 250954 273783 251010 273792
rect 252164 273750 252192 276934
rect 253360 274673 253388 276934
rect 253452 276934 253604 276962
rect 254248 276934 254308 276962
rect 253346 274664 253402 274673
rect 253346 274599 253402 274608
rect 253452 274362 253480 276934
rect 254280 274566 254308 276934
rect 254556 276934 254892 276962
rect 255108 276934 255444 276962
rect 255752 276934 256088 276962
rect 256396 276934 256732 276962
rect 256948 276934 257284 276962
rect 257592 276934 257928 276962
rect 258328 276934 258572 276962
rect 254452 274832 254504 274838
rect 254452 274774 254504 274780
rect 254268 274560 254320 274566
rect 254268 274502 254320 274508
rect 253440 274356 253492 274362
rect 253440 274298 253492 274304
rect 253440 273948 253492 273954
rect 253440 273890 253492 273896
rect 252152 273744 252204 273750
rect 252152 273686 252204 273692
rect 253452 266542 253480 273890
rect 253440 266536 253492 266542
rect 253440 266478 253492 266484
rect 250772 266332 250824 266338
rect 250772 266274 250824 266280
rect 252796 266332 252848 266338
rect 252796 266274 252848 266280
rect 250680 266196 250732 266202
rect 250680 266138 250732 266144
rect 251876 265788 251928 265794
rect 251876 265730 251928 265736
rect 251888 263770 251916 265730
rect 250048 263742 250108 263770
rect 251580 263742 251916 263770
rect 252808 263770 252836 266274
rect 254464 263770 254492 274774
rect 254556 274702 254584 276934
rect 254544 274696 254596 274702
rect 254544 274638 254596 274644
rect 255108 274634 255136 276934
rect 255752 274770 255780 276934
rect 255740 274764 255792 274770
rect 255740 274706 255792 274712
rect 255096 274628 255148 274634
rect 255096 274570 255148 274576
rect 256200 274628 256252 274634
rect 256200 274570 256252 274576
rect 254820 274220 254872 274226
rect 254820 274162 254872 274168
rect 254832 265658 254860 274162
rect 256212 266746 256240 274570
rect 256396 274022 256424 276934
rect 256948 274634 256976 276934
rect 256936 274628 256988 274634
rect 256936 274570 256988 274576
rect 256384 274016 256436 274022
rect 256384 273958 256436 273964
rect 257592 273954 257620 276934
rect 258328 274226 258356 276934
rect 258316 274220 258368 274226
rect 258316 274162 258368 274168
rect 257580 273948 257632 273954
rect 257580 273890 257632 273896
rect 256200 266740 256252 266746
rect 256200 266682 256252 266688
rect 256936 266672 256988 266678
rect 256936 266614 256988 266620
rect 255556 266604 255608 266610
rect 255556 266546 255608 266552
rect 254820 265652 254872 265658
rect 254820 265594 254872 265600
rect 252808 263742 252960 263770
rect 254340 263742 254492 263770
rect 255568 263770 255596 266546
rect 256948 263770 256976 266614
rect 258316 266468 258368 266474
rect 258316 266410 258368 266416
rect 258328 263770 258356 266410
rect 258972 265794 259000 313058
rect 261718 306216 261774 306225
rect 261718 306151 261774 306160
rect 261732 297210 261760 306151
rect 261720 297204 261772 297210
rect 261720 297146 261772 297152
rect 261718 286632 261774 286641
rect 261718 286567 261720 286576
rect 261772 286567 261774 286576
rect 261720 286538 261772 286544
rect 261442 274664 261498 274673
rect 261442 274599 261498 274608
rect 261456 272225 261484 274599
rect 261442 272216 261498 272225
rect 261442 272151 261498 272160
rect 264480 268984 264532 268990
rect 264480 268926 264532 268932
rect 259696 266536 259748 266542
rect 259696 266478 259748 266484
rect 258960 265788 259012 265794
rect 258960 265730 259012 265736
rect 259708 263770 259736 266478
rect 262456 266332 262508 266338
rect 262456 266274 262508 266280
rect 261076 266264 261128 266270
rect 261076 266206 261128 266212
rect 261088 263770 261116 266206
rect 262468 263770 262496 266274
rect 263836 266196 263888 266202
rect 263836 266138 263888 266144
rect 263848 263770 263876 266138
rect 255568 263742 255720 263770
rect 256948 263742 257100 263770
rect 258328 263742 258572 263770
rect 259708 263742 259952 263770
rect 261088 263742 261332 263770
rect 262468 263742 262712 263770
rect 263848 263742 264092 263770
rect 249944 263544 249996 263550
rect 249944 263486 249996 263492
rect 262548 236208 262600 236214
rect 243778 236176 243834 236185
rect 247274 236176 247330 236185
rect 243834 236134 244128 236162
rect 246980 236134 247274 236162
rect 243778 236111 243834 236120
rect 262548 236150 262600 236156
rect 247274 236111 247330 236120
rect 244988 235998 245048 236026
rect 246000 235998 246060 236026
rect 242490 235904 242546 235913
rect 236248 235862 237412 235890
rect 238332 235862 238668 235890
rect 239252 235862 239588 235890
rect 234764 233760 234816 233766
rect 234764 233702 234816 233708
rect 234776 233358 234804 233702
rect 231452 233352 231504 233358
rect 231452 233294 231504 233300
rect 234764 233352 234816 233358
rect 234764 233294 234816 233300
rect 231360 226212 231412 226218
rect 231360 226154 231412 226160
rect 230990 223256 231046 223265
rect 230990 223191 231046 223200
rect 230806 220128 230862 220137
rect 230806 220063 230862 220072
rect 230714 217000 230770 217009
rect 230714 216935 230770 216944
rect 231360 215876 231412 215882
rect 231360 215818 231412 215824
rect 230898 200680 230954 200689
rect 230898 200615 230954 200624
rect 230714 198232 230770 198241
rect 230714 198167 230770 198176
rect 228692 159300 228744 159306
rect 228692 159242 228744 159248
rect 228704 149446 228732 159242
rect 228692 149440 228744 149446
rect 228692 149382 228744 149388
rect 230728 104129 230756 198167
rect 230808 194524 230860 194530
rect 230808 194466 230860 194472
rect 230820 194433 230848 194466
rect 230806 194424 230862 194433
rect 230806 194359 230862 194368
rect 230714 104120 230770 104129
rect 230714 104055 230770 104064
rect 230728 95425 230756 104055
rect 230820 101681 230848 194359
rect 230912 107393 230940 200615
rect 231372 185729 231400 215818
rect 231464 207761 231492 233294
rect 231728 233284 231780 233290
rect 231728 233226 231780 233232
rect 231636 233216 231688 233222
rect 231636 233158 231688 233164
rect 231542 217000 231598 217009
rect 231542 216935 231598 216944
rect 231450 207752 231506 207761
rect 231450 207687 231506 207696
rect 231452 202072 231504 202078
rect 231452 202014 231504 202020
rect 231358 185720 231414 185729
rect 231358 185655 231414 185664
rect 231464 182601 231492 202014
rect 231556 191985 231584 216935
rect 231648 210753 231676 233158
rect 231740 213881 231768 233226
rect 231726 213872 231782 213881
rect 231726 213807 231782 213816
rect 231634 210744 231690 210753
rect 231634 210679 231690 210688
rect 232004 204792 232056 204798
rect 232004 204734 232056 204740
rect 232016 204497 232044 204734
rect 232002 204488 232058 204497
rect 232002 204423 232058 204432
rect 235314 194560 235370 194569
rect 235314 194495 235316 194504
rect 235368 194495 235370 194504
rect 235316 194466 235368 194472
rect 231542 191976 231598 191985
rect 231542 191911 231598 191920
rect 232002 188848 232058 188857
rect 236248 188818 236276 235862
rect 238640 233154 238668 235862
rect 238628 233148 238680 233154
rect 238628 233090 238680 233096
rect 239560 232474 239588 235862
rect 239652 235862 240264 235890
rect 241184 235862 241520 235890
rect 239548 232468 239600 232474
rect 239548 232410 239600 232416
rect 239652 231726 239680 235862
rect 241492 233766 241520 235862
rect 242136 235862 242490 235890
rect 241480 233760 241532 233766
rect 241480 233702 241532 233708
rect 241492 233601 241520 233702
rect 241478 233592 241534 233601
rect 241478 233527 241534 233536
rect 242136 233222 242164 235862
rect 242490 235839 242546 235848
rect 243056 235862 243116 235890
rect 243056 233465 243084 235862
rect 244988 235194 245016 235998
rect 244976 235188 245028 235194
rect 244976 235130 245028 235136
rect 246000 234281 246028 235998
rect 247992 235862 248328 235890
rect 248912 235862 249248 235890
rect 245986 234272 246042 234281
rect 245986 234207 246042 234216
rect 246264 233692 246316 233698
rect 246264 233634 246316 233640
rect 244424 233624 244476 233630
rect 244424 233566 244476 233572
rect 243042 233456 243098 233465
rect 243042 233391 243098 233400
rect 243056 233290 243084 233391
rect 243044 233284 243096 233290
rect 243044 233226 243096 233232
rect 242124 233216 242176 233222
rect 242124 233158 242176 233164
rect 244332 233216 244384 233222
rect 244332 233158 244384 233164
rect 240284 232468 240336 232474
rect 240284 232410 240336 232416
rect 239640 231720 239692 231726
rect 239640 231662 239692 231668
rect 239652 204798 239680 231662
rect 240296 226286 240324 232410
rect 240284 226280 240336 226286
rect 240284 226222 240336 226228
rect 243596 224172 243648 224178
rect 243596 224114 243648 224120
rect 243608 222834 243636 224114
rect 244344 222834 244372 233158
rect 244436 224178 244464 233566
rect 245344 233284 245396 233290
rect 245344 233226 245396 233232
rect 244424 224172 244476 224178
rect 244424 224114 244476 224120
rect 245356 222834 245384 233226
rect 246276 222834 246304 233634
rect 248012 233556 248064 233562
rect 248012 233498 248064 233504
rect 247092 232944 247144 232950
rect 247092 232886 247144 232892
rect 247104 222834 247132 232886
rect 248024 222834 248052 233498
rect 248300 232542 248328 235862
rect 248932 233760 248984 233766
rect 248932 233702 248984 233708
rect 248288 232536 248340 232542
rect 248288 232478 248340 232484
rect 248944 222834 248972 233702
rect 249220 225402 249248 235862
rect 249910 235618 249938 235876
rect 250844 235862 251272 235890
rect 251856 235862 252192 235890
rect 249910 235590 249984 235618
rect 249852 233352 249904 233358
rect 249852 233294 249904 233300
rect 249208 225396 249260 225402
rect 249208 225338 249260 225344
rect 249864 222834 249892 233294
rect 249956 232474 249984 235590
rect 250680 233488 250732 233494
rect 250680 233430 250732 233436
rect 250128 232536 250180 232542
rect 250128 232478 250180 232484
rect 249944 232468 249996 232474
rect 249944 232410 249996 232416
rect 243300 222806 243636 222834
rect 244128 222806 244372 222834
rect 245048 222806 245384 222834
rect 245968 222806 246304 222834
rect 246796 222806 247132 222834
rect 247716 222806 248052 222834
rect 248636 222806 248972 222834
rect 249464 222806 249892 222834
rect 250140 222750 250168 232478
rect 250692 222834 250720 233430
rect 251244 225470 251272 235862
rect 252164 229634 252192 235862
rect 252624 235862 252776 235890
rect 253788 235862 254124 235890
rect 254708 235862 255044 235890
rect 255720 235862 256056 235890
rect 252164 229606 252284 229634
rect 251232 225464 251284 225470
rect 251232 225406 251284 225412
rect 252256 225402 252284 229606
rect 252152 225396 252204 225402
rect 252152 225338 252204 225344
rect 252244 225396 252296 225402
rect 252244 225338 252296 225344
rect 252164 222834 252192 225338
rect 252624 225198 252652 235862
rect 252888 232468 252940 232474
rect 252888 232410 252940 232416
rect 252612 225192 252664 225198
rect 252612 225134 252664 225140
rect 250384 222806 250720 222834
rect 252132 222806 252192 222834
rect 250128 222744 250180 222750
rect 250128 222686 250180 222692
rect 250956 222744 251008 222750
rect 252900 222698 252928 232410
rect 253992 225464 254044 225470
rect 253992 225406 254044 225412
rect 254004 222834 254032 225406
rect 254096 225266 254124 235862
rect 255016 225470 255044 235862
rect 255004 225464 255056 225470
rect 255004 225406 255056 225412
rect 256028 225402 256056 235862
rect 256304 235862 256640 235890
rect 257316 235862 257652 235890
rect 258420 235862 258572 235890
rect 259248 235862 259584 235890
rect 260168 235862 260504 235890
rect 261180 235862 261516 235890
rect 262100 235862 262436 235890
rect 256304 233630 256332 235862
rect 256292 233624 256344 233630
rect 256292 233566 256344 233572
rect 257316 233222 257344 235862
rect 258420 233290 258448 235862
rect 259248 233698 259276 235862
rect 259236 233692 259288 233698
rect 259236 233634 259288 233640
rect 258408 233284 258460 233290
rect 258408 233226 258460 233232
rect 257304 233216 257356 233222
rect 257304 233158 257356 233164
rect 258960 233148 259012 233154
rect 258960 233090 259012 233096
rect 257488 225464 257540 225470
rect 257488 225406 257540 225412
rect 254820 225396 254872 225402
rect 254820 225338 254872 225344
rect 256016 225396 256068 225402
rect 256016 225338 256068 225344
rect 254084 225260 254136 225266
rect 254084 225202 254136 225208
rect 254832 222834 254860 225338
rect 256660 225260 256712 225266
rect 256660 225202 256712 225208
rect 255740 225192 255792 225198
rect 255740 225134 255792 225140
rect 255752 222834 255780 225134
rect 256672 222834 256700 225202
rect 257500 222834 257528 225406
rect 258408 225396 258460 225402
rect 258408 225338 258460 225344
rect 258420 222834 258448 225338
rect 253972 222806 254032 222834
rect 254800 222806 254860 222834
rect 255720 222806 255780 222834
rect 256640 222806 256700 222834
rect 257468 222806 257528 222834
rect 258388 222806 258448 222834
rect 251008 222692 251304 222698
rect 250956 222686 251304 222692
rect 250968 222670 251304 222686
rect 252900 222670 253052 222698
rect 258972 219282 259000 233090
rect 260168 232950 260196 235862
rect 261180 233562 261208 235862
rect 262100 233766 262128 235862
rect 262560 235777 262588 236150
rect 263112 235862 263448 235890
rect 264032 235862 264368 235890
rect 262546 235768 262602 235777
rect 262546 235703 262602 235712
rect 262560 235194 262588 235703
rect 262548 235188 262600 235194
rect 262548 235130 262600 235136
rect 262088 233760 262140 233766
rect 262088 233702 262140 233708
rect 261168 233556 261220 233562
rect 261168 233498 261220 233504
rect 263112 233358 263140 235862
rect 264032 233494 264060 235862
rect 264020 233488 264072 233494
rect 264020 233430 264072 233436
rect 263100 233352 263152 233358
rect 263100 233294 263152 233300
rect 260156 232944 260208 232950
rect 260156 232886 260208 232892
rect 258960 219276 259012 219282
rect 258960 219218 259012 219224
rect 240926 216184 240982 216193
rect 240926 216119 240982 216128
rect 240940 215882 240968 216119
rect 240928 215876 240980 215882
rect 240928 215818 240980 215824
rect 239640 204792 239692 204798
rect 239640 204734 239692 204740
rect 240650 202856 240706 202865
rect 240650 202791 240706 202800
rect 240664 202078 240692 202791
rect 240652 202072 240704 202078
rect 240652 202014 240704 202020
rect 240926 189528 240982 189537
rect 240926 189463 240982 189472
rect 232002 188783 232004 188792
rect 232056 188783 232058 188792
rect 236236 188812 236288 188818
rect 232004 188754 232056 188760
rect 236236 188754 236288 188760
rect 236248 188342 236276 188754
rect 236236 188336 236288 188342
rect 236236 188278 236288 188284
rect 236880 188336 236932 188342
rect 236880 188278 236932 188284
rect 232740 188268 232792 188274
rect 232740 188210 232792 188216
rect 231450 182592 231506 182601
rect 231450 182527 231506 182536
rect 232752 179774 232780 188210
rect 230992 179768 231044 179774
rect 230992 179710 231044 179716
rect 232740 179768 232792 179774
rect 232740 179710 232792 179716
rect 231004 179473 231032 179710
rect 230990 179464 231046 179473
rect 230990 179399 231046 179408
rect 236892 172566 236920 188278
rect 240940 188274 240968 189463
rect 240928 188268 240980 188274
rect 240928 188210 240980 188216
rect 248930 183136 248986 183145
rect 248986 183094 249280 183122
rect 248930 183071 248986 183080
rect 246244 182958 246764 182986
rect 243208 182822 243544 182850
rect 243760 182822 244096 182850
rect 244404 182822 244464 182850
rect 245048 182822 245384 182850
rect 243516 181066 243544 182822
rect 243504 181060 243556 181066
rect 243504 181002 243556 181008
rect 244068 180998 244096 182822
rect 244056 180992 244108 180998
rect 244056 180934 244108 180940
rect 241664 180924 241716 180930
rect 241664 180866 241716 180872
rect 240284 180788 240336 180794
rect 240284 180730 240336 180736
rect 237524 180720 237576 180726
rect 237524 180662 237576 180668
rect 236880 172560 236932 172566
rect 236880 172502 236932 172508
rect 237536 169794 237564 180662
rect 238904 180652 238956 180658
rect 238904 180594 238956 180600
rect 238916 169794 238944 180594
rect 240296 169794 240324 180730
rect 241676 169794 241704 180866
rect 243044 180856 243096 180862
rect 243044 180798 243096 180804
rect 243056 169794 243084 180798
rect 244436 172770 244464 182822
rect 245356 181338 245384 182822
rect 245540 182822 245600 182850
rect 245344 181332 245396 181338
rect 245344 181274 245396 181280
rect 244884 172900 244936 172906
rect 244884 172842 244936 172848
rect 244424 172764 244476 172770
rect 244424 172706 244476 172712
rect 244896 169794 244924 172842
rect 245540 172702 245568 182822
rect 246736 181354 246764 182958
rect 246888 182822 246948 182850
rect 247440 182822 247776 182850
rect 248084 182822 248604 182850
rect 248728 182822 249064 182850
rect 245804 181332 245856 181338
rect 246736 181326 246856 181354
rect 245804 181274 245856 181280
rect 245528 172696 245580 172702
rect 245528 172638 245580 172644
rect 245816 172294 245844 181274
rect 246264 172968 246316 172974
rect 246264 172910 246316 172916
rect 245804 172288 245856 172294
rect 245804 172230 245856 172236
rect 246276 169794 246304 172910
rect 246828 172634 246856 181326
rect 246816 172628 246868 172634
rect 246816 172570 246868 172576
rect 246920 172498 246948 182822
rect 247748 181338 247776 182822
rect 247736 181332 247788 181338
rect 247736 181274 247788 181280
rect 248380 181332 248432 181338
rect 248380 181274 248432 181280
rect 246908 172492 246960 172498
rect 246908 172434 246960 172440
rect 248392 172430 248420 181274
rect 248472 181128 248524 181134
rect 248472 181070 248524 181076
rect 248380 172424 248432 172430
rect 248380 172366 248432 172372
rect 248484 171954 248512 181070
rect 248576 172362 248604 182822
rect 249036 182193 249064 182822
rect 249588 182822 249924 182850
rect 250232 182822 250568 182850
rect 250876 182822 251212 182850
rect 251764 182822 252100 182850
rect 252408 182822 252744 182850
rect 253052 182822 253388 182850
rect 249022 182184 249078 182193
rect 249022 182119 249078 182128
rect 249588 180017 249616 182822
rect 250232 180153 250260 182822
rect 250876 180289 250904 182822
rect 252072 180561 252100 182822
rect 252716 180697 252744 182822
rect 252796 181060 252848 181066
rect 252796 181002 252848 181008
rect 252702 180688 252758 180697
rect 252702 180623 252758 180632
rect 252058 180552 252114 180561
rect 252058 180487 252114 180496
rect 250862 180280 250918 180289
rect 250862 180215 250918 180224
rect 250218 180144 250274 180153
rect 250218 180079 250274 180088
rect 249574 180008 249630 180017
rect 249574 179943 249630 179952
rect 250036 172560 250088 172566
rect 250036 172502 250088 172508
rect 248564 172356 248616 172362
rect 248564 172298 248616 172304
rect 249024 172220 249076 172226
rect 249024 172162 249076 172168
rect 247644 171948 247696 171954
rect 247644 171890 247696 171896
rect 248472 171948 248524 171954
rect 248472 171890 248524 171896
rect 247656 169794 247684 171890
rect 249036 169794 249064 172162
rect 237536 169766 237596 169794
rect 238916 169766 238976 169794
rect 240296 169766 240356 169794
rect 241676 169766 241736 169794
rect 243056 169766 243116 169794
rect 244588 169766 244924 169794
rect 245968 169766 246304 169794
rect 247348 169766 247684 169794
rect 248728 169766 249064 169794
rect 250048 169794 250076 172502
rect 251876 171812 251928 171818
rect 251876 171754 251928 171760
rect 251888 169794 251916 171754
rect 250048 169766 250108 169794
rect 251580 169766 251916 169794
rect 252808 169794 252836 181002
rect 253360 180833 253388 182822
rect 253544 182822 253604 182850
rect 254188 182822 254248 182850
rect 254556 182822 254892 182850
rect 255108 182822 255444 182850
rect 255752 182822 256088 182850
rect 256732 182822 256792 182850
rect 253440 180992 253492 180998
rect 253440 180934 253492 180940
rect 253346 180824 253402 180833
rect 253346 180759 253402 180768
rect 253452 173042 253480 180934
rect 253544 180726 253572 182822
rect 253532 180720 253584 180726
rect 253532 180662 253584 180668
rect 254188 180658 254216 182822
rect 254556 180794 254584 182822
rect 255108 180930 255136 182822
rect 255096 180924 255148 180930
rect 255096 180866 255148 180872
rect 255752 180862 255780 182822
rect 255740 180856 255792 180862
rect 255740 180798 255792 180804
rect 254544 180788 254596 180794
rect 254544 180730 254596 180736
rect 254176 180652 254228 180658
rect 254176 180594 254228 180600
rect 254820 180584 254872 180590
rect 254820 180526 254872 180532
rect 253440 173036 253492 173042
rect 253440 172978 253492 172984
rect 254176 173036 254228 173042
rect 254176 172978 254228 172984
rect 254188 169794 254216 172978
rect 254832 172974 254860 180526
rect 254820 172968 254872 172974
rect 254820 172910 254872 172916
rect 256764 172906 256792 182822
rect 256948 182822 257284 182850
rect 257592 182822 257928 182850
rect 258572 182822 258724 182850
rect 256948 180590 256976 182822
rect 257592 181134 257620 182822
rect 257580 181128 257632 181134
rect 257580 181070 257632 181076
rect 256936 180584 256988 180590
rect 256936 180526 256988 180532
rect 258696 172974 258724 182822
rect 258684 172968 258736 172974
rect 258684 172910 258736 172916
rect 256752 172900 256804 172906
rect 256752 172842 256804 172848
rect 255556 172764 255608 172770
rect 255556 172706 255608 172712
rect 255568 169794 255596 172706
rect 258316 172696 258368 172702
rect 258316 172638 258368 172644
rect 256936 172288 256988 172294
rect 256936 172230 256988 172236
rect 256948 169794 256976 172230
rect 258328 169794 258356 172638
rect 258972 171818 259000 219218
rect 262362 212784 262418 212793
rect 262362 212719 262418 212728
rect 262376 211802 262404 212719
rect 262364 211796 262416 211802
rect 262364 211738 262416 211744
rect 263098 192792 263154 192801
rect 263098 192727 263154 192736
rect 263112 186846 263140 192727
rect 263100 186840 263152 186846
rect 263100 186782 263152 186788
rect 261076 182080 261128 182086
rect 261074 182048 261076 182057
rect 261128 182048 261130 182057
rect 261074 181983 261130 181992
rect 264492 175694 264520 268926
rect 265872 232338 265900 371742
rect 278076 370910 278412 370938
rect 277544 368332 277596 368338
rect 277544 368274 277596 368280
rect 266596 357928 266648 357934
rect 266596 357870 266648 357876
rect 266608 357225 266636 357870
rect 266594 357216 266650 357225
rect 266594 357151 266650 357160
rect 266596 356568 266648 356574
rect 266596 356510 266648 356516
rect 266608 356137 266636 356510
rect 266594 356128 266650 356137
rect 266594 356063 266650 356072
rect 266596 355208 266648 355214
rect 266594 355176 266596 355185
rect 266648 355176 266650 355185
rect 266594 355111 266650 355120
rect 266688 355140 266740 355146
rect 266688 355082 266740 355088
rect 266700 354097 266728 355082
rect 266686 354088 266742 354097
rect 266686 354023 266742 354032
rect 266596 353848 266648 353854
rect 266596 353790 266648 353796
rect 266608 353009 266636 353790
rect 266594 353000 266650 353009
rect 266594 352935 266650 352944
rect 266596 352420 266648 352426
rect 266596 352362 266648 352368
rect 266608 352057 266636 352362
rect 266594 352048 266650 352057
rect 266594 351983 266650 351992
rect 274874 351368 274930 351377
rect 274874 351303 274930 351312
rect 274888 351134 274916 351303
rect 272024 351128 272076 351134
rect 272024 351070 272076 351076
rect 274876 351128 274928 351134
rect 274876 351070 274928 351076
rect 266688 351060 266740 351066
rect 266688 351002 266740 351008
rect 266594 350960 266650 350969
rect 266594 350895 266650 350904
rect 266608 350386 266636 350895
rect 266596 350380 266648 350386
rect 266596 350322 266648 350328
rect 266700 349881 266728 351002
rect 266686 349872 266742 349881
rect 266686 349807 266742 349816
rect 271932 349768 271984 349774
rect 271932 349710 271984 349716
rect 266596 349700 266648 349706
rect 266596 349642 266648 349648
rect 266608 348929 266636 349642
rect 266594 348920 266650 348929
rect 266594 348855 266650 348864
rect 271944 348278 271972 349710
rect 272036 349706 272064 351070
rect 277556 351066 277584 368274
rect 278384 367658 278412 370910
rect 280408 370910 280560 370938
rect 280408 368338 280436 370910
rect 283030 370666 283058 370924
rect 284548 370910 285528 370938
rect 288012 370910 288624 370938
rect 283030 370638 283104 370666
rect 280396 368332 280448 368338
rect 280396 368274 280448 368280
rect 278372 367652 278424 367658
rect 278372 367594 278424 367600
rect 280488 367652 280540 367658
rect 280488 367594 280540 367600
rect 280500 351762 280528 367594
rect 283076 355078 283104 370638
rect 284548 356545 284576 370910
rect 284534 356536 284590 356545
rect 284534 356471 284590 356480
rect 288596 355078 288624 370910
rect 290068 370910 290496 370938
rect 293072 370910 293408 370938
rect 283064 355072 283116 355078
rect 283064 355014 283116 355020
rect 285364 355072 285416 355078
rect 285364 355014 285416 355020
rect 288584 355072 288636 355078
rect 288584 355014 288636 355020
rect 280422 351734 280528 351762
rect 285376 351748 285404 355014
rect 290068 352426 290096 370910
rect 293380 367658 293408 370910
rect 294208 370910 295556 370938
rect 298040 370910 298284 370938
rect 293368 367652 293420 367658
rect 293368 367594 293420 367600
rect 290332 355072 290384 355078
rect 290332 355014 290384 355020
rect 290056 352420 290108 352426
rect 290056 352362 290108 352368
rect 290344 351748 290372 355014
rect 294208 353854 294236 370910
rect 298256 367658 298284 370910
rect 299820 370910 300524 370938
rect 303008 370910 303344 370938
rect 294288 367652 294340 367658
rect 294288 367594 294340 367600
rect 298244 367652 298296 367658
rect 298244 367594 298296 367600
rect 299716 367652 299768 367658
rect 299716 367594 299768 367600
rect 294196 353848 294248 353854
rect 294196 353790 294248 353796
rect 294300 351898 294328 367594
rect 294300 351870 294972 351898
rect 284534 351640 284590 351649
rect 294944 351626 294972 351870
rect 299728 351626 299756 367594
rect 299820 355146 299848 370910
rect 303316 367658 303344 370910
rect 305340 370910 305584 370938
rect 308068 370910 308404 370938
rect 303304 367652 303356 367658
rect 303304 367594 303356 367600
rect 305236 367652 305288 367658
rect 305236 367594 305288 367600
rect 299808 355140 299860 355146
rect 299808 355082 299860 355088
rect 305248 351762 305276 367594
rect 305340 355214 305368 370910
rect 308376 367658 308404 370910
rect 309388 370910 310552 370938
rect 313036 370910 313464 370938
rect 308364 367652 308416 367658
rect 308364 367594 308416 367600
rect 309284 367652 309336 367658
rect 309284 367594 309336 367600
rect 305328 355208 305380 355214
rect 305328 355150 305380 355156
rect 309296 355078 309324 367594
rect 309388 356574 309416 370910
rect 309376 356568 309428 356574
rect 309376 356510 309428 356516
rect 313436 355078 313464 370910
rect 314908 370910 315520 370938
rect 314908 357934 314936 370910
rect 314896 357928 314948 357934
rect 314896 357870 314948 357876
rect 309284 355072 309336 355078
rect 309284 355014 309336 355020
rect 310388 355072 310440 355078
rect 310388 355014 310440 355020
rect 313424 355072 313476 355078
rect 313424 355014 313476 355020
rect 315356 355072 315408 355078
rect 315356 355014 315408 355020
rect 305248 351734 305354 351762
rect 310400 351748 310428 355014
rect 315368 351748 315396 355014
rect 294944 351598 295418 351626
rect 299728 351598 300386 351626
rect 284534 351575 284536 351584
rect 284588 351575 284590 351584
rect 284536 351546 284588 351552
rect 277544 351060 277596 351066
rect 277544 351002 277596 351008
rect 274874 350416 274930 350425
rect 274874 350351 274930 350360
rect 274888 349774 274916 350351
rect 274876 349768 274928 349774
rect 274876 349710 274928 349716
rect 272024 349700 272076 349706
rect 272024 349642 272076 349648
rect 274874 349600 274930 349609
rect 274874 349535 274930 349544
rect 266596 348272 266648 348278
rect 266596 348214 266648 348220
rect 271932 348272 271984 348278
rect 271932 348214 271984 348220
rect 266608 347841 266636 348214
rect 266594 347832 266650 347841
rect 266594 347767 266650 347776
rect 274888 346918 274916 349535
rect 274966 348648 275022 348657
rect 274966 348583 275022 348592
rect 266596 346912 266648 346918
rect 266594 346880 266596 346889
rect 274876 346912 274928 346918
rect 266648 346880 266650 346889
rect 274876 346854 274928 346860
rect 274980 346850 275008 348583
rect 275058 347832 275114 347841
rect 275058 347767 275114 347776
rect 266594 346815 266650 346824
rect 266688 346844 266740 346850
rect 266688 346786 266740 346792
rect 274968 346844 275020 346850
rect 274968 346786 275020 346792
rect 266700 345801 266728 346786
rect 266686 345792 266742 345801
rect 266686 345727 266742 345736
rect 275072 345558 275100 347767
rect 275150 346880 275206 346889
rect 275150 346815 275206 346824
rect 266596 345552 266648 345558
rect 266596 345494 266648 345500
rect 275060 345552 275112 345558
rect 275060 345494 275112 345500
rect 266608 344713 266636 345494
rect 275164 345370 275192 346815
rect 275242 346064 275298 346073
rect 275242 345999 275298 346008
rect 274980 345342 275192 345370
rect 274874 345112 274930 345121
rect 274874 345047 274930 345056
rect 266594 344704 266650 344713
rect 266594 344639 266650 344648
rect 266596 344124 266648 344130
rect 266596 344066 266648 344072
rect 266608 343761 266636 344066
rect 266594 343752 266650 343761
rect 266594 343687 266650 343696
rect 274888 342770 274916 345047
rect 274980 344130 275008 345342
rect 275058 344296 275114 344305
rect 275058 344231 275114 344240
rect 274968 344124 275020 344130
rect 274968 344066 275020 344072
rect 274966 343344 275022 343353
rect 274966 343279 275022 343288
rect 266688 342764 266740 342770
rect 266688 342706 266740 342712
rect 274876 342764 274928 342770
rect 274876 342706 274928 342712
rect 266596 342696 266648 342702
rect 266594 342664 266596 342673
rect 266648 342664 266650 342673
rect 266594 342599 266650 342608
rect 266700 341585 266728 342706
rect 266686 341576 266742 341585
rect 266686 341511 266742 341520
rect 274874 341576 274930 341585
rect 274874 341511 274930 341520
rect 266596 341404 266648 341410
rect 266596 341346 266648 341352
rect 266608 340633 266636 341346
rect 266594 340624 266650 340633
rect 266594 340559 266650 340568
rect 272024 340112 272076 340118
rect 272024 340054 272076 340060
rect 266596 340044 266648 340050
rect 266596 339986 266648 339992
rect 266608 339545 266636 339986
rect 266594 339536 266650 339545
rect 266594 339471 266650 339480
rect 266688 338616 266740 338622
rect 266594 338584 266650 338593
rect 266688 338558 266740 338564
rect 266594 338519 266596 338528
rect 266648 338519 266650 338528
rect 266596 338490 266648 338496
rect 266700 337505 266728 338558
rect 266686 337496 266742 337505
rect 266686 337431 266742 337440
rect 271472 337324 271524 337330
rect 271472 337266 271524 337272
rect 266596 337256 266648 337262
rect 266596 337198 266648 337204
rect 266608 336417 266636 337198
rect 266594 336408 266650 336417
rect 266594 336343 266650 336352
rect 266596 335896 266648 335902
rect 266596 335838 266648 335844
rect 266608 335465 266636 335838
rect 266594 335456 266650 335465
rect 266594 335391 266650 335400
rect 266596 334468 266648 334474
rect 266596 334410 266648 334416
rect 266608 334377 266636 334410
rect 271484 334406 271512 337266
rect 272036 337262 272064 340054
rect 274888 338622 274916 341511
rect 274980 340050 275008 343279
rect 275072 341410 275100 344231
rect 275256 342702 275284 345999
rect 275244 342696 275296 342702
rect 275244 342638 275296 342644
rect 275150 342392 275206 342401
rect 275150 342327 275206 342336
rect 275060 341404 275112 341410
rect 275060 341346 275112 341352
rect 275058 340624 275114 340633
rect 275058 340559 275114 340568
rect 275072 340118 275100 340559
rect 275060 340112 275112 340118
rect 275060 340054 275112 340060
rect 274968 340044 275020 340050
rect 274968 339986 275020 339992
rect 275058 339808 275114 339817
rect 275058 339743 275114 339752
rect 274876 338616 274928 338622
rect 274876 338558 274928 338564
rect 274874 338040 274930 338049
rect 274874 337975 274930 337984
rect 274888 337330 274916 337975
rect 274876 337324 274928 337330
rect 274876 337266 274928 337272
rect 272024 337256 272076 337262
rect 272024 337198 272076 337204
rect 274874 337088 274930 337097
rect 274874 337023 274930 337032
rect 266688 334400 266740 334406
rect 266594 334368 266650 334377
rect 266688 334342 266740 334348
rect 271472 334400 271524 334406
rect 271472 334342 271524 334348
rect 266594 334303 266650 334312
rect 266700 333289 266728 334342
rect 266686 333280 266742 333289
rect 266686 333215 266742 333224
rect 274888 333114 274916 337023
rect 274966 336272 275022 336281
rect 274966 336207 275022 336216
rect 266596 333108 266648 333114
rect 266596 333050 266648 333056
rect 274876 333108 274928 333114
rect 274876 333050 274928 333056
rect 266608 332337 266636 333050
rect 266594 332328 266650 332337
rect 266594 332263 266650 332272
rect 274980 331754 275008 336207
rect 275072 335902 275100 339743
rect 275164 338554 275192 342327
rect 275610 338856 275666 338865
rect 275610 338791 275666 338800
rect 275152 338548 275204 338554
rect 275152 338490 275204 338496
rect 275060 335896 275112 335902
rect 275060 335838 275112 335844
rect 275624 334474 275652 338791
rect 275612 334468 275664 334474
rect 275612 334410 275664 334416
rect 279580 333794 279608 335836
rect 281788 335822 282906 335850
rect 285928 335822 286218 335850
rect 288688 335822 289530 335850
rect 280304 333856 280356 333862
rect 280304 333798 280356 333804
rect 279568 333788 279620 333794
rect 279568 333730 279620 333736
rect 266596 331748 266648 331754
rect 266596 331690 266648 331696
rect 274968 331748 275020 331754
rect 274968 331690 275020 331696
rect 266608 331249 266636 331690
rect 266594 331240 266650 331249
rect 266594 331175 266650 331184
rect 266594 330288 266650 330297
rect 266594 330223 266650 330232
rect 266608 329102 266636 330223
rect 266596 329096 266648 329102
rect 266596 329038 266648 329044
rect 268620 326988 268672 326994
rect 268620 326930 268672 326936
rect 266596 286596 266648 286602
rect 266596 286538 266648 286544
rect 266608 280686 266636 286538
rect 266596 280680 266648 280686
rect 266596 280622 266648 280628
rect 267240 263612 267292 263618
rect 267240 263554 267292 263560
rect 267148 257288 267200 257294
rect 267148 257230 267200 257236
rect 266594 256168 266650 256177
rect 266594 256103 266650 256112
rect 266608 255934 266636 256103
rect 266596 255928 266648 255934
rect 266596 255870 266648 255876
rect 266594 254672 266650 254681
rect 266594 254607 266650 254616
rect 266608 254506 266636 254607
rect 266596 254500 266648 254506
rect 266596 254442 266648 254448
rect 266594 253312 266650 253321
rect 266594 253247 266650 253256
rect 266608 253214 266636 253247
rect 266596 253208 266648 253214
rect 266596 253150 266648 253156
rect 266594 251952 266650 251961
rect 266594 251887 266650 251896
rect 266608 251786 266636 251887
rect 266596 251780 266648 251786
rect 266596 251722 266648 251728
rect 267160 249105 267188 257230
rect 267146 249096 267202 249105
rect 267146 249031 267202 249040
rect 266596 248788 266648 248794
rect 266596 248730 266648 248736
rect 266608 247745 266636 248730
rect 266594 247736 266650 247745
rect 266594 247671 266650 247680
rect 266596 247564 266648 247570
rect 266596 247506 266648 247512
rect 266608 246385 266636 247506
rect 266594 246376 266650 246385
rect 266594 246311 266650 246320
rect 266596 246136 266648 246142
rect 266596 246078 266648 246084
rect 266608 244889 266636 246078
rect 266594 244880 266650 244889
rect 266594 244815 266650 244824
rect 267252 236593 267280 263554
rect 267514 263104 267570 263113
rect 267514 263039 267570 263048
rect 267422 261744 267478 261753
rect 267422 261679 267478 261688
rect 267330 258888 267386 258897
rect 267330 258823 267386 258832
rect 267344 252210 267372 258823
rect 267436 253078 267464 261679
rect 267424 253072 267476 253078
rect 267424 253014 267476 253020
rect 267344 252182 267464 252210
rect 267330 250592 267386 250601
rect 267330 250527 267386 250536
rect 267344 237234 267372 250527
rect 267436 248674 267464 252182
rect 267528 250290 267556 263039
rect 267606 260384 267662 260393
rect 267606 260319 267662 260328
rect 267516 250284 267568 250290
rect 267516 250226 267568 250232
rect 267620 248930 267648 260319
rect 267790 257528 267846 257537
rect 267790 257463 267846 257472
rect 267700 253072 267752 253078
rect 267700 253014 267752 253020
rect 267608 248924 267660 248930
rect 267608 248866 267660 248872
rect 267712 248862 267740 253014
rect 267700 248856 267752 248862
rect 267700 248798 267752 248804
rect 267436 248646 267740 248674
rect 267712 247502 267740 248646
rect 267700 247496 267752 247502
rect 267700 247438 267752 247444
rect 267804 246210 267832 257463
rect 267884 253140 267936 253146
rect 267884 253082 267936 253088
rect 267792 246204 267844 246210
rect 267792 246146 267844 246152
rect 267896 243529 267924 253082
rect 267882 243520 267938 243529
rect 267882 243455 267938 243464
rect 267884 243280 267936 243286
rect 267884 243222 267936 243228
rect 267896 242169 267924 243222
rect 267882 242160 267938 242169
rect 267882 242095 267938 242104
rect 267882 240664 267938 240673
rect 267882 240599 267884 240608
rect 267936 240599 267938 240608
rect 267884 240570 267936 240576
rect 267882 239304 267938 239313
rect 267882 239239 267884 239248
rect 267936 239239 267938 239248
rect 267884 239210 267936 239216
rect 267516 239200 267568 239206
rect 267516 239142 267568 239148
rect 267528 237953 267556 239142
rect 267514 237944 267570 237953
rect 267514 237879 267570 237888
rect 267332 237228 267384 237234
rect 267332 237170 267384 237176
rect 267238 236584 267294 236593
rect 267238 236519 267294 236528
rect 268632 233766 268660 326930
rect 280316 323526 280344 333798
rect 281788 327402 281816 335822
rect 285928 327470 285956 335822
rect 288688 327538 288716 335822
rect 292724 333924 292776 333930
rect 292724 333866 292776 333872
rect 288676 327532 288728 327538
rect 288676 327474 288728 327480
rect 289964 327532 290016 327538
rect 289964 327474 290016 327480
rect 285916 327464 285968 327470
rect 285916 327406 285968 327412
rect 281776 327396 281828 327402
rect 281776 327338 281828 327344
rect 282236 327396 282288 327402
rect 282236 327338 282288 327344
rect 282248 326994 282276 327338
rect 285928 327062 285956 327406
rect 289976 327130 290004 327474
rect 289964 327124 290016 327130
rect 289964 327066 290016 327072
rect 285916 327056 285968 327062
rect 285916 326998 285968 327004
rect 282236 326988 282288 326994
rect 282236 326930 282288 326936
rect 292736 323526 292764 333866
rect 292920 331657 292948 335836
rect 296232 333153 296260 335836
rect 296218 333144 296274 333153
rect 296218 333079 296274 333088
rect 299544 331754 299572 335836
rect 302870 335822 303160 335850
rect 299532 331748 299584 331754
rect 299532 331690 299584 331696
rect 292906 331648 292962 331657
rect 292906 331583 292962 331592
rect 292920 330841 292948 331583
rect 299544 331521 299572 331690
rect 299530 331512 299586 331521
rect 299530 331447 299586 331456
rect 292906 330832 292962 330841
rect 292906 330767 292962 330776
rect 303132 328966 303160 335822
rect 305144 333992 305196 333998
rect 305144 333934 305196 333940
rect 302476 328960 302528 328966
rect 302476 328902 302528 328908
rect 303120 328960 303172 328966
rect 303120 328902 303172 328908
rect 302488 327606 302516 328902
rect 302476 327600 302528 327606
rect 302476 327542 302528 327548
rect 305156 323526 305184 333934
rect 306260 330394 306288 335836
rect 309572 333862 309600 335836
rect 312884 333930 312912 335836
rect 316196 333998 316224 335836
rect 316184 333992 316236 333998
rect 316184 333934 316236 333940
rect 312872 333924 312924 333930
rect 312872 333866 312924 333872
rect 309560 333856 309612 333862
rect 309560 333798 309612 333804
rect 319048 330394 319076 384759
rect 319126 382104 319182 382113
rect 319126 382039 319182 382048
rect 305236 330388 305288 330394
rect 305236 330330 305288 330336
rect 306248 330388 306300 330394
rect 306248 330330 306300 330336
rect 319036 330388 319088 330394
rect 319036 330330 319088 330336
rect 305248 329034 305276 330330
rect 316552 329096 316604 329102
rect 316552 329038 316604 329044
rect 305236 329028 305288 329034
rect 305236 328970 305288 328976
rect 279108 323520 279160 323526
rect 279108 323462 279160 323468
rect 280304 323520 280356 323526
rect 280304 323462 280356 323468
rect 291528 323520 291580 323526
rect 291528 323462 291580 323468
rect 292724 323520 292776 323526
rect 292724 323462 292776 323468
rect 304040 323520 304092 323526
rect 304040 323462 304092 323468
rect 305144 323520 305196 323526
rect 305144 323462 305196 323468
rect 279120 321692 279148 323462
rect 291540 321692 291568 323462
rect 304052 321692 304080 323462
rect 316564 321692 316592 329038
rect 319140 328966 319168 382039
rect 319218 380200 319274 380209
rect 319218 380135 319274 380144
rect 319232 331754 319260 380135
rect 319310 377480 319366 377489
rect 319310 377415 319366 377424
rect 319324 333153 319352 377415
rect 319402 374760 319458 374769
rect 319402 374695 319458 374704
rect 319310 333144 319366 333153
rect 319310 333079 319366 333088
rect 319324 331822 319352 333079
rect 319312 331816 319364 331822
rect 319312 331758 319364 331764
rect 319220 331748 319272 331754
rect 319220 331690 319272 331696
rect 319232 330462 319260 331690
rect 319416 331657 319444 374695
rect 320138 371904 320194 371913
rect 320138 371839 320194 371848
rect 320152 371806 320180 371839
rect 320140 371800 320192 371806
rect 320140 371742 320192 371748
rect 320598 351368 320654 351377
rect 320598 351303 320654 351312
rect 320612 351134 320640 351303
rect 320600 351128 320652 351134
rect 320600 351070 320652 351076
rect 321610 350416 321666 350425
rect 321610 350351 321666 350360
rect 321624 349774 321652 350351
rect 321612 349768 321664 349774
rect 321612 349710 321664 349716
rect 321702 349600 321758 349609
rect 321702 349535 321758 349544
rect 321610 348648 321666 348657
rect 321610 348583 321666 348592
rect 321624 348346 321652 348583
rect 321716 348482 321744 349535
rect 321704 348476 321756 348482
rect 321704 348418 321756 348424
rect 321612 348340 321664 348346
rect 321612 348282 321664 348288
rect 321058 347832 321114 347841
rect 321058 347767 321114 347776
rect 321072 346986 321100 347767
rect 321060 346980 321112 346986
rect 321060 346922 321112 346928
rect 320414 346880 320470 346889
rect 320414 346815 320470 346824
rect 320428 345694 320456 346815
rect 320506 346064 320562 346073
rect 320506 345999 320562 346008
rect 320416 345688 320468 345694
rect 320416 345630 320468 345636
rect 320520 345626 320548 345999
rect 320508 345620 320560 345626
rect 320508 345562 320560 345568
rect 321058 345112 321114 345121
rect 321058 345047 321114 345056
rect 321072 344674 321100 345047
rect 321060 344668 321112 344674
rect 321060 344610 321112 344616
rect 321612 344396 321664 344402
rect 321612 344338 321664 344344
rect 321624 344305 321652 344338
rect 321610 344296 321666 344305
rect 321610 344231 321666 344240
rect 321610 343344 321666 343353
rect 321610 343279 321666 343288
rect 321624 342906 321652 343279
rect 321612 342900 321664 342906
rect 321612 342842 321664 342848
rect 321058 342392 321114 342401
rect 321058 342327 321114 342336
rect 321072 341478 321100 342327
rect 321610 341576 321666 341585
rect 321610 341511 321612 341520
rect 321664 341511 321666 341520
rect 321612 341482 321664 341488
rect 321060 341472 321112 341478
rect 321060 341414 321112 341420
rect 320598 340624 320654 340633
rect 320598 340559 320654 340568
rect 320612 340118 320640 340559
rect 320600 340112 320652 340118
rect 320600 340054 320652 340060
rect 321242 339808 321298 339817
rect 321242 339743 321298 339752
rect 321256 338690 321284 339743
rect 321610 338856 321666 338865
rect 321610 338791 321612 338800
rect 321664 338791 321666 338800
rect 321612 338762 321664 338768
rect 321244 338684 321296 338690
rect 321244 338626 321296 338632
rect 321610 338040 321666 338049
rect 321610 337975 321666 337984
rect 321624 337330 321652 337975
rect 321612 337324 321664 337330
rect 321612 337266 321664 337272
rect 321426 337088 321482 337097
rect 321426 337023 321482 337032
rect 321440 336106 321468 337023
rect 321610 336272 321666 336281
rect 321610 336207 321666 336216
rect 321428 336100 321480 336106
rect 321428 336042 321480 336048
rect 321624 335970 321652 336207
rect 321612 335964 321664 335970
rect 321612 335906 321664 335912
rect 319402 331648 319458 331657
rect 319402 331583 319458 331592
rect 319416 330530 319444 331583
rect 319404 330524 319456 330530
rect 319404 330466 319456 330472
rect 319220 330456 319272 330462
rect 319220 330398 319272 330404
rect 319128 328960 319180 328966
rect 319128 328902 319180 328908
rect 270274 313560 270330 313569
rect 270274 313495 270330 313504
rect 270288 313122 270316 313495
rect 270276 313116 270328 313122
rect 270276 313058 270328 313064
rect 269356 297204 269408 297210
rect 269356 297146 269408 297152
rect 269368 296841 269396 297146
rect 269354 296832 269410 296841
rect 269354 296767 269410 296776
rect 270276 280680 270328 280686
rect 270276 280622 270328 280628
rect 270288 280249 270316 280622
rect 270274 280240 270330 280249
rect 270274 280175 270330 280184
rect 276452 269670 276480 271916
rect 276440 269664 276492 269670
rect 276440 269606 276492 269612
rect 276452 269505 276480 269606
rect 283536 269534 283564 271916
rect 290712 269670 290740 271916
rect 290700 269664 290752 269670
rect 290700 269606 290752 269612
rect 283524 269528 283576 269534
rect 276438 269496 276494 269505
rect 283524 269470 283576 269476
rect 276438 269431 276494 269440
rect 284536 269052 284588 269058
rect 284536 268994 284588 269000
rect 284548 257772 284576 268994
rect 290712 268990 290740 269606
rect 297796 269058 297824 271916
rect 297784 269052 297836 269058
rect 297784 268994 297836 269000
rect 290700 268984 290752 268990
rect 290700 268926 290752 268932
rect 304972 268310 305000 271916
rect 303764 268304 303816 268310
rect 303764 268246 303816 268252
rect 304960 268304 305012 268310
rect 304960 268246 305012 268252
rect 303776 261306 303804 268246
rect 312056 264094 312084 271916
rect 310756 264088 310808 264094
rect 310756 264030 310808 264036
rect 312044 264088 312096 264094
rect 312044 264030 312096 264036
rect 310768 263618 310796 264030
rect 310756 263612 310808 263618
rect 310756 263554 310808 263560
rect 297876 261300 297928 261306
rect 297876 261242 297928 261248
rect 303764 261300 303816 261306
rect 303764 261242 303816 261248
rect 297888 257772 297916 261242
rect 319232 260694 319260 271916
rect 311216 260688 311268 260694
rect 311216 260630 311268 260636
rect 319220 260688 319272 260694
rect 319220 260630 319272 260636
rect 311228 257772 311256 260630
rect 321244 258444 321296 258450
rect 321244 258386 321296 258392
rect 321256 257401 321284 258386
rect 274874 257392 274930 257401
rect 274874 257327 274930 257336
rect 321242 257392 321298 257401
rect 321242 257327 321298 257336
rect 274888 257294 274916 257327
rect 274876 257288 274928 257294
rect 274876 257230 274928 257236
rect 321060 257220 321112 257226
rect 321060 257162 321112 257168
rect 321072 256449 321100 257162
rect 275058 256440 275114 256449
rect 275058 256375 275114 256384
rect 321058 256440 321114 256449
rect 321058 256375 321114 256384
rect 274414 254672 274470 254681
rect 274414 254607 274470 254616
rect 272760 254500 272812 254506
rect 272760 254442 272812 254448
rect 272772 244782 272800 254442
rect 274232 253208 274284 253214
rect 274232 253150 274284 253156
rect 272852 251780 272904 251786
rect 272852 251722 272904 251728
rect 272760 244776 272812 244782
rect 272760 244718 272812 244724
rect 272864 243422 272892 251722
rect 274138 250320 274194 250329
rect 274138 250255 274194 250264
rect 272852 243416 272904 243422
rect 272852 243358 272904 243364
rect 274152 239206 274180 250255
rect 274244 243121 274272 253150
rect 274322 252904 274378 252913
rect 274322 252839 274378 252848
rect 274336 243286 274364 252839
rect 274428 246142 274456 254607
rect 274874 253856 274930 253865
rect 274874 253791 274930 253800
rect 274888 253146 274916 253791
rect 274876 253140 274928 253146
rect 274876 253082 274928 253088
rect 274876 250284 274928 250290
rect 274876 250226 274928 250232
rect 274888 250057 274916 250226
rect 274874 250048 274930 250057
rect 274874 249983 274930 249992
rect 274968 248924 275020 248930
rect 274968 248866 275020 248872
rect 274876 248856 274928 248862
rect 274874 248824 274876 248833
rect 274928 248824 274930 248833
rect 274874 248759 274930 248768
rect 274980 248289 275008 248866
rect 275072 248794 275100 256375
rect 275704 255928 275756 255934
rect 275704 255870 275756 255876
rect 275610 252088 275666 252097
rect 275610 252023 275666 252032
rect 275518 251136 275574 251145
rect 275518 251071 275574 251080
rect 275060 248788 275112 248794
rect 275060 248730 275112 248736
rect 274966 248280 275022 248289
rect 274966 248215 275022 248224
rect 274876 247496 274928 247502
rect 274876 247438 274928 247444
rect 274888 247337 274916 247438
rect 274874 247328 274930 247337
rect 274874 247263 274930 247272
rect 274876 246204 274928 246210
rect 274876 246146 274928 246152
rect 274416 246136 274468 246142
rect 274888 246113 274916 246146
rect 274416 246078 274468 246084
rect 274874 246104 274930 246113
rect 274874 246039 274930 246048
rect 274876 244776 274928 244782
rect 274874 244744 274876 244753
rect 274928 244744 274930 244753
rect 274874 244679 274930 244688
rect 274324 243280 274376 243286
rect 274324 243222 274376 243228
rect 274230 243112 274286 243121
rect 274230 243047 274286 243056
rect 275532 239274 275560 251071
rect 275624 240634 275652 252023
rect 275716 245569 275744 255870
rect 320692 255860 320744 255866
rect 320692 255802 320744 255808
rect 275886 255624 275942 255633
rect 275886 255559 275942 255568
rect 275900 247570 275928 255559
rect 320704 254681 320732 255802
rect 320876 255656 320928 255662
rect 320874 255624 320876 255633
rect 320928 255624 320930 255633
rect 320874 255559 320930 255568
rect 320690 254672 320746 254681
rect 320690 254607 320746 254616
rect 321610 253856 321666 253865
rect 321610 253791 321666 253800
rect 321624 253690 321652 253791
rect 321612 253684 321664 253690
rect 321612 253626 321664 253632
rect 321612 253072 321664 253078
rect 321612 253014 321664 253020
rect 321624 252913 321652 253014
rect 321610 252904 321666 252913
rect 321610 252839 321666 252848
rect 321610 252088 321666 252097
rect 321610 252023 321612 252032
rect 321664 252023 321666 252032
rect 321612 251994 321664 252000
rect 320598 251136 320654 251145
rect 320598 251071 320654 251080
rect 320612 250630 320640 251071
rect 320600 250624 320652 250630
rect 320600 250566 320652 250572
rect 321058 250320 321114 250329
rect 321058 250255 321114 250264
rect 321072 249542 321100 250255
rect 321060 249536 321112 249542
rect 321060 249478 321112 249484
rect 321610 249368 321666 249377
rect 321610 249303 321666 249312
rect 321624 249134 321652 249303
rect 321612 249128 321664 249134
rect 321612 249070 321664 249076
rect 321610 248416 321666 248425
rect 321610 248351 321666 248360
rect 321624 247706 321652 248351
rect 321612 247700 321664 247706
rect 321612 247642 321664 247648
rect 321794 247600 321850 247609
rect 275888 247564 275940 247570
rect 321794 247535 321796 247544
rect 275888 247506 275940 247512
rect 321848 247535 321850 247544
rect 321796 247506 321848 247512
rect 321808 247475 321836 247506
rect 321242 246648 321298 246657
rect 321242 246583 321298 246592
rect 321256 246278 321284 246583
rect 321244 246272 321296 246278
rect 321244 246214 321296 246220
rect 321610 245832 321666 245841
rect 321610 245767 321666 245776
rect 275702 245560 275758 245569
rect 275702 245495 275758 245504
rect 321624 244850 321652 245767
rect 321704 244912 321756 244918
rect 321702 244880 321704 244889
rect 321756 244880 321758 244889
rect 321612 244844 321664 244850
rect 321702 244815 321758 244824
rect 321612 244786 321664 244792
rect 321610 244064 321666 244073
rect 321610 243999 321666 244008
rect 321624 243490 321652 243999
rect 321612 243484 321664 243490
rect 321612 243426 321664 243432
rect 275796 243416 275848 243422
rect 275796 243358 275848 243364
rect 275808 242985 275836 243358
rect 321610 243112 321666 243121
rect 321610 243047 321666 243056
rect 275794 242976 275850 242985
rect 275794 242911 275850 242920
rect 320506 242296 320562 242305
rect 321624 242266 321652 243047
rect 320506 242231 320562 242240
rect 321612 242260 321664 242266
rect 320520 242130 320548 242231
rect 321612 242202 321664 242208
rect 320508 242124 320560 242130
rect 320508 242066 320560 242072
rect 275612 240628 275664 240634
rect 275612 240570 275664 240576
rect 279672 239342 279700 241860
rect 283260 239449 283288 241860
rect 283246 239440 283302 239449
rect 283246 239375 283302 239384
rect 279660 239336 279712 239342
rect 279660 239278 279712 239284
rect 280304 239336 280356 239342
rect 280304 239278 280356 239284
rect 275520 239268 275572 239274
rect 275520 239210 275572 239216
rect 274140 239200 274192 239206
rect 274140 239142 274192 239148
rect 268620 233760 268672 233766
rect 268620 233702 268672 233708
rect 265860 232332 265912 232338
rect 265860 232274 265912 232280
rect 279108 230292 279160 230298
rect 279108 230234 279160 230240
rect 279120 227716 279148 230234
rect 280316 227646 280344 239278
rect 286940 238594 286968 241860
rect 290528 239721 290556 241860
rect 290514 239712 290570 239721
rect 290514 239647 290570 239656
rect 294208 238662 294236 241860
rect 294196 238656 294248 238662
rect 294196 238598 294248 238604
rect 286928 238588 286980 238594
rect 286928 238530 286980 238536
rect 286940 238361 286968 238530
rect 286926 238352 286982 238361
rect 286926 238287 286982 238296
rect 297796 238066 297824 241860
rect 297704 238038 297824 238066
rect 297704 236350 297732 238038
rect 297692 236344 297744 236350
rect 297692 236286 297744 236292
rect 297704 235874 297732 236286
rect 297692 235868 297744 235874
rect 297692 235810 297744 235816
rect 301476 234961 301504 241860
rect 305064 241738 305092 241860
rect 308744 241738 308772 241860
rect 312332 241738 312360 241860
rect 316026 241846 316132 241874
rect 305064 241710 305184 241738
rect 305156 240401 305184 241710
rect 308008 241710 308772 241738
rect 312148 241710 312360 241738
rect 305142 240392 305198 240401
rect 305142 240327 305198 240336
rect 301462 234952 301518 234961
rect 301462 234887 301518 234896
rect 302014 234952 302070 234961
rect 302014 234887 302070 234896
rect 302028 234446 302056 234887
rect 302016 234440 302068 234446
rect 302016 234382 302068 234388
rect 304040 230428 304092 230434
rect 304040 230370 304092 230376
rect 291528 230360 291580 230366
rect 291528 230302 291580 230308
rect 291540 227716 291568 230302
rect 304052 227716 304080 230370
rect 305156 227714 305184 240327
rect 308008 230298 308036 241710
rect 312148 230366 312176 241710
rect 316104 239886 316132 241846
rect 314896 239880 314948 239886
rect 314896 239822 314948 239828
rect 316092 239880 316144 239886
rect 316092 239822 316144 239828
rect 314908 230434 314936 239822
rect 316276 237228 316328 237234
rect 316276 237170 316328 237176
rect 316288 236622 316316 237170
rect 316276 236616 316328 236622
rect 316276 236558 316328 236564
rect 314896 230428 314948 230434
rect 314896 230370 314948 230376
rect 312136 230360 312188 230366
rect 312136 230302 312188 230308
rect 307996 230292 308048 230298
rect 307996 230234 308048 230240
rect 316288 227730 316316 236558
rect 305144 227708 305196 227714
rect 316288 227702 316578 227730
rect 305144 227650 305196 227656
rect 280304 227640 280356 227646
rect 280304 227582 280356 227588
rect 273954 226656 274010 226665
rect 273954 226591 274010 226600
rect 272942 219584 272998 219593
rect 272942 219519 272998 219528
rect 272956 219282 272984 219519
rect 272944 219276 272996 219282
rect 272944 219218 272996 219224
rect 268620 211796 268672 211802
rect 268620 211738 268672 211744
rect 268632 207518 268660 211738
rect 268620 207512 268672 207518
rect 268620 207454 268672 207460
rect 272944 207512 272996 207518
rect 272944 207454 272996 207460
rect 272956 202865 272984 207454
rect 272942 202856 272998 202865
rect 272942 202791 272998 202800
rect 273968 188970 273996 226591
rect 273876 188942 273996 188970
rect 272944 186840 272996 186846
rect 272944 186782 272996 186788
rect 272956 186273 272984 186782
rect 272942 186264 272998 186273
rect 272942 186199 272998 186208
rect 267516 182080 267568 182086
rect 267516 182022 267568 182028
rect 267528 181241 267556 182022
rect 267514 181232 267570 181241
rect 267514 181167 267570 181176
rect 273876 178550 273904 188942
rect 273864 178544 273916 178550
rect 273864 178486 273916 178492
rect 276256 178544 276308 178550
rect 276256 178486 276308 178492
rect 276268 178226 276296 178486
rect 276268 178212 276466 178226
rect 276268 178198 276480 178212
rect 276452 175830 276480 178198
rect 276440 175824 276492 175830
rect 276440 175766 276492 175772
rect 283536 175762 283564 177940
rect 283524 175756 283576 175762
rect 283524 175698 283576 175704
rect 290712 175694 290740 177940
rect 264480 175688 264532 175694
rect 264480 175630 264532 175636
rect 290700 175688 290752 175694
rect 290700 175630 290752 175636
rect 297796 175150 297824 177940
rect 285824 175144 285876 175150
rect 285824 175086 285876 175092
rect 297784 175144 297836 175150
rect 297784 175086 297836 175092
rect 259696 172628 259748 172634
rect 259696 172570 259748 172576
rect 258960 171812 259012 171818
rect 258960 171754 259012 171760
rect 259708 169794 259736 172570
rect 261168 172492 261220 172498
rect 261168 172434 261220 172440
rect 261180 169794 261208 172434
rect 262456 172424 262508 172430
rect 262456 172366 262508 172372
rect 262468 169794 262496 172366
rect 263836 172356 263888 172362
rect 263836 172298 263888 172304
rect 263848 169794 263876 172298
rect 252808 169766 252960 169794
rect 254188 169766 254340 169794
rect 255568 169766 255720 169794
rect 256948 169766 257100 169794
rect 258328 169766 258572 169794
rect 259708 169766 259952 169794
rect 261180 169766 261332 169794
rect 262468 169766 262712 169794
rect 263848 169766 264092 169794
rect 267240 169568 267292 169574
rect 267240 169510 267292 169516
rect 233474 169128 233530 169137
rect 233474 169063 233530 169072
rect 233488 168962 233516 169063
rect 233476 168956 233528 168962
rect 233476 168898 233528 168904
rect 233474 167768 233530 167777
rect 233474 167703 233530 167712
rect 233488 167602 233516 167703
rect 233476 167596 233528 167602
rect 233476 167538 233528 167544
rect 233474 166408 233530 166417
rect 233474 166343 233530 166352
rect 233488 166242 233516 166343
rect 233476 166236 233528 166242
rect 233476 166178 233528 166184
rect 233474 164912 233530 164921
rect 233474 164847 233530 164856
rect 267146 164912 267202 164921
rect 267146 164847 267202 164856
rect 233488 164814 233516 164847
rect 233476 164808 233528 164814
rect 233476 164750 233528 164756
rect 233474 163552 233530 163561
rect 231452 163516 231504 163522
rect 233474 163487 233530 163496
rect 231452 163458 231504 163464
rect 231360 159300 231412 159306
rect 231360 159242 231412 159248
rect 231372 149174 231400 159242
rect 231464 155090 231492 163458
rect 233488 163454 233516 163487
rect 233476 163448 233528 163454
rect 233476 163390 233528 163396
rect 233474 162192 233530 162201
rect 233474 162127 233476 162136
rect 233528 162127 233530 162136
rect 267054 162192 267110 162201
rect 267054 162127 267110 162136
rect 233476 162098 233528 162104
rect 234580 162088 234632 162094
rect 234580 162030 234632 162036
rect 232738 160696 232794 160705
rect 232738 160631 232794 160640
rect 234304 160660 234356 160666
rect 231452 155084 231504 155090
rect 231452 155026 231504 155032
rect 232752 150874 232780 160631
rect 234304 160602 234356 160608
rect 233474 159336 233530 159345
rect 233474 159271 233476 159280
rect 233528 159271 233530 159280
rect 233476 159242 233528 159248
rect 234118 157976 234174 157985
rect 234118 157911 234174 157920
rect 233476 157192 233528 157198
rect 233476 157134 233528 157140
rect 233488 156625 233516 157134
rect 233474 156616 233530 156625
rect 233474 156551 233530 156560
rect 233474 155120 233530 155129
rect 233474 155055 233476 155064
rect 233528 155055 233530 155064
rect 233476 155026 233528 155032
rect 233476 150936 233528 150942
rect 233474 150904 233476 150913
rect 233528 150904 233530 150913
rect 232740 150868 232792 150874
rect 233474 150839 233530 150848
rect 232740 150810 232792 150816
rect 234132 149582 234160 157911
rect 234316 152409 234344 160602
rect 234592 153769 234620 162030
rect 266594 160696 266650 160705
rect 266594 160631 266596 160640
rect 266648 160631 266650 160640
rect 266596 160602 266648 160608
rect 266596 159368 266648 159374
rect 266594 159336 266596 159345
rect 266648 159336 266650 159345
rect 266594 159271 266650 159280
rect 266596 158008 266648 158014
rect 266594 157976 266596 157985
rect 266648 157976 266650 157985
rect 266594 157911 266650 157920
rect 266964 157940 267016 157946
rect 266964 157882 267016 157888
rect 266594 155120 266650 155129
rect 266594 155055 266650 155064
rect 266688 155084 266740 155090
rect 266608 154954 266636 155055
rect 266688 155026 266740 155032
rect 266596 154948 266648 154954
rect 266596 154890 266648 154896
rect 266700 153769 266728 155026
rect 234578 153760 234634 153769
rect 234578 153695 234634 153704
rect 266686 153760 266742 153769
rect 266686 153695 266742 153704
rect 266596 153588 266648 153594
rect 266596 153530 266648 153536
rect 266608 152409 266636 153530
rect 234302 152400 234358 152409
rect 234302 152335 234358 152344
rect 266594 152400 266650 152409
rect 266594 152335 266650 152344
rect 266596 150936 266648 150942
rect 266594 150904 266596 150913
rect 266648 150904 266650 150913
rect 266594 150839 266650 150848
rect 234120 149576 234172 149582
rect 233474 149544 233530 149553
rect 266596 149576 266648 149582
rect 234120 149518 234172 149524
rect 266594 149544 266596 149553
rect 266648 149544 266650 149553
rect 233474 149479 233530 149488
rect 266594 149479 266650 149488
rect 233488 149446 233516 149479
rect 233476 149440 233528 149446
rect 233476 149382 233528 149388
rect 231360 149168 231412 149174
rect 231360 149110 231412 149116
rect 233476 148216 233528 148222
rect 233474 148184 233476 148193
rect 266976 148193 267004 157882
rect 267068 155838 267096 162127
rect 267056 155832 267108 155838
rect 267056 155774 267108 155780
rect 267160 153730 267188 164847
rect 267148 153724 267200 153730
rect 267148 153666 267200 153672
rect 233528 148184 233530 148193
rect 233474 148119 233530 148128
rect 266962 148184 267018 148193
rect 266962 148119 267018 148128
rect 233476 146788 233528 146794
rect 233476 146730 233528 146736
rect 233488 146697 233516 146730
rect 233474 146688 233530 146697
rect 233474 146623 233530 146632
rect 233476 145428 233528 145434
rect 233476 145370 233528 145376
rect 266780 145428 266832 145434
rect 266780 145370 266832 145376
rect 233488 145337 233516 145370
rect 266792 145337 266820 145370
rect 233474 145328 233530 145337
rect 233474 145263 233530 145272
rect 266778 145328 266834 145337
rect 266778 145263 266834 145272
rect 230992 144884 231044 144890
rect 230992 144826 231044 144832
rect 231004 143161 231032 144826
rect 233476 144068 233528 144074
rect 233476 144010 233528 144016
rect 233488 143977 233516 144010
rect 233474 143968 233530 143977
rect 233474 143903 233530 143912
rect 230990 143152 231046 143161
rect 230990 143087 231046 143096
rect 231004 132961 231032 143087
rect 267252 142617 267280 169510
rect 267422 169128 267478 169137
rect 267422 169063 267478 169072
rect 267330 156616 267386 156625
rect 267330 156551 267386 156560
rect 267238 142608 267294 142617
rect 267238 142543 267294 142552
rect 242490 142200 242546 142209
rect 242196 142158 242490 142186
rect 242490 142135 242546 142144
rect 246814 142200 246870 142209
rect 246870 142158 246980 142186
rect 246814 142135 246870 142144
rect 231360 142096 231412 142102
rect 231360 142038 231412 142044
rect 233474 142064 233530 142073
rect 231268 140600 231320 140606
rect 231268 140542 231320 140548
rect 231082 140024 231138 140033
rect 231082 139959 231138 139968
rect 230990 132952 231046 132961
rect 230990 132887 231046 132896
rect 230992 132848 231044 132854
rect 230992 132790 231044 132796
rect 231004 120449 231032 132790
rect 231096 126025 231124 139959
rect 231280 130270 231308 140542
rect 231372 139761 231400 142038
rect 233474 141999 233476 142008
rect 233528 141999 233530 142008
rect 233476 141970 233528 141976
rect 236248 141886 237412 141914
rect 238332 141886 238668 141914
rect 239252 141886 239588 141914
rect 231450 140568 231506 140577
rect 231450 140503 231506 140512
rect 231358 139752 231414 139761
rect 231358 139687 231414 139696
rect 231372 138673 231400 139687
rect 231358 138664 231414 138673
rect 231358 138599 231414 138608
rect 231464 132854 231492 140503
rect 232002 138664 232058 138673
rect 232002 138599 232058 138608
rect 231452 132848 231504 132854
rect 231452 132790 231504 132796
rect 231360 131352 231412 131358
rect 231360 131294 231412 131300
rect 231268 130264 231320 130270
rect 231268 130206 231320 130212
rect 231280 129833 231308 130206
rect 231266 129824 231322 129833
rect 231266 129759 231322 129768
rect 231082 126016 231138 126025
rect 231082 125951 231138 125960
rect 230990 120440 231046 120449
rect 230990 120375 231046 120384
rect 230898 107384 230954 107393
rect 230898 107319 230954 107328
rect 230806 101672 230862 101681
rect 230806 101607 230862 101616
rect 231372 98281 231400 131294
rect 232016 122625 232044 138599
rect 236248 134418 236276 141886
rect 238640 139246 238668 141886
rect 239560 139858 239588 141886
rect 239652 141886 240264 141914
rect 241184 141886 241520 141914
rect 239548 139852 239600 139858
rect 239548 139794 239600 139800
rect 238628 139240 238680 139246
rect 238628 139182 238680 139188
rect 239652 136474 239680 141886
rect 241492 139314 241520 141886
rect 242504 139654 242532 142135
rect 243410 142064 243466 142073
rect 243056 142022 243410 142050
rect 243056 140577 243084 142022
rect 267344 142034 267372 156551
rect 267436 156450 267464 169063
rect 267606 167768 267662 167777
rect 267606 167703 267662 167712
rect 267514 166408 267570 166417
rect 267514 166343 267570 166352
rect 267424 156444 267476 156450
rect 267424 156386 267476 156392
rect 267528 153662 267556 166343
rect 267620 155022 267648 167703
rect 285836 166310 285864 175086
rect 304972 174470 305000 177940
rect 300360 174464 300412 174470
rect 300360 174406 300412 174412
rect 304960 174464 305012 174470
rect 304960 174406 305012 174412
rect 300372 166854 300400 174406
rect 312056 170254 312084 177940
rect 312044 170248 312096 170254
rect 312044 170190 312096 170196
rect 312056 169574 312084 170190
rect 312044 169568 312096 169574
rect 312044 169510 312096 169516
rect 319232 166854 319260 177940
rect 297876 166848 297928 166854
rect 297876 166790 297928 166796
rect 300360 166848 300412 166854
rect 300360 166790 300412 166796
rect 311216 166848 311268 166854
rect 311216 166790 311268 166796
rect 319220 166848 319272 166854
rect 319220 166790 319272 166796
rect 284536 166304 284588 166310
rect 284536 166246 284588 166252
rect 285824 166304 285876 166310
rect 285824 166246 285876 166252
rect 284548 163796 284576 166246
rect 297888 163796 297916 166790
rect 311228 163796 311256 166790
rect 267882 163552 267938 163561
rect 267882 163487 267938 163496
rect 321612 163516 321664 163522
rect 267700 155832 267752 155838
rect 267700 155774 267752 155780
rect 267608 155016 267660 155022
rect 267608 154958 267660 154964
rect 267516 153656 267568 153662
rect 267516 153598 267568 153604
rect 267712 150874 267740 155774
rect 267792 155152 267844 155158
rect 267792 155094 267844 155100
rect 267700 150868 267752 150874
rect 267700 150810 267752 150816
rect 267804 143977 267832 155094
rect 267896 152370 267924 163487
rect 321612 163458 321664 163464
rect 272852 163448 272904 163454
rect 274876 163448 274928 163454
rect 272852 163390 272904 163396
rect 274874 163416 274876 163425
rect 321624 163425 321652 163458
rect 274928 163416 274930 163425
rect 270000 160660 270052 160666
rect 270000 160602 270052 160608
rect 267884 152364 267936 152370
rect 267884 152306 267936 152312
rect 270012 150806 270040 160602
rect 272760 159300 272812 159306
rect 272760 159242 272812 159248
rect 271380 158008 271432 158014
rect 271380 157950 271432 157956
rect 270000 150800 270052 150806
rect 270000 150742 270052 150748
rect 271392 149514 271420 157950
rect 272772 149582 272800 159242
rect 272864 154954 272892 163390
rect 274874 163351 274930 163360
rect 321610 163416 321666 163425
rect 321610 163351 321666 163360
rect 275058 162464 275114 162473
rect 275058 162399 275114 162408
rect 321610 162464 321666 162473
rect 321610 162399 321612 162408
rect 272944 161136 272996 161142
rect 272944 161078 272996 161084
rect 272852 154948 272904 154954
rect 272852 154890 272904 154896
rect 272956 153594 272984 161078
rect 274874 158928 274930 158937
rect 274874 158863 274930 158872
rect 274888 157946 274916 158863
rect 274876 157940 274928 157946
rect 274876 157882 274928 157888
rect 274876 156444 274928 156450
rect 274876 156386 274928 156392
rect 274888 156081 274916 156386
rect 274966 156344 275022 156353
rect 274966 156279 275022 156288
rect 274874 156072 274930 156081
rect 274874 156007 274930 156016
rect 274980 155158 275008 156279
rect 274968 155152 275020 155158
rect 274968 155094 275020 155100
rect 275072 155090 275100 162399
rect 321664 162399 321666 162408
rect 321612 162370 321664 162376
rect 275150 161648 275206 161657
rect 321610 161648 321666 161657
rect 275150 161583 275206 161592
rect 321060 161612 321112 161618
rect 275164 161142 275192 161583
rect 321610 161583 321666 161592
rect 321060 161554 321112 161560
rect 275152 161136 275204 161142
rect 275152 161078 275204 161084
rect 321072 160705 321100 161554
rect 321624 161482 321652 161583
rect 321612 161476 321664 161482
rect 321612 161418 321664 161424
rect 275794 160696 275850 160705
rect 275794 160631 275850 160640
rect 321058 160696 321114 160705
rect 321058 160631 321114 160640
rect 275150 159880 275206 159889
rect 275150 159815 275206 159824
rect 275164 159306 275192 159815
rect 275704 159368 275756 159374
rect 275704 159310 275756 159316
rect 275152 159300 275204 159306
rect 275152 159242 275204 159248
rect 275518 158112 275574 158121
rect 275518 158047 275574 158056
rect 275060 155084 275112 155090
rect 275060 155026 275112 155032
rect 274876 155016 274928 155022
rect 274874 154984 274876 154993
rect 274928 154984 274930 154993
rect 274874 154919 274930 154928
rect 274968 153724 275020 153730
rect 274968 153666 275020 153672
rect 274876 153656 274928 153662
rect 274874 153624 274876 153633
rect 274928 153624 274930 153633
rect 272944 153588 272996 153594
rect 274874 153559 274930 153568
rect 272944 153530 272996 153536
rect 274980 153361 275008 153666
rect 274966 153352 275022 153361
rect 274966 153287 275022 153296
rect 274876 152364 274928 152370
rect 274876 152306 274928 152312
rect 274888 152137 274916 152306
rect 274874 152128 274930 152137
rect 274874 152063 274930 152072
rect 274874 150904 274930 150913
rect 274874 150839 274876 150848
rect 274928 150839 274930 150848
rect 274876 150810 274928 150816
rect 274968 150800 275020 150806
rect 274968 150742 275020 150748
rect 274980 150641 275008 150742
rect 274966 150632 275022 150641
rect 274966 150567 275022 150576
rect 272760 149576 272812 149582
rect 272760 149518 272812 149524
rect 271380 149508 271432 149514
rect 271380 149450 271432 149456
rect 274876 149508 274928 149514
rect 274876 149450 274928 149456
rect 274888 148873 274916 149450
rect 274874 148864 274930 148873
rect 274874 148799 274930 148808
rect 275532 146794 275560 158047
rect 275610 157160 275666 157169
rect 275610 157095 275666 157104
rect 267884 146788 267936 146794
rect 267884 146730 267936 146736
rect 275520 146788 275572 146794
rect 275520 146730 275572 146736
rect 267896 146697 267924 146730
rect 267882 146688 267938 146697
rect 267882 146623 267938 146632
rect 275624 145434 275652 157095
rect 275716 149553 275744 159310
rect 275808 150942 275836 160631
rect 320598 159880 320654 159889
rect 320598 159815 320654 159824
rect 320612 159374 320640 159815
rect 320600 159368 320652 159374
rect 320600 159310 320652 159316
rect 321058 158928 321114 158937
rect 321058 158863 321114 158872
rect 321072 158014 321100 158863
rect 321612 158212 321664 158218
rect 321612 158154 321664 158160
rect 321624 158121 321652 158154
rect 321610 158112 321666 158121
rect 321610 158047 321666 158056
rect 321060 158008 321112 158014
rect 321060 157950 321112 157956
rect 321612 157192 321664 157198
rect 321610 157160 321612 157169
rect 321664 157160 321666 157169
rect 321610 157095 321666 157104
rect 321058 156344 321114 156353
rect 321058 156279 321114 156288
rect 321072 155430 321100 156279
rect 321060 155424 321112 155430
rect 321060 155366 321112 155372
rect 321610 155392 321666 155401
rect 321610 155327 321666 155336
rect 321624 155158 321652 155327
rect 321612 155152 321664 155158
rect 321612 155094 321664 155100
rect 320874 154440 320930 154449
rect 320874 154375 320930 154384
rect 320888 153798 320916 154375
rect 320876 153792 320928 153798
rect 320876 153734 320928 153740
rect 321610 153624 321666 153633
rect 321610 153559 321666 153568
rect 320506 152672 320562 152681
rect 320506 152607 320562 152616
rect 320520 152438 320548 152607
rect 321624 152506 321652 153559
rect 321612 152500 321664 152506
rect 321612 152442 321664 152448
rect 320508 152432 320560 152438
rect 320508 152374 320560 152380
rect 320782 151856 320838 151865
rect 320782 151791 320838 151800
rect 320796 151418 320824 151791
rect 320784 151412 320836 151418
rect 320784 151354 320836 151360
rect 275796 150936 275848 150942
rect 275796 150878 275848 150884
rect 321702 150904 321758 150913
rect 321758 150862 321836 150890
rect 321702 150839 321758 150848
rect 321610 150088 321666 150097
rect 321610 150023 321666 150032
rect 321624 149650 321652 150023
rect 321612 149644 321664 149650
rect 321612 149586 321664 149592
rect 275702 149544 275758 149553
rect 275702 149479 275758 149488
rect 321058 149136 321114 149145
rect 321058 149071 321114 149080
rect 321072 148290 321100 149071
rect 321612 148420 321664 148426
rect 321612 148362 321664 148368
rect 321624 148329 321652 148362
rect 321610 148320 321666 148329
rect 321060 148284 321112 148290
rect 321610 148255 321666 148264
rect 321060 148226 321112 148232
rect 321808 148222 321836 150862
rect 321796 148216 321848 148222
rect 321796 148158 321848 148164
rect 279672 145434 279700 147884
rect 283260 147762 283288 147884
rect 286940 147762 286968 147884
rect 283168 147734 283288 147762
rect 285928 147734 286968 147762
rect 275612 145428 275664 145434
rect 275612 145370 275664 145376
rect 279660 145428 279712 145434
rect 279660 145370 279712 145376
rect 280304 144748 280356 144754
rect 280304 144690 280356 144696
rect 267790 143968 267846 143977
rect 267790 143903 267846 143912
rect 243410 141999 243466 142008
rect 267332 142028 267384 142034
rect 267332 141970 267384 141976
rect 243792 141886 244128 141914
rect 245048 141886 245384 141914
rect 246060 141886 246212 141914
rect 247992 141886 248512 141914
rect 248912 141886 249248 141914
rect 243042 140568 243098 140577
rect 243042 140503 243098 140512
rect 243792 139761 243820 141886
rect 243778 139752 243834 139761
rect 243778 139687 243834 139696
rect 244332 139716 244384 139722
rect 244332 139658 244384 139664
rect 242492 139648 242544 139654
rect 242492 139590 242544 139596
rect 241480 139308 241532 139314
rect 241480 139250 241532 139256
rect 239100 136446 239680 136474
rect 236236 134412 236288 134418
rect 236236 134354 236288 134360
rect 236236 124824 236288 124830
rect 236236 124766 236288 124772
rect 232002 122616 232058 122625
rect 232002 122551 232058 122560
rect 231452 122036 231504 122042
rect 231452 121978 231504 121984
rect 231358 98272 231414 98281
rect 231358 98207 231414 98216
rect 230714 95416 230770 95425
rect 230714 95351 230770 95360
rect 230728 94881 230756 95351
rect 230714 94872 230770 94881
rect 230714 94807 230770 94816
rect 231464 92297 231492 121978
rect 236248 115106 236276 124766
rect 236236 115100 236288 115106
rect 236236 115042 236288 115048
rect 239100 110958 239128 136446
rect 244344 130338 244372 139658
rect 245356 139625 245384 141886
rect 246184 139897 246212 141886
rect 246170 139888 246226 139897
rect 246170 139823 246226 139832
rect 246446 139888 246502 139897
rect 246446 139823 246502 139832
rect 245342 139616 245398 139625
rect 245342 139551 245398 139560
rect 244424 139376 244476 139382
rect 244424 139318 244476 139324
rect 243596 130332 243648 130338
rect 243596 130274 243648 130280
rect 244332 130332 244384 130338
rect 244332 130274 244384 130280
rect 243608 128722 243636 130274
rect 244436 128722 244464 139318
rect 245804 138900 245856 138906
rect 245804 138842 245856 138848
rect 245816 131630 245844 138842
rect 245344 131624 245396 131630
rect 245344 131566 245396 131572
rect 245804 131624 245856 131630
rect 245804 131566 245856 131572
rect 245356 128722 245384 131566
rect 246264 130604 246316 130610
rect 246264 130546 246316 130552
rect 246276 128722 246304 130546
rect 246460 130270 246488 139823
rect 247092 139784 247144 139790
rect 247092 139726 247144 139732
rect 247104 130610 247132 139726
rect 247184 138968 247236 138974
rect 247184 138910 247236 138916
rect 247092 130604 247144 130610
rect 247092 130546 247144 130552
rect 246448 130264 246500 130270
rect 246446 130232 246448 130241
rect 246500 130232 246502 130241
rect 246446 130167 246502 130176
rect 247196 128722 247224 138910
rect 248012 131624 248064 131630
rect 248012 131566 248064 131572
rect 248024 128722 248052 131566
rect 248484 131426 248512 141886
rect 249116 139648 249168 139654
rect 249116 139590 249168 139596
rect 248564 139444 248616 139450
rect 248564 139386 248616 139392
rect 248576 131630 248604 139386
rect 249128 138537 249156 139590
rect 249220 139518 249248 141886
rect 249864 141886 249924 141914
rect 250844 141886 251180 141914
rect 251856 141886 252192 141914
rect 249864 139586 249892 141886
rect 249852 139580 249904 139586
rect 249852 139522 249904 139528
rect 249208 139512 249260 139518
rect 249208 139454 249260 139460
rect 249668 139308 249720 139314
rect 249668 139250 249720 139256
rect 249852 139308 249904 139314
rect 249852 139250 249904 139256
rect 249114 138528 249170 138537
rect 249114 138463 249170 138472
rect 249128 137313 249156 138463
rect 249114 137304 249170 137313
rect 249114 137239 249170 137248
rect 249680 134321 249708 139250
rect 249666 134312 249722 134321
rect 249666 134247 249722 134256
rect 249680 133097 249708 134247
rect 249666 133088 249722 133097
rect 249666 133023 249722 133032
rect 248564 131624 248616 131630
rect 248564 131566 248616 131572
rect 248472 131420 248524 131426
rect 248472 131362 248524 131368
rect 248932 130332 248984 130338
rect 248932 130274 248984 130280
rect 248944 128722 248972 130274
rect 249864 128722 249892 139250
rect 249944 139172 249996 139178
rect 249944 139114 249996 139120
rect 249956 130338 249984 139114
rect 251152 139042 251180 141886
rect 251324 139648 251376 139654
rect 251324 139590 251376 139596
rect 251140 139036 251192 139042
rect 251140 138978 251192 138984
rect 251336 131630 251364 139590
rect 252060 139512 252112 139518
rect 252060 139454 252112 139460
rect 250680 131624 250732 131630
rect 250680 131566 250732 131572
rect 251324 131624 251376 131630
rect 251324 131566 251376 131572
rect 249944 130332 249996 130338
rect 249944 130274 249996 130280
rect 250692 128722 250720 131566
rect 250956 131420 251008 131426
rect 250956 131362 251008 131368
rect 243300 128694 243636 128722
rect 244128 128694 244464 128722
rect 245048 128694 245384 128722
rect 245968 128694 246304 128722
rect 246796 128694 247224 128722
rect 247716 128694 248052 128722
rect 248636 128694 248972 128722
rect 249464 128694 249892 128722
rect 250384 128694 250720 128722
rect 250968 128722 250996 131362
rect 252072 128994 252100 139454
rect 252164 139110 252192 141886
rect 252716 141886 252776 141914
rect 253788 141886 253940 141914
rect 254708 141886 255044 141914
rect 255720 141886 256056 141914
rect 252152 139104 252204 139110
rect 252152 139046 252204 139052
rect 252716 138634 252744 141886
rect 253072 139580 253124 139586
rect 253072 139522 253124 139528
rect 252704 138628 252756 138634
rect 252704 138570 252756 138576
rect 252072 128966 252146 128994
rect 250968 128694 251304 128722
rect 252118 128708 252146 128966
rect 253084 128722 253112 139522
rect 253912 138838 253940 141886
rect 255016 139586 255044 141886
rect 255004 139580 255056 139586
rect 255004 139522 255056 139528
rect 256028 139518 256056 141886
rect 256304 141886 256640 141914
rect 257316 141886 257652 141914
rect 258328 141886 258572 141914
rect 259248 141886 259584 141914
rect 260168 141886 260504 141914
rect 261180 141886 261516 141914
rect 262100 141886 262436 141914
rect 263112 141886 263448 141914
rect 264124 141886 264368 141914
rect 256304 139722 256332 141886
rect 256292 139716 256344 139722
rect 256292 139658 256344 139664
rect 256016 139512 256068 139518
rect 256016 139454 256068 139460
rect 257316 139382 257344 141886
rect 257488 139580 257540 139586
rect 257488 139522 257540 139528
rect 257304 139376 257356 139382
rect 257304 139318 257356 139324
rect 254176 139104 254228 139110
rect 254176 139046 254228 139052
rect 253992 139036 254044 139042
rect 253992 138978 254044 138984
rect 253900 138832 253952 138838
rect 253900 138774 253952 138780
rect 254004 128722 254032 138978
rect 253052 128694 253112 128722
rect 253972 128694 254032 128722
rect 254188 128586 254216 139046
rect 256660 138832 256712 138838
rect 256660 138774 256712 138780
rect 254820 138628 254872 138634
rect 254820 138570 254872 138576
rect 254832 130338 254860 138570
rect 254820 130332 254872 130338
rect 254820 130274 254872 130280
rect 255556 130332 255608 130338
rect 255556 130274 255608 130280
rect 255568 128722 255596 130274
rect 256672 128722 256700 138774
rect 257500 128722 257528 139522
rect 258328 139450 258356 141886
rect 259248 139790 259276 141886
rect 260168 139926 260196 141886
rect 260156 139920 260208 139926
rect 260156 139862 260208 139868
rect 259236 139784 259288 139790
rect 259236 139726 259288 139732
rect 258684 139512 258736 139518
rect 258684 139454 258736 139460
rect 258316 139444 258368 139450
rect 258316 139386 258368 139392
rect 258696 128722 258724 139454
rect 261180 139314 261208 141886
rect 261168 139308 261220 139314
rect 261168 139250 261220 139256
rect 262100 139110 262128 141886
rect 263112 139178 263140 141886
rect 264124 139654 264152 141886
rect 264112 139648 264164 139654
rect 264112 139590 264164 139596
rect 264480 139240 264532 139246
rect 264480 139182 264532 139188
rect 263100 139172 263152 139178
rect 263100 139114 263152 139120
rect 262088 139104 262140 139110
rect 262088 139046 262140 139052
rect 258960 131284 259012 131290
rect 258960 131226 259012 131232
rect 255568 128694 255720 128722
rect 256640 128694 256700 128722
rect 257468 128694 257528 128722
rect 258388 128694 258724 128722
rect 254188 128558 254800 128586
rect 240374 122208 240430 122217
rect 240374 122143 240430 122152
rect 240388 122042 240416 122143
rect 240376 122036 240428 122042
rect 240376 121978 240428 121984
rect 231636 110952 231688 110958
rect 231634 110920 231636 110929
rect 239088 110952 239140 110958
rect 231688 110920 231690 110929
rect 239088 110894 239140 110900
rect 240100 110952 240152 110958
rect 240100 110894 240152 110900
rect 231634 110855 231690 110864
rect 240112 109841 240140 110894
rect 240098 109832 240154 109841
rect 240098 109767 240154 109776
rect 240374 108880 240430 108889
rect 240374 108815 240430 108824
rect 240388 108238 240416 108815
rect 231544 108232 231596 108238
rect 231544 108174 231596 108180
rect 240376 108232 240428 108238
rect 240376 108174 240428 108180
rect 231450 92288 231506 92297
rect 231450 92223 231506 92232
rect 231556 88897 231584 108174
rect 236236 105512 236288 105518
rect 236236 105454 236288 105460
rect 236248 95794 236276 105454
rect 236236 95788 236288 95794
rect 236236 95730 236288 95736
rect 237248 95788 237300 95794
rect 237248 95730 237300 95736
rect 231820 95040 231872 95046
rect 231818 95008 231820 95017
rect 231872 95008 231874 95017
rect 231818 94943 231874 94952
rect 232740 94428 232792 94434
rect 232740 94370 232792 94376
rect 231542 88888 231598 88897
rect 231542 88823 231598 88832
rect 232752 85934 232780 94370
rect 230992 85928 231044 85934
rect 230992 85870 231044 85876
rect 232740 85928 232792 85934
rect 232740 85870 232792 85876
rect 231004 85769 231032 85870
rect 230990 85760 231046 85769
rect 230990 85695 231046 85704
rect 233476 76408 233528 76414
rect 233476 76350 233528 76356
rect 233488 75297 233516 76350
rect 237260 75818 237288 95730
rect 240374 95552 240430 95561
rect 240374 95487 240430 95496
rect 240388 94434 240416 95487
rect 240376 94428 240428 94434
rect 240376 94370 240428 94376
rect 248930 89160 248986 89169
rect 248986 89118 249280 89146
rect 248930 89095 248986 89104
rect 243208 88846 243452 88874
rect 243760 88846 244004 88874
rect 244404 88846 244464 88874
rect 245048 88846 245384 88874
rect 245600 88846 245844 88874
rect 246244 88846 246580 88874
rect 246888 88846 247224 88874
rect 247440 88846 247776 88874
rect 248084 88846 248512 88874
rect 248728 88846 249064 88874
rect 243424 87430 243452 88846
rect 243412 87424 243464 87430
rect 243412 87366 243464 87372
rect 243976 87226 244004 88846
rect 243964 87220 244016 87226
rect 243964 87162 244016 87168
rect 243044 87152 243096 87158
rect 243044 87094 243096 87100
rect 241664 87016 241716 87022
rect 241664 86958 241716 86964
rect 240284 86880 240336 86886
rect 240284 86822 240336 86828
rect 238904 86812 238956 86818
rect 238904 86754 238956 86760
rect 238916 75818 238944 86754
rect 240296 75818 240324 86822
rect 241676 75818 241704 86958
rect 242582 85896 242638 85905
rect 242582 85831 242638 85840
rect 242596 76521 242624 85831
rect 242582 76512 242638 76521
rect 242582 76447 242638 76456
rect 243056 75818 243084 87094
rect 244436 87090 244464 88846
rect 244424 87084 244476 87090
rect 244424 87026 244476 87032
rect 245356 86954 245384 88846
rect 245344 86948 245396 86954
rect 245344 86890 245396 86896
rect 244884 78856 244936 78862
rect 244884 78798 244936 78804
rect 244896 75818 244924 78798
rect 245816 78794 245844 88846
rect 246552 86138 246580 88846
rect 246540 86132 246592 86138
rect 246540 86074 246592 86080
rect 247092 86132 247144 86138
rect 247092 86074 247144 86080
rect 245804 78788 245856 78794
rect 245804 78730 245856 78736
rect 247104 78726 247132 86074
rect 247092 78720 247144 78726
rect 247092 78662 247144 78668
rect 247196 78590 247224 88846
rect 247748 86138 247776 88846
rect 247736 86132 247788 86138
rect 247736 86074 247788 86080
rect 247644 78924 247696 78930
rect 247644 78866 247696 78872
rect 247184 78584 247236 78590
rect 247184 78526 247236 78532
rect 246264 78176 246316 78182
rect 246264 78118 246316 78124
rect 246276 75818 246304 78118
rect 247656 75818 247684 78866
rect 248484 78522 248512 88846
rect 249036 87362 249064 88846
rect 249128 88489 249156 89118
rect 252164 88982 252408 89010
rect 249574 88888 249630 88897
rect 249630 88846 249924 88874
rect 250568 88846 250904 88874
rect 251212 88846 251364 88874
rect 251764 88846 252100 88874
rect 249574 88823 249630 88832
rect 249114 88480 249170 88489
rect 249114 88415 249170 88424
rect 250772 87424 250824 87430
rect 250772 87366 250824 87372
rect 249024 87356 249076 87362
rect 249024 87298 249076 87304
rect 250680 86268 250732 86274
rect 250680 86210 250732 86216
rect 248564 86132 248616 86138
rect 248564 86074 248616 86080
rect 248576 78658 248604 86074
rect 250404 79128 250456 79134
rect 250404 79070 250456 79076
rect 248564 78652 248616 78658
rect 248564 78594 248616 78600
rect 248472 78516 248524 78522
rect 248472 78458 248524 78464
rect 249024 77972 249076 77978
rect 249024 77914 249076 77920
rect 249036 75818 249064 77914
rect 250416 75818 250444 79070
rect 250692 78182 250720 86210
rect 250784 79202 250812 87366
rect 250876 86721 250904 88846
rect 251336 87566 251364 88846
rect 251324 87560 251376 87566
rect 251324 87502 251376 87508
rect 252072 86857 252100 88846
rect 252164 88081 252192 88982
rect 253052 88846 253112 88874
rect 252150 88072 252206 88081
rect 252150 88007 252206 88016
rect 252058 86848 252114 86857
rect 252058 86783 252114 86792
rect 250862 86712 250918 86721
rect 250862 86647 250918 86656
rect 252164 86177 252192 88007
rect 252980 87220 253032 87226
rect 252980 87162 253032 87168
rect 252150 86168 252206 86177
rect 252150 86103 252206 86112
rect 250772 79196 250824 79202
rect 250772 79138 250824 79144
rect 251416 79196 251468 79202
rect 251416 79138 251468 79144
rect 250680 78176 250732 78182
rect 250680 78118 250732 78124
rect 237260 75790 237596 75818
rect 238916 75790 238976 75818
rect 240296 75790 240356 75818
rect 241676 75790 241736 75818
rect 243056 75790 243116 75818
rect 244588 75790 244924 75818
rect 245968 75790 246304 75818
rect 247348 75790 247684 75818
rect 248728 75790 249064 75818
rect 250108 75790 250444 75818
rect 251428 75818 251456 79138
rect 252992 76090 253020 87162
rect 253084 86993 253112 88846
rect 253268 88846 253604 88874
rect 254248 88846 254308 88874
rect 253070 86984 253126 86993
rect 253070 86919 253126 86928
rect 253268 86818 253296 88846
rect 253532 87084 253584 87090
rect 253532 87026 253584 87032
rect 253256 86812 253308 86818
rect 253256 86754 253308 86760
rect 253440 86200 253492 86206
rect 253440 86142 253492 86148
rect 253452 77978 253480 86142
rect 253544 79202 253572 87026
rect 254280 86886 254308 88846
rect 254556 88846 254892 88874
rect 255108 88846 255444 88874
rect 255752 88846 256088 88874
rect 256396 88846 256732 88874
rect 256948 88846 257284 88874
rect 257684 88846 257928 88874
rect 258420 88846 258572 88874
rect 254556 87022 254584 88846
rect 255108 87158 255136 88846
rect 255096 87152 255148 87158
rect 255096 87094 255148 87100
rect 254544 87016 254596 87022
rect 254544 86958 254596 86964
rect 255556 86948 255608 86954
rect 255556 86890 255608 86896
rect 254268 86880 254320 86886
rect 254268 86822 254320 86828
rect 254820 86132 254872 86138
rect 254820 86074 254872 86080
rect 253532 79196 253584 79202
rect 253532 79138 253584 79144
rect 254176 79196 254228 79202
rect 254176 79138 254228 79144
rect 253440 77972 253492 77978
rect 253440 77914 253492 77920
rect 252946 76062 253020 76090
rect 251428 75790 251580 75818
rect 252946 75804 252974 76062
rect 254188 75818 254216 79138
rect 254832 78862 254860 86074
rect 254820 78856 254872 78862
rect 254820 78798 254872 78804
rect 255568 75818 255596 86890
rect 255752 86138 255780 88846
rect 256396 86274 256424 88846
rect 256384 86268 256436 86274
rect 256384 86210 256436 86216
rect 256948 86138 256976 88846
rect 257580 86540 257632 86546
rect 257580 86482 257632 86488
rect 255740 86132 255792 86138
rect 255740 86074 255792 86080
rect 256200 86132 256252 86138
rect 256200 86074 256252 86080
rect 256936 86132 256988 86138
rect 256936 86074 256988 86080
rect 256212 78930 256240 86074
rect 257592 79134 257620 86482
rect 257684 86206 257712 88846
rect 258420 86546 258448 88846
rect 258972 87362 259000 131226
rect 264492 125306 264520 139182
rect 280316 136186 280344 144690
rect 279108 136180 279160 136186
rect 279108 136122 279160 136128
rect 280304 136180 280356 136186
rect 280304 136122 280356 136128
rect 279120 133740 279148 136122
rect 283168 134321 283196 147734
rect 285928 138537 285956 147734
rect 290528 142481 290556 147884
rect 292724 144816 292776 144822
rect 292724 144758 292776 144764
rect 290514 142472 290570 142481
rect 290514 142407 290570 142416
rect 290974 142472 291030 142481
rect 290974 142407 291030 142416
rect 290988 142102 291016 142407
rect 290976 142096 291028 142102
rect 290976 142038 291028 142044
rect 285914 138528 285970 138537
rect 285914 138463 285970 138472
rect 287202 138528 287258 138537
rect 287202 138463 287258 138472
rect 287216 137886 287244 138463
rect 287204 137880 287256 137886
rect 287204 137822 287256 137828
rect 292736 136322 292764 144758
rect 294208 144657 294236 147884
rect 294194 144648 294250 144657
rect 294194 144583 294250 144592
rect 297796 143394 297824 147884
rect 301476 147762 301504 147884
rect 301108 147734 301504 147762
rect 297784 143388 297836 143394
rect 297784 143330 297836 143336
rect 297796 143161 297824 143330
rect 297782 143152 297838 143161
rect 297782 143087 297838 143096
rect 301108 141121 301136 147734
rect 303854 143832 303910 143841
rect 303854 143767 303910 143776
rect 303868 143462 303896 143767
rect 305064 143462 305092 147884
rect 308744 144754 308772 147884
rect 312332 144822 312360 147884
rect 312320 144816 312372 144822
rect 312320 144758 312372 144764
rect 308732 144748 308784 144754
rect 308732 144690 308784 144696
rect 316012 144210 316040 147884
rect 310020 144204 310072 144210
rect 310020 144146 310072 144152
rect 316000 144204 316052 144210
rect 316000 144146 316052 144152
rect 303856 143456 303908 143462
rect 303856 143398 303908 143404
rect 305052 143456 305104 143462
rect 305052 143398 305104 143404
rect 301094 141112 301150 141121
rect 301094 141047 301150 141056
rect 302014 141112 302070 141121
rect 302014 141047 302070 141056
rect 302028 140606 302056 141047
rect 302016 140600 302068 140606
rect 302016 140542 302068 140548
rect 310032 136458 310060 144146
rect 316276 142028 316328 142034
rect 316276 141970 316328 141976
rect 316288 141354 316316 141970
rect 316276 141348 316328 141354
rect 316276 141290 316328 141296
rect 304040 136452 304092 136458
rect 304040 136394 304092 136400
rect 310020 136452 310072 136458
rect 310020 136394 310072 136400
rect 291528 136316 291580 136322
rect 291528 136258 291580 136264
rect 292724 136316 292776 136322
rect 292724 136258 292776 136264
rect 283154 134312 283210 134321
rect 283154 134247 283210 134256
rect 283168 133738 283196 134247
rect 291540 133740 291568 136258
rect 304052 133740 304080 136394
rect 316288 133754 316316 141290
rect 283156 133732 283208 133738
rect 316288 133726 316578 133754
rect 283156 133674 283208 133680
rect 270366 125472 270422 125481
rect 270366 125407 270422 125416
rect 270380 125306 270408 125407
rect 263836 125300 263888 125306
rect 263836 125242 263888 125248
rect 264480 125300 264532 125306
rect 264480 125242 264532 125248
rect 270368 125300 270420 125306
rect 270368 125242 270420 125248
rect 260338 122616 260394 122625
rect 260338 122551 260394 122560
rect 260064 87560 260116 87566
rect 260062 87528 260064 87537
rect 260352 87537 260380 122551
rect 261166 118808 261222 118817
rect 261166 118743 261222 118752
rect 261180 117962 261208 118743
rect 261168 117956 261220 117962
rect 261168 117898 261220 117904
rect 263098 98816 263154 98825
rect 263098 98751 263154 98760
rect 263112 93006 263140 98751
rect 263100 93000 263152 93006
rect 263100 92942 263152 92948
rect 260116 87528 260118 87537
rect 260062 87463 260118 87472
rect 260338 87528 260394 87537
rect 260338 87463 260394 87472
rect 258960 87356 259012 87362
rect 258960 87298 259012 87304
rect 258408 86540 258460 86546
rect 258408 86482 258460 86488
rect 257672 86200 257724 86206
rect 257672 86142 257724 86148
rect 257580 79128 257632 79134
rect 257580 79070 257632 79076
rect 256200 78924 256252 78930
rect 256200 78866 256252 78872
rect 256936 78788 256988 78794
rect 256936 78730 256988 78736
rect 256948 75818 256976 78730
rect 258408 78720 258460 78726
rect 258408 78662 258460 78668
rect 258420 75818 258448 78662
rect 261076 78652 261128 78658
rect 261076 78594 261128 78600
rect 259696 78584 259748 78590
rect 259696 78526 259748 78532
rect 259708 75818 259736 78526
rect 261088 75818 261116 78594
rect 262456 78516 262508 78522
rect 262456 78458 262508 78464
rect 262468 75818 262496 78458
rect 263848 75818 263876 125242
rect 268620 117956 268672 117962
rect 268620 117898 268672 117904
rect 268632 108889 268660 117898
rect 268618 108880 268674 108889
rect 268618 108815 268674 108824
rect 270368 93000 270420 93006
rect 270368 92942 270420 92948
rect 270380 92297 270408 92942
rect 270366 92288 270422 92297
rect 270366 92223 270422 92232
rect 276268 83814 276466 83842
rect 283444 83814 283550 83842
rect 290344 83814 290726 83842
rect 297520 83814 297810 83842
rect 304880 83814 304986 83842
rect 311872 83814 312070 83842
rect 319140 83814 319246 83842
rect 276268 81990 276296 83814
rect 276256 81984 276308 81990
rect 276256 81926 276308 81932
rect 283444 81922 283472 83814
rect 283432 81916 283484 81922
rect 283432 81858 283484 81864
rect 283444 81310 283472 81858
rect 290344 81854 290372 83814
rect 290332 81848 290384 81854
rect 290332 81790 290384 81796
rect 297520 81378 297548 83814
rect 304880 83706 304908 83814
rect 304880 83678 305092 83706
rect 285824 81372 285876 81378
rect 285824 81314 285876 81320
rect 297508 81372 297560 81378
rect 297508 81314 297560 81320
rect 283432 81304 283484 81310
rect 283432 81246 283484 81252
rect 266596 76408 266648 76414
rect 266596 76350 266648 76356
rect 254188 75790 254340 75818
rect 255568 75790 255720 75818
rect 256948 75790 257100 75818
rect 258420 75790 258572 75818
rect 259708 75790 259952 75818
rect 261088 75790 261332 75818
rect 262468 75790 262712 75818
rect 263848 75790 264092 75818
rect 249206 75560 249262 75569
rect 249206 75495 249262 75504
rect 249220 75462 249248 75495
rect 249208 75456 249260 75462
rect 249208 75398 249260 75404
rect 266608 75297 266636 76350
rect 233474 75288 233530 75297
rect 233474 75223 233530 75232
rect 266594 75288 266650 75297
rect 266594 75223 266650 75232
rect 267422 74200 267478 74209
rect 267422 74135 267478 74144
rect 233934 73928 233990 73937
rect 233934 73863 233990 73872
rect 233474 72568 233530 72577
rect 233474 72503 233530 72512
rect 233488 72402 233516 72503
rect 230164 72396 230216 72402
rect 230164 72338 230216 72344
rect 233476 72396 233528 72402
rect 233476 72338 233528 72344
rect 229888 69608 229940 69614
rect 229888 69550 229940 69556
rect 229900 66418 229928 69550
rect 230176 69478 230204 72338
rect 233474 71480 233530 71489
rect 233474 71415 233530 71424
rect 230164 69472 230216 69478
rect 230164 69414 230216 69420
rect 233488 68186 233516 71415
rect 233750 71072 233806 71081
rect 233750 71007 233806 71016
rect 233566 69712 233622 69721
rect 233566 69647 233622 69656
rect 233580 69614 233608 69647
rect 233568 69608 233620 69614
rect 233568 69550 233620 69556
rect 233658 68352 233714 68361
rect 233658 68287 233714 68296
rect 233476 68180 233528 68186
rect 233476 68122 233528 68128
rect 233566 67264 233622 67273
rect 233566 67199 233622 67208
rect 233474 66992 233530 67001
rect 233474 66927 233530 66936
rect 233488 66826 233516 66927
rect 230072 66820 230124 66826
rect 230072 66762 230124 66768
rect 233476 66820 233528 66826
rect 233476 66762 233528 66768
rect 229888 66412 229940 66418
rect 229888 66354 229940 66360
rect 229428 65460 229480 65466
rect 229428 65402 229480 65408
rect 229440 62406 229468 65402
rect 230084 64038 230112 66762
rect 233474 65496 233530 65505
rect 233474 65431 233476 65440
rect 233528 65431 233530 65440
rect 233476 65402 233528 65408
rect 233580 65398 233608 67199
rect 233568 65392 233620 65398
rect 233568 65334 233620 65340
rect 233672 65330 233700 68287
rect 233764 66758 233792 71007
rect 233948 69546 233976 73863
rect 264480 73756 264532 73762
rect 264480 73698 264532 73704
rect 233936 69540 233988 69546
rect 233936 69482 233988 69488
rect 233752 66752 233804 66758
rect 233752 66694 233804 66700
rect 233660 65324 233712 65330
rect 233660 65266 233712 65272
rect 234578 64544 234634 64553
rect 234578 64479 234634 64488
rect 230072 64032 230124 64038
rect 230072 63974 230124 63980
rect 233474 63184 233530 63193
rect 233474 63119 233530 63128
rect 233488 62678 233516 63119
rect 233566 62776 233622 62785
rect 233566 62711 233622 62720
rect 230164 62672 230216 62678
rect 230164 62614 230216 62620
rect 233476 62672 233528 62678
rect 233476 62614 233528 62620
rect 229428 62400 229480 62406
rect 229428 62342 229480 62348
rect 230176 61114 230204 62614
rect 233474 61416 233530 61425
rect 233474 61351 233530 61360
rect 230164 61108 230216 61114
rect 230164 61050 230216 61056
rect 233488 59822 233516 61351
rect 233580 59890 233608 62711
rect 234592 62610 234620 64479
rect 234580 62604 234632 62610
rect 234580 62546 234632 62552
rect 233658 60056 233714 60065
rect 233658 59991 233714 60000
rect 233568 59884 233620 59890
rect 233568 59826 233620 59832
rect 233476 59816 233528 59822
rect 233476 59758 233528 59764
rect 233566 58968 233622 58977
rect 233566 58903 233622 58912
rect 233474 58696 233530 58705
rect 230348 58660 230400 58666
rect 233580 58666 233608 58903
rect 233474 58631 233530 58640
rect 233568 58660 233620 58666
rect 230348 58602 230400 58608
rect 230360 56966 230388 58602
rect 233488 58598 233516 58631
rect 233568 58602 233620 58608
rect 230624 58592 230676 58598
rect 230624 58534 230676 58540
rect 233476 58592 233528 58598
rect 233476 58534 233528 58540
rect 230348 56960 230400 56966
rect 230348 56902 230400 56908
rect 230636 56694 230664 58534
rect 233672 58530 233700 59991
rect 233660 58524 233712 58530
rect 233660 58466 233712 58472
rect 233474 57200 233530 57209
rect 233474 57135 233530 57144
rect 230624 56688 230676 56694
rect 230624 56630 230676 56636
rect 233488 55742 233516 57135
rect 234394 55976 234450 55985
rect 234394 55911 234450 55920
rect 233476 55736 233528 55742
rect 233476 55678 233528 55684
rect 233474 55296 233530 55305
rect 233474 55231 233530 55240
rect 233488 55062 233516 55231
rect 233476 55056 233528 55062
rect 233476 54998 233528 55004
rect 233474 54480 233530 54489
rect 233474 54415 233476 54424
rect 233528 54415 233530 54424
rect 233476 54386 233528 54392
rect 234408 54382 234436 55911
rect 234396 54376 234448 54382
rect 234396 54318 234448 54324
rect 233476 53696 233528 53702
rect 233476 53638 233528 53644
rect 233488 53537 233516 53638
rect 233474 53528 233530 53537
rect 233474 53463 233530 53472
rect 228600 51588 228652 51594
rect 228600 51530 228652 51536
rect 233566 50808 233622 50817
rect 233566 50743 233622 50752
rect 233474 50400 233530 50409
rect 233580 50370 233608 50743
rect 233474 50335 233530 50344
rect 233568 50364 233620 50370
rect 233488 50302 233516 50335
rect 233568 50306 233620 50312
rect 233476 50296 233528 50302
rect 233476 50238 233528 50244
rect 233474 49040 233530 49049
rect 233474 48975 233530 48984
rect 233488 48942 233516 48975
rect 233476 48936 233528 48942
rect 233476 48878 233528 48884
rect 264492 48097 264520 73698
rect 266594 73248 266650 73257
rect 266594 73183 266650 73192
rect 266608 72402 266636 73183
rect 266596 72396 266648 72402
rect 266596 72338 266648 72344
rect 266686 72160 266742 72169
rect 266686 72095 266742 72104
rect 266594 71072 266650 71081
rect 266700 71042 266728 72095
rect 266594 71007 266650 71016
rect 266688 71036 266740 71042
rect 266608 70974 266636 71007
rect 266688 70978 266740 70984
rect 266596 70968 266648 70974
rect 266596 70910 266648 70916
rect 266594 70120 266650 70129
rect 266594 70055 266650 70064
rect 266608 69614 266636 70055
rect 266596 69608 266648 69614
rect 266596 69550 266648 69556
rect 267436 69546 267464 74135
rect 285836 72402 285864 81314
rect 305064 73762 305092 83678
rect 311872 80170 311900 83814
rect 319140 80630 319168 83814
rect 316920 80624 316972 80630
rect 316920 80566 316972 80572
rect 319128 80624 319180 80630
rect 319128 80566 319180 80572
rect 311872 80142 312084 80170
rect 312056 76414 312084 80142
rect 312044 76408 312096 76414
rect 312044 76350 312096 76356
rect 304868 73756 304920 73762
rect 304868 73698 304920 73704
rect 305052 73756 305104 73762
rect 305052 73698 305104 73704
rect 304880 72402 304908 73698
rect 316932 72538 316960 80566
rect 311216 72532 311268 72538
rect 311216 72474 311268 72480
rect 316920 72532 316972 72538
rect 316920 72474 316972 72480
rect 274968 72396 275020 72402
rect 274968 72338 275020 72344
rect 284536 72396 284588 72402
rect 284536 72338 284588 72344
rect 285824 72396 285876 72402
rect 285824 72338 285876 72344
rect 297876 72396 297928 72402
rect 297876 72338 297928 72344
rect 304868 72396 304920 72402
rect 304868 72338 304920 72344
rect 274784 71036 274836 71042
rect 274784 70978 274836 70984
rect 274692 70968 274744 70974
rect 274692 70910 274744 70916
rect 270552 69608 270604 69614
rect 270552 69550 270604 69556
rect 267424 69540 267476 69546
rect 267424 69482 267476 69488
rect 266594 69032 266650 69041
rect 266594 68967 266650 68976
rect 266608 68254 266636 68967
rect 266596 68248 266648 68254
rect 266596 68190 266648 68196
rect 266686 67944 266742 67953
rect 266686 67879 266742 67888
rect 266594 66992 266650 67001
rect 266594 66927 266650 66936
rect 266608 66826 266636 66927
rect 266700 66894 266728 67879
rect 267240 67568 267292 67574
rect 267240 67510 267292 67516
rect 266688 66888 266740 66894
rect 266688 66830 266740 66836
rect 266596 66820 266648 66826
rect 266596 66762 266648 66768
rect 266594 65904 266650 65913
rect 266594 65839 266650 65848
rect 266608 65466 266636 65839
rect 266596 65460 266648 65466
rect 266596 65402 266648 65408
rect 266594 64952 266650 64961
rect 266594 64887 266650 64896
rect 266608 64106 266636 64887
rect 266596 64100 266648 64106
rect 266596 64042 266648 64048
rect 266686 63864 266742 63873
rect 266686 63799 266742 63808
rect 266594 62776 266650 62785
rect 266700 62746 266728 63799
rect 266594 62711 266650 62720
rect 266688 62740 266740 62746
rect 266608 62678 266636 62711
rect 266688 62682 266740 62688
rect 266596 62672 266648 62678
rect 266596 62614 266648 62620
rect 266594 61824 266650 61833
rect 266594 61759 266650 61768
rect 266608 61318 266636 61759
rect 266596 61312 266648 61318
rect 266596 61254 266648 61260
rect 266594 60736 266650 60745
rect 266594 60671 266650 60680
rect 266608 59958 266636 60671
rect 266596 59952 266648 59958
rect 266596 59894 266648 59900
rect 266686 59648 266742 59657
rect 266686 59583 266742 59592
rect 266594 58696 266650 58705
rect 266594 58631 266596 58640
rect 266648 58631 266650 58640
rect 266596 58602 266648 58608
rect 266700 58598 266728 59583
rect 266688 58592 266740 58598
rect 266688 58534 266740 58540
rect 266594 57608 266650 57617
rect 266594 57543 266650 57552
rect 266608 57170 266636 57543
rect 266596 57164 266648 57170
rect 266596 57106 266648 57112
rect 266594 56656 266650 56665
rect 266594 56591 266650 56600
rect 266608 55810 266636 56591
rect 266596 55804 266648 55810
rect 266596 55746 266648 55752
rect 267252 55577 267280 67510
rect 270564 66758 270592 69550
rect 272668 68248 272720 68254
rect 272668 68190 272720 68196
rect 272484 66888 272536 66894
rect 272484 66830 272536 66836
rect 270552 66752 270604 66758
rect 270552 66694 270604 66700
rect 272496 65398 272524 66830
rect 272484 65392 272536 65398
rect 272484 65334 272536 65340
rect 272680 65330 272708 68190
rect 272760 66820 272812 66826
rect 272760 66762 272812 66768
rect 272668 65324 272720 65330
rect 272668 65266 272720 65272
rect 272772 63630 272800 66762
rect 274704 66729 274732 70910
rect 274796 67681 274824 70978
rect 274876 69540 274928 69546
rect 274876 69482 274928 69488
rect 274888 69449 274916 69482
rect 274874 69440 274930 69449
rect 274874 69375 274930 69384
rect 274980 68497 275008 72338
rect 284548 69820 284576 72338
rect 297888 69820 297916 72338
rect 311228 69820 311256 72474
rect 321610 69440 321666 69449
rect 321610 69375 321666 69384
rect 321624 68594 321652 69375
rect 321612 68588 321664 68594
rect 321612 68530 321664 68536
rect 274966 68488 275022 68497
rect 274966 68423 275022 68432
rect 321610 68488 321666 68497
rect 321610 68423 321666 68432
rect 321624 68390 321652 68423
rect 321612 68384 321664 68390
rect 321612 68326 321664 68332
rect 274782 67672 274838 67681
rect 320506 67672 320562 67681
rect 274782 67607 274838 67616
rect 317392 67630 317604 67658
rect 274876 66752 274928 66758
rect 274690 66720 274746 66729
rect 274876 66694 274928 66700
rect 274690 66655 274746 66664
rect 274888 65913 274916 66694
rect 274874 65904 274930 65913
rect 274874 65839 274930 65848
rect 274968 65460 275020 65466
rect 274968 65402 275020 65408
rect 274876 65392 274928 65398
rect 274876 65334 274928 65340
rect 274888 64145 274916 65334
rect 274874 64136 274930 64145
rect 273036 64100 273088 64106
rect 274874 64071 274930 64080
rect 273036 64042 273088 64048
rect 272760 63624 272812 63630
rect 272760 63566 272812 63572
rect 272760 62740 272812 62746
rect 272760 62682 272812 62688
rect 272668 61312 272720 61318
rect 272668 61254 272720 61260
rect 272680 59890 272708 61254
rect 272772 61250 272800 62682
rect 273048 62610 273076 64042
rect 274876 63624 274928 63630
rect 274876 63566 274928 63572
rect 274888 63193 274916 63566
rect 274874 63184 274930 63193
rect 274874 63119 274930 63128
rect 273036 62604 273088 62610
rect 273036 62546 273088 62552
rect 274876 62604 274928 62610
rect 274876 62546 274928 62552
rect 274888 61425 274916 62546
rect 274980 62377 275008 65402
rect 275060 65324 275112 65330
rect 275060 65266 275112 65272
rect 275072 64961 275100 65266
rect 275058 64952 275114 64961
rect 275058 64887 275114 64896
rect 275060 62672 275112 62678
rect 275060 62614 275112 62620
rect 274966 62368 275022 62377
rect 274966 62303 275022 62312
rect 274874 61416 274930 61425
rect 274874 61351 274930 61360
rect 272760 61244 272812 61250
rect 272760 61186 272812 61192
rect 274876 61244 274928 61250
rect 274876 61186 274928 61192
rect 274888 60473 274916 61186
rect 274874 60464 274930 60473
rect 274874 60399 274930 60408
rect 274968 59952 275020 59958
rect 274968 59894 275020 59900
rect 272668 59884 272720 59890
rect 272668 59826 272720 59832
rect 274876 59884 274928 59890
rect 274876 59826 274928 59832
rect 274888 58705 274916 59826
rect 274874 58696 274930 58705
rect 272576 58660 272628 58666
rect 274874 58631 274930 58640
rect 272576 58602 272628 58608
rect 272588 57034 272616 58602
rect 272760 58592 272812 58598
rect 272760 58534 272812 58540
rect 272772 57102 272800 58534
rect 274980 57889 275008 59894
rect 275072 59657 275100 62614
rect 275058 59648 275114 59657
rect 275058 59583 275114 59592
rect 274966 57880 275022 57889
rect 274966 57815 275022 57824
rect 274968 57164 275020 57170
rect 274968 57106 275020 57112
rect 272760 57096 272812 57102
rect 272760 57038 272812 57044
rect 274876 57096 274928 57102
rect 274876 57038 274928 57044
rect 272576 57028 272628 57034
rect 272576 56970 272628 56976
rect 274888 56937 274916 57038
rect 274874 56928 274930 56937
rect 274874 56863 274930 56872
rect 273404 55804 273456 55810
rect 273404 55746 273456 55752
rect 267238 55568 267294 55577
rect 267238 55503 267294 55512
rect 266594 54480 266650 54489
rect 266594 54415 266596 54424
rect 266648 54415 266650 54424
rect 266596 54386 266648 54392
rect 273416 54382 273444 55746
rect 274980 55169 275008 57106
rect 275060 57028 275112 57034
rect 275060 56970 275112 56976
rect 275072 56121 275100 56970
rect 275058 56112 275114 56121
rect 275058 56047 275114 56056
rect 274966 55160 275022 55169
rect 274966 55095 275022 55104
rect 317392 55010 317420 67630
rect 317576 67574 317604 67630
rect 320506 67607 320562 67616
rect 317564 67568 317616 67574
rect 317564 67510 317616 67516
rect 320520 67234 320548 67607
rect 320508 67228 320560 67234
rect 320508 67170 320560 67176
rect 321060 66888 321112 66894
rect 321060 66830 321112 66836
rect 321072 63193 321100 66830
rect 321426 66720 321482 66729
rect 321426 66655 321482 66664
rect 321440 65738 321468 66655
rect 321610 65904 321666 65913
rect 321610 65839 321612 65848
rect 321664 65839 321666 65848
rect 321612 65810 321664 65816
rect 321428 65732 321480 65738
rect 321428 65674 321480 65680
rect 321704 65460 321756 65466
rect 321704 65402 321756 65408
rect 321428 65120 321480 65126
rect 321428 65062 321480 65068
rect 321440 64145 321468 65062
rect 321610 64952 321666 64961
rect 321610 64887 321666 64896
rect 321624 64786 321652 64887
rect 321612 64780 321664 64786
rect 321612 64722 321664 64728
rect 321426 64136 321482 64145
rect 321426 64071 321482 64080
rect 321058 63184 321114 63193
rect 321058 63119 321114 63128
rect 321244 62400 321296 62406
rect 321716 62377 321744 65402
rect 321244 62342 321296 62348
rect 321702 62368 321758 62377
rect 321256 61425 321284 62342
rect 321702 62303 321758 62312
rect 321242 61416 321298 61425
rect 321242 61351 321298 61360
rect 321060 61312 321112 61318
rect 321060 61254 321112 61260
rect 320876 61040 320928 61046
rect 320876 60982 320928 60988
rect 320888 60473 320916 60982
rect 320874 60464 320930 60473
rect 320874 60399 320930 60408
rect 321072 58705 321100 61254
rect 321610 59648 321666 59657
rect 321610 59583 321666 59592
rect 321624 58802 321652 59583
rect 321612 58796 321664 58802
rect 321612 58738 321664 58744
rect 321058 58696 321114 58705
rect 321058 58631 321114 58640
rect 320874 57880 320930 57889
rect 320874 57815 320930 57824
rect 320888 57238 320916 57815
rect 320876 57232 320928 57238
rect 320876 57174 320928 57180
rect 321058 56928 321114 56937
rect 321058 56863 321114 56872
rect 321072 56082 321100 56863
rect 321612 56348 321664 56354
rect 321612 56290 321664 56296
rect 321624 56121 321652 56290
rect 321610 56112 321666 56121
rect 321060 56076 321112 56082
rect 321610 56047 321666 56056
rect 321060 56018 321112 56024
rect 321610 55160 321666 55169
rect 321610 55095 321666 55104
rect 317472 55056 317524 55062
rect 317392 55004 317472 55010
rect 317392 54998 317524 55004
rect 317392 54982 317512 54998
rect 321624 54994 321652 55095
rect 321612 54988 321664 54994
rect 273404 54376 273456 54382
rect 274876 54376 274928 54382
rect 273404 54318 273456 54324
rect 274874 54344 274876 54353
rect 274928 54344 274930 54353
rect 274874 54279 274930 54288
rect 266596 53696 266648 53702
rect 266596 53638 266648 53644
rect 266608 53537 266636 53638
rect 266594 53528 266650 53537
rect 266594 53463 266650 53472
rect 279028 51594 279056 53908
rect 279016 51588 279068 51594
rect 279016 51530 279068 51536
rect 266686 51352 266742 51361
rect 266686 51287 266742 51296
rect 266594 50400 266650 50409
rect 266700 50370 266728 51287
rect 280304 50908 280356 50914
rect 280304 50850 280356 50856
rect 266594 50335 266650 50344
rect 266688 50364 266740 50370
rect 266608 50302 266636 50335
rect 266688 50306 266740 50312
rect 266596 50296 266648 50302
rect 266596 50238 266648 50244
rect 274966 49992 275022 50001
rect 274966 49927 275022 49936
rect 274980 49622 275008 49927
rect 274968 49616 275020 49622
rect 274968 49558 275020 49564
rect 275612 49616 275664 49622
rect 275612 49558 275664 49564
rect 275060 49548 275112 49554
rect 275060 49490 275112 49496
rect 275072 49321 275100 49490
rect 266594 49312 266650 49321
rect 266594 49247 266650 49256
rect 275058 49312 275114 49321
rect 275058 49247 275114 49256
rect 266608 48942 266636 49247
rect 266596 48936 266648 48942
rect 266596 48878 266648 48884
rect 266594 48360 266650 48369
rect 266594 48295 266650 48304
rect 241110 48088 241166 48097
rect 262914 48088 262970 48097
rect 241166 48046 241460 48074
rect 241110 48023 241166 48032
rect 264478 48088 264534 48097
rect 262970 48046 263264 48074
rect 262914 48023 262970 48032
rect 264478 48023 264534 48032
rect 244882 47952 244938 47961
rect 238424 47910 238668 47938
rect 244588 47910 244882 47938
rect 233474 47816 233530 47825
rect 233474 47751 233530 47760
rect 233488 47514 233516 47751
rect 233476 47508 233528 47514
rect 233476 47450 233528 47456
rect 238640 45950 238668 47910
rect 253990 47952 254046 47961
rect 247716 47910 248052 47938
rect 250844 47910 251180 47938
rect 253880 47910 253990 47938
rect 244882 47887 244938 47896
rect 248024 47281 248052 47910
rect 248010 47272 248066 47281
rect 248010 47207 248066 47216
rect 238628 45944 238680 45950
rect 238628 45886 238680 45892
rect 251152 45785 251180 47910
rect 253990 47887 254046 47896
rect 256948 47910 257008 47938
rect 260136 47910 260380 47938
rect 256948 46057 256976 47910
rect 260352 46601 260380 47910
rect 266608 47514 266636 48295
rect 266596 47508 266648 47514
rect 266596 47450 266648 47456
rect 260338 46592 260394 46601
rect 260338 46527 260394 46536
rect 256934 46048 256990 46057
rect 256934 45983 256990 45992
rect 263190 46048 263246 46057
rect 263190 45983 263246 45992
rect 256948 45882 256976 45983
rect 263204 45882 263232 45983
rect 256936 45876 256988 45882
rect 256936 45818 256988 45824
rect 263192 45876 263244 45882
rect 263192 45818 263244 45824
rect 251138 45776 251194 45785
rect 251138 45711 251194 45720
rect 263204 44794 263232 45818
rect 263192 44788 263244 44794
rect 263192 44730 263244 44736
rect 223540 37104 223592 37110
rect 223540 37046 223592 37052
rect 223000 35126 223120 35154
rect 223000 34746 223028 35126
rect 222554 34718 223028 34746
rect 190078 34582 190644 34610
rect 182324 33024 182376 33030
rect 182324 32966 182376 32972
rect 182230 26056 182286 26065
rect 182230 25991 182286 26000
rect 181862 23336 181918 23345
rect 181862 23271 181918 23280
rect 182336 20761 182364 32966
rect 275624 23345 275652 49558
rect 275888 49548 275940 49554
rect 275888 49490 275940 49496
rect 275796 48188 275848 48194
rect 275796 48130 275848 48136
rect 275808 47961 275836 48130
rect 275794 47952 275850 47961
rect 275794 47887 275850 47896
rect 275900 47802 275928 49490
rect 276072 48188 276124 48194
rect 276072 48130 276124 48136
rect 275808 47774 275928 47802
rect 275808 33681 275836 47774
rect 275888 46760 275940 46766
rect 275888 46702 275940 46708
rect 275900 46601 275928 46702
rect 275886 46592 275942 46601
rect 275886 46527 275942 46536
rect 275794 33672 275850 33681
rect 275794 33607 275850 33616
rect 275900 30825 275928 46527
rect 275980 45400 276032 45406
rect 275980 45342 276032 45348
rect 275992 44794 276020 45342
rect 275980 44788 276032 44794
rect 275980 44730 276032 44736
rect 275886 30816 275942 30825
rect 275886 30751 275942 30760
rect 275992 28105 276020 44730
rect 275978 28096 276034 28105
rect 275978 28031 276034 28040
rect 276084 26065 276112 48130
rect 280316 37382 280344 50850
rect 281328 50681 281356 53908
rect 281314 50672 281370 50681
rect 281314 50607 281370 50616
rect 283720 48097 283748 53908
rect 285928 53894 286034 53922
rect 288320 53894 288426 53922
rect 284444 50976 284496 50982
rect 284444 50918 284496 50924
rect 283706 48088 283762 48097
rect 283706 48023 283762 48032
rect 281592 47508 281644 47514
rect 281592 47450 281644 47456
rect 279108 37376 279160 37382
rect 279108 37318 279160 37324
rect 280304 37376 280356 37382
rect 280304 37318 280356 37324
rect 279120 34732 279148 37318
rect 281604 34732 281632 47450
rect 283720 45882 283748 48023
rect 283708 45876 283760 45882
rect 283708 45818 283760 45824
rect 284456 34746 284484 50918
rect 285928 47417 285956 53894
rect 288320 50234 288348 53894
rect 289964 51044 290016 51050
rect 289964 50986 290016 50992
rect 288308 50228 288360 50234
rect 288308 50170 288360 50176
rect 288320 49622 288348 50170
rect 288308 49616 288360 49622
rect 288308 49558 288360 49564
rect 286560 48936 286612 48942
rect 286560 48878 286612 48884
rect 285914 47408 285970 47417
rect 285914 47343 285916 47352
rect 285968 47343 285970 47352
rect 285916 47314 285968 47320
rect 284102 34718 284484 34746
rect 286572 34732 286600 48878
rect 289976 37790 290004 50986
rect 290712 48194 290740 53908
rect 291528 50296 291580 50302
rect 291528 50238 291580 50244
rect 290700 48188 290752 48194
rect 290700 48130 290752 48136
rect 289044 37784 289096 37790
rect 289044 37726 289096 37732
rect 289964 37784 290016 37790
rect 289964 37726 290016 37732
rect 289056 34732 289084 37726
rect 291540 34732 291568 50238
rect 293104 45406 293132 53908
rect 294104 51112 294156 51118
rect 294104 51054 294156 51060
rect 293092 45400 293144 45406
rect 293092 45342 293144 45348
rect 294116 34732 294144 51054
rect 295496 47446 295524 53908
rect 296588 50364 296640 50370
rect 296588 50306 296640 50312
rect 294196 47440 294248 47446
rect 294196 47382 294248 47388
rect 295484 47440 295536 47446
rect 295484 47382 295536 47388
rect 294208 46766 294236 47382
rect 294196 46760 294248 46766
rect 294196 46702 294248 46708
rect 296600 34732 296628 50306
rect 297796 49554 297824 53908
rect 299624 51180 299676 51186
rect 299624 51122 299676 51128
rect 297784 49548 297836 49554
rect 297784 49490 297836 49496
rect 299636 34610 299664 51122
rect 300188 50914 300216 53908
rect 302488 50982 302516 53908
rect 304880 51050 304908 53908
rect 306984 53696 307036 53702
rect 306984 53638 307036 53644
rect 306996 53401 307024 53638
rect 306982 53392 307038 53401
rect 306982 53327 307038 53336
rect 307272 51118 307300 53908
rect 309572 51186 309600 53908
rect 309560 51180 309612 51186
rect 309560 51122 309612 51128
rect 307260 51112 307312 51118
rect 307260 51054 307312 51060
rect 304868 51044 304920 51050
rect 304868 50986 304920 50992
rect 302476 50976 302528 50982
rect 302476 50918 302528 50924
rect 311964 50914 311992 53908
rect 300176 50908 300228 50914
rect 300176 50850 300228 50856
rect 305144 50908 305196 50914
rect 305144 50850 305196 50856
rect 311952 50908 312004 50914
rect 311952 50850 312004 50856
rect 301554 39112 301610 39121
rect 301554 39047 301610 39056
rect 301568 34732 301596 39047
rect 305156 37790 305184 50850
rect 314264 50438 314292 53908
rect 316288 53894 316670 53922
rect 310020 50432 310072 50438
rect 310020 50374 310072 50380
rect 314252 50432 314304 50438
rect 314252 50374 314304 50380
rect 310032 37790 310060 50374
rect 304040 37784 304092 37790
rect 304040 37726 304092 37732
rect 305144 37784 305196 37790
rect 309100 37784 309152 37790
rect 305144 37726 305196 37732
rect 306614 37752 306670 37761
rect 304052 34732 304080 37726
rect 309100 37726 309152 37732
rect 310020 37784 310072 37790
rect 310020 37726 310072 37732
rect 306614 37687 306670 37696
rect 306628 34732 306656 37687
rect 309112 34732 309140 37726
rect 311584 36560 311636 36566
rect 311584 36502 311636 36508
rect 311596 34732 311624 36502
rect 316288 36498 316316 53894
rect 317392 44674 317420 54982
rect 321612 54930 321664 54936
rect 317472 54444 317524 54450
rect 317472 54386 317524 54392
rect 317116 44646 317420 44674
rect 314068 36492 314120 36498
rect 314068 36434 314120 36440
rect 316276 36492 316328 36498
rect 316276 36434 316328 36440
rect 314080 34732 314108 36434
rect 317116 35154 317144 44646
rect 317484 36566 317512 54386
rect 320968 54376 321020 54382
rect 320966 54344 320968 54353
rect 321020 54344 321022 54353
rect 320966 54279 321022 54288
rect 317472 36560 317524 36566
rect 317472 36502 317524 36508
rect 317024 35126 317144 35154
rect 317024 34746 317052 35126
rect 316578 34718 317052 34746
rect 299098 34582 299664 34610
rect 276164 33092 276216 33098
rect 276164 33034 276216 33040
rect 276070 26056 276126 26065
rect 276070 25991 276126 26000
rect 275610 23336 275666 23345
rect 275610 23271 275666 23280
rect 276176 20761 276204 33034
rect 88482 20752 88538 20761
rect 88482 20687 88538 20696
rect 182322 20752 182378 20761
rect 182322 20687 182378 20696
rect 276162 20752 276218 20761
rect 276162 20687 276218 20696
rect 92420 18942 92664 18970
rect 92636 16846 92664 18942
rect 97052 18942 97388 18970
rect 102356 18942 102416 18970
rect 92624 16840 92676 16846
rect 92624 16782 92676 16788
rect 80756 16772 80808 16778
rect 80756 16714 80808 16720
rect 67876 16704 67928 16710
rect 67876 16646 67928 16652
rect 54996 16636 55048 16642
rect 54996 16578 55048 16584
rect 29236 16568 29288 16574
rect 29236 16510 29288 16516
rect 16356 16432 16408 16438
rect 16356 16374 16408 16380
rect 12676 14256 12728 14262
rect 12674 14224 12676 14233
rect 16080 14256 16132 14262
rect 12728 14224 12730 14233
rect 16080 14198 16132 14204
rect 12674 14159 12730 14168
rect 16368 9304 16396 16374
rect 29248 9304 29276 16510
rect 42116 16500 42168 16506
rect 42116 16442 42168 16448
rect 42128 9304 42156 16442
rect 55008 9304 55036 16578
rect 67888 9304 67916 16646
rect 80768 9304 80796 16714
rect 97052 16098 97080 18942
rect 102388 16778 102416 18942
rect 107080 18942 107416 18970
rect 112048 18942 112384 18970
rect 117016 18942 117352 18970
rect 122076 18942 122412 18970
rect 127228 18942 127380 18970
rect 105136 16840 105188 16846
rect 105136 16782 105188 16788
rect 102376 16772 102428 16778
rect 102376 16714 102428 16720
rect 95476 16092 95528 16098
rect 95476 16034 95528 16040
rect 97040 16092 97092 16098
rect 97040 16034 97092 16040
rect 95488 12630 95516 16034
rect 93636 12624 93688 12630
rect 93636 12566 93688 12572
rect 95476 12624 95528 12630
rect 95476 12566 95528 12572
rect 93648 9304 93676 12566
rect 105148 12358 105176 16782
rect 107080 16710 107108 18942
rect 107068 16704 107120 16710
rect 107068 16646 107120 16652
rect 112048 16642 112076 18942
rect 112036 16636 112088 16642
rect 112036 16578 112088 16584
rect 117016 16506 117044 18942
rect 122076 16574 122104 18942
rect 122064 16568 122116 16574
rect 122064 16510 122116 16516
rect 117004 16500 117056 16506
rect 117004 16442 117056 16448
rect 119396 16500 119448 16506
rect 119396 16442 119448 16448
rect 105136 12352 105188 12358
rect 105136 12294 105188 12300
rect 106516 12352 106568 12358
rect 106516 12294 106568 12300
rect 106528 9304 106556 12294
rect 119408 9304 119436 16442
rect 127228 16438 127256 18942
rect 186384 17118 186412 18956
rect 191352 17118 191380 18956
rect 185176 17112 185228 17118
rect 185176 17054 185228 17060
rect 186372 17112 186424 17118
rect 186372 17054 186424 17060
rect 191340 17112 191392 17118
rect 191340 17054 191392 17060
rect 192076 17112 192128 17118
rect 192076 17054 192128 17060
rect 170916 16704 170968 16710
rect 170916 16646 170968 16652
rect 158036 16636 158088 16642
rect 158036 16578 158088 16584
rect 145156 16568 145208 16574
rect 145156 16510 145208 16516
rect 127216 16432 127268 16438
rect 127216 16374 127268 16380
rect 132276 16432 132328 16438
rect 132276 16374 132328 16380
rect 132288 9304 132316 16374
rect 145168 9304 145196 16510
rect 158048 9304 158076 16578
rect 170928 9304 170956 16646
rect 183796 12352 183848 12358
rect 183796 12294 183848 12300
rect 183808 9304 183836 12294
rect 185188 12290 185216 17054
rect 185176 12284 185228 12290
rect 185176 12226 185228 12232
rect 192088 12154 192116 17054
rect 196320 17050 196348 18956
rect 194560 17044 194612 17050
rect 194560 16986 194612 16992
rect 196308 17044 196360 17050
rect 196308 16986 196360 16992
rect 194572 12358 194600 16986
rect 201380 16710 201408 18956
rect 201368 16704 201420 16710
rect 201368 16646 201420 16652
rect 206348 16642 206376 18956
rect 206336 16636 206388 16642
rect 206336 16578 206388 16584
rect 211316 16574 211344 18956
rect 211304 16568 211356 16574
rect 211304 16510 211356 16516
rect 216376 16438 216404 18956
rect 221344 16506 221372 18956
rect 273956 16704 274008 16710
rect 273956 16646 274008 16652
rect 261076 16636 261128 16642
rect 261076 16578 261128 16584
rect 248196 16568 248248 16574
rect 248196 16510 248248 16516
rect 221332 16500 221384 16506
rect 221332 16442 221384 16448
rect 235316 16500 235368 16506
rect 235316 16442 235368 16448
rect 216364 16432 216416 16438
rect 216364 16374 216416 16380
rect 222436 16432 222488 16438
rect 222436 16374 222488 16380
rect 194560 12352 194612 12358
rect 194560 12294 194612 12300
rect 209556 12284 209608 12290
rect 209556 12226 209608 12232
rect 192076 12148 192128 12154
rect 192076 12090 192128 12096
rect 196676 12148 196728 12154
rect 196676 12090 196728 12096
rect 196688 9304 196716 12090
rect 209568 9304 209596 12226
rect 222448 9304 222476 16374
rect 235328 9304 235356 16442
rect 248208 9304 248236 16510
rect 261088 9304 261116 16578
rect 273968 9304 273996 16646
rect 280408 12290 280436 18956
rect 285376 16778 285404 18956
rect 290344 17118 290372 18956
rect 288676 17112 288728 17118
rect 288676 17054 288728 17060
rect 290332 17112 290384 17118
rect 290332 17054 290384 17060
rect 285364 16772 285416 16778
rect 285364 16714 285416 16720
rect 288688 12426 288716 17054
rect 295404 16710 295432 18956
rect 299716 16772 299768 16778
rect 299716 16714 299768 16720
rect 295392 16704 295444 16710
rect 295392 16646 295444 16652
rect 286836 12420 286888 12426
rect 286836 12362 286888 12368
rect 288676 12420 288728 12426
rect 288676 12362 288728 12368
rect 280396 12284 280448 12290
rect 280396 12226 280448 12232
rect 286848 9304 286876 12362
rect 299728 9304 299756 16714
rect 300372 16642 300400 18956
rect 300360 16636 300412 16642
rect 300360 16578 300412 16584
rect 305340 16574 305368 18956
rect 305328 16568 305380 16574
rect 305328 16510 305380 16516
rect 310400 16506 310428 18956
rect 310388 16500 310440 16506
rect 310388 16442 310440 16448
rect 315368 16438 315396 18956
rect 315356 16432 315408 16438
rect 315356 16374 315408 16380
rect 322544 12290 322572 388470
rect 323820 371800 323872 371806
rect 323820 371742 323872 371748
rect 323176 346980 323228 346986
rect 323176 346922 323228 346928
rect 323188 345558 323216 346922
rect 323268 345688 323320 345694
rect 323268 345630 323320 345636
rect 323176 345552 323228 345558
rect 323176 345494 323228 345500
rect 323176 344668 323228 344674
rect 323176 344610 323228 344616
rect 323188 342770 323216 344610
rect 323280 344130 323308 345630
rect 323268 344124 323320 344130
rect 323268 344066 323320 344072
rect 323176 342764 323228 342770
rect 323176 342706 323228 342712
rect 322624 333788 322676 333794
rect 322624 333730 322676 333736
rect 322636 233698 322664 333730
rect 323176 244912 323228 244918
rect 323176 244854 323228 244860
rect 323188 243422 323216 244854
rect 323176 243416 323228 243422
rect 323176 243358 323228 243364
rect 322624 233692 322676 233698
rect 322624 233634 322676 233640
rect 323832 233630 323860 371742
rect 328420 357928 328472 357934
rect 328420 357870 328472 357876
rect 328432 357497 328460 357870
rect 328418 357488 328474 357497
rect 328418 357423 328474 357432
rect 328328 356568 328380 356574
rect 328328 356510 328380 356516
rect 328340 356137 328368 356510
rect 328326 356128 328382 356137
rect 328326 356063 328382 356072
rect 328420 355208 328472 355214
rect 328418 355176 328420 355185
rect 328472 355176 328474 355185
rect 328418 355111 328474 355120
rect 328512 355140 328564 355146
rect 328512 355082 328564 355088
rect 328524 354641 328552 355082
rect 328510 354632 328566 354641
rect 328510 354567 328566 354576
rect 328052 353848 328104 353854
rect 328052 353790 328104 353796
rect 328064 353417 328092 353790
rect 328050 353408 328106 353417
rect 328050 353343 328106 353352
rect 328512 352420 328564 352426
rect 328512 352362 328564 352368
rect 328524 352329 328552 352362
rect 328510 352320 328566 352329
rect 328510 352255 328566 352264
rect 328144 351128 328196 351134
rect 328144 351070 328196 351076
rect 327868 351060 327920 351066
rect 327868 351002 327920 351008
rect 327498 350960 327554 350969
rect 327498 350895 327554 350904
rect 327512 350386 327540 350895
rect 327880 350425 327908 351002
rect 327866 350416 327922 350425
rect 327500 350380 327552 350386
rect 327866 350351 327922 350360
rect 327500 350322 327552 350328
rect 328156 349609 328184 351070
rect 328328 349768 328380 349774
rect 328328 349710 328380 349716
rect 328142 349600 328198 349609
rect 328142 349535 328198 349544
rect 327224 348476 327276 348482
rect 327224 348418 327276 348424
rect 327132 348340 327184 348346
rect 327132 348282 327184 348288
rect 327144 346481 327172 348282
rect 327236 346889 327264 348418
rect 328340 348249 328368 349710
rect 328326 348240 328382 348249
rect 328326 348175 328382 348184
rect 327222 346880 327278 346889
rect 327222 346815 327278 346824
rect 327130 346472 327186 346481
rect 327130 346407 327186 346416
rect 327040 345620 327092 345626
rect 327040 345562 327092 345568
rect 326856 344396 326908 344402
rect 326856 344338 326908 344344
rect 326868 341313 326896 344338
rect 327052 342673 327080 345562
rect 328052 345552 328104 345558
rect 328052 345494 328104 345500
rect 328064 345121 328092 345494
rect 328050 345112 328106 345121
rect 328050 345047 328106 345056
rect 328512 344124 328564 344130
rect 328512 344066 328564 344072
rect 328524 344033 328552 344066
rect 328510 344024 328566 344033
rect 328510 343959 328566 343968
rect 327132 342900 327184 342906
rect 327132 342842 327184 342848
rect 327038 342664 327094 342673
rect 327038 342599 327094 342608
rect 327040 341540 327092 341546
rect 327040 341482 327092 341488
rect 326854 341304 326910 341313
rect 326854 341239 326910 341248
rect 326948 340112 327000 340118
rect 326948 340054 327000 340060
rect 326672 338820 326724 338826
rect 326672 338762 326724 338768
rect 326684 334377 326712 338762
rect 326960 337097 326988 340054
rect 327052 338185 327080 341482
rect 327144 339953 327172 342842
rect 328052 342764 328104 342770
rect 328052 342706 328104 342712
rect 328064 342129 328092 342706
rect 328050 342120 328106 342129
rect 328050 342055 328106 342064
rect 327224 341472 327276 341478
rect 327224 341414 327276 341420
rect 327130 339944 327186 339953
rect 327130 339879 327186 339888
rect 327132 338684 327184 338690
rect 327132 338626 327184 338632
rect 327038 338176 327094 338185
rect 327038 338111 327094 338120
rect 327040 337324 327092 337330
rect 327040 337266 327092 337272
rect 326946 337088 327002 337097
rect 326946 337023 327002 337032
rect 326670 334368 326726 334377
rect 326670 334303 326726 334312
rect 327052 333969 327080 337266
rect 327144 335873 327172 338626
rect 327236 338593 327264 341414
rect 327222 338584 327278 338593
rect 327222 338519 327278 338528
rect 327316 336100 327368 336106
rect 327316 336042 327368 336048
rect 327224 335964 327276 335970
rect 327224 335906 327276 335912
rect 327130 335864 327186 335873
rect 327130 335799 327186 335808
rect 327038 333960 327094 333969
rect 327038 333895 327094 333904
rect 325384 331816 325436 331822
rect 325384 331758 325436 331764
rect 324648 330456 324700 330462
rect 324648 330398 324700 330404
rect 324556 327056 324608 327062
rect 324556 326998 324608 327004
rect 324568 326897 324596 326998
rect 324554 326888 324610 326897
rect 324554 326823 324610 326832
rect 324568 301601 324596 326823
rect 324660 315201 324688 330398
rect 325200 329028 325252 329034
rect 325200 328970 325252 328976
rect 324740 323520 324792 323526
rect 324740 323462 324792 323468
rect 324752 320369 324780 323462
rect 324832 320732 324884 320738
rect 324832 320674 324884 320680
rect 324738 320360 324794 320369
rect 324738 320295 324794 320304
rect 324844 317241 324872 320674
rect 324830 317232 324886 317241
rect 324830 317167 324886 317176
rect 324646 315192 324702 315201
rect 324646 315127 324702 315136
rect 324660 314113 324688 315127
rect 324646 314104 324702 314113
rect 324646 314039 324702 314048
rect 324738 308256 324794 308265
rect 324738 308191 324794 308200
rect 324554 301592 324610 301601
rect 324554 301527 324610 301536
rect 324646 298464 324702 298473
rect 324646 298399 324702 298408
rect 324554 282824 324610 282833
rect 324554 282759 324556 282768
rect 324608 282759 324610 282768
rect 324556 282730 324608 282736
rect 324556 258648 324608 258654
rect 324556 258590 324608 258596
rect 324568 255662 324596 258590
rect 324556 255656 324608 255662
rect 324556 255598 324608 255604
rect 324556 234440 324608 234446
rect 324556 234382 324608 234388
rect 324568 233834 324596 234382
rect 324556 233828 324608 233834
rect 324556 233770 324608 233776
rect 323820 233624 323872 233630
rect 323820 233566 323872 233572
rect 324660 231726 324688 298399
rect 324752 250329 324780 308191
rect 325212 293441 325240 328970
rect 325292 327124 325344 327130
rect 325292 327066 325344 327072
rect 325304 324886 325332 327066
rect 325292 324880 325344 324886
rect 325292 324822 325344 324828
rect 325304 304729 325332 324822
rect 325396 319378 325424 331758
rect 327236 331657 327264 335906
rect 327328 333017 327356 336042
rect 327314 333008 327370 333017
rect 327314 332943 327370 332952
rect 327222 331648 327278 331657
rect 327222 331583 327278 331592
rect 325568 330524 325620 330530
rect 325568 330466 325620 330472
rect 325476 326988 325528 326994
rect 325476 326930 325528 326936
rect 325384 319372 325436 319378
rect 325384 319314 325436 319320
rect 325396 310985 325424 319314
rect 325488 316658 325516 326930
rect 325580 322166 325608 330466
rect 325752 330388 325804 330394
rect 325752 330330 325804 330336
rect 325660 328960 325712 328966
rect 325660 328902 325712 328908
rect 325568 322160 325620 322166
rect 325568 322102 325620 322108
rect 325476 316652 325528 316658
rect 325476 316594 325528 316600
rect 325382 310976 325438 310985
rect 325382 310911 325438 310920
rect 325384 309716 325436 309722
rect 325384 309658 325436 309664
rect 325290 304720 325346 304729
rect 325290 304655 325346 304664
rect 324830 293432 324886 293441
rect 324830 293367 324886 293376
rect 325198 293432 325254 293441
rect 325198 293367 325254 293376
rect 324738 250320 324794 250329
rect 324738 250255 324794 250264
rect 324740 233828 324792 233834
rect 324740 233770 324792 233776
rect 324648 231720 324700 231726
rect 324648 231662 324700 231668
rect 324660 229686 324688 231662
rect 324648 229680 324700 229686
rect 324648 229622 324700 229628
rect 322992 227708 323044 227714
rect 322992 227650 323044 227656
rect 323004 227034 323032 227650
rect 322992 227028 323044 227034
rect 322992 226970 323044 226976
rect 323004 226393 323032 226970
rect 322990 226384 323046 226393
rect 322990 226319 323046 226328
rect 324556 225736 324608 225742
rect 324556 225678 324608 225684
rect 322624 224172 322676 224178
rect 322624 224114 322676 224120
rect 322636 45950 322664 224114
rect 323820 222880 323872 222886
rect 323820 222822 323872 222828
rect 322716 222812 322768 222818
rect 322716 222754 322768 222760
rect 322728 131358 322756 222754
rect 322900 221384 322952 221390
rect 322900 221326 322952 221332
rect 322808 220500 322860 220506
rect 322808 220442 322860 220448
rect 322820 139858 322848 220442
rect 322912 145434 322940 221326
rect 323176 152432 323228 152438
rect 323176 152374 323228 152380
rect 323188 150942 323216 152374
rect 323268 151412 323320 151418
rect 323268 151354 323320 151360
rect 323176 150936 323228 150942
rect 323176 150878 323228 150884
rect 323280 149582 323308 151354
rect 323268 149576 323320 149582
rect 323268 149518 323320 149524
rect 322900 145428 322952 145434
rect 322900 145370 322952 145376
rect 322808 139852 322860 139858
rect 322808 139794 322860 139800
rect 322716 131352 322768 131358
rect 322716 131294 322768 131300
rect 323176 130332 323228 130338
rect 323176 130274 323228 130280
rect 323188 124121 323216 130274
rect 323174 124112 323230 124121
rect 323174 124047 323230 124056
rect 323188 122965 323216 124047
rect 323174 122956 323230 122965
rect 323174 122891 323230 122900
rect 323832 51594 323860 222822
rect 324568 220137 324596 225678
rect 324752 223265 324780 233770
rect 324738 223256 324794 223265
rect 324738 223191 324794 223200
rect 324554 220128 324610 220137
rect 324554 220063 324610 220072
rect 324844 198785 324872 293367
rect 325290 285952 325346 285961
rect 325290 285887 325346 285896
rect 325200 283536 325252 283542
rect 325200 283478 325252 283484
rect 325212 273449 325240 283478
rect 325198 273440 325254 273449
rect 325198 273375 325254 273384
rect 325198 239032 325254 239041
rect 325198 238967 325254 238976
rect 325212 238662 325240 238967
rect 325200 238656 325252 238662
rect 325200 238598 325252 238604
rect 325212 224246 325240 238598
rect 325200 224240 325252 224246
rect 325200 224182 325252 224188
rect 325200 221452 325252 221458
rect 325200 221394 325252 221400
rect 324830 198776 324886 198785
rect 324830 198711 324886 198720
rect 324556 188948 324608 188954
rect 324556 188890 324608 188896
rect 324568 188857 324596 188890
rect 324554 188848 324610 188857
rect 324554 188783 324610 188792
rect 324556 179496 324608 179502
rect 324554 179464 324556 179473
rect 324608 179464 324610 179473
rect 324554 179399 324610 179408
rect 324648 143456 324700 143462
rect 324648 143398 324700 143404
rect 324556 133732 324608 133738
rect 324556 133674 324608 133680
rect 324568 133126 324596 133674
rect 324556 133120 324608 133126
rect 324556 133062 324608 133068
rect 324568 120018 324596 133062
rect 324660 132417 324688 143398
rect 324832 140600 324884 140606
rect 324832 140542 324884 140548
rect 324740 137880 324792 137886
rect 324740 137822 324792 137828
rect 324646 132408 324702 132417
rect 324646 132343 324702 132352
rect 324660 132310 324688 132343
rect 324648 132304 324700 132310
rect 324648 132246 324700 132252
rect 324752 131698 324780 137822
rect 324844 133058 324872 140542
rect 324832 133052 324884 133058
rect 324832 132994 324884 133000
rect 324740 131692 324792 131698
rect 324740 131634 324792 131640
rect 324476 119990 324596 120018
rect 324476 119746 324504 119990
rect 324556 119928 324608 119934
rect 324554 119896 324556 119905
rect 324608 119896 324610 119905
rect 324554 119831 324610 119840
rect 324476 119718 324596 119746
rect 324568 113649 324596 119718
rect 324554 113640 324610 113649
rect 324554 113575 324610 113584
rect 324646 106840 324702 106849
rect 324646 106775 324702 106784
rect 324554 104120 324610 104129
rect 324554 104055 324610 104064
rect 324568 94473 324596 104055
rect 324660 101001 324688 106775
rect 324646 100992 324702 101001
rect 324646 100927 324702 100936
rect 325212 98281 325240 221394
rect 325304 220642 325332 285887
rect 325396 279705 325424 309658
rect 325488 298473 325516 316594
rect 325580 308265 325608 322102
rect 325672 320738 325700 328902
rect 325764 323526 325792 330330
rect 328418 330288 328474 330297
rect 328418 330223 328474 330232
rect 328432 329102 328460 330223
rect 348120 329974 348870 330002
rect 330088 329838 331298 329866
rect 331468 329838 332034 329866
rect 328420 329096 328472 329102
rect 328420 329038 328472 329044
rect 326580 326920 326632 326926
rect 326580 326862 326632 326868
rect 325752 323520 325804 323526
rect 325752 323462 325804 323468
rect 325660 320732 325712 320738
rect 325660 320674 325712 320680
rect 325566 308256 325622 308265
rect 325566 308191 325622 308200
rect 325474 298464 325530 298473
rect 325474 298399 325530 298408
rect 325476 295912 325528 295918
rect 325476 295854 325528 295860
rect 325382 279696 325438 279705
rect 325382 279631 325438 279640
rect 325488 276577 325516 295854
rect 325474 276568 325530 276577
rect 325474 276503 325530 276512
rect 325568 238588 325620 238594
rect 325568 238530 325620 238536
rect 325384 235868 325436 235874
rect 325384 235810 325436 235816
rect 325396 225742 325424 235810
rect 325580 231046 325608 238530
rect 325658 234408 325714 234417
rect 325658 234343 325714 234352
rect 325568 231040 325620 231046
rect 325568 230982 325620 230988
rect 325476 229680 325528 229686
rect 325476 229622 325528 229628
rect 325384 225736 325436 225742
rect 325384 225678 325436 225684
rect 325382 224344 325438 224353
rect 325382 224279 325384 224288
rect 325436 224279 325438 224288
rect 325384 224250 325436 224256
rect 325292 220636 325344 220642
rect 325292 220578 325344 220584
rect 325384 220568 325436 220574
rect 325384 220510 325436 220516
rect 325292 215876 325344 215882
rect 325292 215818 325344 215824
rect 325304 185729 325332 215818
rect 325396 191985 325424 220510
rect 325488 204497 325516 229622
rect 325580 210753 325608 230982
rect 325672 224382 325700 234343
rect 326592 232270 326620 326862
rect 330088 282794 330116 329838
rect 331468 320194 331496 329838
rect 332848 320262 332876 329852
rect 333676 327402 333704 329852
rect 334320 329838 334426 329866
rect 332928 327396 332980 327402
rect 332928 327338 332980 327344
rect 333664 327396 333716 327402
rect 333664 327338 333716 327344
rect 334216 327396 334268 327402
rect 334216 327338 334268 327344
rect 332836 320256 332888 320262
rect 332836 320198 332888 320204
rect 331456 320188 331508 320194
rect 331456 320130 331508 320136
rect 332940 319990 332968 327338
rect 334228 320330 334256 327338
rect 334216 320324 334268 320330
rect 334216 320266 334268 320272
rect 334320 320058 334348 329838
rect 335240 327402 335268 329852
rect 335608 329838 336082 329866
rect 335228 327396 335280 327402
rect 335228 327338 335280 327344
rect 335608 320398 335636 329838
rect 336804 326926 336832 329852
rect 336988 329838 337646 329866
rect 338368 329838 338474 329866
rect 335688 326920 335740 326926
rect 335688 326862 335740 326868
rect 336792 326920 336844 326926
rect 336792 326862 336844 326868
rect 335596 320392 335648 320398
rect 335596 320334 335648 320340
rect 335700 320126 335728 326862
rect 336988 320534 337016 329838
rect 337160 327532 337212 327538
rect 337160 327474 337212 327480
rect 337068 326580 337120 326586
rect 337068 326522 337120 326528
rect 336976 320528 337028 320534
rect 336976 320470 337028 320476
rect 335688 320120 335740 320126
rect 335688 320062 335740 320068
rect 334308 320052 334360 320058
rect 334308 319994 334360 320000
rect 332928 319984 332980 319990
rect 332928 319926 332980 319932
rect 337080 316810 337108 326522
rect 337172 320670 337200 327474
rect 337160 320664 337212 320670
rect 337160 320606 337212 320612
rect 337528 320664 337580 320670
rect 337528 320606 337580 320612
rect 337540 316810 337568 320606
rect 338368 320466 338396 329838
rect 338632 327464 338684 327470
rect 339196 327441 339224 329852
rect 339920 327600 339972 327606
rect 339920 327542 339972 327548
rect 338632 327406 338684 327412
rect 339182 327432 339238 327441
rect 338540 326988 338592 326994
rect 338540 326930 338592 326936
rect 338356 320460 338408 320466
rect 338356 320402 338408 320408
rect 338552 319650 338580 326930
rect 338540 319644 338592 319650
rect 338540 319586 338592 319592
rect 338644 316810 338672 327406
rect 339182 327367 339238 327376
rect 339552 327328 339604 327334
rect 339552 327270 339604 327276
rect 339564 320670 339592 327270
rect 339932 327146 339960 327542
rect 340024 327441 340052 329852
rect 340010 327432 340066 327441
rect 340010 327367 340066 327376
rect 339932 327118 340052 327146
rect 339920 327056 339972 327062
rect 339920 326998 339972 327004
rect 339932 320670 339960 326998
rect 339276 320664 339328 320670
rect 339276 320606 339328 320612
rect 339552 320664 339604 320670
rect 339552 320606 339604 320612
rect 339920 320664 339972 320670
rect 339920 320606 339972 320612
rect 339288 316810 339316 320606
rect 339552 319644 339604 319650
rect 339552 319586 339604 319592
rect 337080 316782 337232 316810
rect 337540 316782 337784 316810
rect 338428 316782 338672 316810
rect 339072 316782 339316 316810
rect 339564 316810 339592 319586
rect 340024 316810 340052 327118
rect 340852 326858 340880 329852
rect 341484 327396 341536 327402
rect 341484 327338 341536 327344
rect 341208 327124 341260 327130
rect 341208 327066 341260 327072
rect 340840 326852 340892 326858
rect 340840 326794 340892 326800
rect 340564 320664 340616 320670
rect 340564 320606 340616 320612
rect 340576 316810 340604 320606
rect 341220 319378 341248 327066
rect 341208 319372 341260 319378
rect 341208 319314 341260 319320
rect 341496 317082 341524 327338
rect 341588 326790 341616 329852
rect 342416 327198 342444 329852
rect 342496 327668 342548 327674
rect 342496 327610 342548 327616
rect 342404 327192 342456 327198
rect 342404 327134 342456 327140
rect 342508 326897 342536 327610
rect 342494 326888 342550 326897
rect 342494 326823 342550 326832
rect 341576 326784 341628 326790
rect 341576 326726 341628 326732
rect 341760 319372 341812 319378
rect 341760 319314 341812 319320
rect 341450 317054 341524 317082
rect 339564 316782 339624 316810
rect 340024 316782 340268 316810
rect 340576 316782 340912 316810
rect 341450 316796 341478 317054
rect 341772 316810 341800 319314
rect 342508 318170 342536 326823
rect 343244 326654 343272 329852
rect 343980 326722 344008 329852
rect 344808 327266 344836 329852
rect 344796 327260 344848 327266
rect 344796 327202 344848 327208
rect 343968 326716 344020 326722
rect 343968 326658 344020 326664
rect 343232 326648 343284 326654
rect 343232 326590 343284 326596
rect 345636 326518 345664 329852
rect 346464 327674 346492 329852
rect 346452 327668 346504 327674
rect 346452 327610 346504 327616
rect 345624 326512 345676 326518
rect 345624 326454 345676 326460
rect 347200 324886 347228 329852
rect 343876 324880 343928 324886
rect 343876 324822 343928 324828
rect 347188 324880 347240 324886
rect 347188 324822 347240 324828
rect 342508 318142 343088 318170
rect 343060 316810 343088 318142
rect 343888 316810 343916 324822
rect 347004 323520 347056 323526
rect 347004 323462 347056 323468
rect 344336 323452 344388 323458
rect 344336 323394 344388 323400
rect 344348 322166 344376 323394
rect 344336 322160 344388 322166
rect 344336 322102 344388 322108
rect 344348 316810 344376 322102
rect 346452 322092 346504 322098
rect 346452 322034 346504 322040
rect 346464 320738 346492 322034
rect 346452 320732 346504 320738
rect 346452 320674 346504 320680
rect 346084 320596 346136 320602
rect 346084 320538 346136 320544
rect 345164 319372 345216 319378
rect 345164 319314 345216 319320
rect 345176 316810 345204 319314
rect 341772 316782 342108 316810
rect 343060 316782 343304 316810
rect 343888 316782 343948 316810
rect 344348 316782 344592 316810
rect 345176 316782 345236 316810
rect 345622 316688 345678 316697
rect 342752 316658 343088 316674
rect 342752 316652 343100 316658
rect 342752 316646 343048 316652
rect 346096 316674 346124 320538
rect 346464 317082 346492 320674
rect 346418 317054 346492 317082
rect 346418 316796 346446 317054
rect 347016 316810 347044 323462
rect 348028 323458 348056 329852
rect 348016 323452 348068 323458
rect 348016 323394 348068 323400
rect 348120 323338 348148 329974
rect 348028 323310 348148 323338
rect 349408 329838 349606 329866
rect 348028 320346 348056 323310
rect 349408 320602 349436 329838
rect 350420 322098 350448 329852
rect 351248 323526 351276 329852
rect 351984 327334 352012 329852
rect 352812 327538 352840 329852
rect 352800 327532 352852 327538
rect 352800 327474 352852 327480
rect 353640 327470 353668 329852
rect 353628 327464 353680 327470
rect 353628 327406 353680 327412
rect 351972 327328 352024 327334
rect 351972 327270 352024 327276
rect 354376 326926 354404 329852
rect 355204 326994 355232 329852
rect 356032 327606 356060 329852
rect 356020 327600 356072 327606
rect 356020 327542 356072 327548
rect 355560 327192 355612 327198
rect 355560 327134 355612 327140
rect 355192 326988 355244 326994
rect 355192 326930 355244 326936
rect 354364 326920 354416 326926
rect 354364 326862 354416 326868
rect 354180 326784 354232 326790
rect 354180 326726 354232 326732
rect 352892 325220 352944 325226
rect 352892 325162 352944 325168
rect 352904 324857 352932 325162
rect 352890 324848 352946 324857
rect 352890 324783 352946 324792
rect 353074 324848 353130 324857
rect 353074 324783 353130 324792
rect 351236 323520 351288 323526
rect 351236 323462 351288 323468
rect 350408 322092 350460 322098
rect 350408 322034 350460 322040
rect 349396 320596 349448 320602
rect 349396 320538 349448 320544
rect 351604 320528 351656 320534
rect 351604 320470 351656 320476
rect 350684 320392 350736 320398
rect 348028 320318 348148 320346
rect 350684 320334 350736 320340
rect 348016 320256 348068 320262
rect 348120 320233 348148 320318
rect 349764 320324 349816 320330
rect 349764 320266 349816 320272
rect 348016 320198 348068 320204
rect 348106 320224 348162 320233
rect 347280 320188 347332 320194
rect 347280 320130 347332 320136
rect 347292 316810 347320 320130
rect 348028 316810 348056 320198
rect 348106 320159 348162 320168
rect 348120 319378 348148 320159
rect 349396 320052 349448 320058
rect 349396 319994 349448 320000
rect 348568 319984 348620 319990
rect 348568 319926 348620 319932
rect 348108 319372 348160 319378
rect 348108 319314 348160 319320
rect 348580 316810 348608 319926
rect 349408 316810 349436 319994
rect 349776 316810 349804 320266
rect 350696 316810 350724 320334
rect 350960 320120 351012 320126
rect 350960 320062 351012 320068
rect 350972 316810 351000 320062
rect 351616 316810 351644 320470
rect 352248 320460 352300 320466
rect 352248 320402 352300 320408
rect 352260 316810 352288 320402
rect 347016 316782 347076 316810
rect 347292 316782 347628 316810
rect 348028 316782 348272 316810
rect 348580 316782 348916 316810
rect 349408 316782 349468 316810
rect 349776 316782 350112 316810
rect 350696 316782 350756 316810
rect 350972 316782 351308 316810
rect 351616 316782 351952 316810
rect 352260 316782 352596 316810
rect 345678 316646 346124 316674
rect 345622 316623 345678 316632
rect 343048 316594 343100 316600
rect 353088 315230 353116 324783
rect 352892 315224 352944 315230
rect 352892 315166 352944 315172
rect 353076 315224 353128 315230
rect 353076 315166 353128 315172
rect 334214 309752 334270 309761
rect 334214 309687 334216 309696
rect 334268 309687 334270 309696
rect 334216 309658 334268 309664
rect 352904 306934 352932 315166
rect 352708 306928 352760 306934
rect 352708 306870 352760 306876
rect 352892 306928 352944 306934
rect 352892 306870 352944 306876
rect 334214 296288 334270 296297
rect 334214 296223 334270 296232
rect 334228 295918 334256 296223
rect 334216 295912 334268 295918
rect 334216 295854 334268 295860
rect 352720 291770 352748 306870
rect 354192 295850 354220 326726
rect 354916 306248 354968 306254
rect 354916 306190 354968 306196
rect 353536 295844 353588 295850
rect 353536 295786 353588 295792
rect 354180 295844 354232 295850
rect 354180 295786 354232 295792
rect 353548 295170 353576 295786
rect 353536 295164 353588 295170
rect 353536 295106 353588 295112
rect 352708 291764 352760 291770
rect 352708 291706 352760 291712
rect 334214 283640 334270 283649
rect 334214 283575 334270 283584
rect 334228 283542 334256 283575
rect 334216 283536 334268 283542
rect 334216 283478 334268 283484
rect 330076 282788 330128 282794
rect 330076 282730 330128 282736
rect 327316 264088 327368 264094
rect 327316 264030 327368 264036
rect 327328 263657 327356 264030
rect 327314 263648 327370 263657
rect 330088 263634 330116 282730
rect 352984 279388 353036 279394
rect 352984 279330 353036 279336
rect 337324 276934 337660 276962
rect 337632 274974 337660 276934
rect 338138 276690 338166 276948
rect 338980 276934 339316 276962
rect 339808 276934 340144 276962
rect 340636 276934 340880 276962
rect 341464 276934 341800 276962
rect 342292 276934 342444 276962
rect 343212 276934 343548 276962
rect 344040 276934 344376 276962
rect 344868 276934 345204 276962
rect 338138 276662 338212 276690
rect 337620 274968 337672 274974
rect 337620 274910 337672 274916
rect 334124 274832 334176 274838
rect 334124 274774 334176 274780
rect 332744 274560 332796 274566
rect 332744 274502 332796 274508
rect 332756 263770 332784 274502
rect 334136 266882 334164 274774
rect 336884 274764 336936 274770
rect 336884 274706 336936 274712
rect 335412 274696 335464 274702
rect 335412 274638 335464 274644
rect 335424 266882 335452 274638
rect 335504 274628 335556 274634
rect 335504 274570 335556 274576
rect 333388 266876 333440 266882
rect 333388 266818 333440 266824
rect 334124 266876 334176 266882
rect 334124 266818 334176 266824
rect 334400 266876 334452 266882
rect 334400 266818 334452 266824
rect 335412 266876 335464 266882
rect 335412 266818 335464 266824
rect 332402 263742 332784 263770
rect 333400 263756 333428 266818
rect 334412 263756 334440 266818
rect 335516 263756 335544 274570
rect 336896 263770 336924 274706
rect 338184 273818 338212 276662
rect 339092 274968 339144 274974
rect 339092 274910 339144 274916
rect 338264 274900 338316 274906
rect 338264 274842 338316 274848
rect 338172 273812 338224 273818
rect 338172 273754 338224 273760
rect 338276 266882 338304 274842
rect 339000 273812 339052 273818
rect 339000 273754 339052 273760
rect 337528 266876 337580 266882
rect 337528 266818 337580 266824
rect 338264 266876 338316 266882
rect 338264 266818 338316 266824
rect 336542 263742 336924 263770
rect 337540 263756 337568 266818
rect 338540 266196 338592 266202
rect 338540 266138 338592 266144
rect 338552 263756 338580 266138
rect 339012 265726 339040 273754
rect 339000 265720 339052 265726
rect 339000 265662 339052 265668
rect 339104 265590 339132 274910
rect 339288 273886 339316 276934
rect 339644 275036 339696 275042
rect 339644 274978 339696 274984
rect 339276 273880 339328 273886
rect 339276 273822 339328 273828
rect 339092 265584 339144 265590
rect 339092 265526 339144 265532
rect 339656 263756 339684 274978
rect 340116 273818 340144 276934
rect 340104 273812 340156 273818
rect 340104 273754 340156 273760
rect 340852 266270 340880 276934
rect 341024 274968 341076 274974
rect 341024 274910 341076 274916
rect 340932 273812 340984 273818
rect 340932 273754 340984 273760
rect 340840 266264 340892 266270
rect 340840 266206 340892 266212
rect 340944 265658 340972 273754
rect 340932 265652 340984 265658
rect 340932 265594 340984 265600
rect 341036 263770 341064 274910
rect 341772 274294 341800 276934
rect 341760 274288 341812 274294
rect 341760 274230 341812 274236
rect 342416 273886 342444 276934
rect 343520 273954 343548 276934
rect 344348 274022 344376 276934
rect 345176 274498 345204 276934
rect 345360 276934 345696 276962
rect 346188 276934 346524 276962
rect 347016 276934 347352 276962
rect 348120 276934 348272 276962
rect 348764 276934 349100 276962
rect 349592 276934 349928 276962
rect 350420 276934 350756 276962
rect 351248 276934 351584 276962
rect 352168 276934 352412 276962
rect 345360 274566 345388 276934
rect 346188 274838 346216 276934
rect 346176 274832 346228 274838
rect 346176 274774 346228 274780
rect 347016 274702 347044 276934
rect 347004 274696 347056 274702
rect 347004 274638 347056 274644
rect 348120 274634 348148 276934
rect 348764 274770 348792 276934
rect 349592 274906 349620 276934
rect 349580 274900 349632 274906
rect 349580 274842 349632 274848
rect 348752 274764 348804 274770
rect 348752 274706 348804 274712
rect 348108 274628 348160 274634
rect 348108 274570 348160 274576
rect 345348 274560 345400 274566
rect 345348 274502 345400 274508
rect 345164 274492 345216 274498
rect 345164 274434 345216 274440
rect 344612 274288 344664 274294
rect 344612 274230 344664 274236
rect 344336 274016 344388 274022
rect 344336 273958 344388 273964
rect 343508 273948 343560 273954
rect 343508 273890 343560 273896
rect 341852 273880 341904 273886
rect 341852 273822 341904 273828
rect 342404 273880 342456 273886
rect 342404 273822 342456 273828
rect 344520 273880 344572 273886
rect 344520 273822 344572 273828
rect 341864 266474 341892 273822
rect 344532 266814 344560 273822
rect 344520 266808 344572 266814
rect 344520 266750 344572 266756
rect 344624 266542 344652 274230
rect 347372 274016 347424 274022
rect 347372 273958 347424 273964
rect 347280 273948 347332 273954
rect 347280 273890 347332 273896
rect 347292 266882 347320 273890
rect 347280 266876 347332 266882
rect 347280 266818 347332 266824
rect 344612 266536 344664 266542
rect 344612 266478 344664 266484
rect 346820 266536 346872 266542
rect 346820 266478 346872 266484
rect 341852 266468 341904 266474
rect 341852 266410 341904 266416
rect 343784 266468 343836 266474
rect 343784 266410 343836 266416
rect 342680 265720 342732 265726
rect 342680 265662 342732 265668
rect 341668 265584 341720 265590
rect 341668 265526 341720 265532
rect 340682 263742 341064 263770
rect 341680 263756 341708 265526
rect 342692 263756 342720 265662
rect 343796 263756 343824 266410
rect 345808 266264 345860 266270
rect 345808 266206 345860 266212
rect 344796 265652 344848 265658
rect 344796 265594 344848 265600
rect 344808 263756 344836 265594
rect 345820 263756 345848 266206
rect 346832 263756 346860 266478
rect 347384 266338 347412 273958
rect 350420 273818 350448 276934
rect 351248 275042 351276 276934
rect 351236 275036 351288 275042
rect 351236 274978 351288 274984
rect 352168 274974 352196 276934
rect 352156 274968 352208 274974
rect 352156 274910 352208 274916
rect 348660 273812 348712 273818
rect 348660 273754 348712 273760
rect 350408 273812 350460 273818
rect 350408 273754 350460 273760
rect 347924 266808 347976 266814
rect 347924 266750 347976 266756
rect 347372 266332 347424 266338
rect 347372 266274 347424 266280
rect 347936 263756 347964 266750
rect 348672 266202 348700 273754
rect 352996 272458 353024 279330
rect 352800 272452 352852 272458
rect 352800 272394 352852 272400
rect 352984 272452 353036 272458
rect 352984 272394 353036 272400
rect 348936 266876 348988 266882
rect 348936 266818 348988 266824
rect 348660 266196 348712 266202
rect 348660 266138 348712 266144
rect 348948 263756 348976 266818
rect 352062 266776 352118 266785
rect 352062 266711 352118 266720
rect 350958 266640 351014 266649
rect 350958 266575 351014 266584
rect 349948 266332 350000 266338
rect 349948 266274 350000 266280
rect 349960 263756 349988 266274
rect 350972 263756 351000 266575
rect 352076 263756 352104 266711
rect 352812 263770 352840 272394
rect 353548 263770 353576 295106
rect 353720 285508 353772 285514
rect 353720 285450 353772 285456
rect 353732 285281 353760 285450
rect 353718 285272 353774 285281
rect 353718 285207 353774 285216
rect 354928 267902 354956 306190
rect 355572 300678 355600 327134
rect 356768 327062 356796 329852
rect 357596 327402 357624 329852
rect 357584 327396 357636 327402
rect 357584 327338 357636 327344
rect 358320 327260 358372 327266
rect 358320 327202 358372 327208
rect 356756 327056 356808 327062
rect 356756 326998 356808 327004
rect 356940 326716 356992 326722
rect 356940 326658 356992 326664
rect 355652 326648 355704 326654
rect 355652 326590 355704 326596
rect 355664 306254 355692 326590
rect 356202 314104 356258 314113
rect 356202 314039 356258 314048
rect 356216 313802 356244 314039
rect 356204 313796 356256 313802
rect 356204 313738 356256 313744
rect 356952 310334 356980 326658
rect 358332 315910 358360 327202
rect 358424 327130 358452 329852
rect 358412 327124 358464 327130
rect 358412 327066 358464 327072
rect 357676 315904 357728 315910
rect 357676 315846 357728 315852
rect 358320 315904 358372 315910
rect 358320 315846 358372 315852
rect 356940 310328 356992 310334
rect 356940 310270 356992 310276
rect 356952 309722 356980 310270
rect 356296 309716 356348 309722
rect 356296 309658 356348 309664
rect 356940 309716 356992 309722
rect 356940 309658 356992 309664
rect 356202 308664 356258 308673
rect 356202 308599 356258 308608
rect 356216 308294 356244 308599
rect 356204 308288 356256 308294
rect 356204 308230 356256 308236
rect 355652 306248 355704 306254
rect 355652 306190 355704 306196
rect 356202 304176 356258 304185
rect 356202 304111 356204 304120
rect 356256 304111 356258 304120
rect 356204 304082 356256 304088
rect 355560 300672 355612 300678
rect 355560 300614 355612 300620
rect 355572 300066 355600 300614
rect 355008 300060 355060 300066
rect 355008 300002 355060 300008
rect 355560 300060 355612 300066
rect 355560 300002 355612 300008
rect 354916 267896 354968 267902
rect 354916 267838 354968 267844
rect 355020 263770 355048 300002
rect 356202 298872 356258 298881
rect 356202 298807 356258 298816
rect 356216 298638 356244 298807
rect 356204 298632 356256 298638
rect 356204 298574 356256 298580
rect 356202 293840 356258 293849
rect 356202 293775 356204 293784
rect 356256 293775 356258 293784
rect 356204 293746 356256 293752
rect 356202 289080 356258 289089
rect 356202 289015 356258 289024
rect 356216 288982 356244 289015
rect 356204 288976 356256 288982
rect 356204 288918 356256 288924
rect 356202 283776 356258 283785
rect 356202 283711 356258 283720
rect 356216 283474 356244 283711
rect 356204 283468 356256 283474
rect 356204 283410 356256 283416
rect 356202 279424 356258 279433
rect 356202 279359 356258 279368
rect 356216 279326 356244 279359
rect 356204 279320 356256 279326
rect 356204 279262 356256 279268
rect 355836 267896 355888 267902
rect 355836 267838 355888 267844
rect 356308 267850 356336 309658
rect 355848 263770 355876 267838
rect 356308 267822 356704 267850
rect 352812 263742 353102 263770
rect 353548 263742 354114 263770
rect 355020 263742 355126 263770
rect 355848 263742 356230 263770
rect 356676 263634 356704 267822
rect 357688 263770 357716 315846
rect 357688 263742 358254 263770
rect 330088 263606 331390 263634
rect 356676 263606 357242 263634
rect 358332 263618 358452 263634
rect 358332 263612 358464 263618
rect 358332 263606 358412 263612
rect 327314 263583 327370 263592
rect 327222 261744 327278 261753
rect 327222 261679 327278 261688
rect 326762 260384 326818 260393
rect 326762 260319 326818 260328
rect 326776 257226 326804 260319
rect 327236 258450 327264 261679
rect 328418 258888 328474 258897
rect 328418 258823 328474 258832
rect 328432 258654 328460 258823
rect 328420 258648 328472 258654
rect 328420 258590 328472 258596
rect 327224 258444 327276 258450
rect 327224 258386 327276 258392
rect 327222 257528 327278 257537
rect 327222 257463 327278 257472
rect 326764 257220 326816 257226
rect 326764 257162 326816 257168
rect 327236 255866 327264 257463
rect 328050 256168 328106 256177
rect 328050 256103 328106 256112
rect 327224 255860 327276 255866
rect 327224 255802 327276 255808
rect 328064 253690 328092 256103
rect 328418 254672 328474 254681
rect 328418 254607 328474 254616
rect 328052 253684 328104 253690
rect 328052 253626 328104 253632
rect 327222 253312 327278 253321
rect 327222 253247 327278 253256
rect 327236 252058 327264 253247
rect 328432 253078 328460 254607
rect 328420 253072 328472 253078
rect 328420 253014 328472 253020
rect 327224 252052 327276 252058
rect 327224 251994 327276 252000
rect 327130 251952 327186 251961
rect 327130 251887 327186 251896
rect 327144 250630 327172 251887
rect 327132 250624 327184 250630
rect 327132 250566 327184 250572
rect 327222 250592 327278 250601
rect 327222 250527 327278 250536
rect 327236 249542 327264 250527
rect 327224 249536 327276 249542
rect 327224 249478 327276 249484
rect 328420 249128 328472 249134
rect 328418 249096 328420 249105
rect 328472 249096 328474 249105
rect 328418 249031 328474 249040
rect 328418 247736 328474 247745
rect 328418 247671 328420 247680
rect 328472 247671 328474 247680
rect 328420 247642 328472 247648
rect 328420 247564 328472 247570
rect 328420 247506 328472 247512
rect 328432 246929 328460 247506
rect 328418 246920 328474 246929
rect 328418 246855 328474 246864
rect 327868 246204 327920 246210
rect 327868 246146 327920 246152
rect 327880 245569 327908 246146
rect 327866 245560 327922 245569
rect 327866 245495 327922 245504
rect 327868 244776 327920 244782
rect 327868 244718 327920 244724
rect 327880 244073 327908 244718
rect 327866 244064 327922 244073
rect 327866 243999 327922 244008
rect 327040 243484 327092 243490
rect 327040 243426 327092 243432
rect 327052 240673 327080 243426
rect 327868 243416 327920 243422
rect 327868 243358 327920 243364
rect 327880 242713 327908 243358
rect 327866 242704 327922 242713
rect 327866 242639 327922 242648
rect 327224 242260 327276 242266
rect 327224 242202 327276 242208
rect 327132 242124 327184 242130
rect 327132 242066 327184 242072
rect 327038 240664 327094 240673
rect 327038 240599 327094 240608
rect 327144 238633 327172 242066
rect 327236 239313 327264 242202
rect 327222 239304 327278 239313
rect 327222 239239 327278 239248
rect 327130 238624 327186 238633
rect 327130 238559 327186 238568
rect 328420 236616 328472 236622
rect 328418 236584 328420 236593
rect 328472 236584 328474 236593
rect 328418 236519 328474 236528
rect 330088 235862 331390 235890
rect 332402 235862 332784 235890
rect 326580 232264 326632 232270
rect 326580 232206 326632 232212
rect 325660 224376 325712 224382
rect 325660 224318 325712 224324
rect 325566 210744 325622 210753
rect 325566 210679 325622 210688
rect 325672 207625 325700 224318
rect 325752 224308 325804 224314
rect 325752 224250 325804 224256
rect 325764 213881 325792 224250
rect 325844 224240 325896 224246
rect 325844 224182 325896 224188
rect 325856 216737 325884 224182
rect 325842 216728 325898 216737
rect 325842 216663 325898 216672
rect 325750 213872 325806 213881
rect 325750 213807 325806 213816
rect 325658 207616 325714 207625
rect 325658 207551 325714 207560
rect 325474 204488 325530 204497
rect 325474 204423 325530 204432
rect 325476 202072 325528 202078
rect 325476 202014 325528 202020
rect 325382 191976 325438 191985
rect 325382 191911 325438 191920
rect 325290 185720 325346 185729
rect 325290 185655 325346 185664
rect 325488 182601 325516 202014
rect 330088 188954 330116 235862
rect 332756 224858 332784 235862
rect 333400 232474 333428 235876
rect 334412 232474 334440 235876
rect 333388 232468 333440 232474
rect 333388 232410 333440 232416
rect 334124 232468 334176 232474
rect 334124 232410 334176 232416
rect 334400 232468 334452 232474
rect 334400 232410 334452 232416
rect 335412 232468 335464 232474
rect 335412 232410 335464 232416
rect 334136 224994 334164 232410
rect 335424 225130 335452 232410
rect 335412 225124 335464 225130
rect 335412 225066 335464 225072
rect 334124 224988 334176 224994
rect 334124 224930 334176 224936
rect 335516 224926 335544 235876
rect 336542 235862 336924 235890
rect 337554 235862 338304 235890
rect 335504 224920 335556 224926
rect 335504 224862 335556 224868
rect 332744 224852 332796 224858
rect 332744 224794 332796 224800
rect 336896 224518 336924 235862
rect 337160 225396 337212 225402
rect 337160 225338 337212 225344
rect 336884 224512 336936 224518
rect 336884 224454 336936 224460
rect 337172 222834 337200 225338
rect 337712 225056 337764 225062
rect 337712 224998 337764 225004
rect 337724 222834 337752 224998
rect 338276 224654 338304 235862
rect 338552 232474 338580 235876
rect 339564 235862 339670 235890
rect 340682 235862 340880 235890
rect 339000 232536 339052 232542
rect 339000 232478 339052 232484
rect 338540 232468 338592 232474
rect 338540 232410 338592 232416
rect 338356 225464 338408 225470
rect 338356 225406 338408 225412
rect 338264 224648 338316 224654
rect 338264 224590 338316 224596
rect 338368 222834 338396 225406
rect 339012 225402 339040 232478
rect 339564 226778 339592 235862
rect 339644 232468 339696 232474
rect 339644 232410 339696 232416
rect 339656 230366 339684 232410
rect 339644 230360 339696 230366
rect 339644 230302 339696 230308
rect 339564 226750 339684 226778
rect 339000 225396 339052 225402
rect 339000 225338 339052 225344
rect 339552 225260 339604 225266
rect 339552 225202 339604 225208
rect 339000 225192 339052 225198
rect 339000 225134 339052 225140
rect 339012 222834 339040 225134
rect 339564 222834 339592 225202
rect 339656 224586 339684 226750
rect 340196 225396 340248 225402
rect 340196 225338 340248 225344
rect 339644 224580 339696 224586
rect 339644 224522 339696 224528
rect 340208 222834 340236 225338
rect 340852 224858 340880 235862
rect 341024 233352 341076 233358
rect 341024 233294 341076 233300
rect 340932 233012 340984 233018
rect 340932 232954 340984 232960
rect 340840 224852 340892 224858
rect 340840 224794 340892 224800
rect 340944 223106 340972 232954
rect 341036 225402 341064 233294
rect 341680 232542 341708 235876
rect 342600 235862 342706 235890
rect 343520 235862 343810 235890
rect 341668 232536 341720 232542
rect 341668 232478 341720 232484
rect 341392 225464 341444 225470
rect 341392 225406 341444 225412
rect 341024 225396 341076 225402
rect 341024 225338 341076 225344
rect 341298 224888 341354 224897
rect 341298 224823 341300 224832
rect 341352 224823 341354 224832
rect 341300 224794 341352 224800
rect 340898 223078 340972 223106
rect 337172 222806 337232 222834
rect 337724 222806 337784 222834
rect 338368 222806 338428 222834
rect 339012 222806 339072 222834
rect 339564 222806 339624 222834
rect 340208 222806 340268 222834
rect 340898 222820 340926 223078
rect 341404 222834 341432 225406
rect 342036 225396 342088 225402
rect 342036 225338 342088 225344
rect 342048 222834 342076 225338
rect 342600 225062 342628 235862
rect 342864 232536 342916 232542
rect 342864 232478 342916 232484
rect 342588 225056 342640 225062
rect 342588 224998 342640 225004
rect 342680 225056 342732 225062
rect 342680 224998 342732 225004
rect 342692 224897 342720 224998
rect 342678 224888 342734 224897
rect 342678 224823 342734 224832
rect 342876 224790 342904 232478
rect 342956 232468 343008 232474
rect 342956 232410 343008 232416
rect 342968 225198 342996 232410
rect 343048 229680 343100 229686
rect 343048 229622 343100 229628
rect 342956 225192 343008 225198
rect 342956 225134 343008 225140
rect 343060 225010 343088 229622
rect 343520 225266 343548 235862
rect 344808 232474 344836 235876
rect 345440 233828 345492 233834
rect 345440 233770 345492 233776
rect 344796 232468 344848 232474
rect 344796 232410 344848 232416
rect 345164 231720 345216 231726
rect 345164 231662 345216 231668
rect 345176 231046 345204 231662
rect 343968 231040 344020 231046
rect 343968 230982 344020 230988
rect 345164 231040 345216 231046
rect 345164 230982 345216 230988
rect 343784 230292 343836 230298
rect 343784 230234 343836 230240
rect 343796 229686 343824 230234
rect 343784 229680 343836 229686
rect 343784 229622 343836 229628
rect 343508 225260 343560 225266
rect 343508 225202 343560 225208
rect 342968 224982 343088 225010
rect 342864 224784 342916 224790
rect 342864 224726 342916 224732
rect 341404 222806 341464 222834
rect 342048 222806 342108 222834
rect 342968 222698 342996 224982
rect 343048 224784 343100 224790
rect 343048 224726 343100 224732
rect 343060 224382 343088 224726
rect 343048 224376 343100 224382
rect 343048 224318 343100 224324
rect 343060 222834 343088 224318
rect 343980 223106 344008 230982
rect 345452 229090 345480 233770
rect 345820 232542 345848 235876
rect 346544 234440 346596 234446
rect 346544 234382 346596 234388
rect 346556 233834 346584 234382
rect 346544 233828 346596 233834
rect 346544 233770 346596 233776
rect 346832 233358 346860 235876
rect 346820 233352 346872 233358
rect 346820 233294 346872 233300
rect 347936 233018 347964 235876
rect 347924 233012 347976 233018
rect 347924 232954 347976 232960
rect 345808 232536 345860 232542
rect 345808 232478 345860 232484
rect 346728 232536 346780 232542
rect 346728 232478 346780 232484
rect 346636 232468 346688 232474
rect 346636 232410 346688 232416
rect 345452 229062 345940 229090
rect 345716 225736 345768 225742
rect 345716 225678 345768 225684
rect 345728 225441 345756 225678
rect 345714 225432 345770 225441
rect 345714 225367 345770 225376
rect 344244 224308 344296 224314
rect 344244 224250 344296 224256
rect 343934 223078 344008 223106
rect 343060 222806 343304 222834
rect 343934 222820 343962 223078
rect 344256 222834 344284 224250
rect 345164 224240 345216 224246
rect 345164 224182 345216 224188
rect 345176 222834 345204 224182
rect 345728 222834 345756 225367
rect 344256 222806 344592 222834
rect 345176 222806 345236 222834
rect 345728 222806 345788 222834
rect 342752 222670 342996 222698
rect 345912 222698 345940 229062
rect 346648 225470 346676 232410
rect 346636 225464 346688 225470
rect 346636 225406 346688 225412
rect 346740 225402 346768 232478
rect 348948 232474 348976 235876
rect 349960 232542 349988 235876
rect 349948 232536 350000 232542
rect 350972 232513 351000 235876
rect 352076 232513 352104 235876
rect 352720 235862 353102 235890
rect 353548 235862 354114 235890
rect 355020 235862 355126 235890
rect 355848 235862 356230 235890
rect 356308 235862 357242 235890
rect 357688 235862 358254 235890
rect 349948 232478 350000 232484
rect 350958 232504 351014 232513
rect 348936 232468 348988 232474
rect 350958 232439 351014 232448
rect 352062 232504 352118 232513
rect 352062 232439 352118 232448
rect 348936 232410 348988 232416
rect 347004 227708 347056 227714
rect 347004 227650 347056 227656
rect 347016 227034 347044 227650
rect 347004 227028 347056 227034
rect 347004 226970 347056 226976
rect 346728 225396 346780 225402
rect 346728 225338 346780 225344
rect 347016 222834 347044 226970
rect 351604 225260 351656 225266
rect 351604 225202 351656 225208
rect 348568 225124 348620 225130
rect 348568 225066 348620 225072
rect 348016 224988 348068 224994
rect 348016 224930 348068 224936
rect 347280 224444 347332 224450
rect 347280 224386 347332 224392
rect 347292 222834 347320 224386
rect 348028 222834 348056 224930
rect 348580 222834 348608 225066
rect 349396 224920 349448 224926
rect 349396 224862 349448 224868
rect 349408 222834 349436 224862
rect 350684 224648 350736 224654
rect 350684 224590 350736 224596
rect 349764 224512 349816 224518
rect 349764 224454 349816 224460
rect 349776 222834 349804 224454
rect 350696 223106 350724 224590
rect 350696 223078 350770 223106
rect 347016 222806 347076 222834
rect 347292 222806 347628 222834
rect 348028 222806 348272 222834
rect 348580 222806 348916 222834
rect 349408 222806 349468 222834
rect 349776 222806 350112 222834
rect 350742 222820 350770 223078
rect 351282 223084 351334 223090
rect 351282 223026 351334 223032
rect 351294 222820 351322 223026
rect 351616 222834 351644 225202
rect 352248 225192 352300 225198
rect 352248 225134 352300 225140
rect 352260 222834 352288 225134
rect 351616 222806 351952 222834
rect 352260 222806 352596 222834
rect 345912 222670 346432 222698
rect 334214 216184 334270 216193
rect 334214 216119 334270 216128
rect 334228 215882 334256 216119
rect 334216 215876 334268 215882
rect 334216 215818 334268 215824
rect 334214 202856 334270 202865
rect 334214 202791 334270 202800
rect 334228 202078 334256 202791
rect 334216 202072 334268 202078
rect 334216 202014 334268 202020
rect 352720 195822 352748 235862
rect 352892 233080 352944 233086
rect 352892 233022 352944 233028
rect 352800 218664 352852 218670
rect 352800 218606 352852 218612
rect 352708 195816 352760 195822
rect 352708 195758 352760 195764
rect 334214 189528 334270 189537
rect 334214 189463 334270 189472
rect 330076 188948 330128 188954
rect 330076 188890 330128 188896
rect 326580 188268 326632 188274
rect 326580 188210 326632 188216
rect 325474 182592 325530 182601
rect 325474 182527 325530 182536
rect 326592 179502 326620 188210
rect 326580 179496 326632 179502
rect 326580 179438 326632 179444
rect 328420 170248 328472 170254
rect 328420 170190 328472 170196
rect 328432 169137 328460 170190
rect 330088 169930 330116 188890
rect 334228 188274 334256 189463
rect 334216 188268 334268 188274
rect 334216 188210 334268 188216
rect 337324 182822 337660 182850
rect 338152 182822 338304 182850
rect 338980 182822 339592 182850
rect 339808 182822 340144 182850
rect 340636 182822 340880 182850
rect 341464 182822 341708 182850
rect 342292 182822 342444 182850
rect 343212 182822 343548 182850
rect 344040 182822 344376 182850
rect 344868 182822 345020 182850
rect 337632 181338 337660 182822
rect 337620 181332 337672 181338
rect 337620 181274 337672 181280
rect 338276 181270 338304 182822
rect 338264 181264 338316 181270
rect 338264 181206 338316 181212
rect 334124 181060 334176 181066
rect 334124 181002 334176 181008
rect 332744 180720 332796 180726
rect 332744 180662 332796 180668
rect 330088 169902 330852 169930
rect 330824 169658 330852 169902
rect 332756 169794 332784 180662
rect 334136 173042 334164 181002
rect 335504 180992 335556 180998
rect 335504 180934 335556 180940
rect 335412 180652 335464 180658
rect 335412 180594 335464 180600
rect 333388 173036 333440 173042
rect 333388 172978 333440 172984
rect 334124 173036 334176 173042
rect 334124 172978 334176 172984
rect 332402 169766 332784 169794
rect 333400 169780 333428 172978
rect 334400 172900 334452 172906
rect 334400 172842 334452 172848
rect 334412 169780 334440 172842
rect 335424 169794 335452 180594
rect 335516 172906 335544 180934
rect 336884 180924 336936 180930
rect 336884 180866 336936 180872
rect 335504 172900 335556 172906
rect 335504 172842 335556 172848
rect 336896 169794 336924 180866
rect 338264 180856 338316 180862
rect 338264 180798 338316 180804
rect 335424 169766 335530 169794
rect 336542 169766 336924 169794
rect 338276 169658 338304 180798
rect 339564 172906 339592 182822
rect 339644 181128 339696 181134
rect 339644 181070 339696 181076
rect 339552 172900 339604 172906
rect 339552 172842 339604 172848
rect 338540 171948 338592 171954
rect 338540 171890 338592 171896
rect 338552 169780 338580 171890
rect 339656 169780 339684 181070
rect 340116 180386 340144 182822
rect 340104 180380 340156 180386
rect 340104 180322 340156 180328
rect 340852 180046 340880 182822
rect 341116 181332 341168 181338
rect 341116 181274 341168 181280
rect 340932 180788 340984 180794
rect 340932 180730 340984 180736
rect 340840 180040 340892 180046
rect 340840 179982 340892 179988
rect 340944 169794 340972 180730
rect 341024 180380 341076 180386
rect 341024 180322 341076 180328
rect 341036 172974 341064 180322
rect 341024 172968 341076 172974
rect 341024 172910 341076 172916
rect 340682 169766 340972 169794
rect 330824 169630 331390 169658
rect 337554 169630 338304 169658
rect 341128 169658 341156 181274
rect 341680 180250 341708 182822
rect 341760 181264 341812 181270
rect 341760 181206 341812 181212
rect 341668 180244 341720 180250
rect 341668 180186 341720 180192
rect 341772 173042 341800 181206
rect 342416 179978 342444 182822
rect 343520 181270 343548 182822
rect 343508 181264 343560 181270
rect 343508 181206 343560 181212
rect 344348 181202 344376 182822
rect 344992 181338 345020 182822
rect 345452 182822 345696 182850
rect 346188 182822 346524 182850
rect 347016 182822 347352 182850
rect 348028 182822 348272 182850
rect 348764 182822 349100 182850
rect 349592 182822 349928 182850
rect 350420 182822 350756 182850
rect 351248 182822 351584 182850
rect 352168 182822 352412 182850
rect 344980 181332 345032 181338
rect 344980 181274 345032 181280
rect 344336 181196 344388 181202
rect 344336 181138 344388 181144
rect 345452 180726 345480 182822
rect 346188 181066 346216 182822
rect 346176 181060 346228 181066
rect 346176 181002 346228 181008
rect 347016 180998 347044 182822
rect 347280 181264 347332 181270
rect 347280 181206 347332 181212
rect 347004 180992 347056 180998
rect 347004 180934 347056 180940
rect 345440 180720 345492 180726
rect 345440 180662 345492 180668
rect 345992 180244 346044 180250
rect 345992 180186 346044 180192
rect 345256 180040 345308 180046
rect 345256 179982 345308 179988
rect 342404 179972 342456 179978
rect 342404 179914 342456 179920
rect 341760 173036 341812 173042
rect 341760 172978 341812 172984
rect 342680 173036 342732 173042
rect 342680 172978 342732 172984
rect 342692 169780 342720 172978
rect 344796 172968 344848 172974
rect 344796 172910 344848 172916
rect 343784 172900 343836 172906
rect 343784 172842 343836 172848
rect 343796 169780 343824 172842
rect 344808 169780 344836 172910
rect 345268 169658 345296 179982
rect 345900 179972 345952 179978
rect 345900 179914 345952 179920
rect 345912 172974 345940 179914
rect 346004 173042 346032 180186
rect 345992 173036 346044 173042
rect 345992 172978 346044 172984
rect 346820 173036 346872 173042
rect 346820 172978 346872 172984
rect 345900 172968 345952 172974
rect 345900 172910 345952 172916
rect 346832 169780 346860 172978
rect 347292 171954 347320 181206
rect 348028 180658 348056 182822
rect 348108 181196 348160 181202
rect 348108 181138 348160 181144
rect 348016 180652 348068 180658
rect 348016 180594 348068 180600
rect 348120 180538 348148 181138
rect 348764 180930 348792 182822
rect 348752 180924 348804 180930
rect 348752 180866 348804 180872
rect 349592 180862 349620 182822
rect 350420 181270 350448 182822
rect 350408 181264 350460 181270
rect 350408 181206 350460 181212
rect 351248 181134 351276 182822
rect 351236 181128 351288 181134
rect 351236 181070 351288 181076
rect 349580 180856 349632 180862
rect 349580 180798 349632 180804
rect 349396 180788 349448 180794
rect 349396 180730 349448 180736
rect 348028 180510 348148 180538
rect 347924 172968 347976 172974
rect 347924 172910 347976 172916
rect 347280 171948 347332 171954
rect 347280 171890 347332 171896
rect 347936 169780 347964 172910
rect 348028 169658 348056 180510
rect 349408 169658 349436 180730
rect 352168 180590 352196 182822
rect 352156 180584 352208 180590
rect 352156 180526 352208 180532
rect 350958 172936 351014 172945
rect 350958 172871 351014 172880
rect 352062 172936 352118 172945
rect 352062 172871 352118 172880
rect 350972 169780 351000 172871
rect 352076 169780 352104 172871
rect 352720 169794 352748 195758
rect 352812 186250 352840 218606
rect 352904 218534 352932 233022
rect 353076 227640 353128 227646
rect 353076 227582 353128 227588
rect 352892 218528 352944 218534
rect 352892 218470 352944 218476
rect 352984 217236 353036 217242
rect 352984 217178 353036 217184
rect 352892 191668 352944 191674
rect 352892 191610 352944 191616
rect 352904 191441 352932 191610
rect 352890 191432 352946 191441
rect 352890 191367 352946 191376
rect 352812 186222 352932 186250
rect 352800 186160 352852 186166
rect 352800 186102 352852 186108
rect 352812 184097 352840 186102
rect 352798 184088 352854 184097
rect 352798 184023 352854 184032
rect 352904 182193 352932 186222
rect 352890 182184 352946 182193
rect 352890 182119 352946 182128
rect 352996 182057 353024 217178
rect 353088 214454 353116 227582
rect 353260 226280 353312 226286
rect 353260 226222 353312 226228
rect 353168 226212 353220 226218
rect 353168 226154 353220 226160
rect 353180 215814 353208 226154
rect 353168 215808 353220 215814
rect 353168 215750 353220 215756
rect 353272 215746 353300 226222
rect 353352 226144 353404 226150
rect 353352 226086 353404 226092
rect 353364 217174 353392 226086
rect 353444 220636 353496 220642
rect 353444 220578 353496 220584
rect 353352 217168 353404 217174
rect 353352 217110 353404 217116
rect 353260 215740 353312 215746
rect 353260 215682 353312 215688
rect 353076 214448 353128 214454
rect 353076 214390 353128 214396
rect 353456 213094 353484 220578
rect 353444 213088 353496 213094
rect 353444 213030 353496 213036
rect 353548 201330 353576 235862
rect 354916 232060 354968 232066
rect 354916 232002 354968 232008
rect 354928 210986 354956 232002
rect 354916 210980 354968 210986
rect 354916 210922 354968 210928
rect 353536 201324 353588 201330
rect 353536 201266 353588 201272
rect 352982 182048 353038 182057
rect 352982 181983 353038 181992
rect 352720 169766 353102 169794
rect 353548 169658 353576 201266
rect 354928 175150 354956 210922
rect 355020 206838 355048 235862
rect 355848 232066 355876 235862
rect 355836 232060 355888 232066
rect 355836 232002 355888 232008
rect 355098 220264 355154 220273
rect 355098 220199 355154 220208
rect 355112 214046 355140 220199
rect 356308 215921 356336 235862
rect 357688 222041 357716 235862
rect 357674 222032 357730 222041
rect 357674 221967 357730 221976
rect 356294 215912 356350 215921
rect 356294 215847 356350 215856
rect 356202 215232 356258 215241
rect 356202 215167 356258 215176
rect 356216 214114 356244 215167
rect 356204 214108 356256 214114
rect 356204 214050 356256 214056
rect 355100 214040 355152 214046
rect 355100 213982 355152 213988
rect 356018 210200 356074 210209
rect 356018 210135 356074 210144
rect 356032 209626 356060 210135
rect 356020 209620 356072 209626
rect 356020 209562 356072 209568
rect 355008 206832 355060 206838
rect 355008 206774 355060 206780
rect 354916 175144 354968 175150
rect 354916 175086 354968 175092
rect 355020 169794 355048 206774
rect 356202 205304 356258 205313
rect 356202 205239 356258 205248
rect 356216 204798 356244 205239
rect 356204 204792 356256 204798
rect 356204 204734 356256 204740
rect 355926 200272 355982 200281
rect 355926 200207 355982 200216
rect 355940 199290 355968 200207
rect 355928 199284 355980 199290
rect 355928 199226 355980 199232
rect 356202 195240 356258 195249
rect 356202 195175 356258 195184
rect 356216 195142 356244 195175
rect 356204 195136 356256 195142
rect 356204 195078 356256 195084
rect 355190 190208 355246 190217
rect 355190 190143 355246 190152
rect 355204 189634 355232 190143
rect 355192 189628 355244 189634
rect 355192 189570 355244 189576
rect 356202 185312 356258 185321
rect 356202 185247 356258 185256
rect 356216 184058 356244 185247
rect 356204 184052 356256 184058
rect 356204 183994 356256 184000
rect 355836 175144 355888 175150
rect 355836 175086 355888 175092
rect 355848 169794 355876 175086
rect 356308 169794 356336 215847
rect 355020 169766 355126 169794
rect 355848 169766 356230 169794
rect 356308 169766 356796 169794
rect 356768 169658 356796 169766
rect 357688 169658 357716 221967
rect 358332 215678 358360 263606
rect 358412 263554 358464 263560
rect 358412 263476 358464 263482
rect 358412 263418 358464 263424
rect 358424 217106 358452 263418
rect 358412 217100 358464 217106
rect 358412 217042 358464 217048
rect 358320 215672 358372 215678
rect 358320 215614 358372 215620
rect 341128 169630 341694 169658
rect 345268 169630 345834 169658
rect 348028 169630 348962 169658
rect 349408 169630 349974 169658
rect 353548 169630 354114 169658
rect 356768 169630 357242 169658
rect 357688 169630 358254 169658
rect 328418 169128 328474 169137
rect 328418 169063 328474 169072
rect 327222 167768 327278 167777
rect 327222 167703 327278 167712
rect 327236 163522 327264 167703
rect 327498 166408 327554 166417
rect 327498 166343 327554 166352
rect 327224 163516 327276 163522
rect 327224 163458 327276 163464
rect 327222 163416 327278 163425
rect 327222 163351 327278 163360
rect 327236 161618 327264 163351
rect 327512 162434 327540 166343
rect 328418 164912 328474 164921
rect 328418 164847 328474 164856
rect 327500 162428 327552 162434
rect 327500 162370 327552 162376
rect 327314 162192 327370 162201
rect 327314 162127 327370 162136
rect 327224 161612 327276 161618
rect 327224 161554 327276 161560
rect 327328 159374 327356 162127
rect 328432 161482 328460 164847
rect 328420 161476 328472 161482
rect 328420 161418 328472 161424
rect 327406 160696 327462 160705
rect 327406 160631 327462 160640
rect 327316 159368 327368 159374
rect 327222 159336 327278 159345
rect 327316 159310 327368 159316
rect 327222 159271 327278 159280
rect 327236 158218 327264 159271
rect 327224 158212 327276 158218
rect 327224 158154 327276 158160
rect 327420 158014 327448 160631
rect 327408 158008 327460 158014
rect 327222 157976 327278 157985
rect 327408 157950 327460 157956
rect 327222 157911 327278 157920
rect 327236 157198 327264 157911
rect 327224 157192 327276 157198
rect 327224 157134 327276 157140
rect 327222 156616 327278 156625
rect 327222 156551 327278 156560
rect 327236 155430 327264 156551
rect 327224 155424 327276 155430
rect 327224 155366 327276 155372
rect 328418 155120 328474 155129
rect 328418 155055 328420 155064
rect 328472 155055 328474 155064
rect 328420 155026 328472 155032
rect 328420 153792 328472 153798
rect 328418 153760 328420 153769
rect 328472 153760 328474 153769
rect 328418 153695 328474 153704
rect 328236 152500 328288 152506
rect 328236 152442 328288 152448
rect 328248 152409 328276 152442
rect 328234 152400 328290 152409
rect 328234 152335 328290 152344
rect 328420 150936 328472 150942
rect 328418 150904 328420 150913
rect 328472 150904 328474 150913
rect 328418 150839 328474 150848
rect 327224 149644 327276 149650
rect 327224 149586 327276 149592
rect 327236 146697 327264 149586
rect 328420 149576 328472 149582
rect 328418 149544 328420 149553
rect 328472 149544 328474 149553
rect 328418 149479 328474 149488
rect 328328 148420 328380 148426
rect 328328 148362 328380 148368
rect 327222 146688 327278 146697
rect 327222 146623 327278 146632
rect 328340 143977 328368 148362
rect 328512 148284 328564 148290
rect 328512 148226 328564 148232
rect 328420 148216 328472 148222
rect 328418 148184 328420 148193
rect 328472 148184 328474 148193
rect 328418 148119 328474 148128
rect 328524 145337 328552 148226
rect 328510 145328 328566 145337
rect 328510 145263 328566 145272
rect 328326 143968 328382 143977
rect 328326 143903 328382 143912
rect 325384 143388 325436 143394
rect 325384 143330 325436 143336
rect 325396 134486 325424 143330
rect 325936 142096 325988 142102
rect 325936 142038 325988 142044
rect 328418 142064 328474 142073
rect 325948 137206 325976 142038
rect 328418 141999 328474 142008
rect 328432 141354 328460 141999
rect 330088 141886 331390 141914
rect 332402 141886 332784 141914
rect 328420 141348 328472 141354
rect 328420 141290 328472 141296
rect 325936 137200 325988 137206
rect 325936 137142 325988 137148
rect 326580 137200 326632 137206
rect 326580 137142 326632 137148
rect 325384 134480 325436 134486
rect 325384 134422 325436 134428
rect 325292 130400 325344 130406
rect 325292 130342 325344 130348
rect 325304 110929 325332 130342
rect 325396 126025 325424 134422
rect 325476 133052 325528 133058
rect 325476 132994 325528 133000
rect 325488 129833 325516 132994
rect 325568 131692 325620 131698
rect 325568 131634 325620 131640
rect 325474 129824 325530 129833
rect 325474 129759 325530 129768
rect 325580 126954 325608 131634
rect 325488 126926 325608 126954
rect 325382 126016 325438 126025
rect 325382 125951 325438 125960
rect 325384 122036 325436 122042
rect 325384 121978 325436 121984
rect 325290 110920 325346 110929
rect 325290 110855 325346 110864
rect 325290 100448 325346 100457
rect 325290 100383 325346 100392
rect 325198 98272 325254 98281
rect 325198 98207 325254 98216
rect 324554 94464 324610 94473
rect 324554 94399 324610 94408
rect 324556 85792 324608 85798
rect 324556 85734 324608 85740
rect 324568 85633 324596 85734
rect 324554 85624 324610 85633
rect 324554 85559 324610 85568
rect 324556 55804 324608 55810
rect 324556 55746 324608 55752
rect 324568 54382 324596 55746
rect 324556 54376 324608 54382
rect 324556 54318 324608 54324
rect 323820 51588 323872 51594
rect 323820 51530 323872 51536
rect 322624 45944 322676 45950
rect 322624 45886 322676 45892
rect 324556 45400 324608 45406
rect 324556 45342 324608 45348
rect 312596 12284 312648 12290
rect 312596 12226 312648 12232
rect 322532 12284 322584 12290
rect 322532 12226 322584 12232
rect 312608 9304 312636 12226
rect 324568 12170 324596 45342
rect 325304 12426 325332 100383
rect 325396 92297 325424 121978
rect 325488 117321 325516 126926
rect 326592 119934 326620 137142
rect 326580 119928 326632 119934
rect 326580 119870 326632 119876
rect 325474 117312 325530 117321
rect 325474 117247 325530 117256
rect 325476 108232 325528 108238
rect 325476 108174 325528 108180
rect 325488 102610 325516 108174
rect 325488 102582 325608 102610
rect 325382 92288 325438 92297
rect 325382 92223 325438 92232
rect 325580 88897 325608 102582
rect 325842 94736 325898 94745
rect 325842 94671 325844 94680
rect 325896 94671 325898 94680
rect 325844 94642 325896 94648
rect 325566 88888 325622 88897
rect 325566 88823 325622 88832
rect 326592 87498 326620 119870
rect 330088 94706 330116 141886
rect 332756 131086 332784 141886
rect 333400 139586 333428 141900
rect 334412 139586 334440 141900
rect 335424 141886 335530 141914
rect 336542 141886 336924 141914
rect 337554 141886 338212 141914
rect 333388 139580 333440 139586
rect 333388 139522 333440 139528
rect 334124 139580 334176 139586
rect 334124 139522 334176 139528
rect 334400 139580 334452 139586
rect 334400 139522 334452 139528
rect 334136 131154 334164 139522
rect 334124 131148 334176 131154
rect 334124 131090 334176 131096
rect 332744 131080 332796 131086
rect 332744 131022 332796 131028
rect 335424 131018 335452 141886
rect 335504 139580 335556 139586
rect 335504 139522 335556 139528
rect 335516 131358 335544 139522
rect 335504 131352 335556 131358
rect 335504 131294 335556 131300
rect 336896 131222 336924 141886
rect 338080 138696 338132 138702
rect 338080 138638 338132 138644
rect 336884 131216 336936 131222
rect 336884 131158 336936 131164
rect 335412 131012 335464 131018
rect 335412 130954 335464 130960
rect 338092 130338 338120 138638
rect 338184 131494 338212 141886
rect 338552 139314 338580 141900
rect 339472 141886 339670 141914
rect 340682 141886 340880 141914
rect 338540 139308 338592 139314
rect 338540 139250 338592 139256
rect 338264 138628 338316 138634
rect 338264 138570 338316 138576
rect 338172 131488 338224 131494
rect 338172 131430 338224 131436
rect 337528 130332 337580 130338
rect 337528 130274 337580 130280
rect 338080 130332 338132 130338
rect 338080 130274 338132 130280
rect 337540 128722 337568 130274
rect 338276 130082 338304 138570
rect 339472 131766 339500 141886
rect 339552 139308 339604 139314
rect 339552 139250 339604 139256
rect 339460 131760 339512 131766
rect 339460 131702 339512 131708
rect 339564 131562 339592 139250
rect 339736 131760 339788 131766
rect 339736 131702 339788 131708
rect 339552 131556 339604 131562
rect 339552 131498 339604 131504
rect 339748 130898 339776 131702
rect 340852 131086 340880 141886
rect 340932 138900 340984 138906
rect 340932 138842 340984 138848
rect 340840 131080 340892 131086
rect 340840 131022 340892 131028
rect 339656 130870 339776 130898
rect 339656 130746 339684 130870
rect 339644 130740 339696 130746
rect 339644 130682 339696 130688
rect 339552 130604 339604 130610
rect 339552 130546 339604 130552
rect 339368 130536 339420 130542
rect 339368 130478 339420 130484
rect 338724 130468 338776 130474
rect 338724 130410 338776 130416
rect 338184 130054 338304 130082
rect 338184 128722 338212 130054
rect 338736 128722 338764 130410
rect 339380 128722 339408 130478
rect 337232 128694 337568 128722
rect 337784 128694 338212 128722
rect 338428 128694 338764 128722
rect 339072 128694 339408 128722
rect 339564 128722 339592 130546
rect 340564 130332 340616 130338
rect 340564 130274 340616 130280
rect 340576 128722 340604 130274
rect 340944 128994 340972 138842
rect 341024 138832 341076 138838
rect 341024 138774 341076 138780
rect 341036 130338 341064 138774
rect 341680 138702 341708 141900
rect 341668 138696 341720 138702
rect 341668 138638 341720 138644
rect 342692 138634 342720 141900
rect 342784 141886 343810 141914
rect 343888 141886 344822 141914
rect 342680 138628 342732 138634
rect 342680 138570 342732 138576
rect 342404 131420 342456 131426
rect 342404 131362 342456 131368
rect 341760 130672 341812 130678
rect 341760 130614 341812 130620
rect 341024 130332 341076 130338
rect 341024 130274 341076 130280
rect 339564 128694 339624 128722
rect 340268 128694 340604 128722
rect 340898 128966 340972 128994
rect 340898 128708 340926 128966
rect 341772 128722 341800 130614
rect 342416 128722 342444 131362
rect 342496 130808 342548 130814
rect 342496 130750 342548 130756
rect 341464 128694 341800 128722
rect 342108 128694 342444 128722
rect 342508 128722 342536 130750
rect 342784 130474 342812 141886
rect 343324 133732 343376 133738
rect 343324 133674 343376 133680
rect 343336 133126 343364 133674
rect 343324 133120 343376 133126
rect 343324 133062 343376 133068
rect 342772 130468 342824 130474
rect 342772 130410 342824 130416
rect 343336 128994 343364 133062
rect 343888 130542 343916 141886
rect 345820 138634 345848 141900
rect 345900 138900 345952 138906
rect 345900 138842 345952 138848
rect 344520 138628 344572 138634
rect 344520 138570 344572 138576
rect 345808 138628 345860 138634
rect 345808 138570 345860 138576
rect 343968 137880 344020 137886
rect 343968 137822 344020 137828
rect 343980 137206 344008 137822
rect 343968 137200 344020 137206
rect 343968 137142 344020 137148
rect 343980 135522 344008 137142
rect 343980 135494 344192 135522
rect 343968 132372 344020 132378
rect 343968 132314 344020 132320
rect 343980 131698 344008 132314
rect 343968 131692 344020 131698
rect 343968 131634 344020 131640
rect 343876 130536 343928 130542
rect 343876 130478 343928 130484
rect 343980 128994 344008 131634
rect 343290 128966 343364 128994
rect 343934 128966 344008 128994
rect 342508 128694 342752 128722
rect 343290 128708 343318 128966
rect 343934 128708 343962 128966
rect 344164 128722 344192 135494
rect 344532 130610 344560 138570
rect 345716 134480 345768 134486
rect 345716 134422 345768 134428
rect 344520 130604 344572 130610
rect 344520 130546 344572 130552
rect 344888 130264 344940 130270
rect 344888 130206 344940 130212
rect 344900 128722 344928 130206
rect 345728 128722 345756 134422
rect 345912 131426 345940 138842
rect 346832 138702 346860 141900
rect 347936 138838 347964 141900
rect 347924 138832 347976 138838
rect 347924 138774 347976 138780
rect 346820 138696 346872 138702
rect 346820 138638 346872 138644
rect 348948 138634 348976 141900
rect 349960 138906 349988 141900
rect 350972 139625 351000 141900
rect 352076 139625 352104 141900
rect 352720 141886 353102 141914
rect 353548 141886 354114 141914
rect 355020 141886 355126 141914
rect 355848 141886 356230 141914
rect 356308 141886 357242 141914
rect 357688 141886 358254 141914
rect 350958 139616 351014 139625
rect 350958 139551 351014 139560
rect 352062 139616 352118 139625
rect 352062 139551 352118 139560
rect 349948 138900 350000 138906
rect 349948 138842 350000 138848
rect 345992 138628 346044 138634
rect 345992 138570 346044 138576
rect 348936 138628 348988 138634
rect 348936 138570 348988 138576
rect 345900 131420 345952 131426
rect 345900 131362 345952 131368
rect 346004 130678 346032 138570
rect 346544 135092 346596 135098
rect 346544 135034 346596 135040
rect 346556 134486 346584 135034
rect 346544 134480 346596 134486
rect 346544 134422 346596 134428
rect 346544 133800 346596 133806
rect 346544 133742 346596 133748
rect 346556 133058 346584 133742
rect 346360 133052 346412 133058
rect 346360 132994 346412 133000
rect 346544 133052 346596 133058
rect 346544 132994 346596 133000
rect 345992 130672 346044 130678
rect 345992 130614 346044 130620
rect 346372 128722 346400 132994
rect 347004 132304 347056 132310
rect 347004 132246 347056 132252
rect 347016 131698 347044 132246
rect 347004 131692 347056 131698
rect 347004 131634 347056 131640
rect 347016 128722 347044 131634
rect 350960 131556 351012 131562
rect 350960 131498 351012 131504
rect 350408 131488 350460 131494
rect 350408 131430 350460 131436
rect 348568 131352 348620 131358
rect 348568 131294 348620 131300
rect 348016 131148 348068 131154
rect 348016 131090 348068 131096
rect 347280 130876 347332 130882
rect 347280 130818 347332 130824
rect 347292 128722 347320 130818
rect 348028 128722 348056 131090
rect 348580 128722 348608 131294
rect 349764 131216 349816 131222
rect 349764 131158 349816 131164
rect 349396 131012 349448 131018
rect 349396 130954 349448 130960
rect 349408 128722 349436 130954
rect 349776 128722 349804 131158
rect 350420 128722 350448 131430
rect 350972 128722 351000 131498
rect 352248 131080 352300 131086
rect 352248 131022 352300 131028
rect 351604 130740 351656 130746
rect 351604 130682 351656 130688
rect 351616 128722 351644 130682
rect 352260 128722 352288 131022
rect 344164 128694 344592 128722
rect 344900 128694 345236 128722
rect 345728 128694 345788 128722
rect 346372 128694 346432 128722
rect 347016 128694 347076 128722
rect 347292 128694 347628 128722
rect 348028 128694 348272 128722
rect 348580 128694 348916 128722
rect 349408 128694 349468 128722
rect 349776 128694 350112 128722
rect 350420 128694 350756 128722
rect 350972 128694 351308 128722
rect 351616 128694 351952 128722
rect 352260 128694 352596 128722
rect 334214 122208 334270 122217
rect 334214 122143 334270 122152
rect 334228 122042 334256 122143
rect 334216 122036 334268 122042
rect 334216 121978 334268 121984
rect 334214 108880 334270 108889
rect 334214 108815 334270 108824
rect 334228 108238 334256 108815
rect 334216 108232 334268 108238
rect 334216 108174 334268 108180
rect 352720 101982 352748 141886
rect 353548 107490 353576 141886
rect 354916 132304 354968 132310
rect 354916 132246 354968 132252
rect 354928 117146 354956 132246
rect 354916 117140 354968 117146
rect 354916 117082 354968 117088
rect 353536 107484 353588 107490
rect 353536 107426 353588 107432
rect 352798 105208 352854 105217
rect 352798 105143 352854 105152
rect 352708 101976 352760 101982
rect 352708 101918 352760 101924
rect 334214 95552 334270 95561
rect 334214 95487 334270 95496
rect 330076 94700 330128 94706
rect 330076 94642 330128 94648
rect 326672 94428 326724 94434
rect 326672 94370 326724 94376
rect 326580 87492 326632 87498
rect 326580 87434 326632 87440
rect 326684 85798 326712 94370
rect 327224 87492 327276 87498
rect 327224 87434 327276 87440
rect 326672 85792 326724 85798
rect 326672 85734 326724 85740
rect 327038 73928 327094 73937
rect 327038 73863 327094 73872
rect 326854 71072 326910 71081
rect 326854 71007 326910 71016
rect 326868 65738 326896 71007
rect 326946 69576 327002 69585
rect 326946 69511 327002 69520
rect 326960 65874 326988 69511
rect 327052 68594 327080 73863
rect 327130 71480 327186 71489
rect 327130 71415 327186 71424
rect 327040 68588 327092 68594
rect 327040 68530 327092 68536
rect 327038 68352 327094 68361
rect 327038 68287 327094 68296
rect 326948 65868 327000 65874
rect 326948 65810 327000 65816
rect 326856 65732 326908 65738
rect 326856 65674 326908 65680
rect 327052 64786 327080 68287
rect 327144 67234 327172 71415
rect 327132 67228 327184 67234
rect 327132 67170 327184 67176
rect 327040 64780 327092 64786
rect 327040 64722 327092 64728
rect 327236 50234 327264 87434
rect 328420 76408 328472 76414
rect 328420 76350 328472 76356
rect 328432 75297 328460 76350
rect 330088 75954 330116 94642
rect 334228 94434 334256 95487
rect 334216 94428 334268 94434
rect 334216 94370 334268 94376
rect 337324 88846 337660 88874
rect 338152 88846 338304 88874
rect 338980 88846 339592 88874
rect 339808 88846 340144 88874
rect 340636 88846 340972 88874
rect 341464 88846 341708 88874
rect 342292 88846 342444 88874
rect 343212 88846 343548 88874
rect 344040 88846 344376 88874
rect 344868 88846 345020 88874
rect 334124 87084 334176 87090
rect 334124 87026 334176 87032
rect 332744 86812 332796 86818
rect 332744 86754 332796 86760
rect 330088 75926 330852 75954
rect 330824 75682 330852 75926
rect 332756 75818 332784 86754
rect 334136 79202 334164 87026
rect 335412 86948 335464 86954
rect 335412 86890 335464 86896
rect 335424 79202 335452 86890
rect 335504 86880 335556 86886
rect 335504 86822 335556 86828
rect 333388 79196 333440 79202
rect 333388 79138 333440 79144
rect 334124 79196 334176 79202
rect 334124 79138 334176 79144
rect 334400 79196 334452 79202
rect 334400 79138 334452 79144
rect 335412 79196 335464 79202
rect 335412 79138 335464 79144
rect 332402 75790 332784 75818
rect 333400 75804 333428 79138
rect 334412 75804 334440 79138
rect 335516 75804 335544 86822
rect 336884 86676 336936 86682
rect 336884 86618 336936 86624
rect 336896 75818 336924 86618
rect 337632 86206 337660 88846
rect 338080 87152 338132 87158
rect 338080 87094 338132 87100
rect 337620 86200 337672 86206
rect 337620 86142 337672 86148
rect 338092 85202 338120 87094
rect 338276 86138 338304 88846
rect 339092 86200 339144 86206
rect 339092 86142 339144 86148
rect 338264 86132 338316 86138
rect 338264 86074 338316 86080
rect 339000 86132 339052 86138
rect 339000 86074 339052 86080
rect 338092 85174 338304 85202
rect 338276 79066 338304 85174
rect 339012 79134 339040 86074
rect 339000 79128 339052 79134
rect 339000 79070 339052 79076
rect 337528 79060 337580 79066
rect 337528 79002 337580 79008
rect 338264 79060 338316 79066
rect 338264 79002 338316 79008
rect 336542 75790 336924 75818
rect 337540 75804 337568 79002
rect 339104 78794 339132 86142
rect 339564 79202 339592 88846
rect 339644 87016 339696 87022
rect 339644 86958 339696 86964
rect 339552 79196 339604 79202
rect 339552 79138 339604 79144
rect 339092 78788 339144 78794
rect 339092 78730 339144 78736
rect 338540 78516 338592 78522
rect 338540 78458 338592 78464
rect 338552 75804 338580 78458
rect 339656 75804 339684 86958
rect 340116 86206 340144 88846
rect 340104 86200 340156 86206
rect 340104 86142 340156 86148
rect 340944 86138 340972 88846
rect 341024 87288 341076 87294
rect 341024 87230 341076 87236
rect 340932 86132 340984 86138
rect 340932 86074 340984 86080
rect 341036 75818 341064 87230
rect 341680 86274 341708 88846
rect 341668 86268 341720 86274
rect 341668 86210 341720 86216
rect 342416 86206 342444 88846
rect 341760 86200 341812 86206
rect 341760 86142 341812 86148
rect 342404 86200 342456 86206
rect 342404 86142 342456 86148
rect 341772 78998 341800 86142
rect 343520 86138 343548 88846
rect 344348 87226 344376 88846
rect 344992 87362 345020 88846
rect 345452 88846 345696 88874
rect 346188 88846 346524 88874
rect 347016 88846 347352 88874
rect 348028 88846 348272 88874
rect 348764 88846 349100 88874
rect 349592 88846 349928 88874
rect 350052 88846 350756 88874
rect 351248 88846 351584 88874
rect 352168 88846 352412 88874
rect 344980 87356 345032 87362
rect 344980 87298 345032 87304
rect 344336 87220 344388 87226
rect 344336 87162 344388 87168
rect 345452 86818 345480 88846
rect 346188 87090 346216 88846
rect 346176 87084 346228 87090
rect 346176 87026 346228 87032
rect 345440 86812 345492 86818
rect 345440 86754 345492 86760
rect 347016 86750 347044 88846
rect 347280 87220 347332 87226
rect 347280 87162 347332 87168
rect 347004 86744 347056 86750
rect 347004 86686 347056 86692
rect 344612 86268 344664 86274
rect 344612 86210 344664 86216
rect 341852 86132 341904 86138
rect 341852 86074 341904 86080
rect 343508 86132 343560 86138
rect 343508 86074 343560 86080
rect 344520 86132 344572 86138
rect 344520 86074 344572 86080
rect 341864 79066 341892 86074
rect 343784 79196 343836 79202
rect 343784 79138 343836 79144
rect 342680 79128 342732 79134
rect 342680 79070 342732 79076
rect 341852 79060 341904 79066
rect 341852 79002 341904 79008
rect 341760 78992 341812 78998
rect 341760 78934 341812 78940
rect 341668 78788 341720 78794
rect 341668 78730 341720 78736
rect 340682 75790 341064 75818
rect 341680 75804 341708 78730
rect 342692 75804 342720 79070
rect 343796 75804 343824 79138
rect 344532 78590 344560 86074
rect 344624 79134 344652 86210
rect 344704 86200 344756 86206
rect 344704 86142 344756 86148
rect 344716 79202 344744 86142
rect 347292 79202 347320 87162
rect 348028 86886 348056 88846
rect 348764 87022 348792 88846
rect 349592 87158 349620 88846
rect 349580 87152 349632 87158
rect 349580 87094 349632 87100
rect 348752 87016 348804 87022
rect 348752 86958 348804 86964
rect 348016 86880 348068 86886
rect 348016 86822 348068 86828
rect 350052 86154 350080 88846
rect 351248 86954 351276 88846
rect 352168 87294 352196 88846
rect 352156 87288 352208 87294
rect 352156 87230 352208 87236
rect 351236 86948 351288 86954
rect 351236 86890 351288 86896
rect 349500 86126 350080 86154
rect 344704 79196 344756 79202
rect 344704 79138 344756 79144
rect 347280 79196 347332 79202
rect 347280 79138 347332 79144
rect 344612 79128 344664 79134
rect 344612 79070 344664 79076
rect 346820 79128 346872 79134
rect 346820 79070 346872 79076
rect 347924 79128 347976 79134
rect 347924 79070 347976 79076
rect 345808 79060 345860 79066
rect 345808 79002 345860 79008
rect 344796 78992 344848 78998
rect 344796 78934 344848 78940
rect 344520 78584 344572 78590
rect 344520 78526 344572 78532
rect 344808 75804 344836 78934
rect 345820 75804 345848 79002
rect 346832 75804 346860 79070
rect 347936 75804 347964 79070
rect 348936 78584 348988 78590
rect 348936 78526 348988 78532
rect 348948 75804 348976 78526
rect 349500 78522 349528 86126
rect 349948 79196 350000 79202
rect 349948 79138 350000 79144
rect 349488 78516 349540 78522
rect 349488 78458 349540 78464
rect 349960 75804 349988 79138
rect 350958 77872 351014 77881
rect 350958 77807 351014 77816
rect 352062 77872 352118 77881
rect 352062 77807 352118 77816
rect 350972 75804 351000 77807
rect 352076 75804 352104 77807
rect 352720 75818 352748 101918
rect 352812 97834 352840 105143
rect 352800 97828 352852 97834
rect 352800 97770 352852 97776
rect 352812 97601 352840 97770
rect 352798 97592 352854 97601
rect 352798 97527 352854 97536
rect 352800 92320 352852 92326
rect 352800 92262 352852 92268
rect 352812 90121 352840 92262
rect 352798 90112 352854 90121
rect 352798 90047 352854 90056
rect 352720 75790 353102 75818
rect 353548 75682 353576 107426
rect 354928 84098 354956 117082
rect 355020 112998 355048 141886
rect 355848 132310 355876 141886
rect 355836 132304 355888 132310
rect 355836 132246 355888 132252
rect 356202 126288 356258 126297
rect 356202 126223 356258 126232
rect 356216 126122 356244 126223
rect 356204 126116 356256 126122
rect 356204 126058 356256 126064
rect 356308 122654 356336 141886
rect 357688 126802 357716 141886
rect 357676 126796 357728 126802
rect 357676 126738 357728 126744
rect 356296 122648 356348 122654
rect 356296 122590 356348 122596
rect 356202 121256 356258 121265
rect 356202 121191 356258 121200
rect 356216 120614 356244 121191
rect 356204 120608 356256 120614
rect 356204 120550 356256 120556
rect 356202 116224 356258 116233
rect 356202 116159 356258 116168
rect 356216 115106 356244 116159
rect 356204 115100 356256 115106
rect 356204 115042 356256 115048
rect 355008 112992 355060 112998
rect 355008 112934 355060 112940
rect 354916 84092 354968 84098
rect 354916 84034 354968 84040
rect 355020 75818 355048 112934
rect 356202 111328 356258 111337
rect 356202 111263 356258 111272
rect 356216 110958 356244 111263
rect 356204 110952 356256 110958
rect 356204 110894 356256 110900
rect 356202 106296 356258 106305
rect 356202 106231 356258 106240
rect 356216 105450 356244 106231
rect 356204 105444 356256 105450
rect 356204 105386 356256 105392
rect 356202 101264 356258 101273
rect 356202 101199 356258 101208
rect 356216 100622 356244 101199
rect 356204 100616 356256 100622
rect 356204 100558 356256 100564
rect 356202 96232 356258 96241
rect 356202 96167 356258 96176
rect 356216 95794 356244 96167
rect 356204 95788 356256 95794
rect 356204 95730 356256 95736
rect 356202 91336 356258 91345
rect 356202 91271 356258 91280
rect 356216 90218 356244 91271
rect 356204 90212 356256 90218
rect 356204 90154 356256 90160
rect 355836 84092 355888 84098
rect 355836 84034 355888 84040
rect 355848 75818 355876 84034
rect 355020 75790 355126 75818
rect 355848 75790 356230 75818
rect 356308 75682 356336 122590
rect 357688 75682 357716 126738
rect 330824 75654 331390 75682
rect 353548 75654 354114 75682
rect 356308 75654 357242 75682
rect 357688 75654 358254 75682
rect 328418 75288 328474 75297
rect 328418 75223 328474 75232
rect 327866 72568 327922 72577
rect 327866 72503 327922 72512
rect 327880 68390 327908 72503
rect 327868 68384 327920 68390
rect 327868 68326 327920 68332
rect 327682 67264 327738 67273
rect 327682 67199 327738 67208
rect 327696 65126 327724 67199
rect 328418 66992 328474 67001
rect 328418 66927 328474 66936
rect 328432 66894 328460 66927
rect 328420 66888 328472 66894
rect 328420 66830 328472 66836
rect 328418 65904 328474 65913
rect 328418 65839 328474 65848
rect 328432 65466 328460 65839
rect 328420 65460 328472 65466
rect 328420 65402 328472 65408
rect 327684 65120 327736 65126
rect 327684 65062 327736 65068
rect 327314 64544 327370 64553
rect 327314 64479 327370 64488
rect 327328 62406 327356 64479
rect 328050 63184 328106 63193
rect 328050 63119 328106 63128
rect 327316 62400 327368 62406
rect 327316 62342 327368 62348
rect 328064 61046 328092 63119
rect 328326 62776 328382 62785
rect 328326 62711 328382 62720
rect 328052 61040 328104 61046
rect 328052 60982 328104 60988
rect 328340 58802 328368 62711
rect 328510 61552 328566 61561
rect 328510 61487 328566 61496
rect 328524 61318 328552 61487
rect 328512 61312 328564 61318
rect 328512 61254 328564 61260
rect 328418 60056 328474 60065
rect 328418 59991 328474 60000
rect 328328 58796 328380 58802
rect 328328 58738 328380 58744
rect 327682 58696 327738 58705
rect 327682 58631 327738 58640
rect 327696 56354 327724 58631
rect 328432 57238 328460 59991
rect 328510 58968 328566 58977
rect 328510 58903 328566 58912
rect 328420 57232 328472 57238
rect 328326 57200 328382 57209
rect 328420 57174 328472 57180
rect 328326 57135 328382 57144
rect 327684 56348 327736 56354
rect 327684 56290 327736 56296
rect 327498 56248 327554 56257
rect 327498 56183 327554 56192
rect 327512 55810 327540 56183
rect 327500 55804 327552 55810
rect 327500 55746 327552 55752
rect 328340 54994 328368 57135
rect 328524 56082 328552 58903
rect 328512 56076 328564 56082
rect 328512 56018 328564 56024
rect 328510 55296 328566 55305
rect 328510 55231 328566 55240
rect 328524 55062 328552 55231
rect 358516 55062 358544 388674
rect 362460 388460 362512 388466
rect 362460 388402 362512 388408
rect 360802 262288 360858 262297
rect 360802 262223 360858 262232
rect 360816 262054 360844 262223
rect 360436 262048 360488 262054
rect 360436 261990 360488 261996
rect 360804 262048 360856 262054
rect 360804 261990 360856 261996
rect 360448 227714 360476 261990
rect 360528 259328 360580 259334
rect 360528 259270 360580 259276
rect 360540 259169 360568 259270
rect 360526 259160 360582 259169
rect 360526 259095 360582 259104
rect 360540 234446 360568 259095
rect 360620 257220 360672 257226
rect 360620 257162 360672 257168
rect 360632 256041 360660 257162
rect 360618 256032 360674 256041
rect 360618 255967 360674 255976
rect 361172 253072 361224 253078
rect 361172 253014 361224 253020
rect 361184 252913 361212 253014
rect 361170 252904 361226 252913
rect 361170 252839 361226 252848
rect 361448 250284 361500 250290
rect 361448 250226 361500 250232
rect 361460 249785 361488 250226
rect 361446 249776 361502 249785
rect 361446 249711 361502 249720
rect 360710 246648 360766 246657
rect 360710 246583 360766 246592
rect 360618 243520 360674 243529
rect 360618 243455 360674 243464
rect 360528 234440 360580 234446
rect 360528 234382 360580 234388
rect 360436 227708 360488 227714
rect 360436 227650 360488 227656
rect 360632 224790 360660 243455
rect 360724 231726 360752 246583
rect 360802 240392 360858 240401
rect 360802 240327 360858 240336
rect 360712 231720 360764 231726
rect 360712 231662 360764 231668
rect 360816 230298 360844 240327
rect 361170 237400 361226 237409
rect 361170 237335 361226 237344
rect 360804 230292 360856 230298
rect 360804 230234 360856 230240
rect 360620 224784 360672 224790
rect 360620 224726 360672 224732
rect 361080 221520 361132 221526
rect 361080 221462 361132 221468
rect 359700 220024 359752 220030
rect 359700 219966 359752 219972
rect 359712 181338 359740 219966
rect 359700 181332 359752 181338
rect 359700 181274 359752 181280
rect 360434 168312 360490 168321
rect 360434 168247 360490 168256
rect 360448 142034 360476 168247
rect 360526 165184 360582 165193
rect 360526 165119 360582 165128
rect 360436 142028 360488 142034
rect 360436 141970 360488 141976
rect 360540 133806 360568 165119
rect 360618 162056 360674 162065
rect 360618 161991 360674 162000
rect 360632 135098 360660 161991
rect 360710 158928 360766 158937
rect 360710 158863 360766 158872
rect 360620 135092 360672 135098
rect 360620 135034 360672 135040
rect 360724 134418 360752 158863
rect 360894 155800 360950 155809
rect 360894 155735 360950 155744
rect 360802 152672 360858 152681
rect 360802 152607 360858 152616
rect 360712 134412 360764 134418
rect 360712 134354 360764 134360
rect 360528 133800 360580 133806
rect 360528 133742 360580 133748
rect 360816 132378 360844 152607
rect 360908 137886 360936 155735
rect 360986 149544 361042 149553
rect 360986 149479 361042 149488
rect 360896 137880 360948 137886
rect 360896 137822 360948 137828
rect 361000 133738 361028 149479
rect 361092 143433 361120 221462
rect 361184 214318 361212 237335
rect 361172 214312 361224 214318
rect 361172 214254 361224 214260
rect 361170 168312 361226 168321
rect 361170 168247 361226 168256
rect 361184 168214 361212 168247
rect 361172 168208 361224 168214
rect 361172 168150 361224 168156
rect 361724 165488 361776 165494
rect 361724 165430 361776 165436
rect 361736 165193 361764 165430
rect 361722 165184 361778 165193
rect 361722 165119 361778 165128
rect 361724 162700 361776 162706
rect 361724 162642 361776 162648
rect 361736 162065 361764 162642
rect 361722 162056 361778 162065
rect 361722 161991 361778 162000
rect 361722 158928 361778 158937
rect 361722 158863 361778 158872
rect 361736 158558 361764 158863
rect 361724 158552 361776 158558
rect 361724 158494 361776 158500
rect 361722 155800 361778 155809
rect 361722 155735 361724 155744
rect 361776 155735 361778 155744
rect 361724 155706 361776 155712
rect 361170 146416 361226 146425
rect 361170 146351 361226 146360
rect 361078 143424 361134 143433
rect 361078 143359 361134 143368
rect 361080 142028 361132 142034
rect 361080 141970 361132 141976
rect 360988 133732 361040 133738
rect 360988 133674 361040 133680
rect 360804 132372 360856 132378
rect 360804 132314 360856 132320
rect 361092 131698 361120 141970
rect 360436 131692 360488 131698
rect 360436 131634 360488 131640
rect 361080 131692 361132 131698
rect 361080 131634 361132 131640
rect 360448 119882 360476 131634
rect 361184 130950 361212 146351
rect 361172 130944 361224 130950
rect 361172 130886 361224 130892
rect 360620 124824 360672 124830
rect 360620 124766 360672 124772
rect 360356 119854 360476 119882
rect 360356 117894 360384 119854
rect 360632 117894 360660 124766
rect 360344 117888 360396 117894
rect 360344 117830 360396 117836
rect 360436 117888 360488 117894
rect 360436 117830 360488 117836
rect 360620 117888 360672 117894
rect 360620 117830 360672 117836
rect 360252 117820 360304 117826
rect 360252 117762 360304 117768
rect 360264 98530 360292 117762
rect 360264 98502 360384 98530
rect 360356 88874 360384 98502
rect 360172 88846 360384 88874
rect 360172 87430 360200 88846
rect 359700 87424 359752 87430
rect 359700 87366 359752 87372
rect 360160 87424 360212 87430
rect 360448 87401 360476 117830
rect 360160 87366 360212 87372
rect 360434 87392 360490 87401
rect 328512 55056 328564 55062
rect 328512 54998 328564 55004
rect 358504 55056 358556 55062
rect 358504 54998 358556 55004
rect 328328 54988 328380 54994
rect 328328 54930 328380 54936
rect 328418 54480 328474 54489
rect 328418 54415 328420 54424
rect 328472 54415 328474 54424
rect 328420 54386 328472 54392
rect 328420 53696 328472 53702
rect 328420 53638 328472 53644
rect 328432 53537 328460 53638
rect 328418 53528 328474 53537
rect 328418 53463 328474 53472
rect 327682 50944 327738 50953
rect 327682 50879 327738 50888
rect 327696 50370 327724 50879
rect 328418 50400 328474 50409
rect 327684 50364 327736 50370
rect 328418 50335 328474 50344
rect 327684 50306 327736 50312
rect 328432 50302 328460 50335
rect 328420 50296 328472 50302
rect 328420 50238 328472 50244
rect 327224 50228 327276 50234
rect 327224 50170 327276 50176
rect 327236 50001 327264 50170
rect 327222 49992 327278 50001
rect 327222 49927 327278 49936
rect 328510 49040 328566 49049
rect 328510 48975 328566 48984
rect 328524 48942 328552 48975
rect 359712 48942 359740 87366
rect 360434 87327 360490 87336
rect 328512 48936 328564 48942
rect 328512 48878 328564 48884
rect 359700 48936 359752 48942
rect 359700 48878 359752 48884
rect 357150 48194 357348 48210
rect 357150 48188 357360 48194
rect 357150 48182 357308 48188
rect 357308 48130 357360 48136
rect 328050 47952 328106 47961
rect 328050 47887 328106 47896
rect 328064 47514 328092 47887
rect 328052 47508 328104 47514
rect 328052 47450 328104 47456
rect 332664 45814 332692 47924
rect 336160 45882 336188 47924
rect 339656 47378 339684 47924
rect 339644 47372 339696 47378
rect 339644 47314 339696 47320
rect 338356 45944 338408 45950
rect 338356 45886 338408 45892
rect 336148 45876 336200 45882
rect 336148 45818 336200 45824
rect 332652 45808 332704 45814
rect 332652 45750 332704 45756
rect 338368 45377 338396 45886
rect 339656 45474 339684 47314
rect 343152 45950 343180 47924
rect 346648 46057 346676 47924
rect 346634 46048 346690 46057
rect 346634 45983 346690 45992
rect 350144 45950 350172 47924
rect 353640 47446 353668 47924
rect 353628 47440 353680 47446
rect 353628 47382 353680 47388
rect 343140 45944 343192 45950
rect 343140 45886 343192 45892
rect 350132 45944 350184 45950
rect 350132 45886 350184 45892
rect 339644 45468 339696 45474
rect 339644 45410 339696 45416
rect 350144 45406 350172 45886
rect 350776 45468 350828 45474
rect 350776 45410 350828 45416
rect 350132 45400 350184 45406
rect 338354 45368 338410 45377
rect 350132 45342 350184 45348
rect 338354 45303 338410 45312
rect 325292 12420 325344 12426
rect 325292 12362 325344 12368
rect 324568 12142 325516 12170
rect 325488 9304 325516 12142
rect 338368 9304 338396 45303
rect 350788 9434 350816 45410
rect 362472 12358 362500 388402
rect 363840 326920 363892 326926
rect 363840 326862 363892 326868
rect 363852 235126 363880 326862
rect 365312 274492 365364 274498
rect 365312 274434 365364 274440
rect 363840 235120 363892 235126
rect 363840 235062 363892 235068
rect 363840 222948 363892 222954
rect 363840 222890 363892 222896
rect 363852 87362 363880 222890
rect 365220 218732 365272 218738
rect 365220 218674 365272 218680
rect 365232 138770 365260 218674
rect 365324 213978 365352 274434
rect 368636 239954 368664 396206
rect 395132 395198 395160 396206
rect 395120 395192 395172 395198
rect 395120 395134 395172 395140
rect 421628 393158 421656 396344
rect 421616 393152 421668 393158
rect 421616 393094 421668 393100
rect 429434 390672 429490 390681
rect 429434 390607 429490 390616
rect 429448 389758 429476 390607
rect 429436 389752 429488 389758
rect 429436 389694 429488 389700
rect 395212 385604 395264 385610
rect 395212 385546 395264 385552
rect 395224 378690 395252 385546
rect 395224 378662 395344 378690
rect 395316 366366 395344 378662
rect 429436 378668 429488 378674
rect 429436 378610 429488 378616
rect 429448 378577 429476 378610
rect 429434 378568 429490 378577
rect 429434 378503 429490 378512
rect 429436 367584 429488 367590
rect 429436 367526 429488 367532
rect 429448 366473 429476 367526
rect 429434 366464 429490 366473
rect 429434 366399 429490 366408
rect 395304 366360 395356 366366
rect 395304 366302 395356 366308
rect 395212 365000 395264 365006
rect 395264 364948 395344 364954
rect 395212 364942 395344 364948
rect 395224 364926 395344 364942
rect 395316 363510 395344 364926
rect 395304 363504 395356 363510
rect 395304 363446 395356 363452
rect 429434 354360 429490 354369
rect 429434 354295 429490 354304
rect 429448 353922 429476 354295
rect 390704 353916 390756 353922
rect 390704 353858 390756 353864
rect 429436 353916 429488 353922
rect 429436 353858 429488 353864
rect 369912 274492 369964 274498
rect 369912 274434 369964 274440
rect 369544 263408 369596 263414
rect 369544 263350 369596 263356
rect 368624 239948 368676 239954
rect 368624 239890 368676 239896
rect 369174 236584 369230 236593
rect 369174 236519 369230 236528
rect 368716 235120 368768 235126
rect 368716 235062 368768 235068
rect 368728 234145 368756 235062
rect 368714 234136 368770 234145
rect 368714 234071 368770 234080
rect 368900 233760 368952 233766
rect 368714 233728 368770 233737
rect 368900 233702 368952 233708
rect 368714 233663 368716 233672
rect 368768 233663 368770 233672
rect 368716 233634 368768 233640
rect 368808 233624 368860 233630
rect 368808 233566 368860 233572
rect 368820 233465 368848 233566
rect 368806 233456 368862 233465
rect 368806 233391 368862 233400
rect 368912 233057 368940 233702
rect 368898 233048 368954 233057
rect 368898 232983 368954 232992
rect 368900 232400 368952 232406
rect 368900 232342 368952 232348
rect 368716 232332 368768 232338
rect 368716 232274 368768 232280
rect 368728 232241 368756 232274
rect 368808 232264 368860 232270
rect 368714 232232 368770 232241
rect 368808 232206 368860 232212
rect 368714 232167 368770 232176
rect 368820 231833 368848 232206
rect 368806 231824 368862 231833
rect 368806 231759 368862 231768
rect 368912 231425 368940 232342
rect 368898 231416 368954 231425
rect 368898 231351 368954 231360
rect 368806 231008 368862 231017
rect 368806 230943 368862 230952
rect 368900 230972 368952 230978
rect 368716 230904 368768 230910
rect 368716 230846 368768 230852
rect 368728 230609 368756 230846
rect 368820 230842 368848 230943
rect 368900 230914 368952 230920
rect 368808 230836 368860 230842
rect 368808 230778 368860 230784
rect 368714 230600 368770 230609
rect 368714 230535 368770 230544
rect 368912 230201 368940 230914
rect 368898 230192 368954 230201
rect 368898 230127 368954 230136
rect 368716 229612 368768 229618
rect 368716 229554 368768 229560
rect 368728 229521 368756 229554
rect 368714 229512 368770 229521
rect 368714 229447 368770 229456
rect 368806 229104 368862 229113
rect 368806 229039 368862 229048
rect 368714 228696 368770 228705
rect 368714 228631 368770 228640
rect 368728 228462 368756 228631
rect 368716 228456 368768 228462
rect 368716 228398 368768 228404
rect 368820 228394 368848 229039
rect 368808 228388 368860 228394
rect 368808 228330 368860 228336
rect 368716 228320 368768 228326
rect 368714 228288 368716 228297
rect 368768 228288 368770 228297
rect 368714 228223 368770 228232
rect 369084 227572 369136 227578
rect 369084 227514 369136 227520
rect 368806 227472 368862 227481
rect 368806 227407 368862 227416
rect 368714 227064 368770 227073
rect 368714 226999 368770 227008
rect 368728 226898 368756 226999
rect 368820 226966 368848 227407
rect 368808 226960 368860 226966
rect 368808 226902 368860 226908
rect 368716 226892 368768 226898
rect 368716 226834 368768 226840
rect 368990 226520 369046 226529
rect 368990 226455 369046 226464
rect 368898 226384 368954 226393
rect 368898 226319 368954 226328
rect 368806 225976 368862 225985
rect 368806 225911 368862 225920
rect 368820 225674 368848 225911
rect 368808 225668 368860 225674
rect 368808 225610 368860 225616
rect 368716 225600 368768 225606
rect 368714 225568 368716 225577
rect 368768 225568 368770 225577
rect 368912 225538 368940 226319
rect 368714 225503 368770 225512
rect 368900 225532 368952 225538
rect 368900 225474 368952 225480
rect 368716 225328 368768 225334
rect 368716 225270 368768 225276
rect 368728 224761 368756 225270
rect 368806 225160 368862 225169
rect 368806 225095 368862 225104
rect 368714 224752 368770 224761
rect 368714 224687 368770 224696
rect 368820 224178 368848 225095
rect 368808 224172 368860 224178
rect 368808 224114 368860 224120
rect 368806 223936 368862 223945
rect 368806 223871 368862 223880
rect 368714 223256 368770 223265
rect 368714 223191 368770 223200
rect 368728 222886 368756 223191
rect 368716 222880 368768 222886
rect 368716 222822 368768 222828
rect 368820 222818 368848 223871
rect 369004 223650 369032 226455
rect 369096 223770 369124 227514
rect 369084 223764 369136 223770
rect 369084 223706 369136 223712
rect 369004 223622 369124 223650
rect 368990 223528 369046 223537
rect 368990 223463 369046 223472
rect 368900 222948 368952 222954
rect 368900 222890 368952 222896
rect 368912 222857 368940 222890
rect 368898 222848 368954 222857
rect 368808 222812 368860 222818
rect 368898 222783 368954 222792
rect 368808 222754 368860 222760
rect 368806 222440 368862 222449
rect 368806 222375 368862 222384
rect 368714 221624 368770 221633
rect 368714 221559 368770 221568
rect 368728 221390 368756 221559
rect 368820 221458 368848 222375
rect 368898 222032 368954 222041
rect 368898 221967 368954 221976
rect 368912 221526 368940 221967
rect 368900 221520 368952 221526
rect 368900 221462 368952 221468
rect 368808 221452 368860 221458
rect 368808 221394 368860 221400
rect 368716 221384 368768 221390
rect 368716 221326 368768 221332
rect 368898 221216 368954 221225
rect 368898 221151 368954 221160
rect 368806 220808 368862 220817
rect 368806 220743 368862 220752
rect 368820 220574 368848 220743
rect 368808 220568 368860 220574
rect 368808 220510 368860 220516
rect 368716 220500 368768 220506
rect 368716 220442 368768 220448
rect 368728 220409 368756 220442
rect 368714 220400 368770 220409
rect 368714 220335 368770 220344
rect 368912 220030 368940 221151
rect 368900 220024 368952 220030
rect 368900 219966 368952 219972
rect 368714 219720 368770 219729
rect 368714 219655 368770 219664
rect 368728 218670 368756 219655
rect 368900 219412 368952 219418
rect 368900 219354 368952 219360
rect 368806 218904 368862 218913
rect 368806 218839 368862 218848
rect 368820 218738 368848 218839
rect 368808 218732 368860 218738
rect 368808 218674 368860 218680
rect 368716 218664 368768 218670
rect 368716 218606 368768 218612
rect 368808 218528 368860 218534
rect 368808 218470 368860 218476
rect 368714 218088 368770 218097
rect 368714 218023 368770 218032
rect 368728 217242 368756 218023
rect 368820 217281 368848 218470
rect 368806 217272 368862 217281
rect 368716 217236 368768 217242
rect 368806 217207 368862 217216
rect 368716 217178 368768 217184
rect 368808 217168 368860 217174
rect 368808 217110 368860 217116
rect 368716 217100 368768 217106
rect 368716 217042 368768 217048
rect 368728 216465 368756 217042
rect 368714 216456 368770 216465
rect 368714 216391 368770 216400
rect 368820 216193 368848 217110
rect 368806 216184 368862 216193
rect 368806 216119 368862 216128
rect 368714 215776 368770 215785
rect 368714 215711 368716 215720
rect 368768 215711 368770 215720
rect 368716 215682 368768 215688
rect 368808 215672 368860 215678
rect 368808 215614 368860 215620
rect 368820 214969 368848 215614
rect 368806 214960 368862 214969
rect 368806 214895 368862 214904
rect 368912 214810 368940 219354
rect 369004 219010 369032 223463
rect 369096 219486 369124 223622
rect 369084 219480 369136 219486
rect 369084 219422 369136 219428
rect 369082 219312 369138 219321
rect 369188 219298 369216 236519
rect 369450 236176 369506 236185
rect 369450 236111 369506 236120
rect 369266 224344 369322 224353
rect 369266 224279 369322 224288
rect 369280 219418 369308 224279
rect 369360 223764 369412 223770
rect 369360 223706 369412 223712
rect 369372 219418 369400 223706
rect 369268 219412 369320 219418
rect 369268 219354 369320 219360
rect 369360 219412 369412 219418
rect 369360 219354 369412 219360
rect 369188 219270 369400 219298
rect 369082 219247 369138 219256
rect 368992 219004 369044 219010
rect 368992 218946 369044 218952
rect 368990 217680 369046 217689
rect 368990 217615 369046 217624
rect 369004 216601 369032 217615
rect 369096 217009 369124 219247
rect 369176 219004 369228 219010
rect 369176 218946 369228 218952
rect 369082 217000 369138 217009
rect 369082 216935 369138 216944
rect 369084 216896 369136 216902
rect 369082 216864 369084 216873
rect 369136 216864 369138 216873
rect 369082 216799 369138 216808
rect 369084 216760 369136 216766
rect 369084 216702 369136 216708
rect 368990 216592 369046 216601
rect 368990 216527 369046 216536
rect 368992 215808 369044 215814
rect 368992 215750 369044 215756
rect 368820 214782 368940 214810
rect 368716 214448 368768 214454
rect 368716 214390 368768 214396
rect 365312 213972 365364 213978
rect 365312 213914 365364 213920
rect 368728 213745 368756 214390
rect 368714 213736 368770 213745
rect 368714 213671 368770 213680
rect 368716 213088 368768 213094
rect 368714 213056 368716 213065
rect 368768 213056 368770 213065
rect 368714 212991 368770 213000
rect 365220 138764 365272 138770
rect 365220 138706 365272 138712
rect 368820 131290 368848 214782
rect 369004 214561 369032 215750
rect 369096 215377 369124 216702
rect 369082 215368 369138 215377
rect 369082 215303 369138 215312
rect 368990 214552 369046 214561
rect 368990 214487 369046 214496
rect 368992 214448 369044 214454
rect 368992 214390 369044 214396
rect 368900 214312 368952 214318
rect 368900 214254 368952 214260
rect 368912 214153 368940 214254
rect 368898 214144 368954 214153
rect 368898 214079 368954 214088
rect 368900 213972 368952 213978
rect 368900 213914 368952 213920
rect 368912 213337 368940 213914
rect 368898 213328 368954 213337
rect 368898 213263 368954 213272
rect 369004 209558 369032 214390
rect 369188 209898 369216 218946
rect 369266 218496 369322 218505
rect 369266 218431 369322 218440
rect 369176 209892 369228 209898
rect 369176 209834 369228 209840
rect 369280 209778 369308 218431
rect 369096 209750 369308 209778
rect 368992 209552 369044 209558
rect 368992 209494 369044 209500
rect 369096 209370 369124 209750
rect 369372 209642 369400 219270
rect 368912 209342 369124 209370
rect 369188 209614 369400 209642
rect 368912 199970 368940 209342
rect 369188 204730 369216 209614
rect 369268 209552 369320 209558
rect 369268 209494 369320 209500
rect 368992 204724 369044 204730
rect 368992 204666 369044 204672
rect 369176 204724 369228 204730
rect 369176 204666 369228 204672
rect 368900 199964 368952 199970
rect 368900 199906 368952 199912
rect 369004 195210 369032 204666
rect 369176 199964 369228 199970
rect 369176 199906 369228 199912
rect 368992 195204 369044 195210
rect 368992 195146 369044 195152
rect 369084 185480 369136 185486
rect 369084 185422 369136 185428
rect 369096 175898 369124 185422
rect 369084 175892 369136 175898
rect 369084 175834 369136 175840
rect 369188 168554 369216 199906
rect 369280 168622 369308 209494
rect 369360 195204 369412 195210
rect 369360 195146 369412 195152
rect 369268 168616 369320 168622
rect 369268 168558 369320 168564
rect 369176 168548 369228 168554
rect 369176 168490 369228 168496
rect 368808 131284 368860 131290
rect 368808 131226 368860 131232
rect 363840 87356 363892 87362
rect 363840 87298 363892 87304
rect 369268 79196 369320 79202
rect 369268 79138 369320 79144
rect 369280 66826 369308 79138
rect 369268 66820 369320 66826
rect 369268 66762 369320 66768
rect 369268 59884 369320 59890
rect 369268 59826 369320 59832
rect 369280 47514 369308 59826
rect 369268 47508 369320 47514
rect 369268 47450 369320 47456
rect 369372 35018 369400 195146
rect 369188 34990 369400 35018
rect 369188 32962 369216 34990
rect 369464 33030 369492 236111
rect 369556 229929 369584 263350
rect 369728 262320 369780 262326
rect 369728 262262 369780 262268
rect 369634 235768 369690 235777
rect 369634 235703 369690 235712
rect 369542 229920 369598 229929
rect 369542 229855 369598 229864
rect 369542 227880 369598 227889
rect 369542 227815 369598 227824
rect 369556 132922 369584 227815
rect 369648 132990 369676 235703
rect 369740 232649 369768 262262
rect 369818 235360 369874 235369
rect 369818 235295 369874 235304
rect 369726 232640 369782 232649
rect 369726 232575 369782 232584
rect 369832 231402 369860 235295
rect 369924 234553 369952 274434
rect 372856 262728 372908 262734
rect 372856 262670 372908 262676
rect 372868 236842 372896 262670
rect 381136 262660 381188 262666
rect 381136 262602 381188 262608
rect 377824 239948 377876 239954
rect 377824 239890 377876 239896
rect 372868 236814 373632 236842
rect 373604 236706 373632 236814
rect 373604 236678 373894 236706
rect 377836 236692 377864 239890
rect 381148 236842 381176 262602
rect 385276 262592 385328 262598
rect 385276 262534 385328 262540
rect 385288 236842 385316 262534
rect 390716 240634 390744 353858
rect 395396 345620 395448 345626
rect 395396 345562 395448 345568
rect 394844 341472 394896 341478
rect 394844 341414 394896 341420
rect 394856 240634 394884 341414
rect 395408 340202 395436 345562
rect 429434 342256 429490 342265
rect 429434 342191 429490 342200
rect 429448 341478 429476 342191
rect 429436 341472 429488 341478
rect 429436 341414 429488 341420
rect 395316 340174 395436 340202
rect 395316 335970 395344 340174
rect 395212 335964 395264 335970
rect 395212 335906 395264 335912
rect 395304 335964 395356 335970
rect 395304 335906 395356 335912
rect 395224 327674 395252 335906
rect 429434 330152 429490 330161
rect 429434 330087 429490 330096
rect 429448 329034 429476 330087
rect 429436 329028 429488 329034
rect 429436 328970 429488 328976
rect 395120 327668 395172 327674
rect 395120 327610 395172 327616
rect 395212 327668 395264 327674
rect 395212 327610 395264 327616
rect 395132 320806 395160 327610
rect 395120 320800 395172 320806
rect 395120 320742 395172 320748
rect 395212 320800 395264 320806
rect 395212 320742 395264 320748
rect 395224 311082 395252 320742
rect 429434 317912 429490 317921
rect 429434 317847 429490 317856
rect 429448 316658 429476 317847
rect 429436 316652 429488 316658
rect 429436 316594 429488 316600
rect 405976 315904 406028 315910
rect 405974 315872 405976 315881
rect 406028 315872 406030 315881
rect 405974 315807 406030 315816
rect 427318 313832 427374 313841
rect 405976 313796 406028 313802
rect 427318 313767 427374 313776
rect 405976 313738 406028 313744
rect 405988 313705 406016 313738
rect 405974 313696 406030 313705
rect 405974 313631 406030 313640
rect 395028 311076 395080 311082
rect 395028 311018 395080 311024
rect 395212 311076 395264 311082
rect 395212 311018 395264 311024
rect 395040 310962 395068 311018
rect 395040 310934 395160 310962
rect 395132 301442 395160 310934
rect 405974 310432 406030 310441
rect 405974 310367 406030 310376
rect 405988 310334 406016 310367
rect 405976 310328 406028 310334
rect 405976 310270 406028 310276
rect 405976 308288 406028 308294
rect 405974 308256 405976 308265
rect 406028 308256 406030 308265
rect 405974 308191 406030 308200
rect 406068 306248 406120 306254
rect 406066 306216 406068 306225
rect 406120 306216 406122 306225
rect 406066 306151 406122 306160
rect 405976 304140 406028 304146
rect 405976 304082 406028 304088
rect 405988 303641 406016 304082
rect 405974 303632 406030 303641
rect 405974 303567 406030 303576
rect 395132 301414 395252 301442
rect 395224 291770 395252 301414
rect 405976 300672 406028 300678
rect 405976 300614 406028 300620
rect 405988 300513 406016 300614
rect 405974 300504 406030 300513
rect 405974 300439 406030 300448
rect 405976 298632 406028 298638
rect 405976 298574 406028 298580
rect 405988 298337 406016 298574
rect 405974 298328 406030 298337
rect 405974 298263 406030 298272
rect 405974 295472 406030 295481
rect 405974 295407 406030 295416
rect 405988 295170 406016 295407
rect 405976 295164 406028 295170
rect 405976 295106 406028 295112
rect 405976 293804 406028 293810
rect 405976 293746 406028 293752
rect 405988 293713 406016 293746
rect 405974 293704 406030 293713
rect 405974 293639 406030 293648
rect 395028 291764 395080 291770
rect 395028 291706 395080 291712
rect 395212 291764 395264 291770
rect 395212 291706 395264 291712
rect 395040 291650 395068 291706
rect 395040 291622 395160 291650
rect 395132 288914 395160 291622
rect 405976 291016 406028 291022
rect 405976 290958 406028 290964
rect 405988 290721 406016 290958
rect 405974 290712 406030 290721
rect 405974 290647 406030 290656
rect 405976 288976 406028 288982
rect 405976 288918 406028 288924
rect 395120 288908 395172 288914
rect 395120 288850 395172 288856
rect 405988 288681 406016 288918
rect 405974 288672 406030 288681
rect 405974 288607 406030 288616
rect 405974 285544 406030 285553
rect 405974 285479 405976 285488
rect 406028 285479 406030 285488
rect 405976 285450 406028 285456
rect 405976 283468 406028 283474
rect 405976 283410 406028 283416
rect 405988 283377 406016 283410
rect 405974 283368 406030 283377
rect 405974 283303 406030 283312
rect 395304 282108 395356 282114
rect 395304 282050 395356 282056
rect 395316 279258 395344 282050
rect 405976 279320 406028 279326
rect 405976 279262 406028 279268
rect 395120 279252 395172 279258
rect 395120 279194 395172 279200
rect 395304 279252 395356 279258
rect 395304 279194 395356 279200
rect 395132 269777 395160 279194
rect 405988 278753 406016 279262
rect 405974 278744 406030 278753
rect 405974 278679 406030 278688
rect 415266 277248 415322 277257
rect 415322 277220 415570 277234
rect 415322 277206 415584 277220
rect 415266 277183 415322 277192
rect 410220 274498 410248 276948
rect 410208 274492 410260 274498
rect 410208 274434 410260 274440
rect 395118 269768 395174 269777
rect 395118 269703 395174 269712
rect 395394 269768 395450 269777
rect 395394 269703 395450 269712
rect 395408 269670 395436 269703
rect 395396 269664 395448 269670
rect 395396 269606 395448 269612
rect 412888 250290 412916 276948
rect 415556 273857 415584 277206
rect 417028 276934 418238 276962
rect 419788 276934 420906 276962
rect 422548 276934 423574 276962
rect 414254 273848 414310 273857
rect 414254 273783 414310 273792
rect 415542 273848 415598 273857
rect 415542 273783 415598 273792
rect 414268 253078 414296 273783
rect 417028 257226 417056 276934
rect 419788 259334 419816 276934
rect 422548 262054 422576 276934
rect 422536 262048 422588 262054
rect 422536 261990 422588 261996
rect 419776 259328 419828 259334
rect 419776 259270 419828 259276
rect 417016 257220 417068 257226
rect 417016 257162 417068 257168
rect 414256 253072 414308 253078
rect 414256 253014 414308 253020
rect 412876 250284 412928 250290
rect 412876 250226 412928 250232
rect 389876 240628 389928 240634
rect 389876 240570 389928 240576
rect 390704 240628 390756 240634
rect 390704 240570 390756 240576
rect 393832 240628 393884 240634
rect 393832 240570 393884 240576
rect 394844 240628 394896 240634
rect 394844 240570 394896 240576
rect 381148 236814 381728 236842
rect 385288 236814 385592 236842
rect 381700 236706 381728 236814
rect 385564 236706 385592 236814
rect 381700 236678 381898 236706
rect 385564 236678 385854 236706
rect 389888 236692 389916 240570
rect 393844 236692 393872 240570
rect 370002 234952 370058 234961
rect 370002 234887 370058 234896
rect 369910 234544 369966 234553
rect 369910 234479 369966 234488
rect 370016 231522 370044 234887
rect 370004 231516 370056 231522
rect 370004 231458 370056 231464
rect 369832 231374 370044 231402
rect 369912 231312 369964 231318
rect 369912 231254 369964 231260
rect 369726 226656 369782 226665
rect 369726 226591 369782 226600
rect 369740 210050 369768 226591
rect 369818 219992 369874 220001
rect 369818 219927 369874 219936
rect 369832 214590 369860 219927
rect 369820 214584 369872 214590
rect 369820 214526 369872 214532
rect 369924 211666 369952 231254
rect 369912 211660 369964 211666
rect 369912 211602 369964 211608
rect 369740 210022 369952 210050
rect 369820 209892 369872 209898
rect 369820 209834 369872 209840
rect 369832 199494 369860 209834
rect 369820 199488 369872 199494
rect 369820 199430 369872 199436
rect 369924 195278 369952 210022
rect 369912 195272 369964 195278
rect 369912 195214 369964 195220
rect 369728 195204 369780 195210
rect 369728 195146 369780 195152
rect 369740 185486 369768 195146
rect 369912 192416 369964 192422
rect 369912 192358 369964 192364
rect 369924 192286 369952 192358
rect 369912 192280 369964 192286
rect 369912 192222 369964 192228
rect 369728 185480 369780 185486
rect 369728 185422 369780 185428
rect 369820 182760 369872 182766
rect 369820 182702 369872 182708
rect 369728 170316 369780 170322
rect 369728 170258 369780 170264
rect 369636 132984 369688 132990
rect 369636 132926 369688 132932
rect 369544 132916 369596 132922
rect 369544 132858 369596 132864
rect 369544 124892 369596 124898
rect 369544 124834 369596 124840
rect 369556 46086 369584 124834
rect 369636 124688 369688 124694
rect 369636 124630 369688 124636
rect 369544 46080 369596 46086
rect 369544 46022 369596 46028
rect 369648 33098 369676 124630
rect 369740 88858 369768 170258
rect 369832 156518 369860 182702
rect 369912 175892 369964 175898
rect 369912 175834 369964 175840
rect 369924 170322 369952 175834
rect 369912 170316 369964 170322
rect 369912 170258 369964 170264
rect 369820 156512 369872 156518
rect 369820 156454 369872 156460
rect 369820 153724 369872 153730
rect 369820 153666 369872 153672
rect 369832 146862 369860 153666
rect 369820 146856 369872 146862
rect 369820 146798 369872 146804
rect 369820 146720 369872 146726
rect 369820 146662 369872 146668
rect 369832 115281 369860 146662
rect 369818 115272 369874 115281
rect 369818 115207 369874 115216
rect 369910 115136 369966 115145
rect 369910 115071 369966 115080
rect 369924 105625 369952 115071
rect 369910 105616 369966 105625
rect 369910 105551 369966 105560
rect 369818 105480 369874 105489
rect 369818 105415 369874 105424
rect 369728 88852 369780 88858
rect 369728 88794 369780 88800
rect 369832 79202 369860 105415
rect 369912 88852 369964 88858
rect 369912 88794 369964 88800
rect 369924 81378 369952 88794
rect 370016 87362 370044 231374
rect 405974 218768 406030 218777
rect 405974 218703 406030 218712
rect 405988 218670 406016 218703
rect 394844 218664 394896 218670
rect 394844 218606 394896 218612
rect 405976 218664 406028 218670
rect 405976 218606 406028 218612
rect 394856 214046 394884 218606
rect 405974 214144 406030 214153
rect 405974 214079 405976 214088
rect 406028 214079 406030 214088
rect 405976 214050 406028 214056
rect 394844 214040 394896 214046
rect 394844 213982 394896 213988
rect 370740 211660 370792 211666
rect 370740 211602 370792 211608
rect 370752 181338 370780 211602
rect 383908 210374 383936 212892
rect 405974 211016 406030 211025
rect 405974 210951 405976 210960
rect 406028 210951 406030 210960
rect 405976 210922 406028 210928
rect 378284 210368 378336 210374
rect 378284 210310 378336 210316
rect 383896 210368 383948 210374
rect 383896 210310 383948 210316
rect 370740 181332 370792 181338
rect 370740 181274 370792 181280
rect 370004 87356 370056 87362
rect 370004 87298 370056 87304
rect 369912 81372 369964 81378
rect 369912 81314 369964 81320
rect 369820 79196 369872 79202
rect 369820 79138 369872 79144
rect 369912 76476 369964 76482
rect 369912 76418 369964 76424
rect 369924 69546 369952 76418
rect 369728 69540 369780 69546
rect 369728 69482 369780 69488
rect 369912 69540 369964 69546
rect 369912 69482 369964 69488
rect 369740 59958 369768 69482
rect 369820 66820 369872 66826
rect 369820 66762 369872 66768
rect 369728 59952 369780 59958
rect 369728 59894 369780 59900
rect 369832 59890 369860 66762
rect 370004 59952 370056 59958
rect 370004 59894 370056 59900
rect 369820 59884 369872 59890
rect 369820 59826 369872 59832
rect 370016 55130 370044 59894
rect 369728 55124 369780 55130
rect 369728 55066 369780 55072
rect 370004 55124 370056 55130
rect 370004 55066 370056 55072
rect 369740 46018 369768 55066
rect 369820 47508 369872 47514
rect 369820 47450 369872 47456
rect 369728 46012 369780 46018
rect 369728 45954 369780 45960
rect 369832 45814 369860 47450
rect 369820 45808 369872 45814
rect 369820 45750 369872 45756
rect 369636 33092 369688 33098
rect 369636 33034 369688 33040
rect 369452 33024 369504 33030
rect 369452 32966 369504 32972
rect 369176 32956 369228 32962
rect 369176 32898 369228 32904
rect 378296 12426 378324 210310
rect 405976 209620 406028 209626
rect 405976 209562 406028 209568
rect 405988 209529 406016 209562
rect 405974 209520 406030 209529
rect 405974 209455 406030 209464
rect 427332 208878 427360 313767
rect 428698 308664 428754 308673
rect 428698 308599 428754 308608
rect 427410 304176 427466 304185
rect 427410 304111 427466 304120
rect 427424 233766 427452 304111
rect 427502 298736 427558 298745
rect 427502 298671 427558 298680
rect 427516 246210 427544 298671
rect 427870 293704 427926 293713
rect 427870 293639 427926 293648
rect 427884 293266 427912 293639
rect 427872 293260 427924 293266
rect 427872 293202 427924 293208
rect 427688 293192 427740 293198
rect 427688 293134 427740 293140
rect 427594 289080 427650 289089
rect 427594 289015 427650 289024
rect 427608 269670 427636 289015
rect 427700 279433 427728 293134
rect 427962 283640 428018 283649
rect 427962 283575 427964 283584
rect 428016 283575 428018 283584
rect 427964 283546 428016 283552
rect 427686 279424 427742 279433
rect 427686 279359 427742 279368
rect 427596 269664 427648 269670
rect 427596 269606 427648 269612
rect 427504 246204 427556 246210
rect 427504 246146 427556 246152
rect 427412 233760 427464 233766
rect 427412 233702 427464 233708
rect 428712 220953 428740 308599
rect 429894 293704 429950 293713
rect 429894 293639 429950 293648
rect 428792 293260 428844 293266
rect 428792 293202 428844 293208
rect 428804 257401 428832 293202
rect 429908 293198 429936 293639
rect 429896 293192 429948 293198
rect 429896 293134 429948 293140
rect 429436 283604 429488 283610
rect 429436 283546 429488 283552
rect 429448 281609 429476 283546
rect 429434 281600 429490 281609
rect 429434 281535 429490 281544
rect 429436 269664 429488 269670
rect 429436 269606 429488 269612
rect 429448 269505 429476 269606
rect 429434 269496 429490 269505
rect 429434 269431 429490 269440
rect 428790 257392 428846 257401
rect 428790 257327 428846 257336
rect 429436 246204 429488 246210
rect 429436 246146 429488 246152
rect 429448 245161 429476 246146
rect 429434 245152 429490 245161
rect 429434 245087 429490 245096
rect 429804 233760 429856 233766
rect 429804 233702 429856 233708
rect 429816 233057 429844 233702
rect 429802 233048 429858 233057
rect 429802 232983 429858 232992
rect 428698 220944 428754 220953
rect 428698 220879 428754 220888
rect 427410 220264 427466 220273
rect 427410 220199 427466 220208
rect 427320 208872 427372 208878
rect 427320 208814 427372 208820
rect 405976 206832 406028 206838
rect 405974 206800 405976 206809
rect 406028 206800 406030 206809
rect 405974 206735 406030 206744
rect 427318 205304 427374 205313
rect 427318 205239 427374 205248
rect 406068 204792 406120 204798
rect 406068 204734 406120 204740
rect 406080 204633 406108 204734
rect 406066 204624 406122 204633
rect 406066 204559 406122 204568
rect 405974 201360 406030 201369
rect 405974 201295 405976 201304
rect 406028 201295 406030 201304
rect 405976 201266 406028 201272
rect 427134 200272 427190 200281
rect 427134 200207 427190 200216
rect 427148 199766 427176 200207
rect 427136 199760 427188 199766
rect 427136 199702 427188 199708
rect 405976 199284 406028 199290
rect 405976 199226 406028 199232
rect 405988 199193 406016 199226
rect 405974 199184 406030 199193
rect 405974 199119 406030 199128
rect 405974 195920 406030 195929
rect 405974 195855 406030 195864
rect 405988 195822 406016 195855
rect 405976 195816 406028 195822
rect 405976 195758 406028 195764
rect 406068 195136 406120 195142
rect 406068 195078 406120 195084
rect 406080 194569 406108 195078
rect 406066 194560 406122 194569
rect 406066 194495 406122 194504
rect 405974 191704 406030 191713
rect 405974 191639 405976 191648
rect 406028 191639 406030 191648
rect 405976 191610 406028 191616
rect 426858 190208 426914 190217
rect 426858 190143 426914 190152
rect 426872 189906 426900 190143
rect 426860 189900 426912 189906
rect 426860 189842 426912 189848
rect 405976 189628 406028 189634
rect 405976 189570 406028 189576
rect 405988 189537 406016 189570
rect 405974 189528 406030 189537
rect 405974 189463 406030 189472
rect 405974 186264 406030 186273
rect 405974 186199 406030 186208
rect 405988 186166 406016 186199
rect 405976 186160 406028 186166
rect 405976 186102 406028 186108
rect 405976 184052 406028 184058
rect 405976 183994 406028 184000
rect 405988 183961 406016 183994
rect 405974 183952 406030 183961
rect 405974 183887 406030 183896
rect 410220 181338 410248 182836
rect 410208 181332 410260 181338
rect 410208 181274 410260 181280
rect 412888 155770 412916 182836
rect 415556 158558 415584 182836
rect 418224 162706 418252 182836
rect 420892 165494 420920 182836
rect 423574 182822 423680 182850
rect 423652 168214 423680 182822
rect 423640 168208 423692 168214
rect 423640 168150 423692 168156
rect 420880 165488 420932 165494
rect 420880 165430 420932 165436
rect 418212 162700 418264 162706
rect 418212 162642 418264 162648
rect 415544 158552 415596 158558
rect 415544 158494 415596 158500
rect 412876 155764 412928 155770
rect 412876 155706 412928 155712
rect 427332 148222 427360 205239
rect 427320 148216 427372 148222
rect 427320 148158 427372 148164
rect 405974 126968 406030 126977
rect 405974 126903 406030 126912
rect 405988 126802 406016 126903
rect 405976 126796 406028 126802
rect 405976 126738 406028 126744
rect 427318 126288 427374 126297
rect 427318 126223 427374 126232
rect 405976 126116 406028 126122
rect 405976 126058 406028 126064
rect 405988 125617 406016 126058
rect 405974 125608 406030 125617
rect 405974 125543 406030 125552
rect 405976 122648 406028 122654
rect 405974 122616 405976 122625
rect 406028 122616 406030 122625
rect 405974 122551 406030 122560
rect 405976 120608 406028 120614
rect 405974 120576 405976 120585
rect 406028 120576 406030 120585
rect 405974 120511 406030 120520
rect 405974 117448 406030 117457
rect 405974 117383 406030 117392
rect 405988 117146 406016 117383
rect 405976 117140 406028 117146
rect 405976 117082 406028 117088
rect 405976 115100 406028 115106
rect 405976 115042 406028 115048
rect 405988 114873 406016 115042
rect 405974 114864 406030 114873
rect 405974 114799 406030 114808
rect 405976 112992 406028 112998
rect 405976 112934 406028 112940
rect 405988 112697 406016 112934
rect 405974 112688 406030 112697
rect 405974 112623 406030 112632
rect 406068 110952 406120 110958
rect 406068 110894 406120 110900
rect 406080 110657 406108 110894
rect 406066 110648 406122 110657
rect 406066 110583 406122 110592
rect 405974 107656 406030 107665
rect 405974 107591 406030 107600
rect 405988 107490 406016 107591
rect 405976 107484 406028 107490
rect 405976 107426 406028 107432
rect 405976 105444 406028 105450
rect 405976 105386 406028 105392
rect 405988 105353 406016 105386
rect 405974 105344 406030 105353
rect 405974 105279 406030 105288
rect 405974 102216 406030 102225
rect 405974 102151 406030 102160
rect 405988 101982 406016 102151
rect 405976 101976 406028 101982
rect 405976 101918 406028 101924
rect 405976 100616 406028 100622
rect 405974 100584 405976 100593
rect 406028 100584 406030 100593
rect 405974 100519 406030 100528
rect 405976 97828 406028 97834
rect 405976 97770 406028 97776
rect 405988 97737 406016 97770
rect 405974 97728 406030 97737
rect 405974 97663 406030 97672
rect 427226 96232 427282 96241
rect 427226 96167 427282 96176
rect 427240 95862 427268 96167
rect 427228 95856 427280 95862
rect 427228 95798 427280 95804
rect 405976 95788 406028 95794
rect 405976 95730 406028 95736
rect 405988 95561 406016 95730
rect 405974 95552 406030 95561
rect 405974 95487 406030 95496
rect 405974 92424 406030 92433
rect 405974 92359 406030 92368
rect 405988 92326 406016 92359
rect 405976 92320 406028 92326
rect 405976 92262 406028 92268
rect 405974 90248 406030 90257
rect 405974 90183 405976 90192
rect 406028 90183 406030 90192
rect 405976 90154 406028 90160
rect 410220 87362 410248 88860
rect 412888 87498 412916 88860
rect 412876 87492 412928 87498
rect 412876 87434 412928 87440
rect 415556 87401 415584 88860
rect 417028 88846 418238 88874
rect 419788 88846 420906 88874
rect 415542 87392 415598 87401
rect 410208 87356 410260 87362
rect 415542 87327 415598 87336
rect 410208 87298 410260 87304
rect 389416 55056 389468 55062
rect 389416 54998 389468 55004
rect 364116 12420 364168 12426
rect 364116 12362 364168 12368
rect 376996 12420 377048 12426
rect 376996 12362 377048 12368
rect 378284 12420 378336 12426
rect 378284 12362 378336 12368
rect 362460 12352 362512 12358
rect 362460 12294 362512 12300
rect 350776 9428 350828 9434
rect 350776 9370 350828 9376
rect 351236 9428 351288 9434
rect 351236 9370 351288 9376
rect 351248 9304 351276 9370
rect 364128 9304 364156 12362
rect 377008 9304 377036 12362
rect 389428 9434 389456 54998
rect 417028 45950 417056 88846
rect 419788 47446 419816 88846
rect 423560 87430 423588 88860
rect 423548 87424 423600 87430
rect 423548 87366 423600 87372
rect 419776 47440 419828 47446
rect 419776 47382 419828 47388
rect 417016 45944 417068 45950
rect 417016 45886 417068 45892
rect 427332 15350 427360 126223
rect 427424 112114 427452 220199
rect 428698 215232 428754 215241
rect 428698 215167 428754 215176
rect 427502 210200 427558 210209
rect 427502 210135 427558 210144
rect 427516 137138 427544 210135
rect 427688 196564 427740 196570
rect 427688 196506 427740 196512
rect 427594 195240 427650 195249
rect 427594 195175 427650 195184
rect 427608 173042 427636 195175
rect 427700 185457 427728 196506
rect 427686 185448 427742 185457
rect 427686 185383 427742 185392
rect 427596 173036 427648 173042
rect 427596 172978 427648 172984
rect 427504 137132 427556 137138
rect 427504 137074 427556 137080
rect 428712 123985 428740 215167
rect 429620 208872 429672 208878
rect 429618 208840 429620 208849
rect 429672 208840 429674 208849
rect 429618 208775 429674 208784
rect 428792 199760 428844 199766
rect 428792 199702 428844 199708
rect 428804 160297 428832 199702
rect 429526 196736 429582 196745
rect 429526 196671 429582 196680
rect 429540 196570 429568 196671
rect 429528 196564 429580 196570
rect 429528 196506 429580 196512
rect 429344 189900 429396 189906
rect 429344 189842 429396 189848
rect 429356 184641 429384 189842
rect 429342 184632 429398 184641
rect 429342 184567 429398 184576
rect 429896 173036 429948 173042
rect 429896 172978 429948 172984
rect 429908 172537 429936 172978
rect 429894 172528 429950 172537
rect 429894 172463 429950 172472
rect 428790 160288 428846 160297
rect 428790 160223 428846 160232
rect 429436 148216 429488 148222
rect 429434 148184 429436 148193
rect 429488 148184 429490 148193
rect 429434 148119 429490 148128
rect 429436 137132 429488 137138
rect 429436 137074 429488 137080
rect 429448 136089 429476 137074
rect 429434 136080 429490 136089
rect 429434 136015 429490 136024
rect 428698 123976 428754 123985
rect 428698 123911 428754 123920
rect 427502 121256 427558 121265
rect 427502 121191 427558 121200
rect 427412 112108 427464 112114
rect 427412 112050 427464 112056
rect 427410 101264 427466 101273
rect 427410 101199 427466 101208
rect 427424 76414 427452 101199
rect 427412 76408 427464 76414
rect 427412 76350 427464 76356
rect 427516 28134 427544 121191
rect 428698 116224 428754 116233
rect 428698 116159 428754 116168
rect 427594 111328 427650 111337
rect 427594 111263 427650 111272
rect 427608 51594 427636 111263
rect 427686 106296 427742 106305
rect 427686 106231 427742 106240
rect 427700 105518 427728 106231
rect 427688 105512 427740 105518
rect 427688 105454 427740 105460
rect 427688 98576 427740 98582
rect 427688 98518 427740 98524
rect 427700 91617 427728 98518
rect 427686 91608 427742 91617
rect 427686 91543 427742 91552
rect 428056 81304 428108 81310
rect 428056 81246 428108 81252
rect 427596 51588 427648 51594
rect 427596 51530 427648 51536
rect 427504 28128 427556 28134
rect 427504 28070 427556 28076
rect 427320 15344 427372 15350
rect 427320 15286 427372 15292
rect 402756 12352 402808 12358
rect 402756 12294 402808 12300
rect 389416 9428 389468 9434
rect 389416 9370 389468 9376
rect 389876 9428 389928 9434
rect 389876 9370 389928 9376
rect 389888 9304 389916 9370
rect 402768 9304 402796 12294
rect 415636 12284 415688 12290
rect 415636 12226 415688 12232
rect 415648 9304 415676 12226
rect 428068 9434 428096 81246
rect 428712 39121 428740 116159
rect 429436 112108 429488 112114
rect 429436 112050 429488 112056
rect 429448 111881 429476 112050
rect 429434 111872 429490 111881
rect 429434 111807 429490 111816
rect 430080 105512 430132 105518
rect 430080 105454 430132 105460
rect 429434 99768 429490 99777
rect 429434 99703 429490 99712
rect 429448 98582 429476 99703
rect 429436 98576 429488 98582
rect 429436 98518 429488 98524
rect 429436 76408 429488 76414
rect 429436 76350 429488 76356
rect 429448 75433 429476 76350
rect 429434 75424 429490 75433
rect 429434 75359 429490 75368
rect 430092 63329 430120 105454
rect 430172 95856 430224 95862
rect 430172 95798 430224 95804
rect 430184 87537 430212 95798
rect 430170 87528 430226 87537
rect 430170 87463 430226 87472
rect 430078 63320 430134 63329
rect 430078 63255 430134 63264
rect 429804 51588 429856 51594
rect 429804 51530 429856 51536
rect 429816 51225 429844 51530
rect 429802 51216 429858 51225
rect 429802 51151 429858 51160
rect 428698 39112 428754 39121
rect 428698 39047 428754 39056
rect 429436 28128 429488 28134
rect 429436 28070 429488 28076
rect 429448 27017 429476 28070
rect 429434 27008 429490 27017
rect 429434 26943 429490 26952
rect 429436 15344 429488 15350
rect 429436 15286 429488 15292
rect 429448 14913 429476 15286
rect 429434 14904 429490 14913
rect 429434 14839 429490 14848
rect 428056 9428 428108 9434
rect 428056 9370 428108 9376
rect 428516 9428 428568 9434
rect 428516 9370 428568 9376
rect 428528 9304 428556 9370
rect 16354 8824 16410 9304
rect 29234 8824 29290 9304
rect 42114 8824 42170 9304
rect 54994 8824 55050 9304
rect 67874 8824 67930 9304
rect 80754 8824 80810 9304
rect 93634 8824 93690 9304
rect 106514 8824 106570 9304
rect 119394 8824 119450 9304
rect 132274 8824 132330 9304
rect 145154 8824 145210 9304
rect 158034 8824 158090 9304
rect 170914 8824 170970 9304
rect 183794 8824 183850 9304
rect 196674 8824 196730 9304
rect 209554 8824 209610 9304
rect 222434 8824 222490 9304
rect 235314 8824 235370 9304
rect 248194 8824 248250 9304
rect 261074 8824 261130 9304
rect 273954 8824 274010 9304
rect 286834 8824 286890 9304
rect 299714 8824 299770 9304
rect 312594 8824 312650 9304
rect 325474 8824 325530 9304
rect 338354 8824 338410 9304
rect 351234 8824 351290 9304
rect 364114 8824 364170 9304
rect 376994 8824 377050 9304
rect 389874 8824 389930 9304
rect 402754 8824 402810 9304
rect 415634 8824 415690 9304
rect 428514 8824 428570 9304
<< via2 >>
rect 13134 391296 13190 391352
rect 13686 380552 13742 380608
rect 13594 369808 13650 369864
rect 13502 359064 13558 359120
rect 13410 348184 13466 348240
rect 13318 337440 13374 337496
rect 14698 326696 14754 326752
rect 13318 315952 13374 316008
rect 13042 272840 13098 272896
rect 38802 315544 38858 315600
rect 16078 313776 16134 313832
rect 13410 305072 13466 305128
rect 13502 294328 13558 294384
rect 13594 261960 13650 262016
rect 13134 251216 13190 251272
rect 13318 240508 13320 240528
rect 13320 240508 13372 240528
rect 13372 240508 13374 240528
rect 13318 240472 13374 240508
rect 12858 229728 12914 229784
rect 13042 218848 13098 218904
rect 13042 208140 13044 208160
rect 13044 208140 13096 208160
rect 13096 208140 13098 208160
rect 13042 208104 13098 208140
rect 13042 197360 13098 197416
rect 13042 186652 13044 186672
rect 13044 186652 13096 186672
rect 13096 186652 13098 186672
rect 13042 186616 13098 186652
rect 13042 175772 13044 175792
rect 13044 175772 13096 175792
rect 13096 175772 13098 175792
rect 13042 175736 13098 175772
rect 12674 154248 12730 154304
rect 38434 313096 38490 313152
rect 38802 310376 38858 310432
rect 16262 308336 16318 308392
rect 16170 293104 16226 293160
rect 16170 219936 16226 219992
rect 16078 184168 16134 184224
rect 13410 164992 13466 165048
rect 13318 143504 13374 143560
rect 13042 132624 13098 132680
rect 16078 126096 16134 126152
rect 13226 121916 13228 121936
rect 13228 121916 13280 121936
rect 13280 121916 13282 121936
rect 13226 121880 13282 121916
rect 12858 111136 12914 111192
rect 12858 100392 12914 100448
rect 13226 89512 13282 89568
rect 13502 78768 13558 78824
rect 13410 68024 13466 68080
rect 13318 57280 13374 57336
rect 13042 46400 13098 46456
rect 12858 35656 12914 35712
rect 12674 24948 12676 24968
rect 12676 24948 12728 24968
rect 12728 24948 12730 24968
rect 12674 24912 12730 24948
rect 38802 308064 38858 308120
rect 38802 305616 38858 305672
rect 16446 304120 16502 304176
rect 16354 298680 16410 298736
rect 16354 214496 16410 214552
rect 16262 195320 16318 195376
rect 16262 120656 16318 120712
rect 38618 303032 38674 303088
rect 38802 300620 38804 300640
rect 38804 300620 38856 300640
rect 38856 300620 38858 300640
rect 38802 300584 38858 300620
rect 38250 298136 38306 298192
rect 38802 295416 38858 295472
rect 18010 293784 18066 293840
rect 18010 293104 18066 293160
rect 38434 293104 38490 293160
rect 38526 290520 38582 290576
rect 17458 289024 17514 289080
rect 38526 288072 38582 288128
rect 38526 285508 38582 285544
rect 38526 285488 38528 285508
rect 38528 285488 38580 285508
rect 38580 285488 38582 285508
rect 17550 283720 17606 283776
rect 38526 283040 38582 283096
rect 38066 280320 38122 280376
rect 51222 308608 51278 308664
rect 50302 300620 50304 300640
rect 50304 300620 50356 300640
rect 50356 300620 50358 300640
rect 50302 300584 50358 300620
rect 53062 326288 53118 326344
rect 54074 326288 54130 326344
rect 55086 326288 55142 326344
rect 56098 326288 56154 326344
rect 55086 315852 55088 315872
rect 55088 315852 55140 315872
rect 55140 315852 55142 315872
rect 55086 315816 55142 315852
rect 51590 313796 51646 313832
rect 51590 313776 51592 313796
rect 51592 313776 51644 313796
rect 51644 313776 51646 313796
rect 54074 310920 54130 310976
rect 55086 308064 55142 308120
rect 54074 306196 54076 306216
rect 54076 306196 54128 306216
rect 54128 306196 54130 306216
rect 54074 306160 54130 306196
rect 51866 304256 51922 304312
rect 73394 304664 73450 304720
rect 55086 300856 55142 300912
rect 51682 298952 51738 299008
rect 52602 293804 52658 293840
rect 52602 293784 52604 293804
rect 52604 293784 52656 293804
rect 52656 293784 52658 293804
rect 54902 292016 54958 292072
rect 18102 279504 18158 279560
rect 38618 278144 38674 278200
rect 54534 289228 54590 289284
rect 74222 314456 74278 314512
rect 74130 311056 74186 311112
rect 74038 290112 74094 290168
rect 54902 289024 54958 289080
rect 74038 288888 74094 288944
rect 51498 287528 51554 287584
rect 51682 287528 51738 287584
rect 52050 283856 52106 283912
rect 74314 308200 74370 308256
rect 75418 299904 75474 299960
rect 75418 298680 75474 298736
rect 74406 296232 74462 296288
rect 74222 293512 74278 293568
rect 74222 291608 74278 291664
rect 75970 296232 76026 296288
rect 75878 293512 75934 293568
rect 74406 289024 74462 289080
rect 74314 288752 74370 288808
rect 74038 279504 74094 279560
rect 74314 279504 74370 279560
rect 52602 279368 52658 279424
rect 74038 278144 74094 278200
rect 53522 266720 53578 266776
rect 54534 266720 54590 266776
rect 55546 266720 55602 266776
rect 56558 266720 56614 266776
rect 73854 263476 73910 263512
rect 73854 263456 73856 263476
rect 73856 263456 73908 263476
rect 73908 263456 73910 263476
rect 49198 262524 49254 262560
rect 49198 262504 49200 262524
rect 49200 262504 49252 262524
rect 49252 262504 49254 262524
rect 46714 259104 46770 259160
rect 46622 255976 46678 256032
rect 46530 252848 46586 252904
rect 46438 249720 46494 249776
rect 47082 237344 47138 237400
rect 17550 209600 17606 209656
rect 16538 208920 16594 208976
rect 17550 208920 17606 208976
rect 16446 204840 16502 204896
rect 38066 219392 38122 219448
rect 38526 216808 38582 216864
rect 38526 214224 38582 214280
rect 17642 199672 17698 199728
rect 17090 189744 17146 189800
rect 38710 211504 38766 211560
rect 38526 209192 38582 209248
rect 38526 206608 38582 206664
rect 38526 204432 38582 204488
rect 38526 201440 38582 201496
rect 38526 199128 38582 199184
rect 38526 196408 38582 196464
rect 38802 194504 38858 194560
rect 38802 191512 38858 191568
rect 38066 189200 38122 189256
rect 38066 186480 38122 186536
rect 38802 184052 38858 184088
rect 38802 184032 38804 184052
rect 38804 184032 38856 184052
rect 38856 184032 38858 184052
rect 16446 115080 16502 115136
rect 16538 111000 16594 111056
rect 18102 106240 18158 106296
rect 17458 101208 17514 101264
rect 18102 96176 18158 96232
rect 17274 91280 17330 91336
rect 46898 165128 46954 165184
rect 46622 162544 46678 162600
rect 46530 158872 46586 158928
rect 46438 155744 46494 155800
rect 51406 210144 51462 210200
rect 51406 206780 51408 206800
rect 51408 206780 51460 206800
rect 51460 206780 51462 206800
rect 51406 206744 51462 206780
rect 51406 205248 51462 205304
rect 53522 232448 53578 232504
rect 54534 232448 54590 232504
rect 56558 230952 56614 231008
rect 55546 229592 55602 229648
rect 53246 221296 53302 221352
rect 51866 220208 51922 220264
rect 51682 215176 51738 215232
rect 54074 210980 54130 211016
rect 54074 210960 54076 210980
rect 54076 210960 54128 210980
rect 54128 210960 54130 210980
rect 74682 235576 74738 235632
rect 74406 235032 74462 235088
rect 74682 234896 74738 234952
rect 72658 210144 72714 210200
rect 73486 210144 73542 210200
rect 51314 195184 51370 195240
rect 51406 185256 51462 185312
rect 51774 200216 51830 200272
rect 51774 190152 51830 190208
rect 55546 172880 55602 172936
rect 53522 171656 53578 171712
rect 54534 171656 54590 171712
rect 56558 172744 56614 172800
rect 73762 206608 73818 206664
rect 73946 204976 74002 205032
rect 73762 199264 73818 199320
rect 73946 199264 74002 199320
rect 73762 189472 73818 189528
rect 74222 230952 74278 231008
rect 74222 221432 74278 221488
rect 74314 220344 74370 220400
rect 74222 213136 74278 213192
rect 74222 204432 74278 204488
rect 74130 203208 74186 203264
rect 75142 233944 75198 234000
rect 80202 357568 80258 357624
rect 80202 356344 80258 356400
rect 80202 354984 80258 355040
rect 79282 354576 79338 354632
rect 80202 353352 80258 353408
rect 80202 352128 80258 352184
rect 87102 351312 87158 351368
rect 80202 350632 80258 350688
rect 79834 350360 79890 350416
rect 87010 350360 87066 350416
rect 86918 349544 86974 349600
rect 78914 349000 78970 349056
rect 78914 347504 78970 347560
rect 79006 346416 79062 346472
rect 78914 346008 78970 346064
rect 87102 348592 87158 348648
rect 87010 347232 87066 347288
rect 78914 344512 78970 344568
rect 78914 343288 78970 343344
rect 78914 342764 78970 342800
rect 78914 342744 78916 342764
rect 78916 342744 78968 342764
rect 78968 342744 78970 342764
rect 78914 341656 78970 341712
rect 78914 340976 78970 341032
rect 78914 339752 78970 339808
rect 80202 338392 80258 338448
rect 78914 337984 78970 338040
rect 80202 336216 80258 336272
rect 80202 335264 80258 335320
rect 80202 334212 80204 334232
rect 80204 334212 80256 334232
rect 80256 334212 80258 334232
rect 80202 334176 80258 334212
rect 78914 333632 78970 333688
rect 80202 332680 80258 332736
rect 80202 330912 80258 330968
rect 78914 329688 78970 329744
rect 81674 313540 81676 313560
rect 81676 313540 81728 313560
rect 81728 313540 81730 313560
rect 81674 313504 81730 313540
rect 81674 296776 81730 296832
rect 84618 284944 84674 285000
rect 84526 284536 84582 284592
rect 84618 281816 84674 281872
rect 84526 281136 84582 281192
rect 81674 280184 81730 280240
rect 131354 384768 131410 384824
rect 96854 355256 96910 355312
rect 96762 351584 96818 351640
rect 87930 346824 87986 346880
rect 88114 346008 88170 346064
rect 87470 345056 87526 345112
rect 87378 343288 87434 343344
rect 87286 341520 87342 341576
rect 88482 344240 88538 344296
rect 87470 342336 87526 342392
rect 87378 339752 87434 339808
rect 87562 340568 87618 340624
rect 87930 338800 87986 338856
rect 87378 337032 87434 337088
rect 87838 336216 87894 336272
rect 88022 337984 88078 338040
rect 95198 333768 95254 333824
rect 131446 382048 131502 382104
rect 131538 380144 131594 380200
rect 131630 377424 131686 377480
rect 131722 374704 131778 374760
rect 131814 372120 131870 372176
rect 131814 351312 131870 351368
rect 131814 350360 131870 350416
rect 131906 349544 131962 349600
rect 131814 348592 131870 348648
rect 132182 347776 132238 347832
rect 131906 346824 131962 346880
rect 131814 346008 131870 346064
rect 132366 345056 132422 345112
rect 131814 344260 131870 344296
rect 131814 344240 131816 344260
rect 131816 344240 131868 344260
rect 131868 344240 131870 344260
rect 131814 343288 131870 343344
rect 131906 342336 131962 342392
rect 131814 341520 131870 341576
rect 131814 340568 131870 340624
rect 131906 339752 131962 339808
rect 131814 338800 131870 338856
rect 131814 337984 131870 338040
rect 131906 337032 131962 337088
rect 131814 336216 131870 336272
rect 77258 263116 77314 263172
rect 79742 261688 79798 261744
rect 79742 260328 79798 260384
rect 79742 258832 79798 258888
rect 80294 257472 80350 257528
rect 79742 256112 79798 256168
rect 87194 258016 87250 258072
rect 131354 257356 131410 257392
rect 131354 257336 131356 257356
rect 131356 257336 131408 257356
rect 131408 257336 131410 257356
rect 87194 256828 87196 256848
rect 87196 256828 87248 256848
rect 87248 256828 87250 256848
rect 87194 256792 87250 256828
rect 87286 255568 87342 255624
rect 87194 255296 87250 255352
rect 79834 254616 79890 254672
rect 79742 253256 79798 253312
rect 131446 255568 131502 255624
rect 131354 254616 131410 254672
rect 87378 254344 87434 254400
rect 131354 253800 131410 253856
rect 87194 252884 87196 252904
rect 87196 252884 87248 252904
rect 87248 252884 87250 252904
rect 87194 252848 87250 252884
rect 131354 252848 131410 252904
rect 87286 252712 87342 252768
rect 79742 251896 79798 251952
rect 87194 251660 87196 251680
rect 87196 251660 87248 251680
rect 87248 251660 87250 251680
rect 87194 251624 87250 251660
rect 79742 250536 79798 250592
rect 87194 250284 87250 250320
rect 87194 250264 87196 250284
rect 87196 250264 87248 250284
rect 87248 250264 87250 250284
rect 87194 249312 87250 249368
rect 77258 249108 77314 249164
rect 87194 248360 87250 248416
rect 131998 250264 132054 250320
rect 132182 251080 132238 251136
rect 132090 249992 132146 250048
rect 131814 248904 131870 248960
rect 131722 248224 131778 248280
rect 77258 247748 77314 247804
rect 88482 247564 88538 247600
rect 88482 247544 88484 247564
rect 88484 247544 88536 247564
rect 88536 247544 88538 247564
rect 87194 246592 87250 246648
rect 77258 246388 77314 246444
rect 87286 245776 87342 245832
rect 78914 245504 78970 245560
rect 87194 244844 87250 244880
rect 87194 244824 87196 244844
rect 87196 244824 87248 244844
rect 87248 244824 87250 244844
rect 78914 244144 78970 244200
rect 131354 245504 131410 245560
rect 131354 244416 131410 244472
rect 87378 244008 87434 244064
rect 87286 243056 87342 243112
rect 80202 242784 80258 242840
rect 87194 242240 87250 242296
rect 78914 240628 78970 240664
rect 78914 240608 78916 240628
rect 78916 240608 78968 240628
rect 78968 240608 78970 240628
rect 79006 239248 79062 239304
rect 131906 242648 131962 242704
rect 98924 241696 98980 241752
rect 95198 239656 95254 239712
rect 91702 239384 91758 239440
rect 79098 238568 79154 238624
rect 102558 238568 102614 238624
rect 78914 236564 78916 236584
rect 78916 236564 78968 236584
rect 78968 236564 78970 236584
rect 78914 236528 78970 236564
rect 109826 235712 109882 235768
rect 132366 256384 132422 256440
rect 133378 252032 133434 252088
rect 132458 247000 132514 247056
rect 132274 246048 132330 246104
rect 132642 243056 132698 243112
rect 139634 357704 139690 357760
rect 174042 357160 174098 357216
rect 139634 356516 139636 356536
rect 139636 356516 139688 356536
rect 139688 356516 139690 356536
rect 139634 356480 139690 356516
rect 173490 356072 173546 356128
rect 139634 355156 139636 355176
rect 139636 355156 139688 355176
rect 139688 355156 139690 355176
rect 139634 355120 139690 355156
rect 174042 355156 174044 355176
rect 174044 355156 174096 355176
rect 174096 355156 174098 355176
rect 174042 355120 174098 355156
rect 139726 354576 139782 354632
rect 173766 354032 173822 354088
rect 139634 353488 139690 353544
rect 174042 352944 174098 353000
rect 139634 352264 139690 352320
rect 174042 351992 174098 352048
rect 182322 351312 182378 351368
rect 139726 350904 139782 350960
rect 173674 350904 173730 350960
rect 139634 350496 139690 350552
rect 180758 349952 180814 350008
rect 173858 349816 173914 349872
rect 139450 349544 139506 349600
rect 172846 348864 172902 348920
rect 139542 348184 139598 348240
rect 190786 359336 190842 359392
rect 191246 351876 191302 351912
rect 191246 351856 191248 351876
rect 191248 351856 191300 351876
rect 191300 351856 191302 351876
rect 341942 393744 341998 393800
rect 225286 384768 225342 384824
rect 225194 382048 225250 382104
rect 180942 349000 180998 349056
rect 180850 348320 180906 348376
rect 174042 347776 174098 347832
rect 180758 347232 180814 347288
rect 139634 346860 139636 346880
rect 139636 346860 139688 346880
rect 139688 346860 139690 346880
rect 139634 346824 139690 346860
rect 174042 346860 174044 346880
rect 174044 346860 174096 346880
rect 174096 346860 174098 346880
rect 174042 346824 174098 346860
rect 139818 346280 139874 346336
rect 173122 345736 173178 345792
rect 139726 345328 139782 345384
rect 139634 344104 139690 344160
rect 139634 342608 139690 342664
rect 139726 342200 139782 342256
rect 139634 341248 139690 341304
rect 136966 332136 137022 332192
rect 137058 330776 137114 330832
rect 137242 328736 137298 328792
rect 137150 328056 137206 328112
rect 137242 320304 137298 320360
rect 137150 317176 137206 317232
rect 137058 314048 137114 314104
rect 136966 310920 137022 310976
rect 172754 341520 172810 341576
rect 139818 339888 139874 339944
rect 139726 338528 139782 338584
rect 181034 346824 181090 346880
rect 182322 346008 182378 346064
rect 180850 345736 180906 345792
rect 181034 345736 181090 345792
rect 173306 344648 173362 344704
rect 180942 344648 180998 344704
rect 173674 343732 173676 343752
rect 173676 343732 173728 343752
rect 173728 343732 173730 343752
rect 173674 343696 173730 343732
rect 173030 342608 173086 342664
rect 172938 340568 172994 340624
rect 139910 338120 139966 338176
rect 139726 336760 139782 336816
rect 139634 335808 139690 335864
rect 139634 334312 139690 334368
rect 139634 333904 139690 333960
rect 139634 332952 139690 333008
rect 173306 335400 173362 335456
rect 182322 344240 182378 344296
rect 181402 343288 181458 343344
rect 182138 342336 182194 342392
rect 181770 341520 181826 341576
rect 181402 340568 181458 340624
rect 181586 339752 181642 339808
rect 173674 339480 173730 339536
rect 174042 338548 174098 338584
rect 182322 338800 182378 338856
rect 174042 338528 174044 338548
rect 174044 338528 174096 338548
rect 174096 338528 174098 338548
rect 173950 337440 174006 337496
rect 180390 337440 180446 337496
rect 173490 336352 173546 336408
rect 173398 334312 173454 334368
rect 181586 337032 181642 337088
rect 180942 336080 180998 336136
rect 173306 333224 173362 333280
rect 172846 332272 172902 332328
rect 139634 331592 139690 331648
rect 173674 331184 173730 331240
rect 140370 330232 140426 330288
rect 172110 330232 172166 330288
rect 158586 330096 158642 330152
rect 159598 330096 159654 330152
rect 137518 307792 137574 307848
rect 136874 304664 136930 304720
rect 137518 304664 137574 304720
rect 136414 301536 136470 301592
rect 136874 284808 136930 284864
rect 136874 282496 136930 282552
rect 136874 282224 136930 282280
rect 75418 217352 75474 217408
rect 74406 211640 74462 211696
rect 74406 205384 74462 205440
rect 74314 200488 74370 200544
rect 74314 191920 74370 191976
rect 74314 190968 74370 191024
rect 74222 187976 74278 188032
rect 74498 187024 74554 187080
rect 74222 186888 74278 186944
rect 74038 185120 74094 185176
rect 74406 181176 74462 181232
rect 73762 179952 73818 180008
rect 72658 169752 72714 169808
rect 74498 179952 74554 180008
rect 74406 171656 74462 171712
rect 73486 169480 73542 169536
rect 49198 168836 49200 168856
rect 49200 168836 49252 168856
rect 49252 168836 49254 168856
rect 49198 168800 49254 168836
rect 47082 143368 47138 143424
rect 38802 127456 38858 127512
rect 38250 125552 38306 125608
rect 38802 122696 38858 122752
rect 38802 120248 38858 120304
rect 38250 117528 38306 117584
rect 38802 114944 38858 115000
rect 38802 112768 38858 112824
rect 38250 110456 38306 110512
rect 38802 107484 38858 107520
rect 38802 107464 38804 107484
rect 38804 107464 38856 107484
rect 38856 107464 38858 107484
rect 38802 105288 38858 105344
rect 38618 102432 38674 102488
rect 38802 100256 38858 100312
rect 38802 97828 38858 97864
rect 38802 97808 38804 97828
rect 38804 97808 38856 97828
rect 38856 97808 38858 97828
rect 38066 95360 38122 95416
rect 37606 92504 37662 92560
rect 51222 126232 51278 126288
rect 51222 116168 51278 116224
rect 53522 139560 53578 139616
rect 54534 139560 54590 139616
rect 55638 132352 55694 132408
rect 55454 131536 55510 131592
rect 74038 141600 74094 141656
rect 74130 141464 74186 141520
rect 74314 141736 74370 141792
rect 54074 127184 54130 127240
rect 53154 122696 53210 122752
rect 74130 122696 74186 122752
rect 52602 121200 52658 121256
rect 73394 120520 73450 120576
rect 73394 119704 73450 119760
rect 54074 117140 54130 117176
rect 54074 117120 54076 117140
rect 54076 117120 54128 117140
rect 54128 117120 54130 117140
rect 52142 113040 52198 113096
rect 52602 111272 52658 111328
rect 38802 90056 38858 90112
rect 52602 106240 52658 106296
rect 52602 101208 52658 101264
rect 52602 96176 52658 96232
rect 52602 91280 52658 91336
rect 53062 79040 53118 79096
rect 54074 79040 54130 79096
rect 55086 78904 55142 78960
rect 56098 79040 56154 79096
rect 73486 116168 73542 116224
rect 72566 88288 72622 88344
rect 73578 112768 73634 112824
rect 73670 109504 73726 109560
rect 73670 108824 73726 108880
rect 73578 86384 73634 86440
rect 74406 126368 74462 126424
rect 74314 120520 74370 120576
rect 74222 105424 74278 105480
rect 74222 105288 74278 105344
rect 74682 94308 74684 94328
rect 74684 94308 74736 94328
rect 74736 94308 74738 94328
rect 74682 94272 74738 94308
rect 81674 219548 81730 219584
rect 81674 219528 81676 219548
rect 81676 219528 81728 219548
rect 81728 219528 81730 219548
rect 81674 202800 81730 202856
rect 81674 186208 81730 186264
rect 79190 169072 79246 169128
rect 77258 167644 77314 167700
rect 77258 166284 77314 166340
rect 77258 164808 77314 164844
rect 77258 164788 77260 164808
rect 77260 164788 77312 164808
rect 77312 164788 77314 164808
rect 77258 163448 77314 163484
rect 77258 163428 77260 163448
rect 77260 163428 77312 163448
rect 77312 163428 77314 163448
rect 87194 164040 87250 164096
rect 87102 163088 87158 163144
rect 77258 162068 77314 162124
rect 87286 161864 87342 161920
rect 87194 161320 87250 161376
rect 87194 160368 87250 160424
rect 81766 159960 81822 160016
rect 79282 159300 79338 159336
rect 79282 159280 79284 159300
rect 79284 159280 79336 159300
rect 79336 159280 79338 159300
rect 87194 158872 87250 158928
rect 87286 158600 87342 158656
rect 79742 157940 79798 157976
rect 79742 157920 79744 157940
rect 79744 157920 79796 157940
rect 79796 157920 79798 157940
rect 87194 157648 87250 157704
rect 77258 156512 77314 156548
rect 77258 156492 77260 156512
rect 77260 156492 77312 156512
rect 77312 156492 77314 156512
rect 87194 156288 87250 156344
rect 87194 155336 87250 155392
rect 79742 155084 79798 155120
rect 79742 155064 79744 155084
rect 79744 155064 79796 155084
rect 79796 155064 79798 155084
rect 87194 154404 87250 154440
rect 87194 154384 87196 154404
rect 87196 154384 87248 154404
rect 87248 154384 87250 154404
rect 81766 153704 81822 153760
rect 87194 153568 87250 153624
rect 87194 152616 87250 152672
rect 81766 152344 81822 152400
rect 88114 151800 88170 151856
rect 79742 150848 79798 150904
rect 87102 150848 87158 150904
rect 79742 148148 79798 148184
rect 79742 148128 79744 148148
rect 79744 148128 79796 148148
rect 79796 148128 79798 148148
rect 81766 149524 81768 149544
rect 81768 149524 81820 149544
rect 81820 149524 81822 149544
rect 81766 149488 81822 149524
rect 87194 150032 87250 150088
rect 87194 149080 87250 149136
rect 80110 146632 80166 146688
rect 87286 148264 87342 148320
rect 79742 145272 79798 145328
rect 79742 143912 79798 143968
rect 77258 142484 77314 142540
rect 82318 141600 82374 141656
rect 77718 141464 77774 141520
rect 98878 145136 98934 145192
rect 95198 144456 95254 144512
rect 109734 143096 109790 143152
rect 106146 142552 106202 142608
rect 131354 163360 131410 163416
rect 131446 161592 131502 161648
rect 131354 160676 131356 160696
rect 131356 160676 131408 160696
rect 131408 160676 131410 160696
rect 131354 160640 131410 160676
rect 131354 159824 131410 159880
rect 131998 162408 132054 162464
rect 131630 152208 131686 152264
rect 131354 150440 131410 150496
rect 132182 158872 132238 158928
rect 132274 157104 132330 157160
rect 132090 156016 132146 156072
rect 131998 155064 132054 155120
rect 131906 153568 131962 153624
rect 131814 149488 131870 149544
rect 131354 148808 131410 148864
rect 132550 158056 132606 158112
rect 132366 156288 132422 156344
rect 132458 150848 132514 150904
rect 132642 153296 132698 153352
rect 81674 125452 81676 125472
rect 81676 125452 81728 125472
rect 81728 125452 81730 125472
rect 81674 125416 81730 125452
rect 73854 91144 73910 91200
rect 73670 86248 73726 86304
rect 73486 86112 73542 86168
rect 73762 86112 73818 86168
rect 72842 85840 72898 85896
rect 72842 76456 72898 76512
rect 78178 110864 78234 110920
rect 78178 109640 78234 109696
rect 81674 108824 81730 108880
rect 81674 92232 81730 92288
rect 78914 75776 78970 75832
rect 78914 73872 78970 73928
rect 78914 72784 78970 72840
rect 78914 71560 78970 71616
rect 80202 71152 80258 71208
rect 78914 69792 78970 69848
rect 78914 68568 78970 68624
rect 78914 67480 78970 67536
rect 78914 66800 78970 66856
rect 78914 65576 78970 65632
rect 78914 64624 78970 64680
rect 78914 63400 78970 63456
rect 78914 62856 78970 62912
rect 78914 61496 78970 61552
rect 78914 60272 78970 60328
rect 78914 57280 78970 57336
rect 78914 56192 78970 56248
rect 87378 69384 87434 69440
rect 131354 69420 131356 69440
rect 131356 69420 131408 69440
rect 131408 69420 131410 69440
rect 131354 69384 131410 69420
rect 87194 68432 87250 68488
rect 131446 68432 131502 68488
rect 87194 67616 87250 67672
rect 132366 67616 132422 67672
rect 87194 66700 87196 66720
rect 87196 66700 87248 66720
rect 87248 66700 87250 66720
rect 87194 66664 87250 66700
rect 131354 66684 131410 66720
rect 131354 66664 131356 66684
rect 131356 66664 131408 66684
rect 131408 66664 131410 66684
rect 87286 65848 87342 65904
rect 132366 65848 132422 65904
rect 87286 64896 87342 64952
rect 131354 64896 131410 64952
rect 87194 64080 87250 64136
rect 131446 64080 131502 64136
rect 87194 63128 87250 63184
rect 132366 63128 132422 63184
rect 87286 62312 87342 62368
rect 87194 61360 87250 61416
rect 87194 60408 87250 60464
rect 80202 59048 80258 59104
rect 80202 58504 80258 58560
rect 131354 62312 131410 62368
rect 131722 61360 131778 61416
rect 131354 60408 131410 60464
rect 87378 59592 87434 59648
rect 132642 59592 132698 59648
rect 87194 58640 87250 58696
rect 132550 58640 132606 58696
rect 87194 57824 87250 57880
rect 132642 57824 132698 57880
rect 87194 56872 87250 56928
rect 87286 56056 87342 56112
rect 79558 55648 79614 55704
rect 78914 54560 78970 54616
rect 87378 55104 87434 55160
rect 132642 56872 132698 56928
rect 132550 56056 132606 56112
rect 132642 55104 132698 55160
rect 134206 55124 134262 55160
rect 134206 55104 134208 55124
rect 134208 55104 134260 55124
rect 134260 55104 134262 55124
rect 87194 54324 87196 54344
rect 87196 54324 87248 54344
rect 87248 54324 87250 54344
rect 87194 54288 87250 54324
rect 78914 53608 78970 53664
rect 79006 50752 79062 50808
rect 78914 50244 78916 50264
rect 78916 50244 78968 50264
rect 78968 50244 78970 50264
rect 78914 50208 78970 50244
rect 87470 49256 87526 49312
rect 78914 49120 78970 49176
rect 67874 48032 67930 48088
rect 74314 48032 74370 48088
rect 87102 48032 87158 48088
rect 88298 48032 88354 48088
rect 72566 47388 72568 47408
rect 72568 47388 72620 47408
rect 72620 47388 72622 47408
rect 72566 47352 72622 47388
rect 74682 47352 74738 47408
rect 64194 45856 64250 45912
rect 88114 33616 88170 33672
rect 88206 30760 88262 30816
rect 88298 28040 88354 28096
rect 93634 50616 93690 50672
rect 102374 51296 102430 51352
rect 105134 49256 105190 49312
rect 105134 48032 105190 48088
rect 107526 50208 107582 50264
rect 106606 47352 106662 47408
rect 109458 50208 109514 50264
rect 109458 47216 109514 47272
rect 118198 53064 118254 53120
rect 113598 47488 113654 47544
rect 118658 44632 118714 44688
rect 132642 54324 132644 54344
rect 132644 54324 132696 54344
rect 132696 54324 132698 54344
rect 132642 54288 132698 54324
rect 137610 298544 137666 298600
rect 137610 285216 137666 285272
rect 137518 273792 137574 273848
rect 136966 238604 136968 238624
rect 136968 238604 137020 238624
rect 137020 238604 137022 238624
rect 136966 238568 137022 238604
rect 136966 235712 137022 235768
rect 136966 235032 137022 235088
rect 137150 233028 137152 233048
rect 137152 233028 137204 233048
rect 137204 233028 137206 233048
rect 137150 232992 137206 233028
rect 137702 279640 137758 279696
rect 138622 278144 138678 278200
rect 137794 276512 137850 276568
rect 138070 273384 138126 273440
rect 161714 328736 161770 328792
rect 160702 328056 160758 328112
rect 201826 333088 201882 333144
rect 201826 332136 201882 332192
rect 205598 331592 205654 331648
rect 208726 328056 208782 328112
rect 212314 333496 212370 333552
rect 225378 380144 225434 380200
rect 319034 384768 319090 384824
rect 225470 377424 225526 377480
rect 225562 374704 225618 374760
rect 225470 333088 225526 333144
rect 225378 331592 225434 331648
rect 225838 372120 225894 372176
rect 233474 357704 233530 357760
rect 233474 356516 233476 356536
rect 233476 356516 233528 356536
rect 233528 356516 233530 356536
rect 233474 356480 233530 356516
rect 233474 355156 233476 355176
rect 233476 355156 233528 355176
rect 233528 355156 233530 355176
rect 233474 355120 233530 355156
rect 233566 354576 233622 354632
rect 233474 353488 233530 353544
rect 233474 352264 233530 352320
rect 226298 351332 226354 351368
rect 226298 351312 226300 351332
rect 226300 351312 226352 351332
rect 226352 351312 226354 351332
rect 226574 350360 226630 350416
rect 226482 349544 226538 349600
rect 226390 348592 226446 348648
rect 233474 350904 233530 350960
rect 233566 350496 233622 350552
rect 233474 349544 233530 349600
rect 226390 347776 226446 347832
rect 226482 346824 226538 346880
rect 226390 346008 226446 346064
rect 226022 345056 226078 345112
rect 226390 344260 226446 344296
rect 226390 344240 226392 344260
rect 226392 344240 226444 344260
rect 226444 344240 226446 344260
rect 226390 343288 226446 343344
rect 226482 342336 226538 342392
rect 226390 341520 226446 341576
rect 233474 348220 233476 348240
rect 233476 348220 233528 348240
rect 233528 348220 233530 348240
rect 233474 348184 233530 348220
rect 233474 346860 233476 346880
rect 233476 346860 233528 346880
rect 233528 346860 233530 346880
rect 233474 346824 233530 346860
rect 233566 346416 233622 346472
rect 233474 345192 233530 345248
rect 233474 343968 233530 344024
rect 233474 342200 233530 342256
rect 233474 341112 233530 341168
rect 226390 340568 226446 340624
rect 225930 339752 225986 339808
rect 226482 338820 226538 338856
rect 226482 338800 226484 338820
rect 226484 338800 226536 338820
rect 226536 338800 226538 338820
rect 225930 337984 225986 338040
rect 225930 337032 225986 337088
rect 226482 336216 226538 336272
rect 234578 342608 234634 342664
rect 233658 339888 233714 339944
rect 233566 338528 233622 338584
rect 233474 337032 233530 337088
rect 175514 313504 175570 313560
rect 145522 310104 145578 310160
rect 145430 296776 145486 296832
rect 145614 283484 145616 283504
rect 145616 283484 145668 283504
rect 145668 283484 145670 283504
rect 145614 283448 145670 283484
rect 138622 269712 138678 269768
rect 142394 263592 142450 263648
rect 159046 274608 159102 274664
rect 157758 274472 157814 274528
rect 158402 274472 158458 274528
rect 157206 274336 157262 274392
rect 156194 263864 156250 263920
rect 167878 306160 167934 306216
rect 175514 296776 175570 296832
rect 168062 286304 168118 286360
rect 175790 280184 175846 280240
rect 139818 263048 139874 263104
rect 138806 259920 138862 259976
rect 138806 250400 138862 250456
rect 139542 248360 139598 248416
rect 138898 244144 138954 244200
rect 140186 238432 140242 238488
rect 140370 261688 140426 261744
rect 140370 260328 140426 260384
rect 140554 258832 140610 258888
rect 140554 257472 140610 257528
rect 140554 256112 140610 256168
rect 140554 254616 140610 254672
rect 140462 253256 140518 253312
rect 140370 250536 140426 250592
rect 140278 237208 140334 237264
rect 140738 251896 140794 251952
rect 140554 249584 140610 249640
rect 140646 246864 140702 246920
rect 140554 245504 140610 245560
rect 140646 242784 140702 242840
rect 140554 240628 140610 240664
rect 140554 240608 140556 240628
rect 140556 240608 140608 240628
rect 140608 240608 140610 240628
rect 140554 239268 140610 239304
rect 140554 239248 140556 239268
rect 140556 239248 140608 239268
rect 140608 239248 140610 239268
rect 173398 263048 173454 263104
rect 172938 253276 172994 253312
rect 172938 253256 172940 253276
rect 172940 253256 172992 253276
rect 172992 253256 172994 253276
rect 173122 250536 173178 250592
rect 173490 261688 173546 261744
rect 173306 249040 173362 249096
rect 173306 247680 173362 247736
rect 173766 260328 173822 260384
rect 173858 258832 173914 258888
rect 173766 254616 173822 254672
rect 173674 251916 173730 251952
rect 173674 251896 173676 251916
rect 173676 251896 173728 251916
rect 173728 251896 173730 251916
rect 173306 244824 173362 244880
rect 173306 243464 173362 243520
rect 172938 242104 172994 242160
rect 173950 257472 174006 257528
rect 173674 246320 173730 246376
rect 173582 240608 173638 240664
rect 174042 256112 174098 256168
rect 173858 239248 173914 239304
rect 142762 238296 142818 238352
rect 174042 237888 174098 237944
rect 172938 236528 172994 236584
rect 147454 236120 147510 236176
rect 137702 234896 137758 234952
rect 139266 234896 139322 234952
rect 137702 226328 137758 226384
rect 137334 223200 137390 223256
rect 137242 220072 137298 220128
rect 137150 216944 137206 217000
rect 137058 213816 137114 213872
rect 136966 210688 137022 210744
rect 136874 204432 136930 204488
rect 136874 200896 136930 200952
rect 136966 141872 137022 141928
rect 136874 139832 136930 139888
rect 136874 132896 136930 132952
rect 137334 141056 137390 141112
rect 137242 134392 137298 134448
rect 137058 125960 137114 126016
rect 136966 123240 137022 123296
rect 136874 120384 136930 120440
rect 136874 113176 136930 113232
rect 136874 110728 136930 110784
rect 137702 216536 137758 216592
rect 138162 208240 138218 208296
rect 138162 207560 138218 207616
rect 137702 191920 137758 191976
rect 137794 188520 137850 188576
rect 137610 185664 137666 185720
rect 145154 216128 145210 216184
rect 148374 236120 148430 236176
rect 148650 235984 148706 236040
rect 148742 235848 148798 235904
rect 147822 235032 147878 235088
rect 152054 234896 152110 234952
rect 149294 233672 149350 233728
rect 150122 233672 150178 233728
rect 149294 232992 149350 233048
rect 153250 233536 153306 233592
rect 145430 202800 145486 202856
rect 145614 189472 145670 189528
rect 137886 182536 137942 182592
rect 138898 179408 138954 179464
rect 148742 179952 148798 180008
rect 148742 173016 148798 173072
rect 154722 181992 154778 182048
rect 155274 181176 155330 181232
rect 157206 180904 157262 180960
rect 158402 181040 158458 181096
rect 157758 180768 157814 180824
rect 156562 180632 156618 180688
rect 155918 179952 155974 180008
rect 159046 180496 159102 180552
rect 167970 212728 168026 212784
rect 169258 192736 169314 192792
rect 139634 164856 139690 164912
rect 139634 163496 139690 163552
rect 139634 162136 139690 162192
rect 139634 159300 139690 159336
rect 139634 159280 139636 159300
rect 139636 159280 139688 159300
rect 139688 159280 139690 159300
rect 139634 155084 139690 155120
rect 139634 155064 139636 155084
rect 139636 155064 139688 155084
rect 139688 155064 139690 155084
rect 139542 153704 139598 153760
rect 138898 148128 138954 148184
rect 139634 146632 139690 146688
rect 139634 145272 139690 145328
rect 139634 143912 139690 143968
rect 140554 169072 140610 169128
rect 140554 167712 140610 167768
rect 140554 166352 140610 166408
rect 140370 156560 140426 156616
rect 140278 142552 140334 142608
rect 140646 160640 140702 160696
rect 140462 150848 140518 150904
rect 140738 157920 140794 157976
rect 140830 152344 140886 152400
rect 140554 149488 140610 149544
rect 147914 142144 147970 142200
rect 150674 142144 150730 142200
rect 167786 142180 167788 142200
rect 167788 142180 167840 142200
rect 167840 142180 167842 142200
rect 167786 142144 167842 142180
rect 147454 142008 147510 142064
rect 137610 140376 137666 140432
rect 141842 139868 141844 139888
rect 141844 139868 141896 139888
rect 141896 139868 141898 139888
rect 141842 139832 141898 139868
rect 137610 129768 137666 129824
rect 137518 98488 137574 98544
rect 137610 92232 137666 92288
rect 137794 104064 137850 104120
rect 137794 95224 137850 95280
rect 138162 94544 138218 94600
rect 144234 122288 144290 122344
rect 149110 141056 149166 141112
rect 152054 141056 152110 141112
rect 148190 139832 148246 139888
rect 167878 118752 167934 118808
rect 147362 113584 147418 113640
rect 147362 112496 147418 112552
rect 143958 108824 144014 108880
rect 168246 98760 168302 98816
rect 144418 95496 144474 95552
rect 137702 88832 137758 88888
rect 138162 85468 138164 85488
rect 138164 85468 138216 85488
rect 138216 85468 138218 85488
rect 138162 85432 138218 85468
rect 155366 89104 155422 89160
rect 155918 87336 155974 87392
rect 156562 86792 156618 86848
rect 157758 87064 157814 87120
rect 158402 86928 158458 86984
rect 157206 86656 157262 86712
rect 159046 87064 159102 87120
rect 218018 268352 218074 268408
rect 182322 257336 182378 257392
rect 182322 256384 182378 256440
rect 181586 255568 181642 255624
rect 181586 252848 181642 252904
rect 181494 249720 181550 249776
rect 225562 255568 225618 255624
rect 182322 254616 182378 254672
rect 181770 253800 181826 253856
rect 225378 253800 225434 253856
rect 181770 252032 181826 252088
rect 182322 251080 182378 251136
rect 182230 250264 182286 250320
rect 181954 248632 182010 248688
rect 181862 248224 181918 248280
rect 182322 247272 182378 247328
rect 181678 246048 181734 246104
rect 181586 245504 181642 245560
rect 182046 244552 182102 244608
rect 225378 250264 225434 250320
rect 225746 252848 225802 252904
rect 230806 333088 230862 333144
rect 233474 335844 233476 335864
rect 233476 335844 233528 335864
rect 233528 335844 233530 335864
rect 233474 335808 233530 335844
rect 230898 332136 230954 332192
rect 230806 330776 230862 330832
rect 233750 338120 233806 338176
rect 233658 334312 233714 334368
rect 233474 333904 233530 333960
rect 233474 332952 233530 333008
rect 233474 331456 233530 331512
rect 233474 330232 233530 330288
rect 251966 330096 252022 330152
rect 252610 330096 252666 330152
rect 230990 328736 231046 328792
rect 231358 320304 231414 320360
rect 231358 317176 231414 317232
rect 230990 314048 231046 314104
rect 230898 310920 230954 310976
rect 230806 307792 230862 307848
rect 230714 298408 230770 298464
rect 230714 289060 230716 289080
rect 230716 289060 230768 289080
rect 230768 289060 230770 289080
rect 230714 289024 230770 289060
rect 231358 285216 231414 285272
rect 226022 251080 226078 251136
rect 225930 249312 225986 249368
rect 225838 248360 225894 248416
rect 225654 247544 225710 247600
rect 225378 244824 225434 244880
rect 225562 244008 225618 244064
rect 181034 243364 181036 243384
rect 181036 243364 181088 243384
rect 181088 243364 181090 243384
rect 181034 243328 181090 243364
rect 180298 242784 180354 242840
rect 189222 239656 189278 239712
rect 192902 236936 192958 236992
rect 200170 238296 200226 238352
rect 211026 239656 211082 239712
rect 207254 234896 207310 234952
rect 219766 237752 219822 237808
rect 222434 240608 222490 240664
rect 222802 240608 222858 240664
rect 226390 257336 226446 257392
rect 226298 256384 226354 256440
rect 226298 254636 226354 254672
rect 226298 254616 226300 254636
rect 226300 254616 226352 254636
rect 226352 254616 226354 254636
rect 227218 252032 227274 252088
rect 226206 246592 226262 246648
rect 226114 245776 226170 245832
rect 226298 243092 226300 243112
rect 226300 243092 226352 243112
rect 226352 243092 226354 243112
rect 226298 243056 226354 243092
rect 226390 242240 226446 242296
rect 230990 238976 231046 239032
rect 230898 238296 230954 238352
rect 179286 219528 179342 219584
rect 178918 202800 178974 202856
rect 178918 186208 178974 186264
rect 173582 169072 173638 169128
rect 173490 167712 173546 167768
rect 173398 166352 173454 166408
rect 172938 164856 172994 164912
rect 173122 163496 173178 163552
rect 173306 156560 173362 156616
rect 173398 153704 173454 153760
rect 173766 162136 173822 162192
rect 173674 159316 173676 159336
rect 173676 159316 173728 159336
rect 173728 159316 173730 159336
rect 173674 159280 173730 159316
rect 173674 157920 173730 157976
rect 173582 155084 173638 155120
rect 173582 155064 173584 155084
rect 173584 155064 173636 155084
rect 173636 155064 173638 155084
rect 173582 152380 173584 152400
rect 173584 152380 173636 152400
rect 173636 152380 173638 152400
rect 173582 152344 173638 152380
rect 174042 160660 174098 160696
rect 174042 160640 174044 160660
rect 174044 160640 174096 160660
rect 174096 160640 174098 160660
rect 173582 150848 173638 150904
rect 172754 149488 172810 149544
rect 173582 148164 173584 148184
rect 173584 148164 173636 148184
rect 173636 148164 173638 148184
rect 173582 148128 173638 148164
rect 173858 146632 173914 146688
rect 173950 145272 174006 145328
rect 174042 143912 174098 143968
rect 173582 142552 173638 142608
rect 175514 125436 175570 125472
rect 175514 125416 175516 125436
rect 175516 125416 175568 125436
rect 175568 125416 175570 125436
rect 174870 108824 174926 108880
rect 175514 92232 175570 92288
rect 182966 174920 183022 174976
rect 218018 175464 218074 175520
rect 181770 163360 181826 163416
rect 181310 162408 181366 162464
rect 180298 160912 180354 160968
rect 181678 159824 181734 159880
rect 181402 158872 181458 158928
rect 181402 153160 181458 153216
rect 182322 160660 182378 160696
rect 182322 160640 182324 160660
rect 182324 160640 182376 160660
rect 182376 160640 182378 160660
rect 182322 158056 182378 158112
rect 181678 149488 181734 149544
rect 182322 157104 182378 157160
rect 182322 156288 182378 156344
rect 182138 156016 182194 156072
rect 182322 154964 182324 154984
rect 182324 154964 182376 154984
rect 182376 154964 182378 154984
rect 182322 154928 182378 154964
rect 182322 153604 182324 153624
rect 182324 153604 182376 153624
rect 182376 153604 182378 153624
rect 182322 153568 182378 153604
rect 182322 152072 182378 152128
rect 182322 150884 182324 150904
rect 182324 150884 182376 150904
rect 182376 150884 182378 150904
rect 182322 150848 182378 150884
rect 182230 150576 182286 150632
rect 181862 148808 181918 148864
rect 192902 144592 192958 144648
rect 189222 144456 189278 144512
rect 196214 140512 196270 140568
rect 203758 143232 203814 143288
rect 207254 141056 207310 141112
rect 207898 141056 207954 141112
rect 219674 142028 219730 142064
rect 219674 142008 219676 142028
rect 219676 142008 219728 142028
rect 219728 142008 219730 142028
rect 225746 160640 225802 160696
rect 225654 152616 225710 152672
rect 226298 163360 226354 163416
rect 226206 162408 226262 162464
rect 226114 159824 226170 159880
rect 226114 157104 226170 157160
rect 226022 155336 226078 155392
rect 225930 154384 225986 154440
rect 225838 153568 225894 153624
rect 225562 150032 225618 150088
rect 225930 148264 225986 148320
rect 226298 161592 226354 161648
rect 226298 158056 226354 158112
rect 226206 151800 226262 151856
rect 227218 158872 227274 158928
rect 226390 156288 226446 156344
rect 226482 150848 226538 150904
rect 226298 149116 226300 149136
rect 226300 149116 226352 149136
rect 226352 149116 226354 149136
rect 226298 149080 226354 149116
rect 177630 114808 177686 114864
rect 177630 105424 177686 105480
rect 182506 83664 182562 83720
rect 155366 75524 155422 75560
rect 155366 75504 155368 75524
rect 155368 75504 155420 75524
rect 155420 75504 155422 75524
rect 139634 75232 139690 75288
rect 173858 75232 173914 75288
rect 172938 74144 172994 74200
rect 139818 73736 139874 73792
rect 139634 72512 139690 72568
rect 139726 71424 139782 71480
rect 139634 68296 139690 68352
rect 140002 71016 140058 71072
rect 139910 69520 139966 69576
rect 139726 67344 139782 67400
rect 139634 67072 139690 67128
rect 139910 65440 139966 65496
rect 139634 64216 139690 64272
rect 139726 63128 139782 63184
rect 139634 61360 139690 61416
rect 139818 62720 139874 62776
rect 139726 60000 139782 60056
rect 139726 58912 139782 58968
rect 139634 58640 139690 58696
rect 139634 57280 139690 57336
rect 139542 55920 139598 55976
rect 139634 54444 139690 54480
rect 139634 54424 139636 54444
rect 139636 54424 139688 54444
rect 139688 54424 139690 54444
rect 139634 53472 139690 53528
rect 173490 73192 173546 73248
rect 173490 72104 173546 72160
rect 173306 71036 173362 71072
rect 173306 71016 173308 71036
rect 173308 71016 173360 71036
rect 173360 71016 173362 71036
rect 173306 70084 173362 70120
rect 173306 70064 173308 70084
rect 173308 70064 173360 70084
rect 173360 70064 173362 70084
rect 173122 68976 173178 69032
rect 173674 67888 173730 67944
rect 173122 64896 173178 64952
rect 173122 61768 173178 61824
rect 172754 56600 172810 56656
rect 174042 66956 174098 66992
rect 174042 66936 174044 66956
rect 174044 66936 174096 66956
rect 174096 66936 174098 66956
rect 174042 65848 174098 65904
rect 173490 63808 173546 63864
rect 174042 62740 174098 62776
rect 174042 62720 174044 62740
rect 174044 62720 174096 62740
rect 174096 62720 174098 62740
rect 173490 60680 173546 60736
rect 174042 59592 174098 59648
rect 174042 58640 174098 58696
rect 173490 57552 173546 57608
rect 182322 69384 182378 69440
rect 226298 69384 226354 69440
rect 181678 68432 181734 68488
rect 226390 68432 226446 68488
rect 181402 67616 181458 67672
rect 226298 67616 226354 67672
rect 181034 66120 181090 66176
rect 181770 65848 181826 65904
rect 180850 65440 180906 65496
rect 181034 65440 181090 65496
rect 182322 64896 182378 64952
rect 181586 64080 181642 64136
rect 182322 63128 182378 63184
rect 182322 62312 182378 62368
rect 181586 61360 181642 61416
rect 181218 60408 181274 60464
rect 182322 59592 182378 59648
rect 181586 58640 181642 58696
rect 182322 57824 182378 57880
rect 182322 56484 182378 56520
rect 182322 56464 182324 56484
rect 182324 56464 182376 56484
rect 182376 56464 182378 56484
rect 181770 56056 181826 56112
rect 173398 55512 173454 55568
rect 174042 54444 174098 54480
rect 174042 54424 174044 54444
rect 174044 54424 174096 54444
rect 174096 54424 174098 54444
rect 181678 55104 181734 55160
rect 226298 66700 226300 66720
rect 226300 66700 226352 66720
rect 226352 66700 226354 66720
rect 226298 66664 226354 66700
rect 226298 65848 226354 65904
rect 226206 64896 226262 64952
rect 225930 64080 225986 64136
rect 225746 63128 225802 63184
rect 226298 62348 226300 62368
rect 226300 62348 226352 62368
rect 226352 62348 226354 62368
rect 226298 62312 226354 62348
rect 225930 61360 225986 61416
rect 226298 60408 226354 60464
rect 226114 59592 226170 59648
rect 226298 58640 226354 58696
rect 226298 57824 226354 57880
rect 226298 56908 226300 56928
rect 226300 56908 226352 56928
rect 226352 56908 226354 56928
rect 226298 56872 226354 56908
rect 225378 56056 225434 56112
rect 225378 55104 225434 55160
rect 182322 54288 182378 54344
rect 174042 53472 174098 53528
rect 142854 51024 142910 51080
rect 139726 50616 139782 50672
rect 139634 50344 139690 50400
rect 140554 48984 140610 49040
rect 140002 48032 140058 48088
rect 147730 48032 147786 48088
rect 153986 48032 154042 48088
rect 160058 47896 160114 47952
rect 163002 47216 163058 47272
rect 167602 48032 167658 48088
rect 166406 47760 166462 47816
rect 168890 47896 168946 47952
rect 168890 45992 168946 46048
rect 165946 45856 166002 45912
rect 163002 45720 163058 45776
rect 173950 51296 174006 51352
rect 174042 50344 174098 50400
rect 173306 49256 173362 49312
rect 181862 49256 181918 49312
rect 174042 48304 174098 48360
rect 169718 44788 169774 44824
rect 169718 44768 169720 44788
rect 169720 44768 169772 44788
rect 169772 44768 169774 44788
rect 88390 26000 88446 26056
rect 88022 23280 88078 23336
rect 182230 47896 182286 47952
rect 182138 46536 182194 46592
rect 181954 33616 182010 33672
rect 182046 30760 182102 30816
rect 182138 28040 182194 28096
rect 187290 50616 187346 50672
rect 191982 50344 192038 50400
rect 199066 50208 199122 50264
rect 203758 49256 203814 49312
rect 212038 53064 212094 53120
rect 207530 39056 207586 39112
rect 212590 43408 212646 43464
rect 226298 54324 226300 54344
rect 226300 54324 226352 54344
rect 226352 54324 226354 54344
rect 226298 54288 226354 54324
rect 230898 226328 230954 226384
rect 232002 304664 232058 304720
rect 232002 301536 232058 301592
rect 231450 279640 231506 279696
rect 231634 282804 231636 282824
rect 231636 282804 231688 282824
rect 231688 282804 231690 282824
rect 231634 282768 231690 282804
rect 231542 276512 231598 276568
rect 236050 289060 236052 289080
rect 236052 289060 236104 289080
rect 236104 289060 236106 289080
rect 236050 289024 236106 289060
rect 246170 316904 246226 316960
rect 253530 328736 253586 328792
rect 240650 310104 240706 310160
rect 240926 296776 240982 296832
rect 240926 283484 240928 283504
rect 240928 283484 240980 283504
rect 240980 283484 240982 283504
rect 240926 283448 240982 283484
rect 232738 274336 232794 274392
rect 231634 273384 231690 273440
rect 233474 263048 233530 263104
rect 233474 261688 233530 261744
rect 233474 260328 233530 260384
rect 233474 258832 233530 258888
rect 233474 257472 233530 257528
rect 233474 256112 233530 256168
rect 232738 254616 232794 254672
rect 232830 251896 232886 251952
rect 233474 250980 233476 251000
rect 233476 250980 233528 251000
rect 233528 250980 233530 251000
rect 233474 250944 233530 250980
rect 233474 249720 233530 249776
rect 234210 253256 234266 253312
rect 233566 248360 233622 248416
rect 233566 244144 233622 244200
rect 234302 246864 234358 246920
rect 234210 245504 234266 245560
rect 234118 242784 234174 242840
rect 233474 240628 233530 240664
rect 233474 240608 233476 240628
rect 233476 240608 233528 240628
rect 233528 240608 233530 240628
rect 233474 239268 233530 239304
rect 233474 239248 233476 239268
rect 233476 239248 233528 239268
rect 233528 239248 233530 239268
rect 233566 238568 233622 238624
rect 233474 237072 233530 237128
rect 231818 234896 231874 234952
rect 247918 274608 247974 274664
rect 247274 273692 247276 273712
rect 247276 273692 247328 273712
rect 247328 273692 247330 273712
rect 247274 273656 247330 273692
rect 250862 274336 250918 274392
rect 252058 274472 252114 274528
rect 250954 273792 251010 273848
rect 253346 274608 253402 274664
rect 261718 306160 261774 306216
rect 261718 286596 261774 286632
rect 261718 286576 261720 286596
rect 261720 286576 261772 286596
rect 261772 286576 261774 286596
rect 261442 274608 261498 274664
rect 261442 272160 261498 272216
rect 243778 236120 243834 236176
rect 247274 236120 247330 236176
rect 230990 223200 231046 223256
rect 230806 220072 230862 220128
rect 230714 216944 230770 217000
rect 230898 200624 230954 200680
rect 230714 198176 230770 198232
rect 230806 194368 230862 194424
rect 230714 104064 230770 104120
rect 231542 216944 231598 217000
rect 231450 207696 231506 207752
rect 231358 185664 231414 185720
rect 231726 213816 231782 213872
rect 231634 210688 231690 210744
rect 232002 204432 232058 204488
rect 235314 194524 235370 194560
rect 235314 194504 235316 194524
rect 235316 194504 235368 194524
rect 235368 194504 235370 194524
rect 231542 191920 231598 191976
rect 232002 188812 232058 188848
rect 241478 233536 241534 233592
rect 242490 235848 242546 235904
rect 245986 234216 246042 234272
rect 243042 233400 243098 233456
rect 262546 235712 262602 235768
rect 240926 216128 240982 216184
rect 240650 202800 240706 202856
rect 240926 189472 240982 189528
rect 232002 188792 232004 188812
rect 232004 188792 232056 188812
rect 232056 188792 232058 188812
rect 231450 182536 231506 182592
rect 230990 179408 231046 179464
rect 248930 183080 248986 183136
rect 249022 182128 249078 182184
rect 252702 180632 252758 180688
rect 252058 180496 252114 180552
rect 250862 180224 250918 180280
rect 250218 180088 250274 180144
rect 249574 179952 249630 180008
rect 253346 180768 253402 180824
rect 262362 212728 262418 212784
rect 263098 192736 263154 192792
rect 261074 182028 261076 182048
rect 261076 182028 261128 182048
rect 261128 182028 261130 182048
rect 261074 181992 261130 182028
rect 266594 357160 266650 357216
rect 266594 356072 266650 356128
rect 266594 355156 266596 355176
rect 266596 355156 266648 355176
rect 266648 355156 266650 355176
rect 266594 355120 266650 355156
rect 266686 354032 266742 354088
rect 266594 352944 266650 353000
rect 266594 351992 266650 352048
rect 274874 351312 274930 351368
rect 266594 350904 266650 350960
rect 266686 349816 266742 349872
rect 266594 348864 266650 348920
rect 284534 356480 284590 356536
rect 284534 351604 284590 351640
rect 284534 351584 284536 351604
rect 284536 351584 284588 351604
rect 284588 351584 284590 351604
rect 274874 350360 274930 350416
rect 274874 349544 274930 349600
rect 266594 347776 266650 347832
rect 274966 348592 275022 348648
rect 266594 346860 266596 346880
rect 266596 346860 266648 346880
rect 266648 346860 266650 346880
rect 266594 346824 266650 346860
rect 275058 347776 275114 347832
rect 266686 345736 266742 345792
rect 275150 346824 275206 346880
rect 275242 346008 275298 346064
rect 274874 345056 274930 345112
rect 266594 344648 266650 344704
rect 266594 343696 266650 343752
rect 275058 344240 275114 344296
rect 274966 343288 275022 343344
rect 266594 342644 266596 342664
rect 266596 342644 266648 342664
rect 266648 342644 266650 342664
rect 266594 342608 266650 342644
rect 266686 341520 266742 341576
rect 274874 341520 274930 341576
rect 266594 340568 266650 340624
rect 266594 339480 266650 339536
rect 266594 338548 266650 338584
rect 266594 338528 266596 338548
rect 266596 338528 266648 338548
rect 266648 338528 266650 338548
rect 266686 337440 266742 337496
rect 266594 336352 266650 336408
rect 266594 335400 266650 335456
rect 275150 342336 275206 342392
rect 275058 340568 275114 340624
rect 275058 339752 275114 339808
rect 274874 337984 274930 338040
rect 274874 337032 274930 337088
rect 266594 334312 266650 334368
rect 266686 333224 266742 333280
rect 274966 336216 275022 336272
rect 266594 332272 266650 332328
rect 275610 338800 275666 338856
rect 266594 331184 266650 331240
rect 266594 330232 266650 330288
rect 266594 256112 266650 256168
rect 266594 254616 266650 254672
rect 266594 253256 266650 253312
rect 266594 251896 266650 251952
rect 267146 249040 267202 249096
rect 266594 247680 266650 247736
rect 266594 246320 266650 246376
rect 266594 244824 266650 244880
rect 267514 263048 267570 263104
rect 267422 261688 267478 261744
rect 267330 258832 267386 258888
rect 267330 250536 267386 250592
rect 267606 260328 267662 260384
rect 267790 257472 267846 257528
rect 267882 243464 267938 243520
rect 267882 242104 267938 242160
rect 267882 240628 267938 240664
rect 267882 240608 267884 240628
rect 267884 240608 267936 240628
rect 267936 240608 267938 240628
rect 267882 239268 267938 239304
rect 267882 239248 267884 239268
rect 267884 239248 267936 239268
rect 267936 239248 267938 239268
rect 267514 237888 267570 237944
rect 267238 236528 267294 236584
rect 296218 333088 296274 333144
rect 292906 331592 292962 331648
rect 299530 331456 299586 331512
rect 292906 330776 292962 330832
rect 319126 382048 319182 382104
rect 319218 380144 319274 380200
rect 319310 377424 319366 377480
rect 319402 374704 319458 374760
rect 319310 333088 319366 333144
rect 320138 371848 320194 371904
rect 320598 351312 320654 351368
rect 321610 350360 321666 350416
rect 321702 349544 321758 349600
rect 321610 348592 321666 348648
rect 321058 347776 321114 347832
rect 320414 346824 320470 346880
rect 320506 346008 320562 346064
rect 321058 345056 321114 345112
rect 321610 344240 321666 344296
rect 321610 343288 321666 343344
rect 321058 342336 321114 342392
rect 321610 341540 321666 341576
rect 321610 341520 321612 341540
rect 321612 341520 321664 341540
rect 321664 341520 321666 341540
rect 320598 340568 320654 340624
rect 321242 339752 321298 339808
rect 321610 338820 321666 338856
rect 321610 338800 321612 338820
rect 321612 338800 321664 338820
rect 321664 338800 321666 338820
rect 321610 337984 321666 338040
rect 321426 337032 321482 337088
rect 321610 336216 321666 336272
rect 319402 331592 319458 331648
rect 270274 313504 270330 313560
rect 269354 296776 269410 296832
rect 270274 280184 270330 280240
rect 276438 269440 276494 269496
rect 274874 257336 274930 257392
rect 321242 257336 321298 257392
rect 275058 256384 275114 256440
rect 321058 256384 321114 256440
rect 274414 254616 274470 254672
rect 274138 250264 274194 250320
rect 274322 252848 274378 252904
rect 274874 253800 274930 253856
rect 274874 249992 274930 250048
rect 274874 248804 274876 248824
rect 274876 248804 274928 248824
rect 274928 248804 274930 248824
rect 274874 248768 274930 248804
rect 275610 252032 275666 252088
rect 275518 251080 275574 251136
rect 274966 248224 275022 248280
rect 274874 247272 274930 247328
rect 274874 246048 274930 246104
rect 274874 244724 274876 244744
rect 274876 244724 274928 244744
rect 274928 244724 274930 244744
rect 274874 244688 274930 244724
rect 274230 243056 274286 243112
rect 275886 255568 275942 255624
rect 320874 255604 320876 255624
rect 320876 255604 320928 255624
rect 320928 255604 320930 255624
rect 320874 255568 320930 255604
rect 320690 254616 320746 254672
rect 321610 253800 321666 253856
rect 321610 252848 321666 252904
rect 321610 252052 321666 252088
rect 321610 252032 321612 252052
rect 321612 252032 321664 252052
rect 321664 252032 321666 252052
rect 320598 251080 320654 251136
rect 321058 250264 321114 250320
rect 321610 249312 321666 249368
rect 321610 248360 321666 248416
rect 321794 247564 321850 247600
rect 321794 247544 321796 247564
rect 321796 247544 321848 247564
rect 321848 247544 321850 247564
rect 321242 246592 321298 246648
rect 321610 245776 321666 245832
rect 275702 245504 275758 245560
rect 321702 244860 321704 244880
rect 321704 244860 321756 244880
rect 321756 244860 321758 244880
rect 321702 244824 321758 244860
rect 321610 244008 321666 244064
rect 321610 243056 321666 243112
rect 275794 242920 275850 242976
rect 320506 242240 320562 242296
rect 283246 239384 283302 239440
rect 290514 239656 290570 239712
rect 286926 238296 286982 238352
rect 305142 240336 305198 240392
rect 301462 234896 301518 234952
rect 302014 234896 302070 234952
rect 273954 226600 274010 226656
rect 272942 219528 272998 219584
rect 272942 202800 272998 202856
rect 272942 186208 272998 186264
rect 267514 181176 267570 181232
rect 233474 169072 233530 169128
rect 233474 167712 233530 167768
rect 233474 166352 233530 166408
rect 233474 164856 233530 164912
rect 267146 164856 267202 164912
rect 233474 163496 233530 163552
rect 233474 162156 233530 162192
rect 233474 162136 233476 162156
rect 233476 162136 233528 162156
rect 233528 162136 233530 162156
rect 267054 162136 267110 162192
rect 232738 160640 232794 160696
rect 233474 159300 233530 159336
rect 233474 159280 233476 159300
rect 233476 159280 233528 159300
rect 233528 159280 233530 159300
rect 234118 157920 234174 157976
rect 233474 156560 233530 156616
rect 233474 155084 233530 155120
rect 233474 155064 233476 155084
rect 233476 155064 233528 155084
rect 233528 155064 233530 155084
rect 233474 150884 233476 150904
rect 233476 150884 233528 150904
rect 233528 150884 233530 150904
rect 233474 150848 233530 150884
rect 266594 160660 266650 160696
rect 266594 160640 266596 160660
rect 266596 160640 266648 160660
rect 266648 160640 266650 160660
rect 266594 159316 266596 159336
rect 266596 159316 266648 159336
rect 266648 159316 266650 159336
rect 266594 159280 266650 159316
rect 266594 157956 266596 157976
rect 266596 157956 266648 157976
rect 266648 157956 266650 157976
rect 266594 157920 266650 157956
rect 266594 155064 266650 155120
rect 234578 153704 234634 153760
rect 266686 153704 266742 153760
rect 234302 152344 234358 152400
rect 266594 152344 266650 152400
rect 266594 150884 266596 150904
rect 266596 150884 266648 150904
rect 266648 150884 266650 150904
rect 266594 150848 266650 150884
rect 233474 149488 233530 149544
rect 266594 149524 266596 149544
rect 266596 149524 266648 149544
rect 266648 149524 266650 149544
rect 266594 149488 266650 149524
rect 233474 148164 233476 148184
rect 233476 148164 233528 148184
rect 233528 148164 233530 148184
rect 233474 148128 233530 148164
rect 266962 148128 267018 148184
rect 233474 146632 233530 146688
rect 233474 145272 233530 145328
rect 266778 145272 266834 145328
rect 233474 143912 233530 143968
rect 230990 143096 231046 143152
rect 267422 169072 267478 169128
rect 267330 156560 267386 156616
rect 267238 142552 267294 142608
rect 242490 142144 242546 142200
rect 246814 142144 246870 142200
rect 231082 139968 231138 140024
rect 230990 132896 231046 132952
rect 233474 142028 233530 142064
rect 233474 142008 233476 142028
rect 233476 142008 233528 142028
rect 233528 142008 233530 142028
rect 231450 140512 231506 140568
rect 231358 139696 231414 139752
rect 231358 138608 231414 138664
rect 232002 138608 232058 138664
rect 231266 129768 231322 129824
rect 231082 125960 231138 126016
rect 230990 120384 231046 120440
rect 230898 107328 230954 107384
rect 230806 101616 230862 101672
rect 243410 142008 243466 142064
rect 267606 167712 267662 167768
rect 267514 166352 267570 166408
rect 267882 163496 267938 163552
rect 274874 163396 274876 163416
rect 274876 163396 274928 163416
rect 274928 163396 274930 163416
rect 274874 163360 274930 163396
rect 321610 163360 321666 163416
rect 275058 162408 275114 162464
rect 321610 162428 321666 162464
rect 321610 162408 321612 162428
rect 321612 162408 321664 162428
rect 321664 162408 321666 162428
rect 274874 158872 274930 158928
rect 274966 156288 275022 156344
rect 274874 156016 274930 156072
rect 275150 161592 275206 161648
rect 321610 161592 321666 161648
rect 275794 160640 275850 160696
rect 321058 160640 321114 160696
rect 275150 159824 275206 159880
rect 275518 158056 275574 158112
rect 274874 154964 274876 154984
rect 274876 154964 274928 154984
rect 274928 154964 274930 154984
rect 274874 154928 274930 154964
rect 274874 153604 274876 153624
rect 274876 153604 274928 153624
rect 274928 153604 274930 153624
rect 274874 153568 274930 153604
rect 274966 153296 275022 153352
rect 274874 152072 274930 152128
rect 274874 150868 274930 150904
rect 274874 150848 274876 150868
rect 274876 150848 274928 150868
rect 274928 150848 274930 150868
rect 274966 150576 275022 150632
rect 274874 148808 274930 148864
rect 275610 157104 275666 157160
rect 267882 146632 267938 146688
rect 320598 159824 320654 159880
rect 321058 158872 321114 158928
rect 321610 158056 321666 158112
rect 321610 157140 321612 157160
rect 321612 157140 321664 157160
rect 321664 157140 321666 157160
rect 321610 157104 321666 157140
rect 321058 156288 321114 156344
rect 321610 155336 321666 155392
rect 320874 154384 320930 154440
rect 321610 153568 321666 153624
rect 320506 152616 320562 152672
rect 320782 151800 320838 151856
rect 321702 150848 321758 150904
rect 321610 150032 321666 150088
rect 275702 149488 275758 149544
rect 321058 149080 321114 149136
rect 321610 148264 321666 148320
rect 267790 143912 267846 143968
rect 243042 140512 243098 140568
rect 243778 139696 243834 139752
rect 232002 122560 232058 122616
rect 231358 98216 231414 98272
rect 230714 95360 230770 95416
rect 230714 94816 230770 94872
rect 246170 139832 246226 139888
rect 246446 139832 246502 139888
rect 245342 139560 245398 139616
rect 246446 130212 246448 130232
rect 246448 130212 246500 130232
rect 246500 130212 246502 130232
rect 246446 130176 246502 130212
rect 249114 138472 249170 138528
rect 249114 137248 249170 137304
rect 249666 134256 249722 134312
rect 249666 133032 249722 133088
rect 240374 122152 240430 122208
rect 231634 110900 231636 110920
rect 231636 110900 231688 110920
rect 231688 110900 231690 110920
rect 231634 110864 231690 110900
rect 240098 109776 240154 109832
rect 240374 108824 240430 108880
rect 231450 92232 231506 92288
rect 231818 94988 231820 95008
rect 231820 94988 231872 95008
rect 231872 94988 231874 95008
rect 231818 94952 231874 94988
rect 231542 88832 231598 88888
rect 230990 85704 231046 85760
rect 240374 95496 240430 95552
rect 248930 89104 248986 89160
rect 242582 85840 242638 85896
rect 242582 76456 242638 76512
rect 249574 88832 249630 88888
rect 249114 88424 249170 88480
rect 252150 88016 252206 88072
rect 252058 86792 252114 86848
rect 250862 86656 250918 86712
rect 252150 86112 252206 86168
rect 253070 86928 253126 86984
rect 290514 142416 290570 142472
rect 290974 142416 291030 142472
rect 285914 138472 285970 138528
rect 287202 138472 287258 138528
rect 294194 144592 294250 144648
rect 297782 143096 297838 143152
rect 303854 143776 303910 143832
rect 301094 141056 301150 141112
rect 302014 141056 302070 141112
rect 283154 134256 283210 134312
rect 270366 125416 270422 125472
rect 260338 122560 260394 122616
rect 261166 118752 261222 118808
rect 263098 98760 263154 98816
rect 260062 87508 260064 87528
rect 260064 87508 260116 87528
rect 260116 87508 260118 87528
rect 260062 87472 260118 87508
rect 260338 87472 260394 87528
rect 268618 108824 268674 108880
rect 270366 92232 270422 92288
rect 249206 75504 249262 75560
rect 233474 75232 233530 75288
rect 266594 75232 266650 75288
rect 267422 74144 267478 74200
rect 233934 73872 233990 73928
rect 233474 72512 233530 72568
rect 233474 71424 233530 71480
rect 233750 71016 233806 71072
rect 233566 69656 233622 69712
rect 233658 68296 233714 68352
rect 233566 67208 233622 67264
rect 233474 66936 233530 66992
rect 233474 65460 233530 65496
rect 233474 65440 233476 65460
rect 233476 65440 233528 65460
rect 233528 65440 233530 65460
rect 234578 64488 234634 64544
rect 233474 63128 233530 63184
rect 233566 62720 233622 62776
rect 233474 61360 233530 61416
rect 233658 60000 233714 60056
rect 233566 58912 233622 58968
rect 233474 58640 233530 58696
rect 233474 57144 233530 57200
rect 234394 55920 234450 55976
rect 233474 55240 233530 55296
rect 233474 54444 233530 54480
rect 233474 54424 233476 54444
rect 233476 54424 233528 54444
rect 233528 54424 233530 54444
rect 233474 53472 233530 53528
rect 233566 50752 233622 50808
rect 233474 50344 233530 50400
rect 233474 48984 233530 49040
rect 266594 73192 266650 73248
rect 266686 72104 266742 72160
rect 266594 71016 266650 71072
rect 266594 70064 266650 70120
rect 266594 68976 266650 69032
rect 266686 67888 266742 67944
rect 266594 66936 266650 66992
rect 266594 65848 266650 65904
rect 266594 64896 266650 64952
rect 266686 63808 266742 63864
rect 266594 62720 266650 62776
rect 266594 61768 266650 61824
rect 266594 60680 266650 60736
rect 266686 59592 266742 59648
rect 266594 58660 266650 58696
rect 266594 58640 266596 58660
rect 266596 58640 266648 58660
rect 266648 58640 266650 58660
rect 266594 57552 266650 57608
rect 266594 56600 266650 56656
rect 274874 69384 274930 69440
rect 321610 69384 321666 69440
rect 274966 68432 275022 68488
rect 321610 68432 321666 68488
rect 274782 67616 274838 67672
rect 274690 66664 274746 66720
rect 274874 65848 274930 65904
rect 274874 64080 274930 64136
rect 274874 63128 274930 63184
rect 275058 64896 275114 64952
rect 274966 62312 275022 62368
rect 274874 61360 274930 61416
rect 274874 60408 274930 60464
rect 274874 58640 274930 58696
rect 275058 59592 275114 59648
rect 274966 57824 275022 57880
rect 274874 56872 274930 56928
rect 267238 55512 267294 55568
rect 266594 54444 266650 54480
rect 266594 54424 266596 54444
rect 266596 54424 266648 54444
rect 266648 54424 266650 54444
rect 275058 56056 275114 56112
rect 274966 55104 275022 55160
rect 320506 67616 320562 67672
rect 321426 66664 321482 66720
rect 321610 65868 321666 65904
rect 321610 65848 321612 65868
rect 321612 65848 321664 65868
rect 321664 65848 321666 65868
rect 321610 64896 321666 64952
rect 321426 64080 321482 64136
rect 321058 63128 321114 63184
rect 321702 62312 321758 62368
rect 321242 61360 321298 61416
rect 320874 60408 320930 60464
rect 321610 59592 321666 59648
rect 321058 58640 321114 58696
rect 320874 57824 320930 57880
rect 321058 56872 321114 56928
rect 321610 56056 321666 56112
rect 321610 55104 321666 55160
rect 274874 54324 274876 54344
rect 274876 54324 274928 54344
rect 274928 54324 274930 54344
rect 274874 54288 274930 54324
rect 266594 53472 266650 53528
rect 266686 51296 266742 51352
rect 266594 50344 266650 50400
rect 274966 49936 275022 49992
rect 266594 49256 266650 49312
rect 275058 49256 275114 49312
rect 266594 48304 266650 48360
rect 241110 48032 241166 48088
rect 262914 48032 262970 48088
rect 264478 48032 264534 48088
rect 233474 47760 233530 47816
rect 244882 47896 244938 47952
rect 248010 47216 248066 47272
rect 253990 47896 254046 47952
rect 260338 46536 260394 46592
rect 256934 45992 256990 46048
rect 263190 45992 263246 46048
rect 251138 45720 251194 45776
rect 182230 26000 182286 26056
rect 181862 23280 181918 23336
rect 275794 47896 275850 47952
rect 275886 46536 275942 46592
rect 275794 33616 275850 33672
rect 275886 30760 275942 30816
rect 275978 28040 276034 28096
rect 281314 50616 281370 50672
rect 283706 48032 283762 48088
rect 285914 47372 285970 47408
rect 285914 47352 285916 47372
rect 285916 47352 285968 47372
rect 285968 47352 285970 47372
rect 306982 53336 307038 53392
rect 301554 39056 301610 39112
rect 306614 37696 306670 37752
rect 320966 54324 320968 54344
rect 320968 54324 321020 54344
rect 321020 54324 321022 54344
rect 320966 54288 321022 54324
rect 276070 26000 276126 26056
rect 275610 23280 275666 23336
rect 88482 20696 88538 20752
rect 182322 20696 182378 20752
rect 276162 20696 276218 20752
rect 12674 14204 12676 14224
rect 12676 14204 12728 14224
rect 12728 14204 12730 14224
rect 12674 14168 12730 14204
rect 328418 357432 328474 357488
rect 328326 356072 328382 356128
rect 328418 355156 328420 355176
rect 328420 355156 328472 355176
rect 328472 355156 328474 355176
rect 328418 355120 328474 355156
rect 328510 354576 328566 354632
rect 328050 353352 328106 353408
rect 328510 352264 328566 352320
rect 327498 350904 327554 350960
rect 327866 350360 327922 350416
rect 328142 349544 328198 349600
rect 328326 348184 328382 348240
rect 327222 346824 327278 346880
rect 327130 346416 327186 346472
rect 328050 345056 328106 345112
rect 328510 343968 328566 344024
rect 327038 342608 327094 342664
rect 326854 341248 326910 341304
rect 328050 342064 328106 342120
rect 327130 339888 327186 339944
rect 327038 338120 327094 338176
rect 326946 337032 327002 337088
rect 326670 334312 326726 334368
rect 327222 338528 327278 338584
rect 327130 335808 327186 335864
rect 327038 333904 327094 333960
rect 324554 326832 324610 326888
rect 324738 320304 324794 320360
rect 324830 317176 324886 317232
rect 324646 315136 324702 315192
rect 324646 314048 324702 314104
rect 324738 308200 324794 308256
rect 324554 301536 324610 301592
rect 324646 298408 324702 298464
rect 324554 282788 324610 282824
rect 324554 282768 324556 282788
rect 324556 282768 324608 282788
rect 324608 282768 324610 282788
rect 327314 332952 327370 333008
rect 327222 331592 327278 331648
rect 325382 310920 325438 310976
rect 325290 304664 325346 304720
rect 324830 293376 324886 293432
rect 325198 293376 325254 293432
rect 324738 250264 324794 250320
rect 322990 226328 323046 226384
rect 323174 124056 323230 124112
rect 323174 122900 323230 122956
rect 324738 223200 324794 223256
rect 324554 220072 324610 220128
rect 325290 285896 325346 285952
rect 325198 273384 325254 273440
rect 325198 238976 325254 239032
rect 324830 198720 324886 198776
rect 324554 188792 324610 188848
rect 324554 179444 324556 179464
rect 324556 179444 324608 179464
rect 324608 179444 324610 179464
rect 324554 179408 324610 179444
rect 324646 132352 324702 132408
rect 324554 119876 324556 119896
rect 324556 119876 324608 119896
rect 324608 119876 324610 119896
rect 324554 119840 324610 119876
rect 324554 113584 324610 113640
rect 324646 106784 324702 106840
rect 324554 104064 324610 104120
rect 324646 100936 324702 100992
rect 328418 330232 328474 330288
rect 325566 308200 325622 308256
rect 325474 298408 325530 298464
rect 325382 279640 325438 279696
rect 325474 276512 325530 276568
rect 325658 234352 325714 234408
rect 325382 224308 325438 224344
rect 325382 224288 325384 224308
rect 325384 224288 325436 224308
rect 325436 224288 325438 224308
rect 339182 327376 339238 327432
rect 340010 327376 340066 327432
rect 342494 326832 342550 326888
rect 345622 316632 345678 316688
rect 352890 324792 352946 324848
rect 353074 324792 353130 324848
rect 348106 320168 348162 320224
rect 334214 309716 334270 309752
rect 334214 309696 334216 309716
rect 334216 309696 334268 309716
rect 334268 309696 334270 309716
rect 334214 296232 334270 296288
rect 334214 283584 334270 283640
rect 327314 263592 327370 263648
rect 352062 266720 352118 266776
rect 350958 266584 351014 266640
rect 353718 285216 353774 285272
rect 356202 314048 356258 314104
rect 356202 308608 356258 308664
rect 356202 304140 356258 304176
rect 356202 304120 356204 304140
rect 356204 304120 356256 304140
rect 356256 304120 356258 304140
rect 356202 298816 356258 298872
rect 356202 293804 356258 293840
rect 356202 293784 356204 293804
rect 356204 293784 356256 293804
rect 356256 293784 356258 293804
rect 356202 289024 356258 289080
rect 356202 283720 356258 283776
rect 356202 279368 356258 279424
rect 327222 261688 327278 261744
rect 326762 260328 326818 260384
rect 328418 258832 328474 258888
rect 327222 257472 327278 257528
rect 328050 256112 328106 256168
rect 328418 254616 328474 254672
rect 327222 253256 327278 253312
rect 327130 251896 327186 251952
rect 327222 250536 327278 250592
rect 328418 249076 328420 249096
rect 328420 249076 328472 249096
rect 328472 249076 328474 249096
rect 328418 249040 328474 249076
rect 328418 247700 328474 247736
rect 328418 247680 328420 247700
rect 328420 247680 328472 247700
rect 328472 247680 328474 247700
rect 328418 246864 328474 246920
rect 327866 245504 327922 245560
rect 327866 244008 327922 244064
rect 327866 242648 327922 242704
rect 327038 240608 327094 240664
rect 327222 239248 327278 239304
rect 327130 238568 327186 238624
rect 328418 236564 328420 236584
rect 328420 236564 328472 236584
rect 328472 236564 328474 236584
rect 328418 236528 328474 236564
rect 325566 210688 325622 210744
rect 325842 216672 325898 216728
rect 325750 213816 325806 213872
rect 325658 207560 325714 207616
rect 325474 204432 325530 204488
rect 325382 191920 325438 191976
rect 325290 185664 325346 185720
rect 341298 224852 341354 224888
rect 341298 224832 341300 224852
rect 341300 224832 341352 224852
rect 341352 224832 341354 224852
rect 342678 224832 342734 224888
rect 345714 225376 345770 225432
rect 350958 232448 351014 232504
rect 352062 232448 352118 232504
rect 334214 216128 334270 216184
rect 334214 202800 334270 202856
rect 334214 189472 334270 189528
rect 325474 182536 325530 182592
rect 350958 172880 351014 172936
rect 352062 172880 352118 172936
rect 352890 191376 352946 191432
rect 352798 184032 352854 184088
rect 352890 182128 352946 182184
rect 352982 181992 353038 182048
rect 355098 220208 355154 220264
rect 357674 221976 357730 222032
rect 356294 215856 356350 215912
rect 356202 215176 356258 215232
rect 356018 210144 356074 210200
rect 356202 205248 356258 205304
rect 355926 200216 355982 200272
rect 356202 195184 356258 195240
rect 355190 190152 355246 190208
rect 356202 185256 356258 185312
rect 328418 169072 328474 169128
rect 327222 167712 327278 167768
rect 327498 166352 327554 166408
rect 327222 163360 327278 163416
rect 328418 164856 328474 164912
rect 327314 162136 327370 162192
rect 327406 160640 327462 160696
rect 327222 159280 327278 159336
rect 327222 157920 327278 157976
rect 327222 156560 327278 156616
rect 328418 155084 328474 155120
rect 328418 155064 328420 155084
rect 328420 155064 328472 155084
rect 328472 155064 328474 155084
rect 328418 153740 328420 153760
rect 328420 153740 328472 153760
rect 328472 153740 328474 153760
rect 328418 153704 328474 153740
rect 328234 152344 328290 152400
rect 328418 150884 328420 150904
rect 328420 150884 328472 150904
rect 328472 150884 328474 150904
rect 328418 150848 328474 150884
rect 328418 149524 328420 149544
rect 328420 149524 328472 149544
rect 328472 149524 328474 149544
rect 328418 149488 328474 149524
rect 327222 146632 327278 146688
rect 328418 148164 328420 148184
rect 328420 148164 328472 148184
rect 328472 148164 328474 148184
rect 328418 148128 328474 148164
rect 328510 145272 328566 145328
rect 328326 143912 328382 143968
rect 328418 142008 328474 142064
rect 325474 129768 325530 129824
rect 325382 125960 325438 126016
rect 325290 110864 325346 110920
rect 325290 100392 325346 100448
rect 325198 98216 325254 98272
rect 324554 94408 324610 94464
rect 324554 85568 324610 85624
rect 325474 117256 325530 117312
rect 325382 92232 325438 92288
rect 325842 94700 325898 94736
rect 325842 94680 325844 94700
rect 325844 94680 325896 94700
rect 325896 94680 325898 94700
rect 325566 88832 325622 88888
rect 350958 139560 351014 139616
rect 352062 139560 352118 139616
rect 334214 122152 334270 122208
rect 334214 108824 334270 108880
rect 352798 105152 352854 105208
rect 334214 95496 334270 95552
rect 327038 73872 327094 73928
rect 326854 71016 326910 71072
rect 326946 69520 327002 69576
rect 327130 71424 327186 71480
rect 327038 68296 327094 68352
rect 350958 77816 351014 77872
rect 352062 77816 352118 77872
rect 352798 97536 352854 97592
rect 352798 90056 352854 90112
rect 356202 126232 356258 126288
rect 356202 121200 356258 121256
rect 356202 116168 356258 116224
rect 356202 111272 356258 111328
rect 356202 106240 356258 106296
rect 356202 101208 356258 101264
rect 356202 96176 356258 96232
rect 356202 91280 356258 91336
rect 328418 75232 328474 75288
rect 327866 72512 327922 72568
rect 327682 67208 327738 67264
rect 328418 66936 328474 66992
rect 328418 65848 328474 65904
rect 327314 64488 327370 64544
rect 328050 63128 328106 63184
rect 328326 62720 328382 62776
rect 328510 61496 328566 61552
rect 328418 60000 328474 60056
rect 327682 58640 327738 58696
rect 328510 58912 328566 58968
rect 328326 57144 328382 57200
rect 327498 56192 327554 56248
rect 328510 55240 328566 55296
rect 360802 262232 360858 262288
rect 360526 259104 360582 259160
rect 360618 255976 360674 256032
rect 361170 252848 361226 252904
rect 361446 249720 361502 249776
rect 360710 246592 360766 246648
rect 360618 243464 360674 243520
rect 360802 240336 360858 240392
rect 361170 237344 361226 237400
rect 360434 168256 360490 168312
rect 360526 165128 360582 165184
rect 360618 162000 360674 162056
rect 360710 158872 360766 158928
rect 360894 155744 360950 155800
rect 360802 152616 360858 152672
rect 360986 149488 361042 149544
rect 361170 168256 361226 168312
rect 361722 165128 361778 165184
rect 361722 162000 361778 162056
rect 361722 158872 361778 158928
rect 361722 155764 361778 155800
rect 361722 155744 361724 155764
rect 361724 155744 361776 155764
rect 361776 155744 361778 155764
rect 361170 146360 361226 146416
rect 361078 143368 361134 143424
rect 328418 54444 328474 54480
rect 328418 54424 328420 54444
rect 328420 54424 328472 54444
rect 328472 54424 328474 54444
rect 328418 53472 328474 53528
rect 327682 50888 327738 50944
rect 328418 50344 328474 50400
rect 327222 49936 327278 49992
rect 328510 48984 328566 49040
rect 360434 87336 360490 87392
rect 328050 47896 328106 47952
rect 346634 45992 346690 46048
rect 338354 45312 338410 45368
rect 429434 390616 429490 390672
rect 429434 378512 429490 378568
rect 429434 366408 429490 366464
rect 429434 354304 429490 354360
rect 369174 236528 369230 236584
rect 368714 234080 368770 234136
rect 368714 233692 368770 233728
rect 368714 233672 368716 233692
rect 368716 233672 368768 233692
rect 368768 233672 368770 233692
rect 368806 233400 368862 233456
rect 368898 232992 368954 233048
rect 368714 232176 368770 232232
rect 368806 231768 368862 231824
rect 368898 231360 368954 231416
rect 368806 230952 368862 231008
rect 368714 230544 368770 230600
rect 368898 230136 368954 230192
rect 368714 229456 368770 229512
rect 368806 229048 368862 229104
rect 368714 228640 368770 228696
rect 368714 228268 368716 228288
rect 368716 228268 368768 228288
rect 368768 228268 368770 228288
rect 368714 228232 368770 228268
rect 368806 227416 368862 227472
rect 368714 227008 368770 227064
rect 368990 226464 369046 226520
rect 368898 226328 368954 226384
rect 368806 225920 368862 225976
rect 368714 225548 368716 225568
rect 368716 225548 368768 225568
rect 368768 225548 368770 225568
rect 368714 225512 368770 225548
rect 368806 225104 368862 225160
rect 368714 224696 368770 224752
rect 368806 223880 368862 223936
rect 368714 223200 368770 223256
rect 368990 223472 369046 223528
rect 368898 222792 368954 222848
rect 368806 222384 368862 222440
rect 368714 221568 368770 221624
rect 368898 221976 368954 222032
rect 368898 221160 368954 221216
rect 368806 220752 368862 220808
rect 368714 220344 368770 220400
rect 368714 219664 368770 219720
rect 368806 218848 368862 218904
rect 368714 218032 368770 218088
rect 368806 217216 368862 217272
rect 368714 216400 368770 216456
rect 368806 216128 368862 216184
rect 368714 215740 368770 215776
rect 368714 215720 368716 215740
rect 368716 215720 368768 215740
rect 368768 215720 368770 215740
rect 368806 214904 368862 214960
rect 369082 219256 369138 219312
rect 369450 236120 369506 236176
rect 369266 224288 369322 224344
rect 368990 217624 369046 217680
rect 369082 216944 369138 217000
rect 369082 216844 369084 216864
rect 369084 216844 369136 216864
rect 369136 216844 369138 216864
rect 369082 216808 369138 216844
rect 368990 216536 369046 216592
rect 368714 213680 368770 213736
rect 368714 213036 368716 213056
rect 368716 213036 368768 213056
rect 368768 213036 368770 213056
rect 368714 213000 368770 213036
rect 369082 215312 369138 215368
rect 368990 214496 369046 214552
rect 368898 214088 368954 214144
rect 368898 213272 368954 213328
rect 369266 218440 369322 218496
rect 369634 235712 369690 235768
rect 369542 229864 369598 229920
rect 369542 227824 369598 227880
rect 369818 235304 369874 235360
rect 369726 232584 369782 232640
rect 429434 342200 429490 342256
rect 429434 330096 429490 330152
rect 429434 317856 429490 317912
rect 405974 315852 405976 315872
rect 405976 315852 406028 315872
rect 406028 315852 406030 315872
rect 405974 315816 406030 315852
rect 427318 313776 427374 313832
rect 405974 313640 406030 313696
rect 405974 310376 406030 310432
rect 405974 308236 405976 308256
rect 405976 308236 406028 308256
rect 406028 308236 406030 308256
rect 405974 308200 406030 308236
rect 406066 306196 406068 306216
rect 406068 306196 406120 306216
rect 406120 306196 406122 306216
rect 406066 306160 406122 306196
rect 405974 303576 406030 303632
rect 405974 300448 406030 300504
rect 405974 298272 406030 298328
rect 405974 295416 406030 295472
rect 405974 293648 406030 293704
rect 405974 290656 406030 290712
rect 405974 288616 406030 288672
rect 405974 285508 406030 285544
rect 405974 285488 405976 285508
rect 405976 285488 406028 285508
rect 406028 285488 406030 285508
rect 405974 283312 406030 283368
rect 405974 278688 406030 278744
rect 415266 277192 415322 277248
rect 395118 269712 395174 269768
rect 395394 269712 395450 269768
rect 414254 273792 414310 273848
rect 415542 273792 415598 273848
rect 370002 234896 370058 234952
rect 369910 234488 369966 234544
rect 369726 226600 369782 226656
rect 369818 219936 369874 219992
rect 369818 115216 369874 115272
rect 369910 115080 369966 115136
rect 369910 105560 369966 105616
rect 369818 105424 369874 105480
rect 405974 218712 406030 218768
rect 405974 214108 406030 214144
rect 405974 214088 405976 214108
rect 405976 214088 406028 214108
rect 406028 214088 406030 214108
rect 405974 210980 406030 211016
rect 405974 210960 405976 210980
rect 405976 210960 406028 210980
rect 406028 210960 406030 210980
rect 405974 209464 406030 209520
rect 428698 308608 428754 308664
rect 427410 304120 427466 304176
rect 427502 298680 427558 298736
rect 427870 293648 427926 293704
rect 427594 289024 427650 289080
rect 427962 283604 428018 283640
rect 427962 283584 427964 283604
rect 427964 283584 428016 283604
rect 428016 283584 428018 283604
rect 427686 279368 427742 279424
rect 429894 293648 429950 293704
rect 429434 281544 429490 281600
rect 429434 269440 429490 269496
rect 428790 257336 428846 257392
rect 429434 245096 429490 245152
rect 429802 232992 429858 233048
rect 428698 220888 428754 220944
rect 427410 220208 427466 220264
rect 405974 206780 405976 206800
rect 405976 206780 406028 206800
rect 406028 206780 406030 206800
rect 405974 206744 406030 206780
rect 427318 205248 427374 205304
rect 406066 204568 406122 204624
rect 405974 201324 406030 201360
rect 405974 201304 405976 201324
rect 405976 201304 406028 201324
rect 406028 201304 406030 201324
rect 427134 200216 427190 200272
rect 405974 199128 406030 199184
rect 405974 195864 406030 195920
rect 406066 194504 406122 194560
rect 405974 191668 406030 191704
rect 405974 191648 405976 191668
rect 405976 191648 406028 191668
rect 406028 191648 406030 191668
rect 426858 190152 426914 190208
rect 405974 189472 406030 189528
rect 405974 186208 406030 186264
rect 405974 183896 406030 183952
rect 405974 126912 406030 126968
rect 427318 126232 427374 126288
rect 405974 125552 406030 125608
rect 405974 122596 405976 122616
rect 405976 122596 406028 122616
rect 406028 122596 406030 122616
rect 405974 122560 406030 122596
rect 405974 120556 405976 120576
rect 405976 120556 406028 120576
rect 406028 120556 406030 120576
rect 405974 120520 406030 120556
rect 405974 117392 406030 117448
rect 405974 114808 406030 114864
rect 405974 112632 406030 112688
rect 406066 110592 406122 110648
rect 405974 107600 406030 107656
rect 405974 105288 406030 105344
rect 405974 102160 406030 102216
rect 405974 100564 405976 100584
rect 405976 100564 406028 100584
rect 406028 100564 406030 100584
rect 405974 100528 406030 100564
rect 405974 97672 406030 97728
rect 427226 96176 427282 96232
rect 405974 95496 406030 95552
rect 405974 92368 406030 92424
rect 405974 90212 406030 90248
rect 405974 90192 405976 90212
rect 405976 90192 406028 90212
rect 406028 90192 406030 90212
rect 415542 87336 415598 87392
rect 428698 215176 428754 215232
rect 427502 210144 427558 210200
rect 427594 195184 427650 195240
rect 427686 185392 427742 185448
rect 429618 208820 429620 208840
rect 429620 208820 429672 208840
rect 429672 208820 429674 208840
rect 429618 208784 429674 208820
rect 429526 196680 429582 196736
rect 429342 184576 429398 184632
rect 429894 172472 429950 172528
rect 428790 160232 428846 160288
rect 429434 148164 429436 148184
rect 429436 148164 429488 148184
rect 429488 148164 429490 148184
rect 429434 148128 429490 148164
rect 429434 136024 429490 136080
rect 428698 123920 428754 123976
rect 427502 121200 427558 121256
rect 427410 101208 427466 101264
rect 428698 116168 428754 116224
rect 427594 111272 427650 111328
rect 427686 106240 427742 106296
rect 427686 91552 427742 91608
rect 429434 111816 429490 111872
rect 429434 99712 429490 99768
rect 429434 75368 429490 75424
rect 430170 87472 430226 87528
rect 430078 63264 430134 63320
rect 429802 51160 429858 51216
rect 428698 39056 428754 39112
rect 429434 26952 429490 27008
rect 429434 14848 429490 14904
<< metal3 >>
rect 341702 393740 341708 393804
rect 341772 393802 341778 393804
rect 341937 393802 342003 393805
rect 341772 393800 342003 393802
rect 341772 393744 341942 393800
rect 341998 393744 342003 393800
rect 341772 393742 342003 393744
rect 341772 393740 341778 393742
rect 341937 393739 342003 393742
rect 9896 391354 10376 391384
rect 13129 391354 13195 391357
rect 9896 391352 13195 391354
rect 9896 391296 13134 391352
rect 13190 391296 13195 391352
rect 9896 391294 13195 391296
rect 9896 391264 10376 391294
rect 13129 391291 13195 391294
rect 429429 390674 429495 390677
rect 434416 390674 434896 390704
rect 429429 390672 434896 390674
rect 429429 390616 429434 390672
rect 429490 390616 434896 390672
rect 429429 390614 434896 390616
rect 429429 390611 429495 390614
rect 434416 390584 434896 390614
rect 128638 384826 128698 385408
rect 131349 384826 131415 384829
rect 128638 384824 131415 384826
rect 128638 384768 131354 384824
rect 131410 384768 131415 384824
rect 128638 384766 131415 384768
rect 222662 384826 222722 385408
rect 225281 384826 225347 384829
rect 222662 384824 225347 384826
rect 222662 384768 225286 384824
rect 225342 384768 225347 384824
rect 222662 384766 225347 384768
rect 316686 384826 316746 385408
rect 319029 384826 319095 384829
rect 316686 384824 319095 384826
rect 316686 384768 319034 384824
rect 319090 384768 319095 384824
rect 316686 384766 319095 384768
rect 131349 384763 131415 384766
rect 225281 384763 225347 384766
rect 319029 384763 319095 384766
rect 128638 382106 128698 382688
rect 131441 382106 131507 382109
rect 128638 382104 131507 382106
rect 128638 382048 131446 382104
rect 131502 382048 131507 382104
rect 128638 382046 131507 382048
rect 222662 382106 222722 382688
rect 225189 382106 225255 382109
rect 222662 382104 225255 382106
rect 222662 382048 225194 382104
rect 225250 382048 225255 382104
rect 222662 382046 225255 382048
rect 316686 382106 316746 382688
rect 319121 382106 319187 382109
rect 316686 382104 319187 382106
rect 316686 382048 319126 382104
rect 319182 382048 319187 382104
rect 316686 382046 319187 382048
rect 131441 382043 131507 382046
rect 225189 382043 225255 382046
rect 319121 382043 319187 382046
rect 9896 380610 10376 380640
rect 13681 380610 13747 380613
rect 9896 380608 13747 380610
rect 9896 380552 13686 380608
rect 13742 380552 13747 380608
rect 9896 380550 13747 380552
rect 9896 380520 10376 380550
rect 13681 380547 13747 380550
rect 131533 380202 131599 380205
rect 225373 380202 225439 380205
rect 319213 380202 319279 380205
rect 128668 380200 131599 380202
rect 128668 380144 131538 380200
rect 131594 380144 131599 380200
rect 128668 380142 131599 380144
rect 222692 380200 225439 380202
rect 222692 380144 225378 380200
rect 225434 380144 225439 380200
rect 222692 380142 225439 380144
rect 316716 380200 319279 380202
rect 316716 380144 319218 380200
rect 319274 380144 319279 380200
rect 316716 380142 319279 380144
rect 131533 380139 131599 380142
rect 225373 380139 225439 380142
rect 319213 380139 319279 380142
rect 429429 378570 429495 378573
rect 434416 378570 434896 378600
rect 429429 378568 434896 378570
rect 429429 378512 429434 378568
rect 429490 378512 434896 378568
rect 429429 378510 434896 378512
rect 429429 378507 429495 378510
rect 434416 378480 434896 378510
rect 131625 377482 131691 377485
rect 225465 377482 225531 377485
rect 319305 377482 319371 377485
rect 128668 377480 131691 377482
rect 128668 377424 131630 377480
rect 131686 377424 131691 377480
rect 128668 377422 131691 377424
rect 222692 377480 225531 377482
rect 222692 377424 225470 377480
rect 225526 377424 225531 377480
rect 222692 377422 225531 377424
rect 316716 377480 319371 377482
rect 316716 377424 319310 377480
rect 319366 377424 319371 377480
rect 316716 377422 319371 377424
rect 131625 377419 131691 377422
rect 225465 377419 225531 377422
rect 319305 377419 319371 377422
rect 131717 374762 131783 374765
rect 225557 374762 225623 374765
rect 319397 374762 319463 374765
rect 128668 374760 131783 374762
rect 128668 374704 131722 374760
rect 131778 374704 131783 374760
rect 128668 374702 131783 374704
rect 222692 374760 225623 374762
rect 222692 374704 225562 374760
rect 225618 374704 225623 374760
rect 222692 374702 225623 374704
rect 316716 374760 319463 374762
rect 316716 374704 319402 374760
rect 319458 374704 319463 374760
rect 316716 374702 319463 374704
rect 131717 374699 131783 374702
rect 225557 374699 225623 374702
rect 319397 374699 319463 374702
rect 131809 372178 131875 372181
rect 225833 372178 225899 372181
rect 128668 372176 131875 372178
rect 128668 372120 131814 372176
rect 131870 372120 131875 372176
rect 128668 372118 131875 372120
rect 222692 372176 225899 372178
rect 222692 372120 225838 372176
rect 225894 372120 225899 372176
rect 222692 372118 225899 372120
rect 131809 372115 131875 372118
rect 225833 372115 225899 372118
rect 316686 371906 316746 372080
rect 320133 371906 320199 371909
rect 316686 371904 320199 371906
rect 316686 371848 320138 371904
rect 320194 371848 320199 371904
rect 316686 371846 320199 371848
rect 320133 371843 320199 371846
rect 9896 369866 10376 369896
rect 13589 369866 13655 369869
rect 9896 369864 13655 369866
rect 9896 369808 13594 369864
rect 13650 369808 13655 369864
rect 9896 369806 13655 369808
rect 9896 369776 10376 369806
rect 13589 369803 13655 369806
rect 429429 366466 429495 366469
rect 434416 366466 434896 366496
rect 429429 366464 434896 366466
rect 429429 366408 429434 366464
rect 429490 366408 434896 366464
rect 429429 366406 434896 366408
rect 429429 366403 429495 366406
rect 434416 366376 434896 366406
rect 190781 359394 190847 359397
rect 191190 359394 191196 359396
rect 190781 359392 191196 359394
rect 190781 359336 190786 359392
rect 190842 359336 191196 359392
rect 190781 359334 191196 359336
rect 190781 359331 190847 359334
rect 191190 359332 191196 359334
rect 191260 359332 191266 359396
rect 9896 359122 10376 359152
rect 13497 359122 13563 359125
rect 9896 359120 13563 359122
rect 9896 359064 13502 359120
rect 13558 359064 13563 359120
rect 9896 359062 13563 359064
rect 9896 359032 10376 359062
rect 13497 359059 13563 359062
rect 139629 357762 139695 357765
rect 233469 357762 233535 357765
rect 139629 357760 143050 357762
rect 139629 357704 139634 357760
rect 139690 357704 143050 357760
rect 139629 357702 143050 357704
rect 139629 357699 139695 357702
rect 80197 357626 80263 357629
rect 76382 357624 80263 357626
rect 76382 357568 80202 357624
rect 80258 357568 80263 357624
rect 76382 357566 80263 357568
rect 76382 357188 76442 357566
rect 80197 357563 80263 357566
rect 142990 357256 143050 357702
rect 233469 357760 237074 357762
rect 233469 357704 233474 357760
rect 233530 357704 237074 357760
rect 233469 357702 237074 357704
rect 233469 357699 233535 357702
rect 237014 357256 237074 357702
rect 328413 357490 328479 357493
rect 328413 357488 331098 357490
rect 328413 357432 328418 357488
rect 328474 357432 331098 357488
rect 328413 357430 331098 357432
rect 328413 357427 328479 357430
rect 331038 357256 331098 357430
rect 174037 357218 174103 357221
rect 266589 357218 266655 357221
rect 170804 357216 174103 357218
rect 170804 357160 174042 357216
rect 174098 357160 174103 357216
rect 170804 357158 174103 357160
rect 264828 357216 266655 357218
rect 264828 357160 266594 357216
rect 266650 357160 266655 357216
rect 264828 357158 266655 357160
rect 174037 357155 174103 357158
rect 266589 357155 266655 357158
rect 139629 356538 139695 356541
rect 233469 356538 233535 356541
rect 284529 356540 284595 356541
rect 284478 356538 284484 356540
rect 139629 356536 143050 356538
rect 139629 356480 139634 356536
rect 139690 356480 143050 356536
rect 139629 356478 143050 356480
rect 139629 356475 139695 356478
rect 80197 356402 80263 356405
rect 76382 356400 80263 356402
rect 76382 356344 80202 356400
rect 80258 356344 80263 356400
rect 76382 356342 80263 356344
rect 76382 356100 76442 356342
rect 80197 356339 80263 356342
rect 142990 356168 143050 356478
rect 233469 356536 237074 356538
rect 233469 356480 233474 356536
rect 233530 356480 237074 356536
rect 233469 356478 237074 356480
rect 284438 356478 284484 356538
rect 284548 356536 284595 356540
rect 284590 356480 284595 356536
rect 233469 356475 233535 356478
rect 237014 356168 237074 356478
rect 284478 356476 284484 356478
rect 284548 356476 284595 356480
rect 284529 356475 284595 356476
rect 173485 356130 173551 356133
rect 266589 356130 266655 356133
rect 170804 356128 173551 356130
rect 170804 356072 173490 356128
rect 173546 356072 173551 356128
rect 170804 356070 173551 356072
rect 264828 356128 266655 356130
rect 264828 356072 266594 356128
rect 266650 356072 266655 356128
rect 264828 356070 266655 356072
rect 173485 356067 173551 356070
rect 266589 356067 266655 356070
rect 328321 356130 328387 356133
rect 328321 356128 331068 356130
rect 328321 356072 328326 356128
rect 328382 356072 331068 356128
rect 328321 356070 331068 356072
rect 328321 356067 328387 356070
rect 96849 355316 96915 355317
rect 96798 355252 96804 355316
rect 96868 355314 96915 355316
rect 96868 355312 96960 355314
rect 96910 355256 96960 355312
rect 96868 355254 96960 355256
rect 96868 355252 96915 355254
rect 96849 355251 96915 355252
rect 139629 355178 139695 355181
rect 174037 355178 174103 355181
rect 139629 355176 143020 355178
rect 76198 355042 76258 355148
rect 139629 355120 139634 355176
rect 139690 355120 143020 355176
rect 139629 355118 143020 355120
rect 170804 355176 174103 355178
rect 170804 355120 174042 355176
rect 174098 355120 174103 355176
rect 170804 355118 174103 355120
rect 139629 355115 139695 355118
rect 174037 355115 174103 355118
rect 233469 355178 233535 355181
rect 266589 355178 266655 355181
rect 233469 355176 237044 355178
rect 233469 355120 233474 355176
rect 233530 355120 237044 355176
rect 233469 355118 237044 355120
rect 264828 355176 266655 355178
rect 264828 355120 266594 355176
rect 266650 355120 266655 355176
rect 264828 355118 266655 355120
rect 233469 355115 233535 355118
rect 266589 355115 266655 355118
rect 328413 355178 328479 355181
rect 328413 355176 331068 355178
rect 328413 355120 328418 355176
rect 328474 355120 331068 355176
rect 328413 355118 331068 355120
rect 328413 355115 328479 355118
rect 80197 355042 80263 355045
rect 76198 355040 80263 355042
rect 76198 354984 80202 355040
rect 80258 354984 80263 355040
rect 76198 354982 80263 354984
rect 80197 354979 80263 354982
rect 79277 354634 79343 354637
rect 76382 354632 79343 354634
rect 76382 354576 79282 354632
rect 79338 354576 79343 354632
rect 76382 354574 79343 354576
rect 76382 354060 76442 354574
rect 79277 354571 79343 354574
rect 139721 354634 139787 354637
rect 233561 354634 233627 354637
rect 328505 354634 328571 354637
rect 139721 354632 143050 354634
rect 139721 354576 139726 354632
rect 139782 354576 143050 354632
rect 139721 354574 143050 354576
rect 139721 354571 139787 354574
rect 142990 354128 143050 354574
rect 233561 354632 237074 354634
rect 233561 354576 233566 354632
rect 233622 354576 237074 354632
rect 233561 354574 237074 354576
rect 233561 354571 233627 354574
rect 237014 354128 237074 354574
rect 328505 354632 331098 354634
rect 328505 354576 328510 354632
rect 328566 354576 331098 354632
rect 328505 354574 331098 354576
rect 328505 354571 328571 354574
rect 331038 354128 331098 354574
rect 429429 354362 429495 354365
rect 434416 354362 434896 354392
rect 429429 354360 434896 354362
rect 429429 354304 429434 354360
rect 429490 354304 434896 354360
rect 429429 354302 434896 354304
rect 429429 354299 429495 354302
rect 434416 354272 434896 354302
rect 173761 354090 173827 354093
rect 266681 354090 266747 354093
rect 170804 354088 173827 354090
rect 170804 354032 173766 354088
rect 173822 354032 173827 354088
rect 170804 354030 173827 354032
rect 264828 354088 266747 354090
rect 264828 354032 266686 354088
rect 266742 354032 266747 354088
rect 264828 354030 266747 354032
rect 173761 354027 173827 354030
rect 266681 354027 266747 354030
rect 139629 353546 139695 353549
rect 233469 353546 233535 353549
rect 139629 353544 143050 353546
rect 139629 353488 139634 353544
rect 139690 353488 143050 353544
rect 139629 353486 143050 353488
rect 139629 353483 139695 353486
rect 80197 353410 80263 353413
rect 76382 353408 80263 353410
rect 76382 353352 80202 353408
rect 80258 353352 80263 353408
rect 76382 353350 80263 353352
rect 76382 352972 76442 353350
rect 80197 353347 80263 353350
rect 142990 353040 143050 353486
rect 233469 353544 237074 353546
rect 233469 353488 233474 353544
rect 233530 353488 237074 353544
rect 233469 353486 237074 353488
rect 233469 353483 233535 353486
rect 237014 353040 237074 353486
rect 328045 353410 328111 353413
rect 328045 353408 331098 353410
rect 328045 353352 328050 353408
rect 328106 353352 331098 353408
rect 328045 353350 331098 353352
rect 328045 353347 328111 353350
rect 331038 353040 331098 353350
rect 174037 353002 174103 353005
rect 266589 353002 266655 353005
rect 170804 353000 174103 353002
rect 170804 352944 174042 353000
rect 174098 352944 174103 353000
rect 170804 352942 174103 352944
rect 264828 353000 266655 353002
rect 264828 352944 266594 353000
rect 266650 352944 266655 353000
rect 264828 352942 266655 352944
rect 174037 352939 174103 352942
rect 266589 352939 266655 352942
rect 139629 352322 139695 352325
rect 233469 352322 233535 352325
rect 328505 352322 328571 352325
rect 139629 352320 143050 352322
rect 139629 352264 139634 352320
rect 139690 352264 143050 352320
rect 139629 352262 143050 352264
rect 139629 352259 139695 352262
rect 80197 352186 80263 352189
rect 76382 352184 80263 352186
rect 76382 352128 80202 352184
rect 80258 352128 80263 352184
rect 76382 352126 80263 352128
rect 76382 352020 76442 352126
rect 80197 352123 80263 352126
rect 142990 352088 143050 352262
rect 233469 352320 237074 352322
rect 233469 352264 233474 352320
rect 233530 352264 237074 352320
rect 233469 352262 237074 352264
rect 233469 352259 233535 352262
rect 237014 352088 237074 352262
rect 328505 352320 331098 352322
rect 328505 352264 328510 352320
rect 328566 352264 331098 352320
rect 328505 352262 331098 352264
rect 328505 352259 328571 352262
rect 331038 352088 331098 352262
rect 174037 352050 174103 352053
rect 266589 352050 266655 352053
rect 170804 352048 174103 352050
rect 170804 351992 174042 352048
rect 174098 351992 174103 352048
rect 170804 351990 174103 351992
rect 264828 352048 266655 352050
rect 264828 351992 266594 352048
rect 266650 351992 266655 352048
rect 264828 351990 266655 351992
rect 174037 351987 174103 351990
rect 266589 351987 266655 351990
rect 191241 351916 191307 351917
rect 191190 351914 191196 351916
rect 191150 351854 191196 351914
rect 191260 351912 191307 351916
rect 191302 351856 191307 351912
rect 191190 351852 191196 351854
rect 191260 351852 191307 351856
rect 191241 351851 191307 351852
rect 96757 351644 96823 351645
rect 284529 351644 284595 351645
rect 96757 351640 96804 351644
rect 96868 351642 96874 351644
rect 284478 351642 284484 351644
rect 96757 351584 96762 351640
rect 96757 351580 96804 351584
rect 96868 351582 96914 351642
rect 284438 351582 284484 351642
rect 284548 351640 284595 351644
rect 284590 351584 284595 351640
rect 96868 351580 96874 351582
rect 284478 351580 284484 351582
rect 284548 351580 284595 351584
rect 96757 351579 96823 351580
rect 284529 351579 284595 351580
rect 87097 351370 87163 351373
rect 131809 351370 131875 351373
rect 87097 351368 90028 351370
rect 87097 351312 87102 351368
rect 87158 351312 90028 351368
rect 87097 351310 90028 351312
rect 129772 351368 131875 351370
rect 129772 351312 131814 351368
rect 131870 351312 131875 351368
rect 129772 351310 131875 351312
rect 87097 351307 87163 351310
rect 131809 351307 131875 351310
rect 182317 351370 182383 351373
rect 226293 351370 226359 351373
rect 182317 351368 184052 351370
rect 182317 351312 182322 351368
rect 182378 351312 184052 351368
rect 182317 351310 184052 351312
rect 223796 351368 226359 351370
rect 223796 351312 226298 351368
rect 226354 351312 226359 351368
rect 223796 351310 226359 351312
rect 182317 351307 182383 351310
rect 226293 351307 226359 351310
rect 274869 351370 274935 351373
rect 320593 351370 320659 351373
rect 274869 351368 278076 351370
rect 274869 351312 274874 351368
rect 274930 351312 278076 351368
rect 274869 351310 278076 351312
rect 317820 351368 320659 351370
rect 317820 351312 320598 351368
rect 320654 351312 320659 351368
rect 317820 351310 320659 351312
rect 274869 351307 274935 351310
rect 320593 351307 320659 351310
rect 139721 350962 139787 350965
rect 173669 350962 173735 350965
rect 139721 350960 143020 350962
rect 76198 350690 76258 350932
rect 139721 350904 139726 350960
rect 139782 350904 143020 350960
rect 139721 350902 143020 350904
rect 170804 350960 173735 350962
rect 170804 350904 173674 350960
rect 173730 350904 173735 350960
rect 170804 350902 173735 350904
rect 139721 350899 139787 350902
rect 173669 350899 173735 350902
rect 233469 350962 233535 350965
rect 266589 350962 266655 350965
rect 233469 350960 237044 350962
rect 233469 350904 233474 350960
rect 233530 350904 237044 350960
rect 233469 350902 237044 350904
rect 264828 350960 266655 350962
rect 264828 350904 266594 350960
rect 266650 350904 266655 350960
rect 264828 350902 266655 350904
rect 233469 350899 233535 350902
rect 266589 350899 266655 350902
rect 327493 350962 327559 350965
rect 327493 350960 331068 350962
rect 327493 350904 327498 350960
rect 327554 350904 331068 350960
rect 327493 350902 331068 350904
rect 327493 350899 327559 350902
rect 80197 350690 80263 350693
rect 76198 350688 80263 350690
rect 76198 350632 80202 350688
rect 80258 350632 80263 350688
rect 76198 350630 80263 350632
rect 80197 350627 80263 350630
rect 139629 350554 139695 350557
rect 233561 350554 233627 350557
rect 139629 350552 143050 350554
rect 139629 350496 139634 350552
rect 139690 350496 143050 350552
rect 139629 350494 143050 350496
rect 139629 350491 139695 350494
rect 79829 350418 79895 350421
rect 76382 350416 79895 350418
rect 76382 350360 79834 350416
rect 79890 350360 79895 350416
rect 76382 350358 79895 350360
rect 76382 349844 76442 350358
rect 79829 350355 79895 350358
rect 87005 350418 87071 350421
rect 131809 350418 131875 350421
rect 87005 350416 90028 350418
rect 87005 350360 87010 350416
rect 87066 350360 90028 350416
rect 87005 350358 90028 350360
rect 129772 350416 131875 350418
rect 129772 350360 131814 350416
rect 131870 350360 131875 350416
rect 129772 350358 131875 350360
rect 87005 350355 87071 350358
rect 131809 350355 131875 350358
rect 142990 349912 143050 350494
rect 233561 350552 237074 350554
rect 233561 350496 233566 350552
rect 233622 350496 237074 350552
rect 233561 350494 237074 350496
rect 233561 350491 233627 350494
rect 226569 350418 226635 350421
rect 223796 350416 226635 350418
rect 180753 350010 180819 350013
rect 184022 350010 184082 350388
rect 223796 350360 226574 350416
rect 226630 350360 226635 350416
rect 223796 350358 226635 350360
rect 226569 350355 226635 350358
rect 180753 350008 184082 350010
rect 180753 349952 180758 350008
rect 180814 349952 184082 350008
rect 180753 349950 184082 349952
rect 180753 349947 180819 349950
rect 237014 349912 237074 350494
rect 274869 350418 274935 350421
rect 321605 350418 321671 350421
rect 274869 350416 278076 350418
rect 274869 350360 274874 350416
rect 274930 350360 278076 350416
rect 274869 350358 278076 350360
rect 317820 350416 321671 350418
rect 317820 350360 321610 350416
rect 321666 350360 321671 350416
rect 317820 350358 321671 350360
rect 274869 350355 274935 350358
rect 321605 350355 321671 350358
rect 327861 350418 327927 350421
rect 327861 350416 331098 350418
rect 327861 350360 327866 350416
rect 327922 350360 331098 350416
rect 327861 350358 331098 350360
rect 327861 350355 327927 350358
rect 331038 349912 331098 350358
rect 173853 349874 173919 349877
rect 266681 349874 266747 349877
rect 170804 349872 173919 349874
rect 170804 349816 173858 349872
rect 173914 349816 173919 349872
rect 170804 349814 173919 349816
rect 264828 349872 266747 349874
rect 264828 349816 266686 349872
rect 266742 349816 266747 349872
rect 264828 349814 266747 349816
rect 173853 349811 173919 349814
rect 266681 349811 266747 349814
rect 86913 349602 86979 349605
rect 131901 349602 131967 349605
rect 86913 349600 90028 349602
rect 86913 349544 86918 349600
rect 86974 349544 90028 349600
rect 86913 349542 90028 349544
rect 129772 349600 131967 349602
rect 129772 349544 131906 349600
rect 131962 349544 131967 349600
rect 129772 349542 131967 349544
rect 86913 349539 86979 349542
rect 131901 349539 131967 349542
rect 139445 349602 139511 349605
rect 226477 349602 226543 349605
rect 139445 349600 143050 349602
rect 139445 349544 139450 349600
rect 139506 349544 143050 349600
rect 223796 349600 226543 349602
rect 139445 349542 143050 349544
rect 139445 349539 139511 349542
rect 78909 349058 78975 349061
rect 76382 349056 78975 349058
rect 76382 349000 78914 349056
rect 78970 349000 78975 349056
rect 76382 348998 78975 349000
rect 76382 348892 76442 348998
rect 78909 348995 78975 348998
rect 142990 348960 143050 349542
rect 180937 349058 181003 349061
rect 184022 349058 184082 349572
rect 223796 349544 226482 349600
rect 226538 349544 226543 349600
rect 223796 349542 226543 349544
rect 226477 349539 226543 349542
rect 233469 349602 233535 349605
rect 274869 349602 274935 349605
rect 321697 349602 321763 349605
rect 233469 349600 237074 349602
rect 233469 349544 233474 349600
rect 233530 349544 237074 349600
rect 233469 349542 237074 349544
rect 233469 349539 233535 349542
rect 180937 349056 184082 349058
rect 180937 349000 180942 349056
rect 180998 349000 184082 349056
rect 180937 348998 184082 349000
rect 180937 348995 181003 348998
rect 237014 348960 237074 349542
rect 274869 349600 278076 349602
rect 274869 349544 274874 349600
rect 274930 349544 278076 349600
rect 274869 349542 278076 349544
rect 317820 349600 321763 349602
rect 317820 349544 321702 349600
rect 321758 349544 321763 349600
rect 317820 349542 321763 349544
rect 274869 349539 274935 349542
rect 321697 349539 321763 349542
rect 328137 349602 328203 349605
rect 328137 349600 331098 349602
rect 328137 349544 328142 349600
rect 328198 349544 331098 349600
rect 328137 349542 331098 349544
rect 328137 349539 328203 349542
rect 331038 348960 331098 349542
rect 172841 348922 172907 348925
rect 266589 348922 266655 348925
rect 170804 348920 172907 348922
rect 170804 348864 172846 348920
rect 172902 348864 172907 348920
rect 170804 348862 172907 348864
rect 264828 348920 266655 348922
rect 264828 348864 266594 348920
rect 266650 348864 266655 348920
rect 264828 348862 266655 348864
rect 172841 348859 172907 348862
rect 266589 348859 266655 348862
rect 87097 348650 87163 348653
rect 131809 348650 131875 348653
rect 226385 348650 226451 348653
rect 87097 348648 90028 348650
rect 87097 348592 87102 348648
rect 87158 348592 90028 348648
rect 87097 348590 90028 348592
rect 129772 348648 131875 348650
rect 129772 348592 131814 348648
rect 131870 348592 131875 348648
rect 223796 348648 226451 348650
rect 129772 348590 131875 348592
rect 87097 348587 87163 348590
rect 131809 348587 131875 348590
rect 180845 348378 180911 348381
rect 184022 348378 184082 348620
rect 223796 348592 226390 348648
rect 226446 348592 226451 348648
rect 223796 348590 226451 348592
rect 226385 348587 226451 348590
rect 274961 348650 275027 348653
rect 321605 348650 321671 348653
rect 274961 348648 278076 348650
rect 274961 348592 274966 348648
rect 275022 348592 278076 348648
rect 274961 348590 278076 348592
rect 317820 348648 321671 348650
rect 317820 348592 321610 348648
rect 321666 348592 321671 348648
rect 317820 348590 321671 348592
rect 274961 348587 275027 348590
rect 321605 348587 321671 348590
rect 180845 348376 184082 348378
rect 180845 348320 180850 348376
rect 180906 348320 184082 348376
rect 180845 348318 184082 348320
rect 180845 348315 180911 348318
rect 9896 348242 10376 348272
rect 13405 348242 13471 348245
rect 9896 348240 13471 348242
rect 9896 348184 13410 348240
rect 13466 348184 13471 348240
rect 9896 348182 13471 348184
rect 9896 348152 10376 348182
rect 13405 348179 13471 348182
rect 139537 348242 139603 348245
rect 233469 348242 233535 348245
rect 328321 348242 328387 348245
rect 139537 348240 143050 348242
rect 139537 348184 139542 348240
rect 139598 348184 143050 348240
rect 139537 348182 143050 348184
rect 139537 348179 139603 348182
rect 142990 347872 143050 348182
rect 233469 348240 237074 348242
rect 233469 348184 233474 348240
rect 233530 348184 237074 348240
rect 233469 348182 237074 348184
rect 233469 348179 233535 348182
rect 237014 347872 237074 348182
rect 328321 348240 331098 348242
rect 328321 348184 328326 348240
rect 328382 348184 331098 348240
rect 328321 348182 331098 348184
rect 328321 348179 328387 348182
rect 331038 347872 331098 348182
rect 132177 347834 132243 347837
rect 174037 347834 174103 347837
rect 226385 347834 226451 347837
rect 266589 347834 266655 347837
rect 129772 347832 132243 347834
rect 76198 347562 76258 347804
rect 78909 347562 78975 347565
rect 76198 347560 78975 347562
rect 76198 347504 78914 347560
rect 78970 347504 78975 347560
rect 76198 347502 78975 347504
rect 78909 347499 78975 347502
rect 87005 347290 87071 347293
rect 89998 347290 90058 347804
rect 129772 347776 132182 347832
rect 132238 347776 132243 347832
rect 129772 347774 132243 347776
rect 170804 347832 174103 347834
rect 170804 347776 174042 347832
rect 174098 347776 174103 347832
rect 223796 347832 226451 347834
rect 170804 347774 174103 347776
rect 132177 347771 132243 347774
rect 174037 347771 174103 347774
rect 87005 347288 90058 347290
rect 87005 347232 87010 347288
rect 87066 347232 90058 347288
rect 87005 347230 90058 347232
rect 180753 347290 180819 347293
rect 184022 347290 184082 347804
rect 223796 347776 226390 347832
rect 226446 347776 226451 347832
rect 223796 347774 226451 347776
rect 264828 347832 266655 347834
rect 264828 347776 266594 347832
rect 266650 347776 266655 347832
rect 264828 347774 266655 347776
rect 226385 347771 226451 347774
rect 266589 347771 266655 347774
rect 275053 347834 275119 347837
rect 321053 347834 321119 347837
rect 275053 347832 278076 347834
rect 275053 347776 275058 347832
rect 275114 347776 278076 347832
rect 275053 347774 278076 347776
rect 317820 347832 321119 347834
rect 317820 347776 321058 347832
rect 321114 347776 321119 347832
rect 317820 347774 321119 347776
rect 275053 347771 275119 347774
rect 321053 347771 321119 347774
rect 180753 347288 184082 347290
rect 180753 347232 180758 347288
rect 180814 347232 184082 347288
rect 180753 347230 184082 347232
rect 87005 347227 87071 347230
rect 180753 347227 180819 347230
rect 87925 346882 87991 346885
rect 131901 346882 131967 346885
rect 87925 346880 90028 346882
rect 76198 346474 76258 346852
rect 87925 346824 87930 346880
rect 87986 346824 90028 346880
rect 87925 346822 90028 346824
rect 129772 346880 131967 346882
rect 129772 346824 131906 346880
rect 131962 346824 131967 346880
rect 129772 346822 131967 346824
rect 87925 346819 87991 346822
rect 131901 346819 131967 346822
rect 139629 346882 139695 346885
rect 174037 346882 174103 346885
rect 139629 346880 143020 346882
rect 139629 346824 139634 346880
rect 139690 346824 143020 346880
rect 139629 346822 143020 346824
rect 170804 346880 174103 346882
rect 170804 346824 174042 346880
rect 174098 346824 174103 346880
rect 170804 346822 174103 346824
rect 139629 346819 139695 346822
rect 174037 346819 174103 346822
rect 181029 346882 181095 346885
rect 226477 346882 226543 346885
rect 181029 346880 184052 346882
rect 181029 346824 181034 346880
rect 181090 346824 184052 346880
rect 181029 346822 184052 346824
rect 223796 346880 226543 346882
rect 223796 346824 226482 346880
rect 226538 346824 226543 346880
rect 223796 346822 226543 346824
rect 181029 346819 181095 346822
rect 226477 346819 226543 346822
rect 233469 346882 233535 346885
rect 266589 346882 266655 346885
rect 233469 346880 237044 346882
rect 233469 346824 233474 346880
rect 233530 346824 237044 346880
rect 233469 346822 237044 346824
rect 264828 346880 266655 346882
rect 264828 346824 266594 346880
rect 266650 346824 266655 346880
rect 264828 346822 266655 346824
rect 233469 346819 233535 346822
rect 266589 346819 266655 346822
rect 275145 346882 275211 346885
rect 320409 346882 320475 346885
rect 275145 346880 278076 346882
rect 275145 346824 275150 346880
rect 275206 346824 278076 346880
rect 275145 346822 278076 346824
rect 317820 346880 320475 346882
rect 317820 346824 320414 346880
rect 320470 346824 320475 346880
rect 317820 346822 320475 346824
rect 275145 346819 275211 346822
rect 320409 346819 320475 346822
rect 327217 346882 327283 346885
rect 327217 346880 331068 346882
rect 327217 346824 327222 346880
rect 327278 346824 331068 346880
rect 327217 346822 331068 346824
rect 327217 346819 327283 346822
rect 79001 346474 79067 346477
rect 76198 346472 79067 346474
rect 76198 346416 79006 346472
rect 79062 346416 79067 346472
rect 76198 346414 79067 346416
rect 79001 346411 79067 346414
rect 233561 346474 233627 346477
rect 327125 346474 327191 346477
rect 233561 346472 237074 346474
rect 233561 346416 233566 346472
rect 233622 346416 237074 346472
rect 233561 346414 237074 346416
rect 233561 346411 233627 346414
rect 139813 346338 139879 346341
rect 139813 346336 143050 346338
rect 139813 346280 139818 346336
rect 139874 346280 143050 346336
rect 139813 346278 143050 346280
rect 139813 346275 139879 346278
rect 78909 346066 78975 346069
rect 76382 346064 78975 346066
rect 76382 346008 78914 346064
rect 78970 346008 78975 346064
rect 76382 346006 78975 346008
rect 76382 345764 76442 346006
rect 78909 346003 78975 346006
rect 88109 346066 88175 346069
rect 131809 346066 131875 346069
rect 88109 346064 90028 346066
rect 88109 346008 88114 346064
rect 88170 346008 90028 346064
rect 88109 346006 90028 346008
rect 129772 346064 131875 346066
rect 129772 346008 131814 346064
rect 131870 346008 131875 346064
rect 129772 346006 131875 346008
rect 88109 346003 88175 346006
rect 131809 346003 131875 346006
rect 142990 345832 143050 346278
rect 182317 346066 182383 346069
rect 226385 346066 226451 346069
rect 182317 346064 184052 346066
rect 182317 346008 182322 346064
rect 182378 346008 184052 346064
rect 182317 346006 184052 346008
rect 223796 346064 226451 346066
rect 223796 346008 226390 346064
rect 226446 346008 226451 346064
rect 223796 346006 226451 346008
rect 182317 346003 182383 346006
rect 226385 346003 226451 346006
rect 237014 345832 237074 346414
rect 327125 346472 331098 346474
rect 327125 346416 327130 346472
rect 327186 346416 331098 346472
rect 327125 346414 331098 346416
rect 327125 346411 327191 346414
rect 275237 346066 275303 346069
rect 320501 346066 320567 346069
rect 275237 346064 278076 346066
rect 275237 346008 275242 346064
rect 275298 346008 278076 346064
rect 275237 346006 278076 346008
rect 317820 346064 320567 346066
rect 317820 346008 320506 346064
rect 320562 346008 320567 346064
rect 317820 346006 320567 346008
rect 275237 346003 275303 346006
rect 320501 346003 320567 346006
rect 331038 345832 331098 346414
rect 173117 345794 173183 345797
rect 170804 345792 173183 345794
rect 170804 345736 173122 345792
rect 173178 345736 173183 345792
rect 170804 345734 173183 345736
rect 173117 345731 173183 345734
rect 180845 345794 180911 345797
rect 181029 345794 181095 345797
rect 266681 345794 266747 345797
rect 180845 345792 181095 345794
rect 180845 345736 180850 345792
rect 180906 345736 181034 345792
rect 181090 345736 181095 345792
rect 180845 345734 181095 345736
rect 264828 345792 266747 345794
rect 264828 345736 266686 345792
rect 266742 345736 266747 345792
rect 264828 345734 266747 345736
rect 180845 345731 180911 345734
rect 181029 345731 181095 345734
rect 266681 345731 266747 345734
rect 139721 345386 139787 345389
rect 139721 345384 143050 345386
rect 139721 345328 139726 345384
rect 139782 345328 143050 345384
rect 139721 345326 143050 345328
rect 139721 345323 139787 345326
rect 87465 345114 87531 345117
rect 132361 345114 132427 345117
rect 87465 345112 90028 345114
rect 87465 345056 87470 345112
rect 87526 345056 90028 345112
rect 87465 345054 90028 345056
rect 129772 345112 132427 345114
rect 129772 345056 132366 345112
rect 132422 345056 132427 345112
rect 129772 345054 132427 345056
rect 87465 345051 87531 345054
rect 132361 345051 132427 345054
rect 142990 344744 143050 345326
rect 233469 345250 233535 345253
rect 233469 345248 237074 345250
rect 233469 345192 233474 345248
rect 233530 345192 237074 345248
rect 233469 345190 237074 345192
rect 233469 345187 233535 345190
rect 226017 345114 226083 345117
rect 223796 345112 226083 345114
rect 173301 344706 173367 344709
rect 170804 344704 173367 344706
rect 76198 344570 76258 344676
rect 170804 344648 173306 344704
rect 173362 344648 173367 344704
rect 170804 344646 173367 344648
rect 173301 344643 173367 344646
rect 180937 344706 181003 344709
rect 184022 344706 184082 345084
rect 223796 345056 226022 345112
rect 226078 345056 226083 345112
rect 223796 345054 226083 345056
rect 226017 345051 226083 345054
rect 237014 344744 237074 345190
rect 274869 345114 274935 345117
rect 321053 345114 321119 345117
rect 274869 345112 278076 345114
rect 274869 345056 274874 345112
rect 274930 345056 278076 345112
rect 274869 345054 278076 345056
rect 317820 345112 321119 345114
rect 317820 345056 321058 345112
rect 321114 345056 321119 345112
rect 317820 345054 321119 345056
rect 274869 345051 274935 345054
rect 321053 345051 321119 345054
rect 328045 345114 328111 345117
rect 328045 345112 331098 345114
rect 328045 345056 328050 345112
rect 328106 345056 331098 345112
rect 328045 345054 331098 345056
rect 328045 345051 328111 345054
rect 331038 344744 331098 345054
rect 266589 344706 266655 344709
rect 180937 344704 184082 344706
rect 180937 344648 180942 344704
rect 180998 344648 184082 344704
rect 180937 344646 184082 344648
rect 264828 344704 266655 344706
rect 264828 344648 266594 344704
rect 266650 344648 266655 344704
rect 264828 344646 266655 344648
rect 180937 344643 181003 344646
rect 266589 344643 266655 344646
rect 78909 344570 78975 344573
rect 76198 344568 78975 344570
rect 76198 344512 78914 344568
rect 78970 344512 78975 344568
rect 76198 344510 78975 344512
rect 78909 344507 78975 344510
rect 88477 344298 88543 344301
rect 131809 344298 131875 344301
rect 88477 344296 90028 344298
rect 88477 344240 88482 344296
rect 88538 344240 90028 344296
rect 88477 344238 90028 344240
rect 129772 344296 131875 344298
rect 129772 344240 131814 344296
rect 131870 344240 131875 344296
rect 129772 344238 131875 344240
rect 88477 344235 88543 344238
rect 131809 344235 131875 344238
rect 182317 344298 182383 344301
rect 226385 344298 226451 344301
rect 182317 344296 184052 344298
rect 182317 344240 182322 344296
rect 182378 344240 184052 344296
rect 182317 344238 184052 344240
rect 223796 344296 226451 344298
rect 223796 344240 226390 344296
rect 226446 344240 226451 344296
rect 223796 344238 226451 344240
rect 182317 344235 182383 344238
rect 226385 344235 226451 344238
rect 275053 344298 275119 344301
rect 321605 344298 321671 344301
rect 275053 344296 278076 344298
rect 275053 344240 275058 344296
rect 275114 344240 278076 344296
rect 275053 344238 278076 344240
rect 317820 344296 321671 344298
rect 317820 344240 321610 344296
rect 321666 344240 321671 344296
rect 317820 344238 321671 344240
rect 275053 344235 275119 344238
rect 321605 344235 321671 344238
rect 139629 344162 139695 344165
rect 139629 344160 143050 344162
rect 139629 344104 139634 344160
rect 139690 344104 143050 344160
rect 139629 344102 143050 344104
rect 139629 344099 139695 344102
rect 142990 343792 143050 344102
rect 233469 344026 233535 344029
rect 328505 344026 328571 344029
rect 233469 344024 237074 344026
rect 233469 343968 233474 344024
rect 233530 343968 237074 344024
rect 233469 343966 237074 343968
rect 233469 343963 233535 343966
rect 237014 343792 237074 343966
rect 328505 344024 331098 344026
rect 328505 343968 328510 344024
rect 328566 343968 331098 344024
rect 328505 343966 331098 343968
rect 328505 343963 328571 343966
rect 331038 343792 331098 343966
rect 173669 343754 173735 343757
rect 266589 343754 266655 343757
rect 170804 343752 173735 343754
rect 76198 343346 76258 343724
rect 170804 343696 173674 343752
rect 173730 343696 173735 343752
rect 170804 343694 173735 343696
rect 264828 343752 266655 343754
rect 264828 343696 266594 343752
rect 266650 343696 266655 343752
rect 264828 343694 266655 343696
rect 173669 343691 173735 343694
rect 266589 343691 266655 343694
rect 78909 343346 78975 343349
rect 76198 343344 78975 343346
rect 76198 343288 78914 343344
rect 78970 343288 78975 343344
rect 76198 343286 78975 343288
rect 78909 343283 78975 343286
rect 87373 343346 87439 343349
rect 131809 343346 131875 343349
rect 87373 343344 90028 343346
rect 87373 343288 87378 343344
rect 87434 343288 90028 343344
rect 87373 343286 90028 343288
rect 129772 343344 131875 343346
rect 129772 343288 131814 343344
rect 131870 343288 131875 343344
rect 129772 343286 131875 343288
rect 87373 343283 87439 343286
rect 131809 343283 131875 343286
rect 181397 343346 181463 343349
rect 226385 343346 226451 343349
rect 181397 343344 184052 343346
rect 181397 343288 181402 343344
rect 181458 343288 184052 343344
rect 181397 343286 184052 343288
rect 223796 343344 226451 343346
rect 223796 343288 226390 343344
rect 226446 343288 226451 343344
rect 223796 343286 226451 343288
rect 181397 343283 181463 343286
rect 226385 343283 226451 343286
rect 274961 343346 275027 343349
rect 321605 343346 321671 343349
rect 274961 343344 278076 343346
rect 274961 343288 274966 343344
rect 275022 343288 278076 343344
rect 274961 343286 278076 343288
rect 317820 343344 321671 343346
rect 317820 343288 321610 343344
rect 321666 343288 321671 343344
rect 317820 343286 321671 343288
rect 274961 343283 275027 343286
rect 321605 343283 321671 343286
rect 78909 342802 78975 342805
rect 76382 342800 78975 342802
rect 76382 342744 78914 342800
rect 78970 342744 78975 342800
rect 76382 342742 78975 342744
rect 76382 342636 76442 342742
rect 78909 342739 78975 342742
rect 139629 342666 139695 342669
rect 173025 342666 173091 342669
rect 139629 342664 143020 342666
rect 139629 342608 139634 342664
rect 139690 342608 143020 342664
rect 139629 342606 143020 342608
rect 170804 342664 173091 342666
rect 170804 342608 173030 342664
rect 173086 342608 173091 342664
rect 170804 342606 173091 342608
rect 139629 342603 139695 342606
rect 173025 342603 173091 342606
rect 234573 342666 234639 342669
rect 266589 342666 266655 342669
rect 234573 342664 237044 342666
rect 234573 342608 234578 342664
rect 234634 342608 237044 342664
rect 234573 342606 237044 342608
rect 264828 342664 266655 342666
rect 264828 342608 266594 342664
rect 266650 342608 266655 342664
rect 264828 342606 266655 342608
rect 234573 342603 234639 342606
rect 266589 342603 266655 342606
rect 327033 342666 327099 342669
rect 327033 342664 331068 342666
rect 327033 342608 327038 342664
rect 327094 342608 331068 342664
rect 327033 342606 331068 342608
rect 327033 342603 327099 342606
rect 87465 342394 87531 342397
rect 131901 342394 131967 342397
rect 87465 342392 90028 342394
rect 87465 342336 87470 342392
rect 87526 342336 90028 342392
rect 87465 342334 90028 342336
rect 129772 342392 131967 342394
rect 129772 342336 131906 342392
rect 131962 342336 131967 342392
rect 129772 342334 131967 342336
rect 87465 342331 87531 342334
rect 131901 342331 131967 342334
rect 182133 342394 182199 342397
rect 226477 342394 226543 342397
rect 182133 342392 184052 342394
rect 182133 342336 182138 342392
rect 182194 342336 184052 342392
rect 182133 342334 184052 342336
rect 223796 342392 226543 342394
rect 223796 342336 226482 342392
rect 226538 342336 226543 342392
rect 223796 342334 226543 342336
rect 182133 342331 182199 342334
rect 226477 342331 226543 342334
rect 275145 342394 275211 342397
rect 321053 342394 321119 342397
rect 275145 342392 278076 342394
rect 275145 342336 275150 342392
rect 275206 342336 278076 342392
rect 275145 342334 278076 342336
rect 317820 342392 321119 342394
rect 317820 342336 321058 342392
rect 321114 342336 321119 342392
rect 317820 342334 321119 342336
rect 275145 342331 275211 342334
rect 321053 342331 321119 342334
rect 139721 342258 139787 342261
rect 233469 342258 233535 342261
rect 429429 342258 429495 342261
rect 434416 342258 434896 342288
rect 139721 342256 143050 342258
rect 139721 342200 139726 342256
rect 139782 342200 143050 342256
rect 139721 342198 143050 342200
rect 139721 342195 139787 342198
rect 78909 341714 78975 341717
rect 76382 341712 78975 341714
rect 76382 341656 78914 341712
rect 78970 341656 78975 341712
rect 76382 341654 78975 341656
rect 76382 341548 76442 341654
rect 78909 341651 78975 341654
rect 142990 341616 143050 342198
rect 233469 342256 237074 342258
rect 233469 342200 233474 342256
rect 233530 342200 237074 342256
rect 233469 342198 237074 342200
rect 233469 342195 233535 342198
rect 237014 341616 237074 342198
rect 429429 342256 434896 342258
rect 429429 342200 429434 342256
rect 429490 342200 434896 342256
rect 429429 342198 434896 342200
rect 429429 342195 429495 342198
rect 434416 342168 434896 342198
rect 328045 342122 328111 342125
rect 328045 342120 331098 342122
rect 328045 342064 328050 342120
rect 328106 342064 331098 342120
rect 328045 342062 331098 342064
rect 328045 342059 328111 342062
rect 331038 341616 331098 342062
rect 87281 341578 87347 341581
rect 131809 341578 131875 341581
rect 172749 341578 172815 341581
rect 87281 341576 90028 341578
rect 87281 341520 87286 341576
rect 87342 341520 90028 341576
rect 87281 341518 90028 341520
rect 129772 341576 131875 341578
rect 129772 341520 131814 341576
rect 131870 341520 131875 341576
rect 129772 341518 131875 341520
rect 170804 341576 172815 341578
rect 170804 341520 172754 341576
rect 172810 341520 172815 341576
rect 170804 341518 172815 341520
rect 87281 341515 87347 341518
rect 131809 341515 131875 341518
rect 172749 341515 172815 341518
rect 181765 341578 181831 341581
rect 226385 341578 226451 341581
rect 266681 341578 266747 341581
rect 181765 341576 184052 341578
rect 181765 341520 181770 341576
rect 181826 341520 184052 341576
rect 181765 341518 184052 341520
rect 223796 341576 226451 341578
rect 223796 341520 226390 341576
rect 226446 341520 226451 341576
rect 223796 341518 226451 341520
rect 264828 341576 266747 341578
rect 264828 341520 266686 341576
rect 266742 341520 266747 341576
rect 264828 341518 266747 341520
rect 181765 341515 181831 341518
rect 226385 341515 226451 341518
rect 266681 341515 266747 341518
rect 274869 341578 274935 341581
rect 321605 341578 321671 341581
rect 274869 341576 278076 341578
rect 274869 341520 274874 341576
rect 274930 341520 278076 341576
rect 274869 341518 278076 341520
rect 317820 341576 321671 341578
rect 317820 341520 321610 341576
rect 321666 341520 321671 341576
rect 317820 341518 321671 341520
rect 274869 341515 274935 341518
rect 321605 341515 321671 341518
rect 139629 341306 139695 341309
rect 326849 341306 326915 341309
rect 139629 341304 143050 341306
rect 139629 341248 139634 341304
rect 139690 341248 143050 341304
rect 139629 341246 143050 341248
rect 139629 341243 139695 341246
rect 78909 341034 78975 341037
rect 76382 341032 78975 341034
rect 76382 340976 78914 341032
rect 78970 340976 78975 341032
rect 76382 340974 78975 340976
rect 76382 340596 76442 340974
rect 78909 340971 78975 340974
rect 142990 340664 143050 341246
rect 326849 341304 331098 341306
rect 326849 341248 326854 341304
rect 326910 341248 331098 341304
rect 326849 341246 331098 341248
rect 326849 341243 326915 341246
rect 233469 341170 233535 341173
rect 233469 341168 237074 341170
rect 233469 341112 233474 341168
rect 233530 341112 237074 341168
rect 233469 341110 237074 341112
rect 233469 341107 233535 341110
rect 237014 340664 237074 341110
rect 331038 340664 331098 341246
rect 87557 340626 87623 340629
rect 131809 340626 131875 340629
rect 172933 340626 172999 340629
rect 87557 340624 90028 340626
rect 87557 340568 87562 340624
rect 87618 340568 90028 340624
rect 87557 340566 90028 340568
rect 129772 340624 131875 340626
rect 129772 340568 131814 340624
rect 131870 340568 131875 340624
rect 129772 340566 131875 340568
rect 170804 340624 172999 340626
rect 170804 340568 172938 340624
rect 172994 340568 172999 340624
rect 170804 340566 172999 340568
rect 87557 340563 87623 340566
rect 131809 340563 131875 340566
rect 172933 340563 172999 340566
rect 181397 340626 181463 340629
rect 226385 340626 226451 340629
rect 266589 340626 266655 340629
rect 181397 340624 184052 340626
rect 181397 340568 181402 340624
rect 181458 340568 184052 340624
rect 181397 340566 184052 340568
rect 223796 340624 226451 340626
rect 223796 340568 226390 340624
rect 226446 340568 226451 340624
rect 223796 340566 226451 340568
rect 264828 340624 266655 340626
rect 264828 340568 266594 340624
rect 266650 340568 266655 340624
rect 264828 340566 266655 340568
rect 181397 340563 181463 340566
rect 226385 340563 226451 340566
rect 266589 340563 266655 340566
rect 275053 340626 275119 340629
rect 320593 340626 320659 340629
rect 275053 340624 278076 340626
rect 275053 340568 275058 340624
rect 275114 340568 278076 340624
rect 275053 340566 278076 340568
rect 317820 340624 320659 340626
rect 317820 340568 320598 340624
rect 320654 340568 320659 340624
rect 317820 340566 320659 340568
rect 275053 340563 275119 340566
rect 320593 340563 320659 340566
rect 139813 339946 139879 339949
rect 233653 339946 233719 339949
rect 327125 339946 327191 339949
rect 139813 339944 143050 339946
rect 139813 339888 139818 339944
rect 139874 339888 143050 339944
rect 139813 339886 143050 339888
rect 139813 339883 139879 339886
rect 78909 339810 78975 339813
rect 76382 339808 78975 339810
rect 76382 339752 78914 339808
rect 78970 339752 78975 339808
rect 76382 339750 78975 339752
rect 76382 339508 76442 339750
rect 78909 339747 78975 339750
rect 87373 339810 87439 339813
rect 131901 339810 131967 339813
rect 87373 339808 90028 339810
rect 87373 339752 87378 339808
rect 87434 339752 90028 339808
rect 87373 339750 90028 339752
rect 129772 339808 131967 339810
rect 129772 339752 131906 339808
rect 131962 339752 131967 339808
rect 129772 339750 131967 339752
rect 87373 339747 87439 339750
rect 131901 339747 131967 339750
rect 142990 339576 143050 339886
rect 233653 339944 237074 339946
rect 233653 339888 233658 339944
rect 233714 339888 237074 339944
rect 233653 339886 237074 339888
rect 233653 339883 233719 339886
rect 181581 339810 181647 339813
rect 225925 339810 225991 339813
rect 181581 339808 184052 339810
rect 181581 339752 181586 339808
rect 181642 339752 184052 339808
rect 181581 339750 184052 339752
rect 223796 339808 225991 339810
rect 223796 339752 225930 339808
rect 225986 339752 225991 339808
rect 223796 339750 225991 339752
rect 181581 339747 181647 339750
rect 225925 339747 225991 339750
rect 237014 339576 237074 339886
rect 327125 339944 331098 339946
rect 327125 339888 327130 339944
rect 327186 339888 331098 339944
rect 327125 339886 331098 339888
rect 327125 339883 327191 339886
rect 275053 339810 275119 339813
rect 321237 339810 321303 339813
rect 275053 339808 278076 339810
rect 275053 339752 275058 339808
rect 275114 339752 278076 339808
rect 275053 339750 278076 339752
rect 317820 339808 321303 339810
rect 317820 339752 321242 339808
rect 321298 339752 321303 339808
rect 317820 339750 321303 339752
rect 275053 339747 275119 339750
rect 321237 339747 321303 339750
rect 331038 339576 331098 339886
rect 173669 339538 173735 339541
rect 266589 339538 266655 339541
rect 170804 339536 173735 339538
rect 170804 339480 173674 339536
rect 173730 339480 173735 339536
rect 170804 339478 173735 339480
rect 264828 339536 266655 339538
rect 264828 339480 266594 339536
rect 266650 339480 266655 339536
rect 264828 339478 266655 339480
rect 173669 339475 173735 339478
rect 266589 339475 266655 339478
rect 87925 338858 87991 338861
rect 131809 338858 131875 338861
rect 87925 338856 90028 338858
rect 87925 338800 87930 338856
rect 87986 338800 90028 338856
rect 87925 338798 90028 338800
rect 129772 338856 131875 338858
rect 129772 338800 131814 338856
rect 131870 338800 131875 338856
rect 129772 338798 131875 338800
rect 87925 338795 87991 338798
rect 131809 338795 131875 338798
rect 182317 338858 182383 338861
rect 226477 338858 226543 338861
rect 182317 338856 184052 338858
rect 182317 338800 182322 338856
rect 182378 338800 184052 338856
rect 182317 338798 184052 338800
rect 223796 338856 226543 338858
rect 223796 338800 226482 338856
rect 226538 338800 226543 338856
rect 223796 338798 226543 338800
rect 182317 338795 182383 338798
rect 226477 338795 226543 338798
rect 275605 338858 275671 338861
rect 321605 338858 321671 338861
rect 275605 338856 278076 338858
rect 275605 338800 275610 338856
rect 275666 338800 278076 338856
rect 275605 338798 278076 338800
rect 317820 338856 321671 338858
rect 317820 338800 321610 338856
rect 321666 338800 321671 338856
rect 317820 338798 321671 338800
rect 275605 338795 275671 338798
rect 321605 338795 321671 338798
rect 139721 338586 139787 338589
rect 174037 338586 174103 338589
rect 139721 338584 143020 338586
rect 76198 338450 76258 338556
rect 139721 338528 139726 338584
rect 139782 338528 143020 338584
rect 139721 338526 143020 338528
rect 170804 338584 174103 338586
rect 170804 338528 174042 338584
rect 174098 338528 174103 338584
rect 170804 338526 174103 338528
rect 139721 338523 139787 338526
rect 174037 338523 174103 338526
rect 233561 338586 233627 338589
rect 266589 338586 266655 338589
rect 233561 338584 237044 338586
rect 233561 338528 233566 338584
rect 233622 338528 237044 338584
rect 233561 338526 237044 338528
rect 264828 338584 266655 338586
rect 264828 338528 266594 338584
rect 266650 338528 266655 338584
rect 264828 338526 266655 338528
rect 233561 338523 233627 338526
rect 266589 338523 266655 338526
rect 327217 338586 327283 338589
rect 327217 338584 331068 338586
rect 327217 338528 327222 338584
rect 327278 338528 331068 338584
rect 327217 338526 331068 338528
rect 327217 338523 327283 338526
rect 80197 338450 80263 338453
rect 76198 338448 80263 338450
rect 76198 338392 80202 338448
rect 80258 338392 80263 338448
rect 76198 338390 80263 338392
rect 80197 338387 80263 338390
rect 139905 338178 139971 338181
rect 233745 338178 233811 338181
rect 327033 338178 327099 338181
rect 139905 338176 143050 338178
rect 139905 338120 139910 338176
rect 139966 338120 143050 338176
rect 139905 338118 143050 338120
rect 139905 338115 139971 338118
rect 78909 338042 78975 338045
rect 76382 338040 78975 338042
rect 76382 337984 78914 338040
rect 78970 337984 78975 338040
rect 76382 337982 78975 337984
rect 9896 337498 10376 337528
rect 13313 337498 13379 337501
rect 9896 337496 13379 337498
rect 9896 337440 13318 337496
rect 13374 337440 13379 337496
rect 76382 337468 76442 337982
rect 78909 337979 78975 337982
rect 88017 338042 88083 338045
rect 131809 338042 131875 338045
rect 88017 338040 90028 338042
rect 88017 337984 88022 338040
rect 88078 337984 90028 338040
rect 88017 337982 90028 337984
rect 129772 338040 131875 338042
rect 129772 337984 131814 338040
rect 131870 337984 131875 338040
rect 129772 337982 131875 337984
rect 88017 337979 88083 337982
rect 131809 337979 131875 337982
rect 142990 337536 143050 338118
rect 233745 338176 237074 338178
rect 233745 338120 233750 338176
rect 233806 338120 237074 338176
rect 233745 338118 237074 338120
rect 233745 338115 233811 338118
rect 225925 338042 225991 338045
rect 223796 338040 225991 338042
rect 173945 337498 174011 337501
rect 170804 337496 174011 337498
rect 9896 337438 13379 337440
rect 170804 337440 173950 337496
rect 174006 337440 174011 337496
rect 170804 337438 174011 337440
rect 9896 337408 10376 337438
rect 13313 337435 13379 337438
rect 173945 337435 174011 337438
rect 180385 337498 180451 337501
rect 184022 337498 184082 338012
rect 223796 337984 225930 338040
rect 225986 337984 225991 338040
rect 223796 337982 225991 337984
rect 225925 337979 225991 337982
rect 237014 337536 237074 338118
rect 327033 338176 331098 338178
rect 327033 338120 327038 338176
rect 327094 338120 331098 338176
rect 327033 338118 331098 338120
rect 327033 338115 327099 338118
rect 274869 338042 274935 338045
rect 321605 338042 321671 338045
rect 274869 338040 278076 338042
rect 274869 337984 274874 338040
rect 274930 337984 278076 338040
rect 274869 337982 278076 337984
rect 317820 338040 321671 338042
rect 317820 337984 321610 338040
rect 321666 337984 321671 338040
rect 317820 337982 321671 337984
rect 274869 337979 274935 337982
rect 321605 337979 321671 337982
rect 331038 337536 331098 338118
rect 266681 337498 266747 337501
rect 180385 337496 184082 337498
rect 180385 337440 180390 337496
rect 180446 337440 184082 337496
rect 180385 337438 184082 337440
rect 264828 337496 266747 337498
rect 264828 337440 266686 337496
rect 266742 337440 266747 337496
rect 264828 337438 266747 337440
rect 180385 337435 180451 337438
rect 266681 337435 266747 337438
rect 87373 337090 87439 337093
rect 131901 337090 131967 337093
rect 87373 337088 90028 337090
rect 87373 337032 87378 337088
rect 87434 337032 90028 337088
rect 87373 337030 90028 337032
rect 129772 337088 131967 337090
rect 129772 337032 131906 337088
rect 131962 337032 131967 337088
rect 129772 337030 131967 337032
rect 87373 337027 87439 337030
rect 131901 337027 131967 337030
rect 181581 337090 181647 337093
rect 225925 337090 225991 337093
rect 181581 337088 184052 337090
rect 181581 337032 181586 337088
rect 181642 337032 184052 337088
rect 181581 337030 184052 337032
rect 223796 337088 225991 337090
rect 223796 337032 225930 337088
rect 225986 337032 225991 337088
rect 223796 337030 225991 337032
rect 181581 337027 181647 337030
rect 225925 337027 225991 337030
rect 233469 337090 233535 337093
rect 274869 337090 274935 337093
rect 321421 337090 321487 337093
rect 233469 337088 237074 337090
rect 233469 337032 233474 337088
rect 233530 337032 237074 337088
rect 233469 337030 237074 337032
rect 233469 337027 233535 337030
rect 139721 336818 139787 336821
rect 139721 336816 143050 336818
rect 139721 336760 139726 336816
rect 139782 336760 143050 336816
rect 139721 336758 143050 336760
rect 139721 336755 139787 336758
rect 142990 336448 143050 336758
rect 237014 336448 237074 337030
rect 274869 337088 278076 337090
rect 274869 337032 274874 337088
rect 274930 337032 278076 337088
rect 274869 337030 278076 337032
rect 317820 337088 321487 337090
rect 317820 337032 321426 337088
rect 321482 337032 321487 337088
rect 317820 337030 321487 337032
rect 274869 337027 274935 337030
rect 321421 337027 321487 337030
rect 326941 337090 327007 337093
rect 326941 337088 331098 337090
rect 326941 337032 326946 337088
rect 327002 337032 331098 337088
rect 326941 337030 331098 337032
rect 326941 337027 327007 337030
rect 331038 336448 331098 337030
rect 173485 336410 173551 336413
rect 266589 336410 266655 336413
rect 170804 336408 173551 336410
rect 76198 336274 76258 336380
rect 170804 336352 173490 336408
rect 173546 336352 173551 336408
rect 170804 336350 173551 336352
rect 264828 336408 266655 336410
rect 264828 336352 266594 336408
rect 266650 336352 266655 336408
rect 264828 336350 266655 336352
rect 173485 336347 173551 336350
rect 266589 336347 266655 336350
rect 80197 336274 80263 336277
rect 76198 336272 80263 336274
rect 76198 336216 80202 336272
rect 80258 336216 80263 336272
rect 76198 336214 80263 336216
rect 80197 336211 80263 336214
rect 87833 336274 87899 336277
rect 131809 336274 131875 336277
rect 226477 336274 226543 336277
rect 87833 336272 90028 336274
rect 87833 336216 87838 336272
rect 87894 336216 90028 336272
rect 87833 336214 90028 336216
rect 129772 336272 131875 336274
rect 129772 336216 131814 336272
rect 131870 336216 131875 336272
rect 223796 336272 226543 336274
rect 129772 336214 131875 336216
rect 87833 336211 87899 336214
rect 131809 336211 131875 336214
rect 180937 336138 181003 336141
rect 184022 336138 184082 336244
rect 223796 336216 226482 336272
rect 226538 336216 226543 336272
rect 223796 336214 226543 336216
rect 226477 336211 226543 336214
rect 274961 336274 275027 336277
rect 321605 336274 321671 336277
rect 274961 336272 278076 336274
rect 274961 336216 274966 336272
rect 275022 336216 278076 336272
rect 274961 336214 278076 336216
rect 317820 336272 321671 336274
rect 317820 336216 321610 336272
rect 321666 336216 321671 336272
rect 317820 336214 321671 336216
rect 274961 336211 275027 336214
rect 321605 336211 321671 336214
rect 180937 336136 184082 336138
rect 180937 336080 180942 336136
rect 180998 336080 184082 336136
rect 180937 336078 184082 336080
rect 180937 336075 181003 336078
rect 139629 335866 139695 335869
rect 233469 335866 233535 335869
rect 327125 335866 327191 335869
rect 139629 335864 143050 335866
rect 139629 335808 139634 335864
rect 139690 335808 143050 335864
rect 139629 335806 143050 335808
rect 139629 335803 139695 335806
rect 142990 335496 143050 335806
rect 233469 335864 237074 335866
rect 233469 335808 233474 335864
rect 233530 335808 237074 335864
rect 233469 335806 237074 335808
rect 233469 335803 233535 335806
rect 237014 335496 237074 335806
rect 327125 335864 331098 335866
rect 327125 335808 327130 335864
rect 327186 335808 331098 335864
rect 327125 335806 331098 335808
rect 327125 335803 327191 335806
rect 331038 335496 331098 335806
rect 173301 335458 173367 335461
rect 266589 335458 266655 335461
rect 170804 335456 173367 335458
rect 76198 335322 76258 335428
rect 170804 335400 173306 335456
rect 173362 335400 173367 335456
rect 170804 335398 173367 335400
rect 264828 335456 266655 335458
rect 264828 335400 266594 335456
rect 266650 335400 266655 335456
rect 264828 335398 266655 335400
rect 173301 335395 173367 335398
rect 266589 335395 266655 335398
rect 80197 335322 80263 335325
rect 76198 335320 80263 335322
rect 76198 335264 80202 335320
rect 80258 335264 80263 335320
rect 76198 335262 80263 335264
rect 80197 335259 80263 335262
rect 139629 334370 139695 334373
rect 173393 334370 173459 334373
rect 139629 334368 143020 334370
rect 76198 334234 76258 334340
rect 139629 334312 139634 334368
rect 139690 334312 143020 334368
rect 139629 334310 143020 334312
rect 170804 334368 173459 334370
rect 170804 334312 173398 334368
rect 173454 334312 173459 334368
rect 170804 334310 173459 334312
rect 139629 334307 139695 334310
rect 173393 334307 173459 334310
rect 233653 334370 233719 334373
rect 266589 334370 266655 334373
rect 233653 334368 237044 334370
rect 233653 334312 233658 334368
rect 233714 334312 237044 334368
rect 233653 334310 237044 334312
rect 264828 334368 266655 334370
rect 264828 334312 266594 334368
rect 266650 334312 266655 334368
rect 264828 334310 266655 334312
rect 233653 334307 233719 334310
rect 266589 334307 266655 334310
rect 326665 334370 326731 334373
rect 326665 334368 331068 334370
rect 326665 334312 326670 334368
rect 326726 334312 331068 334368
rect 326665 334310 331068 334312
rect 326665 334307 326731 334310
rect 80197 334234 80263 334237
rect 76198 334232 80263 334234
rect 76198 334176 80202 334232
rect 80258 334176 80263 334232
rect 76198 334174 80263 334176
rect 80197 334171 80263 334174
rect 139629 333962 139695 333965
rect 233469 333962 233535 333965
rect 327033 333962 327099 333965
rect 139629 333960 143050 333962
rect 139629 333904 139634 333960
rect 139690 333904 143050 333960
rect 139629 333902 143050 333904
rect 139629 333899 139695 333902
rect 95193 333826 95259 333829
rect 104894 333826 104900 333828
rect 95193 333824 104900 333826
rect 95193 333768 95198 333824
rect 95254 333768 104900 333824
rect 95193 333766 104900 333768
rect 95193 333763 95259 333766
rect 104894 333764 104900 333766
rect 104964 333764 104970 333828
rect 78909 333690 78975 333693
rect 76382 333688 78975 333690
rect 76382 333632 78914 333688
rect 78970 333632 78975 333688
rect 76382 333630 78975 333632
rect 76382 333252 76442 333630
rect 78909 333627 78975 333630
rect 142990 333320 143050 333902
rect 233469 333960 237074 333962
rect 233469 333904 233474 333960
rect 233530 333904 237074 333960
rect 233469 333902 237074 333904
rect 233469 333899 233535 333902
rect 212166 333492 212172 333556
rect 212236 333554 212242 333556
rect 212309 333554 212375 333557
rect 212236 333552 212375 333554
rect 212236 333496 212314 333552
rect 212370 333496 212375 333552
rect 212236 333494 212375 333496
rect 212236 333492 212242 333494
rect 212309 333491 212375 333494
rect 237014 333320 237074 333902
rect 327033 333960 331098 333962
rect 327033 333904 327038 333960
rect 327094 333904 331098 333960
rect 327033 333902 331098 333904
rect 327033 333899 327099 333902
rect 331038 333320 331098 333902
rect 173301 333282 173367 333285
rect 266681 333282 266747 333285
rect 170804 333280 173367 333282
rect 170804 333224 173306 333280
rect 173362 333224 173367 333280
rect 170804 333222 173367 333224
rect 264828 333280 266747 333282
rect 264828 333224 266686 333280
rect 266742 333224 266747 333280
rect 264828 333222 266747 333224
rect 173301 333219 173367 333222
rect 266681 333219 266747 333222
rect 201821 333146 201887 333149
rect 225465 333146 225531 333149
rect 230801 333146 230867 333149
rect 201821 333144 230867 333146
rect 201821 333088 201826 333144
rect 201882 333088 225470 333144
rect 225526 333088 230806 333144
rect 230862 333088 230867 333144
rect 201821 333086 230867 333088
rect 201821 333083 201887 333086
rect 225465 333083 225531 333086
rect 230801 333083 230867 333086
rect 295518 333084 295524 333148
rect 295588 333146 295594 333148
rect 296213 333146 296279 333149
rect 319305 333146 319371 333149
rect 295588 333144 319371 333146
rect 295588 333088 296218 333144
rect 296274 333088 319310 333144
rect 319366 333088 319371 333144
rect 295588 333086 319371 333088
rect 295588 333084 295594 333086
rect 296213 333083 296279 333086
rect 319305 333083 319371 333086
rect 139629 333010 139695 333013
rect 233469 333010 233535 333013
rect 327309 333010 327375 333013
rect 139629 333008 143050 333010
rect 139629 332952 139634 333008
rect 139690 332952 143050 333008
rect 139629 332950 143050 332952
rect 139629 332947 139695 332950
rect 80197 332738 80263 332741
rect 76382 332736 80263 332738
rect 76382 332680 80202 332736
rect 80258 332680 80263 332736
rect 76382 332678 80263 332680
rect 76382 332300 76442 332678
rect 80197 332675 80263 332678
rect 142990 332368 143050 332950
rect 233469 333008 237074 333010
rect 233469 332952 233474 333008
rect 233530 332952 237074 333008
rect 233469 332950 237074 332952
rect 233469 332947 233535 332950
rect 237014 332368 237074 332950
rect 327309 333008 331098 333010
rect 327309 332952 327314 333008
rect 327370 332952 331098 333008
rect 327309 332950 331098 332952
rect 327309 332947 327375 332950
rect 331038 332368 331098 332950
rect 172841 332330 172907 332333
rect 266589 332330 266655 332333
rect 170804 332328 172907 332330
rect 170804 332272 172846 332328
rect 172902 332272 172907 332328
rect 170804 332270 172907 332272
rect 264828 332328 266655 332330
rect 264828 332272 266594 332328
rect 266650 332272 266655 332328
rect 264828 332270 266655 332272
rect 172841 332267 172907 332270
rect 266589 332267 266655 332270
rect 136961 332194 137027 332197
rect 137278 332194 137284 332196
rect 136961 332192 137284 332194
rect 136961 332136 136966 332192
rect 137022 332136 137284 332192
rect 136961 332134 137284 332136
rect 136961 332131 137027 332134
rect 137278 332132 137284 332134
rect 137348 332132 137354 332196
rect 201678 332132 201684 332196
rect 201748 332194 201754 332196
rect 201821 332194 201887 332197
rect 201748 332192 201887 332194
rect 201748 332136 201826 332192
rect 201882 332136 201887 332192
rect 201748 332134 201887 332136
rect 201748 332132 201754 332134
rect 201821 332131 201887 332134
rect 230893 332196 230959 332197
rect 230893 332192 230940 332196
rect 231004 332194 231010 332196
rect 230893 332136 230898 332192
rect 230893 332132 230940 332136
rect 231004 332134 231050 332194
rect 231004 332132 231010 332134
rect 230893 332131 230959 332132
rect 139629 331650 139695 331653
rect 139629 331648 143050 331650
rect 139629 331592 139634 331648
rect 139690 331592 143050 331648
rect 139629 331590 143050 331592
rect 139629 331587 139695 331590
rect 142990 331280 143050 331590
rect 204438 331588 204444 331652
rect 204508 331650 204514 331652
rect 205593 331650 205659 331653
rect 225373 331650 225439 331653
rect 230934 331650 230940 331652
rect 204508 331648 230940 331650
rect 204508 331592 205598 331648
rect 205654 331592 225378 331648
rect 225434 331592 230940 331648
rect 204508 331590 230940 331592
rect 204508 331588 204514 331590
rect 205593 331587 205659 331590
rect 225373 331587 225439 331590
rect 230934 331588 230940 331590
rect 231004 331588 231010 331652
rect 292901 331650 292967 331653
rect 319397 331650 319463 331653
rect 292901 331648 319463 331650
rect 292901 331592 292906 331648
rect 292962 331592 319402 331648
rect 319458 331592 319463 331648
rect 292901 331590 319463 331592
rect 292901 331587 292967 331590
rect 319397 331587 319463 331590
rect 327217 331650 327283 331653
rect 327217 331648 331098 331650
rect 327217 331592 327222 331648
rect 327278 331592 331098 331648
rect 327217 331590 331098 331592
rect 327217 331587 327283 331590
rect 233469 331514 233535 331517
rect 233469 331512 237074 331514
rect 233469 331456 233474 331512
rect 233530 331456 237074 331512
rect 233469 331454 237074 331456
rect 233469 331451 233535 331454
rect 237014 331280 237074 331454
rect 299382 331452 299388 331516
rect 299452 331514 299458 331516
rect 299525 331514 299591 331517
rect 299452 331512 299591 331514
rect 299452 331456 299530 331512
rect 299586 331456 299591 331512
rect 299452 331454 299591 331456
rect 299452 331452 299458 331454
rect 299525 331451 299591 331454
rect 331038 331280 331098 331590
rect 173669 331242 173735 331245
rect 266589 331242 266655 331245
rect 170804 331240 173735 331242
rect 76198 330970 76258 331212
rect 170804 331184 173674 331240
rect 173730 331184 173735 331240
rect 170804 331182 173735 331184
rect 264828 331240 266655 331242
rect 264828 331184 266594 331240
rect 266650 331184 266655 331240
rect 264828 331182 266655 331184
rect 173669 331179 173735 331182
rect 266589 331179 266655 331182
rect 80197 330970 80263 330973
rect 76198 330968 80263 330970
rect 76198 330912 80202 330968
rect 80258 330912 80263 330968
rect 76198 330910 80263 330912
rect 80197 330907 80263 330910
rect 137053 330834 137119 330837
rect 137278 330834 137284 330836
rect 137053 330832 137284 330834
rect 137053 330776 137058 330832
rect 137114 330776 137284 330832
rect 137053 330774 137284 330776
rect 137053 330771 137119 330774
rect 137278 330772 137284 330774
rect 137348 330772 137354 330836
rect 230801 330834 230867 330837
rect 231302 330834 231308 330836
rect 230801 330832 231308 330834
rect 230801 330776 230806 330832
rect 230862 330776 231308 330832
rect 230801 330774 231308 330776
rect 230801 330771 230867 330774
rect 231302 330772 231308 330774
rect 231372 330772 231378 330836
rect 292758 330772 292764 330836
rect 292828 330834 292834 330836
rect 292901 330834 292967 330837
rect 292828 330832 292967 330834
rect 292828 330776 292906 330832
rect 292962 330776 292967 330832
rect 292828 330774 292967 330776
rect 292828 330772 292834 330774
rect 292901 330771 292967 330774
rect 140365 330290 140431 330293
rect 172105 330290 172171 330293
rect 140365 330288 143020 330290
rect 76198 329746 76258 330260
rect 140365 330232 140370 330288
rect 140426 330232 143020 330288
rect 140365 330230 143020 330232
rect 170804 330288 172171 330290
rect 170804 330232 172110 330288
rect 172166 330232 172171 330288
rect 170804 330230 172171 330232
rect 140365 330227 140431 330230
rect 172105 330227 172171 330230
rect 233469 330290 233535 330293
rect 266589 330290 266655 330293
rect 233469 330288 237044 330290
rect 233469 330232 233474 330288
rect 233530 330232 237044 330288
rect 233469 330230 237044 330232
rect 264828 330288 266655 330290
rect 264828 330232 266594 330288
rect 266650 330232 266655 330288
rect 264828 330230 266655 330232
rect 233469 330227 233535 330230
rect 266589 330227 266655 330230
rect 328413 330290 328479 330293
rect 328413 330288 331068 330290
rect 328413 330232 328418 330288
rect 328474 330232 331068 330288
rect 328413 330230 331068 330232
rect 328413 330227 328479 330230
rect 158581 330156 158647 330157
rect 159593 330156 159659 330157
rect 251961 330156 252027 330157
rect 158581 330154 158628 330156
rect 158536 330152 158628 330154
rect 158536 330096 158586 330152
rect 158536 330094 158628 330096
rect 158581 330092 158628 330094
rect 158692 330092 158698 330156
rect 159542 330092 159548 330156
rect 159612 330154 159659 330156
rect 159612 330152 159704 330154
rect 159654 330096 159704 330152
rect 159612 330094 159704 330096
rect 159612 330092 159659 330094
rect 251910 330092 251916 330156
rect 251980 330154 252027 330156
rect 252605 330156 252671 330157
rect 252605 330154 252652 330156
rect 251980 330152 252072 330154
rect 252022 330096 252072 330152
rect 251980 330094 252072 330096
rect 252560 330152 252652 330154
rect 252560 330096 252610 330152
rect 252560 330094 252652 330096
rect 251980 330092 252027 330094
rect 158581 330091 158647 330092
rect 159593 330091 159659 330092
rect 251961 330091 252027 330092
rect 252605 330092 252652 330094
rect 252716 330092 252722 330156
rect 429429 330154 429495 330157
rect 434416 330154 434896 330184
rect 429429 330152 434896 330154
rect 429429 330096 429434 330152
rect 429490 330096 434896 330152
rect 429429 330094 434896 330096
rect 252605 330091 252671 330092
rect 429429 330091 429495 330094
rect 434416 330064 434896 330094
rect 78909 329746 78975 329749
rect 76198 329744 78975 329746
rect 76198 329688 78914 329744
rect 78970 329688 78975 329744
rect 76198 329686 78975 329688
rect 78909 329683 78975 329686
rect 137237 328794 137303 328797
rect 161709 328796 161775 328797
rect 230985 328796 231051 328797
rect 137462 328794 137468 328796
rect 137237 328792 137468 328794
rect 137237 328736 137242 328792
rect 137298 328736 137468 328792
rect 137237 328734 137468 328736
rect 137237 328731 137303 328734
rect 137462 328732 137468 328734
rect 137532 328732 137538 328796
rect 161709 328794 161756 328796
rect 161664 328792 161756 328794
rect 161664 328736 161714 328792
rect 161664 328734 161756 328736
rect 161709 328732 161756 328734
rect 161820 328732 161826 328796
rect 230934 328794 230940 328796
rect 230858 328734 230940 328794
rect 231004 328794 231051 328796
rect 231854 328794 231860 328796
rect 231004 328792 231860 328794
rect 231046 328736 231860 328792
rect 230934 328732 230940 328734
rect 231004 328734 231860 328736
rect 231004 328732 231051 328734
rect 231854 328732 231860 328734
rect 231924 328732 231930 328796
rect 253382 328732 253388 328796
rect 253452 328794 253458 328796
rect 253525 328794 253591 328797
rect 253452 328792 253591 328794
rect 253452 328736 253530 328792
rect 253586 328736 253591 328792
rect 253452 328734 253591 328736
rect 253452 328732 253458 328734
rect 161709 328731 161775 328732
rect 230985 328731 231051 328732
rect 253525 328731 253591 328734
rect 137145 328114 137211 328117
rect 160697 328116 160763 328117
rect 208721 328116 208787 328117
rect 137462 328114 137468 328116
rect 137145 328112 137468 328114
rect 137145 328056 137150 328112
rect 137206 328056 137468 328112
rect 137145 328054 137468 328056
rect 137145 328051 137211 328054
rect 137462 328052 137468 328054
rect 137532 328052 137538 328116
rect 160646 328052 160652 328116
rect 160716 328114 160763 328116
rect 160716 328112 160808 328114
rect 160758 328056 160808 328112
rect 160716 328054 160808 328056
rect 160716 328052 160763 328054
rect 208670 328052 208676 328116
rect 208740 328114 208787 328116
rect 208740 328112 208832 328114
rect 208782 328056 208832 328112
rect 208740 328054 208832 328056
rect 208740 328052 208787 328054
rect 160697 328051 160763 328052
rect 208721 328051 208787 328052
rect 339177 327434 339243 327437
rect 339494 327434 339500 327436
rect 339177 327432 339500 327434
rect 339177 327376 339182 327432
rect 339238 327376 339500 327432
rect 339177 327374 339500 327376
rect 339177 327371 339243 327374
rect 339494 327372 339500 327374
rect 339564 327372 339570 327436
rect 340005 327434 340071 327437
rect 340966 327434 340972 327436
rect 340005 327432 340972 327434
rect 340005 327376 340010 327432
rect 340066 327376 340972 327432
rect 340005 327374 340972 327376
rect 340005 327371 340071 327374
rect 340966 327372 340972 327374
rect 341036 327372 341042 327436
rect 324549 326890 324615 326893
rect 336366 326890 336372 326892
rect 324549 326888 336372 326890
rect 324549 326832 324554 326888
rect 324610 326832 336372 326888
rect 324549 326830 336372 326832
rect 324549 326827 324615 326830
rect 336366 326828 336372 326830
rect 336436 326890 336442 326892
rect 342489 326890 342555 326893
rect 336436 326888 342555 326890
rect 336436 326832 342494 326888
rect 342550 326832 342555 326888
rect 336436 326830 342555 326832
rect 336436 326828 336442 326830
rect 342489 326827 342555 326830
rect 9896 326754 10376 326784
rect 14693 326754 14759 326757
rect 9896 326752 14759 326754
rect 9896 326696 14698 326752
rect 14754 326696 14759 326752
rect 9896 326694 14759 326696
rect 9896 326664 10376 326694
rect 14693 326691 14759 326694
rect 52638 326284 52644 326348
rect 52708 326346 52714 326348
rect 53057 326346 53123 326349
rect 52708 326344 53123 326346
rect 52708 326288 53062 326344
rect 53118 326288 53123 326344
rect 52708 326286 53123 326288
rect 52708 326284 52714 326286
rect 53057 326283 53123 326286
rect 54069 326346 54135 326349
rect 55081 326348 55147 326349
rect 54662 326346 54668 326348
rect 54069 326344 54668 326346
rect 54069 326288 54074 326344
rect 54130 326288 54668 326344
rect 54069 326286 54668 326288
rect 54069 326283 54135 326286
rect 54662 326284 54668 326286
rect 54732 326284 54738 326348
rect 55030 326346 55036 326348
rect 54990 326286 55036 326346
rect 55100 326344 55147 326348
rect 55142 326288 55147 326344
rect 55030 326284 55036 326286
rect 55100 326284 55147 326288
rect 55950 326284 55956 326348
rect 56020 326346 56026 326348
rect 56093 326346 56159 326349
rect 56020 326344 56159 326346
rect 56020 326288 56098 326344
rect 56154 326288 56159 326344
rect 56020 326286 56159 326288
rect 56020 326284 56026 326286
rect 55081 326283 55147 326284
rect 56093 326283 56159 326286
rect 352885 324850 352951 324853
rect 353069 324850 353135 324853
rect 352885 324848 353135 324850
rect 352885 324792 352890 324848
rect 352946 324792 353074 324848
rect 353130 324792 353135 324848
rect 352885 324790 353135 324792
rect 352885 324787 352951 324790
rect 353069 324787 353135 324790
rect 137237 320362 137303 320365
rect 231353 320362 231419 320365
rect 324733 320362 324799 320365
rect 134740 320360 137303 320362
rect 134740 320304 137242 320360
rect 137298 320304 137303 320360
rect 134740 320302 137303 320304
rect 228764 320360 231419 320362
rect 228764 320304 231358 320360
rect 231414 320304 231419 320360
rect 228764 320302 231419 320304
rect 322788 320360 324799 320362
rect 322788 320304 324738 320360
rect 324794 320304 324799 320360
rect 322788 320302 324799 320304
rect 137237 320299 137303 320302
rect 231353 320299 231419 320302
rect 324733 320299 324799 320302
rect 348101 320226 348167 320229
rect 353294 320226 353300 320228
rect 348101 320224 353300 320226
rect 348101 320168 348106 320224
rect 348162 320168 353300 320224
rect 348101 320166 353300 320168
rect 348101 320163 348167 320166
rect 353294 320164 353300 320166
rect 353364 320164 353370 320228
rect 429429 317914 429495 317917
rect 434416 317914 434896 317944
rect 429429 317912 434896 317914
rect 429429 317856 429434 317912
rect 429490 317856 434896 317912
rect 429429 317854 434896 317856
rect 429429 317851 429495 317854
rect 434416 317824 434896 317854
rect 137145 317234 137211 317237
rect 231353 317234 231419 317237
rect 324825 317234 324891 317237
rect 134740 317232 137211 317234
rect 134740 317176 137150 317232
rect 137206 317176 137211 317232
rect 134740 317174 137211 317176
rect 228764 317232 231419 317234
rect 228764 317176 231358 317232
rect 231414 317176 231419 317232
rect 228764 317174 231419 317176
rect 322788 317232 324891 317234
rect 322788 317176 324830 317232
rect 324886 317176 324891 317232
rect 322788 317174 324891 317176
rect 137145 317171 137211 317174
rect 231353 317171 231419 317174
rect 324825 317171 324891 317174
rect 246165 316964 246231 316965
rect 246165 316960 246212 316964
rect 246276 316962 246282 316964
rect 246165 316904 246170 316960
rect 246165 316900 246212 316904
rect 246276 316902 246322 316962
rect 246276 316900 246282 316902
rect 246165 316899 246231 316900
rect 345617 316690 345683 316693
rect 345574 316688 345683 316690
rect 345574 316632 345622 316688
rect 345678 316632 345683 316688
rect 345574 316627 345683 316632
rect 345574 316556 345634 316627
rect 345566 316492 345572 316556
rect 345636 316492 345642 316556
rect 9896 316010 10376 316040
rect 13313 316010 13379 316013
rect 9896 316008 13379 316010
rect 9896 315952 13318 316008
rect 13374 315952 13379 316008
rect 9896 315950 13379 315952
rect 9896 315920 10376 315950
rect 13313 315947 13379 315950
rect 55081 315874 55147 315877
rect 55950 315874 55956 315876
rect 55081 315872 55956 315874
rect 55081 315816 55086 315872
rect 55142 315816 55956 315872
rect 55081 315814 55956 315816
rect 55081 315811 55147 315814
rect 55950 315812 55956 315814
rect 56020 315812 56026 315876
rect 405969 315874 406035 315877
rect 405969 315872 409114 315874
rect 405969 315816 405974 315872
rect 406030 315816 409114 315872
rect 405969 315814 409114 315816
rect 405969 315811 406035 315814
rect 38797 315602 38863 315605
rect 35748 315600 38863 315602
rect 35748 315544 38802 315600
rect 38858 315544 38863 315600
rect 409054 315572 409114 315814
rect 35748 315542 38863 315544
rect 38797 315539 38863 315542
rect 355686 315330 355692 315332
rect 345574 315270 355692 315330
rect 324641 315194 324707 315197
rect 345574 315196 345634 315270
rect 355686 315268 355692 315270
rect 355756 315268 355762 315332
rect 345566 315194 345572 315196
rect 324641 315192 345572 315194
rect 324641 315136 324646 315192
rect 324702 315136 345572 315192
rect 324641 315134 345572 315136
rect 324641 315131 324707 315134
rect 345566 315132 345572 315134
rect 345636 315132 345642 315196
rect 70862 314514 70922 315028
rect 340966 314860 340972 314924
rect 341036 314922 341042 314924
rect 351822 314922 351828 314924
rect 341036 314862 351828 314922
rect 341036 314860 341042 314862
rect 351822 314860 351828 314862
rect 351892 314860 351898 314924
rect 339494 314588 339500 314652
rect 339564 314588 339570 314652
rect 352006 314588 352012 314652
rect 352076 314588 352082 314652
rect 74217 314514 74283 314517
rect 70862 314512 74283 314514
rect 70862 314456 74222 314512
rect 74278 314456 74283 314512
rect 70862 314454 74283 314456
rect 339502 314514 339562 314588
rect 352014 314514 352074 314588
rect 339502 314454 352074 314514
rect 74217 314451 74283 314454
rect 16073 313834 16139 313837
rect 19894 313834 19954 314348
rect 16073 313832 19954 313834
rect 16073 313776 16078 313832
rect 16134 313776 19954 313832
rect 16073 313774 19954 313776
rect 51585 313834 51651 313837
rect 55038 313834 55098 314280
rect 137053 314106 137119 314109
rect 230985 314106 231051 314109
rect 324641 314106 324707 314109
rect 134740 314104 137119 314106
rect 134740 314048 137058 314104
rect 137114 314048 137119 314104
rect 134740 314046 137119 314048
rect 228764 314104 231051 314106
rect 228764 314048 230990 314104
rect 231046 314048 231051 314104
rect 228764 314046 231051 314048
rect 322788 314104 324707 314106
rect 322788 314048 324646 314104
rect 324702 314048 324707 314104
rect 322788 314046 324707 314048
rect 352750 314106 352810 314280
rect 356197 314106 356263 314109
rect 352750 314104 356263 314106
rect 352750 314048 356202 314104
rect 356258 314048 356263 314104
rect 352750 314046 356263 314048
rect 137053 314043 137119 314046
rect 230985 314043 231051 314046
rect 324641 314043 324707 314046
rect 356197 314043 356263 314046
rect 51585 313832 55098 313834
rect 51585 313776 51590 313832
rect 51646 313776 55098 313832
rect 51585 313774 55098 313776
rect 424694 313834 424754 314280
rect 427313 313834 427379 313837
rect 424694 313832 427379 313834
rect 424694 313776 427318 313832
rect 427374 313776 427379 313832
rect 424694 313774 427379 313776
rect 16073 313771 16139 313774
rect 51585 313771 51651 313774
rect 427313 313771 427379 313774
rect 405969 313698 406035 313701
rect 405969 313696 409114 313698
rect 405969 313640 405974 313696
rect 406030 313640 409114 313696
rect 405969 313638 409114 313640
rect 405969 313635 406035 313638
rect 81669 313562 81735 313565
rect 175509 313562 175575 313565
rect 270269 313562 270335 313565
rect 81669 313560 85060 313562
rect 81669 313504 81674 313560
rect 81730 313504 85060 313560
rect 81669 313502 85060 313504
rect 175509 313560 178900 313562
rect 175509 313504 175514 313560
rect 175570 313504 178900 313560
rect 175509 313502 178900 313504
rect 270269 313560 272924 313562
rect 270269 313504 270274 313560
rect 270330 313504 272924 313560
rect 270269 313502 272924 313504
rect 81669 313499 81735 313502
rect 175509 313499 175575 313502
rect 270269 313499 270335 313502
rect 38429 313154 38495 313157
rect 35748 313152 38495 313154
rect 35748 313096 38434 313152
rect 38490 313096 38495 313152
rect 409054 313124 409114 313638
rect 35748 313094 38495 313096
rect 38429 313091 38495 313094
rect 70862 311114 70922 311356
rect 74125 311114 74191 311117
rect 70862 311112 74191 311114
rect 70862 311056 74130 311112
rect 74186 311056 74191 311112
rect 70862 311054 74191 311056
rect 74125 311051 74191 311054
rect 54069 310978 54135 310981
rect 54846 310978 54852 310980
rect 54069 310976 54852 310978
rect 54069 310920 54074 310976
rect 54130 310920 54852 310976
rect 54069 310918 54852 310920
rect 54069 310915 54135 310918
rect 54846 310916 54852 310918
rect 54916 310978 54922 310980
rect 55030 310978 55036 310980
rect 54916 310918 55036 310978
rect 54916 310916 54922 310918
rect 55030 310916 55036 310918
rect 55100 310916 55106 310980
rect 136961 310978 137027 310981
rect 230893 310978 230959 310981
rect 325377 310978 325443 310981
rect 134740 310976 137027 310978
rect 134740 310920 136966 310976
rect 137022 310920 137027 310976
rect 134740 310918 137027 310920
rect 228764 310976 230959 310978
rect 228764 310920 230898 310976
rect 230954 310920 230959 310976
rect 228764 310918 230959 310920
rect 322788 310976 325443 310978
rect 322788 310920 325382 310976
rect 325438 310920 325443 310976
rect 322788 310918 325443 310920
rect 136961 310915 137027 310918
rect 230893 310915 230959 310918
rect 325377 310915 325443 310918
rect 35718 310434 35778 310472
rect 38797 310434 38863 310437
rect 35718 310432 38863 310434
rect 35718 310376 38802 310432
rect 38858 310376 38863 310432
rect 35718 310374 38863 310376
rect 38797 310371 38863 310374
rect 405969 310434 406035 310437
rect 408870 310434 408930 310540
rect 405969 310432 408930 310434
rect 405969 310376 405974 310432
rect 406030 310376 408930 310432
rect 405969 310374 408930 310376
rect 405969 310371 406035 310374
rect 148326 310170 148908 310230
rect 242350 310170 242932 310230
rect 145517 310162 145583 310165
rect 148326 310162 148386 310170
rect 145517 310160 148386 310162
rect 145517 310104 145522 310160
rect 145578 310104 148386 310160
rect 145517 310102 148386 310104
rect 240645 310162 240711 310165
rect 242350 310162 242410 310170
rect 240645 310160 242410 310162
rect 240645 310104 240650 310160
rect 240706 310104 242410 310160
rect 240645 310102 242410 310104
rect 145517 310099 145583 310102
rect 240645 310099 240711 310102
rect 334209 309754 334275 309757
rect 336926 309754 336986 310200
rect 334209 309752 336986 309754
rect 334209 309696 334214 309752
rect 334270 309696 336986 309752
rect 334209 309694 336986 309696
rect 334209 309691 334275 309694
rect 16257 308394 16323 308397
rect 19894 308394 19954 309316
rect 51217 308666 51283 308669
rect 55038 308666 55098 309248
rect 51217 308664 55098 308666
rect 51217 308608 51222 308664
rect 51278 308608 55098 308664
rect 51217 308606 55098 308608
rect 352750 308666 352810 309248
rect 356197 308666 356263 308669
rect 352750 308664 356263 308666
rect 352750 308608 356202 308664
rect 356258 308608 356263 308664
rect 352750 308606 356263 308608
rect 424694 308666 424754 309248
rect 428693 308666 428759 308669
rect 424694 308664 428759 308666
rect 424694 308608 428698 308664
rect 428754 308608 428759 308664
rect 424694 308606 428759 308608
rect 51217 308603 51283 308606
rect 356197 308603 356263 308606
rect 428693 308603 428759 308606
rect 16257 308392 19954 308394
rect 16257 308336 16262 308392
rect 16318 308336 19954 308392
rect 16257 308334 19954 308336
rect 16257 308331 16323 308334
rect 55030 308196 55036 308260
rect 55100 308196 55106 308260
rect 73430 308258 73436 308260
rect 70678 308198 73436 308258
rect 55038 308125 55098 308196
rect 38797 308122 38863 308125
rect 35748 308120 38863 308122
rect 35748 308064 38802 308120
rect 38858 308064 38863 308120
rect 35748 308062 38863 308064
rect 55038 308120 55147 308125
rect 55038 308064 55086 308120
rect 55142 308064 55147 308120
rect 55038 308062 55147 308064
rect 38797 308059 38863 308062
rect 55081 308059 55147 308062
rect 70678 307684 70738 308198
rect 73430 308196 73436 308198
rect 73500 308258 73506 308260
rect 74309 308258 74375 308261
rect 324733 308258 324799 308261
rect 325561 308258 325627 308261
rect 73500 308256 74375 308258
rect 73500 308200 74314 308256
rect 74370 308200 74375 308256
rect 73500 308198 74375 308200
rect 73500 308196 73506 308198
rect 74309 308195 74375 308198
rect 322758 308256 325627 308258
rect 322758 308200 324738 308256
rect 324794 308200 325566 308256
rect 325622 308200 325627 308256
rect 322758 308198 325627 308200
rect 137513 307850 137579 307853
rect 230801 307850 230867 307853
rect 134740 307848 137579 307850
rect 134740 307792 137518 307848
rect 137574 307792 137579 307848
rect 134740 307790 137579 307792
rect 228764 307848 230867 307850
rect 228764 307792 230806 307848
rect 230862 307792 230867 307848
rect 322758 307820 322818 308198
rect 324733 308195 324799 308198
rect 325561 308195 325627 308198
rect 405969 308258 406035 308261
rect 405969 308256 409114 308258
rect 405969 308200 405974 308256
rect 406030 308200 409114 308256
rect 405969 308198 409114 308200
rect 405969 308195 406035 308198
rect 409054 308092 409114 308198
rect 228764 307790 230867 307792
rect 137513 307787 137579 307790
rect 230801 307787 230867 307790
rect 54069 306218 54135 306221
rect 54662 306218 54668 306220
rect 54069 306216 54668 306218
rect 54069 306160 54074 306216
rect 54130 306160 54668 306216
rect 54069 306158 54668 306160
rect 54069 306155 54135 306158
rect 54662 306156 54668 306158
rect 54732 306156 54738 306220
rect 164702 306218 164762 306800
rect 167873 306218 167939 306221
rect 164702 306216 167939 306218
rect 164702 306160 167878 306216
rect 167934 306160 167939 306216
rect 164702 306158 167939 306160
rect 258726 306218 258786 306800
rect 261713 306218 261779 306221
rect 258726 306216 261779 306218
rect 258726 306160 261718 306216
rect 261774 306160 261779 306216
rect 258726 306158 261779 306160
rect 167873 306155 167939 306158
rect 261713 306155 261779 306158
rect 406061 306218 406127 306221
rect 406061 306216 409114 306218
rect 406061 306160 406066 306216
rect 406122 306160 409114 306216
rect 406061 306158 409114 306160
rect 406061 306155 406127 306158
rect 38797 305674 38863 305677
rect 35748 305672 38863 305674
rect 35748 305616 38802 305672
rect 38858 305616 38863 305672
rect 409054 305644 409114 306158
rect 429470 305748 429476 305812
rect 429540 305810 429546 305812
rect 434416 305810 434896 305840
rect 429540 305750 434896 305810
rect 429540 305748 429546 305750
rect 434416 305720 434896 305750
rect 35748 305614 38863 305616
rect 38797 305611 38863 305614
rect 9896 305130 10376 305160
rect 13405 305130 13471 305133
rect 9896 305128 13471 305130
rect 9896 305072 13410 305128
rect 13466 305072 13471 305128
rect 9896 305070 13471 305072
rect 9896 305040 10376 305070
rect 13405 305067 13471 305070
rect 73389 304722 73455 304725
rect 136869 304722 136935 304725
rect 137513 304722 137579 304725
rect 231997 304722 232063 304725
rect 325285 304722 325351 304725
rect 70678 304720 73455 304722
rect 70678 304664 73394 304720
rect 73450 304664 73455 304720
rect 70678 304662 73455 304664
rect 134740 304720 137579 304722
rect 134740 304664 136874 304720
rect 136930 304664 137518 304720
rect 137574 304664 137579 304720
rect 134740 304662 137579 304664
rect 228764 304720 232063 304722
rect 228764 304664 232002 304720
rect 232058 304664 232063 304720
rect 228764 304662 232063 304664
rect 322788 304720 325351 304722
rect 322788 304664 325290 304720
rect 325346 304664 325351 304720
rect 322788 304662 325351 304664
rect 51861 304314 51927 304317
rect 51861 304312 55068 304314
rect 16441 304178 16507 304181
rect 19894 304178 19954 304284
rect 51861 304256 51866 304312
rect 51922 304256 55068 304312
rect 51861 304254 55068 304256
rect 51861 304251 51927 304254
rect 16441 304176 19954 304178
rect 16441 304120 16446 304176
rect 16502 304120 19954 304176
rect 70678 304148 70738 304662
rect 73389 304659 73455 304662
rect 136869 304659 136935 304662
rect 137513 304659 137579 304662
rect 231997 304659 232063 304662
rect 325285 304659 325351 304662
rect 352750 304178 352810 304216
rect 356197 304178 356263 304181
rect 352750 304176 356263 304178
rect 16441 304118 19954 304120
rect 352750 304120 356202 304176
rect 356258 304120 356263 304176
rect 352750 304118 356263 304120
rect 424694 304178 424754 304216
rect 427405 304178 427471 304181
rect 424694 304176 427471 304178
rect 424694 304120 427410 304176
rect 427466 304120 427471 304176
rect 424694 304118 427471 304120
rect 16441 304115 16507 304118
rect 356197 304115 356263 304118
rect 427405 304115 427471 304118
rect 405969 303634 406035 303637
rect 405969 303632 409114 303634
rect 405969 303576 405974 303632
rect 406030 303576 409114 303632
rect 405969 303574 409114 303576
rect 405969 303571 406035 303574
rect 38613 303090 38679 303093
rect 35748 303088 38679 303090
rect 35748 303032 38618 303088
rect 38674 303032 38679 303088
rect 409054 303060 409114 303574
rect 35748 303030 38679 303032
rect 38613 303027 38679 303030
rect 136409 301594 136475 301597
rect 231997 301594 232063 301597
rect 324549 301594 324615 301597
rect 134740 301592 136475 301594
rect 134740 301536 136414 301592
rect 136470 301536 136475 301592
rect 134740 301534 136475 301536
rect 228764 301592 232063 301594
rect 228764 301536 232002 301592
rect 232058 301536 232063 301592
rect 228764 301534 232063 301536
rect 322788 301592 324615 301594
rect 322788 301536 324554 301592
rect 324610 301536 324615 301592
rect 322788 301534 324615 301536
rect 136409 301531 136475 301534
rect 231997 301531 232063 301534
rect 324549 301531 324615 301534
rect 55081 300916 55147 300917
rect 55030 300852 55036 300916
rect 55100 300914 55147 300916
rect 55100 300912 55192 300914
rect 55142 300856 55192 300912
rect 55100 300854 55192 300856
rect 55100 300852 55147 300854
rect 55081 300851 55147 300852
rect 38797 300642 38863 300645
rect 35748 300640 38863 300642
rect 35748 300584 38802 300640
rect 38858 300584 38863 300640
rect 35748 300582 38863 300584
rect 38797 300579 38863 300582
rect 50297 300642 50363 300645
rect 52638 300642 52644 300644
rect 50297 300640 52644 300642
rect 50297 300584 50302 300640
rect 50358 300584 52644 300640
rect 50297 300582 52644 300584
rect 50297 300579 50363 300582
rect 52638 300580 52644 300582
rect 52708 300580 52714 300644
rect 405969 300506 406035 300509
rect 408870 300506 408930 300612
rect 405969 300504 408930 300506
rect 70862 300098 70922 300476
rect 405969 300448 405974 300504
rect 406030 300448 408930 300504
rect 405969 300446 408930 300448
rect 405969 300443 406035 300446
rect 70862 300038 73498 300098
rect 73438 299962 73498 300038
rect 75413 299962 75479 299965
rect 73438 299960 75479 299962
rect 73438 299904 75418 299960
rect 75474 299904 75479 299960
rect 73438 299902 75479 299904
rect 75413 299899 75479 299902
rect 16349 298738 16415 298741
rect 19894 298738 19954 299388
rect 51677 299010 51743 299013
rect 55038 299010 55098 299320
rect 51677 299008 55098 299010
rect 51677 298952 51682 299008
rect 51738 298952 55098 299008
rect 51677 298950 55098 298952
rect 51677 298947 51743 298950
rect 352750 298874 352810 299320
rect 356197 298874 356263 298877
rect 352750 298872 356263 298874
rect 352750 298816 356202 298872
rect 356258 298816 356263 298872
rect 352750 298814 356263 298816
rect 356197 298811 356263 298814
rect 16349 298736 19954 298738
rect 16349 298680 16354 298736
rect 16410 298680 19954 298736
rect 16349 298678 19954 298680
rect 16349 298675 16415 298678
rect 74534 298676 74540 298740
rect 74604 298738 74610 298740
rect 75413 298738 75479 298741
rect 74604 298736 75479 298738
rect 74604 298680 75418 298736
rect 75474 298680 75479 298736
rect 74604 298678 75479 298680
rect 424694 298738 424754 299320
rect 427497 298738 427563 298741
rect 424694 298736 427563 298738
rect 424694 298680 427502 298736
rect 427558 298680 427563 298736
rect 424694 298678 427563 298680
rect 74604 298676 74610 298678
rect 75413 298675 75479 298678
rect 427497 298675 427563 298678
rect 137605 298602 137671 298605
rect 134710 298600 137671 298602
rect 134710 298544 137610 298600
rect 137666 298544 137671 298600
rect 134710 298542 137671 298544
rect 38245 298194 38311 298197
rect 134710 298196 134770 298542
rect 137605 298539 137671 298542
rect 230709 298466 230775 298469
rect 324641 298466 324707 298469
rect 325469 298466 325535 298469
rect 228764 298464 230775 298466
rect 228764 298408 230714 298464
rect 230770 298408 230775 298464
rect 228764 298406 230775 298408
rect 322788 298464 325535 298466
rect 322788 298408 324646 298464
rect 324702 298408 325474 298464
rect 325530 298408 325535 298464
rect 322788 298406 325535 298408
rect 230709 298403 230775 298406
rect 324641 298403 324707 298406
rect 325469 298403 325535 298406
rect 405969 298330 406035 298333
rect 405969 298328 409114 298330
rect 405969 298272 405974 298328
rect 406030 298272 409114 298328
rect 405969 298270 409114 298272
rect 405969 298267 406035 298270
rect 35748 298192 38311 298194
rect 35748 298136 38250 298192
rect 38306 298136 38311 298192
rect 35748 298134 38311 298136
rect 38245 298131 38311 298134
rect 134702 298132 134708 298196
rect 134772 298132 134778 298196
rect 409054 298164 409114 298270
rect 148326 296842 148908 296902
rect 242350 296842 242932 296902
rect 81669 296834 81735 296837
rect 145425 296834 145491 296837
rect 148326 296834 148386 296842
rect 81669 296832 85060 296834
rect 70862 296290 70922 296804
rect 81669 296776 81674 296832
rect 81730 296776 85060 296832
rect 81669 296774 85060 296776
rect 145425 296832 148386 296834
rect 145425 296776 145430 296832
rect 145486 296776 148386 296832
rect 145425 296774 148386 296776
rect 175509 296834 175575 296837
rect 240921 296834 240987 296837
rect 242350 296834 242410 296842
rect 175509 296832 178900 296834
rect 175509 296776 175514 296832
rect 175570 296776 178900 296832
rect 175509 296774 178900 296776
rect 240921 296832 242410 296834
rect 240921 296776 240926 296832
rect 240982 296776 242410 296832
rect 240921 296774 242410 296776
rect 269349 296834 269415 296837
rect 269349 296832 272924 296834
rect 269349 296776 269354 296832
rect 269410 296776 272924 296832
rect 269349 296774 272924 296776
rect 81669 296771 81735 296774
rect 145425 296771 145491 296774
rect 175509 296771 175575 296774
rect 240921 296771 240987 296774
rect 269349 296771 269415 296774
rect 74401 296290 74467 296293
rect 75965 296290 76031 296293
rect 70862 296288 76031 296290
rect 70862 296232 74406 296288
rect 74462 296232 75970 296288
rect 76026 296232 76031 296288
rect 70862 296230 76031 296232
rect 74401 296227 74467 296230
rect 75965 296227 76031 296230
rect 334209 296290 334275 296293
rect 336926 296290 336986 296872
rect 334209 296288 336986 296290
rect 334209 296232 334214 296288
rect 334270 296232 336986 296288
rect 334209 296230 336986 296232
rect 334209 296227 334275 296230
rect 35718 295474 35778 295512
rect 38797 295474 38863 295477
rect 35718 295472 38863 295474
rect 35718 295416 38802 295472
rect 38858 295416 38863 295472
rect 35718 295414 38863 295416
rect 38797 295411 38863 295414
rect 322750 295412 322756 295476
rect 322820 295412 322826 295476
rect 405969 295474 406035 295477
rect 408870 295474 408930 295580
rect 405969 295472 408930 295474
rect 405969 295416 405974 295472
rect 406030 295416 408930 295472
rect 405969 295414 408930 295416
rect 136910 295338 136916 295340
rect 134740 295278 136916 295338
rect 136910 295276 136916 295278
rect 136980 295276 136986 295340
rect 230750 295338 230756 295340
rect 228764 295278 230756 295338
rect 230750 295276 230756 295278
rect 230820 295276 230826 295340
rect 322758 295308 322818 295412
rect 405969 295411 406035 295414
rect 9896 294386 10376 294416
rect 13497 294386 13563 294389
rect 9896 294384 13563 294386
rect 9896 294328 13502 294384
rect 13558 294328 13563 294384
rect 9896 294326 13563 294328
rect 9896 294296 10376 294326
rect 13497 294323 13563 294326
rect 18005 293842 18071 293845
rect 19894 293842 19954 294356
rect 18005 293840 19954 293842
rect 18005 293784 18010 293840
rect 18066 293784 19954 293840
rect 18005 293782 19954 293784
rect 52597 293842 52663 293845
rect 55038 293842 55098 294288
rect 52597 293840 55098 293842
rect 52597 293784 52602 293840
rect 52658 293784 55098 293840
rect 52597 293782 55098 293784
rect 352750 293842 352810 294288
rect 356197 293842 356263 293845
rect 352750 293840 356263 293842
rect 352750 293784 356202 293840
rect 356258 293784 356263 293840
rect 352750 293782 356263 293784
rect 18005 293779 18071 293782
rect 52597 293779 52663 293782
rect 356197 293779 356263 293782
rect 405969 293706 406035 293709
rect 424694 293706 424754 294288
rect 427865 293706 427931 293709
rect 405969 293704 409114 293706
rect 405969 293648 405974 293704
rect 406030 293648 409114 293704
rect 405969 293646 409114 293648
rect 424694 293704 427931 293706
rect 424694 293648 427870 293704
rect 427926 293648 427931 293704
rect 424694 293646 427931 293648
rect 405969 293643 406035 293646
rect 74217 293570 74283 293573
rect 75873 293570 75939 293573
rect 70678 293568 75939 293570
rect 70678 293512 74222 293568
rect 74278 293512 75878 293568
rect 75934 293512 75939 293568
rect 70678 293510 75939 293512
rect 16165 293162 16231 293165
rect 18005 293162 18071 293165
rect 38429 293162 38495 293165
rect 16165 293160 18071 293162
rect 16165 293104 16170 293160
rect 16226 293104 18010 293160
rect 18066 293104 18071 293160
rect 16165 293102 18071 293104
rect 35748 293160 38495 293162
rect 35748 293104 38434 293160
rect 38490 293104 38495 293160
rect 70678 293132 70738 293510
rect 74217 293507 74283 293510
rect 75873 293507 75939 293510
rect 322750 293372 322756 293436
rect 322820 293434 322826 293436
rect 324825 293434 324891 293437
rect 325193 293434 325259 293437
rect 322820 293432 325259 293434
rect 322820 293376 324830 293432
rect 324886 293376 325198 293432
rect 325254 293376 325259 293432
rect 322820 293374 325259 293376
rect 322820 293372 322826 293374
rect 324825 293371 324891 293374
rect 325193 293371 325259 293374
rect 409054 293132 409114 293646
rect 427865 293643 427931 293646
rect 429889 293706 429955 293709
rect 434416 293706 434896 293736
rect 429889 293704 434896 293706
rect 429889 293648 429894 293704
rect 429950 293648 434896 293704
rect 429889 293646 434896 293648
rect 429889 293643 429955 293646
rect 434416 293616 434896 293646
rect 35748 293102 38495 293104
rect 16165 293099 16231 293102
rect 18005 293099 18071 293102
rect 38429 293099 38495 293102
rect 137830 292754 137836 292756
rect 134710 292694 137836 292754
rect 134710 292180 134770 292694
rect 137830 292692 137836 292694
rect 137900 292692 137906 292756
rect 322750 292284 322756 292348
rect 322820 292284 322826 292348
rect 229278 292210 229284 292212
rect 228764 292150 229284 292210
rect 229278 292148 229284 292150
rect 229348 292148 229354 292212
rect 322758 292180 322818 292284
rect 54897 292074 54963 292077
rect 55030 292074 55036 292076
rect 54897 292072 55036 292074
rect 54897 292016 54902 292072
rect 54958 292016 55036 292072
rect 54897 292014 55036 292016
rect 54897 292011 54963 292014
rect 55030 292012 55036 292014
rect 55100 292012 55106 292076
rect 165614 291876 165620 291940
rect 165684 291938 165690 291940
rect 178678 291938 178684 291940
rect 165684 291878 178684 291938
rect 165684 291876 165690 291878
rect 178678 291876 178684 291878
rect 178748 291876 178754 291940
rect 259454 291876 259460 291940
rect 259524 291938 259530 291940
rect 272702 291938 272708 291940
rect 259524 291878 272708 291938
rect 259524 291876 259530 291878
rect 272702 291876 272708 291878
rect 272772 291876 272778 291940
rect 74217 291668 74283 291669
rect 74166 291666 74172 291668
rect 74126 291606 74172 291666
rect 74236 291664 74283 291668
rect 74278 291608 74283 291664
rect 74166 291604 74172 291606
rect 74236 291604 74283 291608
rect 74217 291603 74283 291604
rect 229278 291332 229284 291396
rect 229348 291394 229354 291396
rect 231854 291394 231860 291396
rect 229348 291334 231860 291394
rect 229348 291332 229354 291334
rect 231854 291332 231860 291334
rect 231924 291332 231930 291396
rect 258718 291332 258724 291396
rect 258788 291394 258794 291396
rect 263686 291394 263692 291396
rect 258788 291334 263692 291394
rect 258788 291332 258794 291334
rect 263686 291332 263692 291334
rect 263756 291332 263762 291396
rect 405969 290714 406035 290717
rect 405969 290712 409114 290714
rect 405969 290656 405974 290712
rect 406030 290656 409114 290712
rect 405969 290654 409114 290656
rect 405969 290651 406035 290654
rect 38521 290578 38587 290581
rect 35748 290576 38587 290578
rect 35748 290520 38526 290576
rect 38582 290520 38587 290576
rect 409054 290548 409114 290654
rect 35748 290518 38587 290520
rect 38521 290515 38587 290518
rect 74033 290170 74099 290173
rect 70678 290168 74099 290170
rect 70678 290112 74038 290168
rect 74094 290112 74099 290168
rect 70678 290110 74099 290112
rect 70678 289596 70738 290110
rect 74033 290107 74099 290110
rect 228726 289564 228732 289628
rect 228796 289564 228802 289628
rect 322750 289564 322756 289628
rect 322820 289564 322826 289628
rect 137830 289354 137836 289356
rect 17453 289082 17519 289085
rect 19894 289082 19954 289324
rect 134710 289294 137836 289354
rect 54529 289286 54595 289289
rect 54529 289284 55068 289286
rect 54529 289228 54534 289284
rect 54590 289228 55068 289284
rect 54529 289226 55068 289228
rect 54529 289223 54595 289226
rect 54897 289082 54963 289085
rect 74401 289084 74467 289085
rect 17453 289080 19954 289082
rect 17453 289024 17458 289080
rect 17514 289024 19954 289080
rect 17453 289022 19954 289024
rect 54854 289080 54963 289082
rect 54854 289024 54902 289080
rect 54958 289048 54963 289080
rect 55030 289048 55036 289050
rect 54958 289024 55036 289048
rect 17453 289019 17519 289022
rect 54854 288988 55036 289024
rect 55030 288986 55036 288988
rect 55100 288986 55106 289050
rect 74350 289020 74356 289084
rect 74420 289082 74467 289084
rect 74420 289080 74512 289082
rect 74462 289024 74512 289080
rect 134710 289052 134770 289294
rect 137830 289292 137836 289294
rect 137900 289292 137906 289356
rect 228734 289082 228794 289564
rect 230709 289082 230775 289085
rect 228734 289080 230775 289082
rect 228734 289052 230714 289080
rect 74420 289022 74512 289024
rect 228764 289024 230714 289052
rect 230770 289024 230775 289080
rect 228764 289022 230775 289024
rect 74420 289020 74467 289022
rect 74401 289019 74467 289020
rect 230709 289019 230775 289022
rect 236045 289084 236111 289085
rect 236045 289080 236092 289084
rect 236156 289082 236162 289084
rect 236045 289024 236050 289080
rect 236045 289020 236092 289024
rect 236156 289022 236202 289082
rect 322758 289052 322818 289564
rect 352750 289082 352810 289256
rect 356197 289082 356263 289085
rect 352750 289080 356263 289082
rect 352750 289024 356202 289080
rect 356258 289024 356263 289080
rect 352750 289022 356263 289024
rect 424694 289082 424754 289256
rect 427589 289082 427655 289085
rect 424694 289080 427655 289082
rect 424694 289024 427594 289080
rect 427650 289024 427655 289080
rect 424694 289022 427655 289024
rect 236156 289020 236162 289022
rect 236045 289019 236111 289020
rect 356197 289019 356263 289022
rect 427589 289019 427655 289022
rect 74033 288946 74099 288949
rect 74166 288946 74172 288948
rect 74033 288944 74172 288946
rect 74033 288888 74038 288944
rect 74094 288888 74172 288944
rect 74033 288886 74172 288888
rect 74033 288883 74099 288886
rect 74166 288884 74172 288886
rect 74236 288884 74242 288948
rect 74309 288812 74375 288813
rect 74309 288810 74356 288812
rect 74264 288808 74356 288810
rect 74264 288752 74314 288808
rect 74264 288750 74356 288752
rect 74309 288748 74356 288750
rect 74420 288748 74426 288812
rect 74309 288747 74375 288748
rect 405969 288674 406035 288677
rect 405969 288672 409114 288674
rect 405969 288616 405974 288672
rect 406030 288616 409114 288672
rect 405969 288614 409114 288616
rect 405969 288611 406035 288614
rect 38521 288130 38587 288133
rect 35748 288128 38587 288130
rect 35748 288072 38526 288128
rect 38582 288072 38587 288128
rect 409054 288100 409114 288614
rect 35748 288070 38587 288072
rect 38521 288067 38587 288070
rect 51493 287586 51559 287589
rect 51677 287586 51743 287589
rect 51493 287584 51743 287586
rect 51493 287528 51498 287584
rect 51554 287528 51682 287584
rect 51738 287528 51743 287584
rect 51493 287526 51743 287528
rect 51493 287523 51559 287526
rect 51677 287523 51743 287526
rect 54478 287524 54484 287588
rect 54548 287586 54554 287588
rect 55030 287586 55036 287588
rect 54548 287526 55036 287586
rect 54548 287524 54554 287526
rect 55030 287524 55036 287526
rect 55100 287524 55106 287588
rect 164702 286362 164762 286808
rect 258726 286634 258786 286808
rect 261713 286634 261779 286637
rect 258726 286632 261779 286634
rect 258726 286576 261718 286632
rect 261774 286576 261779 286632
rect 258726 286574 261779 286576
rect 261713 286571 261779 286574
rect 168057 286362 168123 286365
rect 164702 286360 168123 286362
rect 164702 286304 168062 286360
rect 168118 286304 168123 286360
rect 164702 286302 168123 286304
rect 168057 286299 168123 286302
rect 325285 285954 325351 285957
rect 322788 285952 325351 285954
rect 35718 285546 35778 285584
rect 38521 285546 38587 285549
rect 35718 285544 38587 285546
rect 35718 285488 38526 285544
rect 38582 285488 38587 285544
rect 35718 285486 38587 285488
rect 38521 285483 38587 285486
rect 70678 285002 70738 285924
rect 322788 285896 325290 285952
rect 325346 285896 325351 285952
rect 322788 285894 325351 285896
rect 325285 285891 325351 285894
rect 134710 285274 134770 285856
rect 137605 285274 137671 285277
rect 134710 285272 137671 285274
rect 134710 285216 137610 285272
rect 137666 285216 137671 285272
rect 134710 285214 137671 285216
rect 228734 285274 228794 285856
rect 405969 285546 406035 285549
rect 408870 285546 408930 285652
rect 405969 285544 408930 285546
rect 405969 285488 405974 285544
rect 406030 285488 408930 285544
rect 405969 285486 408930 285488
rect 405969 285483 406035 285486
rect 231353 285274 231419 285277
rect 353713 285276 353779 285277
rect 228734 285272 231419 285274
rect 228734 285216 231358 285272
rect 231414 285216 231419 285272
rect 228734 285214 231419 285216
rect 137605 285211 137671 285214
rect 231353 285211 231419 285214
rect 353662 285212 353668 285276
rect 353732 285274 353779 285276
rect 353732 285272 353824 285274
rect 353774 285216 353824 285272
rect 353732 285214 353824 285216
rect 353732 285212 353779 285214
rect 353713 285211 353779 285212
rect 84613 285002 84679 285005
rect 70678 285000 84679 285002
rect 70678 284944 84618 285000
rect 84674 284944 84679 285000
rect 70678 284942 84679 284944
rect 84613 284939 84679 284942
rect 136869 284866 136935 284869
rect 138566 284866 138572 284868
rect 136869 284864 138572 284866
rect 136869 284808 136874 284864
rect 136930 284808 138572 284864
rect 136869 284806 138572 284808
rect 136869 284803 136935 284806
rect 138566 284804 138572 284806
rect 138636 284804 138642 284868
rect 84521 284596 84587 284597
rect 84470 284594 84476 284596
rect 84430 284534 84476 284594
rect 84540 284592 84587 284596
rect 84582 284536 84587 284592
rect 84470 284532 84476 284534
rect 84540 284532 84587 284536
rect 84521 284531 84587 284532
rect 17545 283778 17611 283781
rect 19894 283778 19954 284292
rect 52045 283914 52111 283917
rect 55038 283914 55098 284224
rect 52045 283912 55098 283914
rect 52045 283856 52050 283912
rect 52106 283856 55098 283912
rect 52045 283854 55098 283856
rect 52045 283851 52111 283854
rect 17545 283776 19954 283778
rect 17545 283720 17550 283776
rect 17606 283720 19954 283776
rect 17545 283718 19954 283720
rect 352750 283778 352810 284224
rect 356197 283778 356263 283781
rect 352750 283776 356263 283778
rect 352750 283720 356202 283776
rect 356258 283720 356263 283776
rect 352750 283718 356263 283720
rect 17545 283715 17611 283718
rect 356197 283715 356263 283718
rect 9896 283642 10376 283672
rect 13630 283642 13636 283644
rect 9896 283582 13636 283642
rect 9896 283552 10376 283582
rect 13630 283580 13636 283582
rect 13700 283580 13706 283644
rect 334209 283642 334275 283645
rect 424694 283642 424754 284224
rect 427957 283642 428023 283645
rect 334209 283640 336956 283642
rect 334209 283584 334214 283640
rect 334270 283584 336956 283640
rect 334209 283582 336956 283584
rect 424694 283640 428023 283642
rect 424694 283584 427962 283640
rect 428018 283584 428023 283640
rect 424694 283582 428023 283584
rect 334209 283579 334275 283582
rect 427957 283579 428023 283582
rect 148326 283514 148908 283574
rect 242350 283514 242932 283574
rect 145609 283506 145675 283509
rect 148326 283506 148386 283514
rect 145609 283504 148386 283506
rect 145609 283448 145614 283504
rect 145670 283448 148386 283504
rect 145609 283446 148386 283448
rect 240921 283506 240987 283509
rect 242350 283506 242410 283514
rect 240921 283504 242410 283506
rect 240921 283448 240926 283504
rect 240982 283448 242410 283504
rect 240921 283446 242410 283448
rect 145609 283443 145675 283446
rect 240921 283443 240987 283446
rect 405969 283370 406035 283373
rect 405969 283368 409114 283370
rect 405969 283312 405974 283368
rect 406030 283312 409114 283368
rect 405969 283310 409114 283312
rect 405969 283307 406035 283310
rect 38521 283098 38587 283101
rect 35748 283096 38587 283098
rect 35748 283040 38526 283096
rect 38582 283040 38587 283096
rect 409054 283068 409114 283310
rect 35748 283038 38587 283040
rect 38521 283035 38587 283038
rect 73614 282826 73620 282828
rect 70678 282766 73620 282826
rect 70678 282252 70738 282766
rect 73614 282764 73620 282766
rect 73684 282826 73690 282828
rect 84654 282826 84660 282828
rect 73684 282766 84660 282826
rect 73684 282764 73690 282766
rect 84654 282764 84660 282766
rect 84724 282764 84730 282828
rect 231629 282826 231695 282829
rect 324549 282826 324615 282829
rect 228764 282824 231695 282826
rect 228764 282768 231634 282824
rect 231690 282768 231695 282824
rect 228764 282766 231695 282768
rect 322788 282824 324615 282826
rect 322788 282768 324554 282824
rect 324610 282768 324615 282824
rect 322788 282766 324615 282768
rect 231629 282763 231695 282766
rect 324549 282763 324615 282766
rect 134710 282554 134770 282728
rect 136869 282554 136935 282557
rect 134710 282552 136935 282554
rect 134710 282496 136874 282552
rect 136930 282496 136935 282552
rect 134710 282494 136935 282496
rect 136869 282491 136935 282494
rect 136869 282282 136935 282285
rect 137278 282282 137284 282284
rect 136869 282280 137284 282282
rect 136869 282224 136874 282280
rect 136930 282224 137284 282280
rect 136869 282222 137284 282224
rect 136869 282219 136935 282222
rect 137278 282220 137284 282222
rect 137348 282220 137354 282284
rect 84613 281876 84679 281877
rect 84613 281874 84660 281876
rect 84568 281872 84660 281874
rect 84568 281816 84618 281872
rect 84568 281814 84660 281816
rect 84613 281812 84660 281814
rect 84724 281812 84730 281876
rect 84613 281811 84679 281812
rect 429429 281602 429495 281605
rect 434416 281602 434896 281632
rect 429429 281600 434896 281602
rect 429429 281544 429434 281600
rect 429490 281544 434896 281600
rect 429429 281542 434896 281544
rect 429429 281539 429495 281542
rect 434416 281512 434896 281542
rect 84521 281194 84587 281197
rect 84654 281194 84660 281196
rect 84521 281192 84660 281194
rect 84521 281136 84526 281192
rect 84582 281136 84660 281192
rect 84521 281134 84660 281136
rect 84521 281131 84587 281134
rect 84654 281132 84660 281134
rect 84724 281132 84730 281196
rect 35718 280378 35778 280552
rect 38061 280378 38127 280381
rect 35718 280376 38127 280378
rect 35718 280320 38066 280376
rect 38122 280320 38127 280376
rect 35718 280318 38127 280320
rect 38061 280315 38127 280318
rect 81669 280242 81735 280245
rect 175785 280242 175851 280245
rect 270269 280242 270335 280245
rect 81669 280240 85060 280242
rect 81669 280184 81674 280240
rect 81730 280184 85060 280240
rect 81669 280182 85060 280184
rect 175785 280240 178900 280242
rect 175785 280184 175790 280240
rect 175846 280184 178900 280240
rect 175785 280182 178900 280184
rect 270269 280240 272924 280242
rect 270269 280184 270274 280240
rect 270330 280184 272924 280240
rect 270269 280182 272924 280184
rect 81669 280179 81735 280182
rect 175785 280179 175851 280182
rect 270269 280179 270335 280182
rect 137697 279698 137763 279701
rect 231445 279698 231511 279701
rect 325377 279698 325443 279701
rect 134740 279696 137763 279698
rect 134740 279640 137702 279696
rect 137758 279640 137763 279696
rect 134740 279638 137763 279640
rect 228764 279696 231511 279698
rect 228764 279640 231450 279696
rect 231506 279640 231511 279696
rect 228764 279638 231511 279640
rect 322788 279696 325443 279698
rect 322788 279640 325382 279696
rect 325438 279640 325443 279696
rect 322788 279638 325443 279640
rect 137697 279635 137763 279638
rect 231445 279635 231511 279638
rect 325377 279635 325443 279638
rect 352742 279636 352748 279700
rect 352812 279698 352818 279700
rect 408870 279698 408930 280620
rect 352812 279638 408930 279698
rect 352812 279636 352818 279638
rect 18097 279562 18163 279565
rect 74033 279562 74099 279565
rect 74309 279562 74375 279565
rect 18097 279560 20138 279562
rect 18097 279504 18102 279560
rect 18158 279504 20138 279560
rect 18097 279502 20138 279504
rect 18097 279499 18163 279502
rect 20078 279396 20138 279502
rect 74033 279560 74234 279562
rect 74033 279504 74038 279560
rect 74094 279504 74234 279560
rect 74033 279502 74234 279504
rect 74033 279499 74099 279502
rect 52597 279426 52663 279429
rect 74174 279428 74234 279502
rect 74309 279560 74418 279562
rect 74309 279504 74314 279560
rect 74370 279504 74418 279560
rect 74309 279499 74418 279504
rect 74358 279428 74418 279499
rect 52597 279424 55068 279426
rect 52597 279368 52602 279424
rect 52658 279368 55068 279424
rect 52597 279366 55068 279368
rect 52597 279363 52663 279366
rect 74166 279364 74172 279428
rect 74236 279364 74242 279428
rect 74350 279364 74356 279428
rect 74420 279364 74426 279428
rect 356197 279426 356263 279429
rect 427681 279426 427747 279429
rect 352780 279424 356263 279426
rect 352780 279368 356202 279424
rect 356258 279368 356263 279424
rect 352780 279366 356263 279368
rect 424724 279424 427747 279426
rect 424724 279368 427686 279424
rect 427742 279368 427747 279424
rect 424724 279366 427747 279368
rect 356197 279363 356263 279366
rect 427681 279363 427747 279366
rect 54662 279228 54668 279292
rect 54732 279228 54738 279292
rect 54670 279020 54730 279228
rect 54662 278956 54668 279020
rect 54732 278956 54738 279020
rect 405969 278746 406035 278749
rect 405969 278744 409114 278746
rect 38613 278202 38679 278205
rect 35748 278200 38679 278202
rect 35748 278144 38618 278200
rect 38674 278144 38679 278200
rect 35748 278142 38679 278144
rect 70862 278202 70922 278716
rect 405969 278688 405974 278744
rect 406030 278688 409114 278744
rect 405969 278686 409114 278688
rect 405969 278683 406035 278686
rect 74033 278202 74099 278205
rect 138617 278204 138683 278205
rect 138566 278202 138572 278204
rect 70862 278200 74099 278202
rect 70862 278144 74038 278200
rect 74094 278144 74099 278200
rect 70862 278142 74099 278144
rect 138526 278142 138572 278202
rect 138636 278200 138683 278204
rect 138678 278144 138683 278200
rect 409054 278172 409114 278686
rect 38613 278139 38679 278142
rect 74033 278139 74099 278142
rect 138566 278140 138572 278142
rect 138636 278140 138683 278144
rect 138617 278139 138683 278140
rect 415118 277188 415124 277252
rect 415188 277250 415194 277252
rect 415261 277250 415327 277253
rect 415188 277248 415327 277250
rect 415188 277192 415266 277248
rect 415322 277192 415327 277248
rect 415188 277190 415327 277192
rect 415188 277188 415194 277190
rect 415261 277187 415327 277190
rect 137789 276570 137855 276573
rect 231537 276570 231603 276573
rect 325469 276570 325535 276573
rect 134740 276568 137855 276570
rect 134740 276512 137794 276568
rect 137850 276512 137855 276568
rect 134740 276510 137855 276512
rect 228764 276568 231603 276570
rect 228764 276512 231542 276568
rect 231598 276512 231603 276568
rect 228764 276510 231603 276512
rect 322788 276568 325535 276570
rect 322788 276512 325474 276568
rect 325530 276512 325535 276568
rect 322788 276510 325535 276512
rect 137789 276507 137855 276510
rect 231537 276507 231603 276510
rect 325469 276507 325535 276510
rect 159041 274666 159107 274669
rect 247913 274668 247979 274669
rect 167822 274666 167828 274668
rect 159041 274664 167828 274666
rect 159041 274608 159046 274664
rect 159102 274608 167828 274664
rect 159041 274606 167828 274608
rect 159041 274603 159107 274606
rect 167822 274604 167828 274606
rect 167892 274604 167898 274668
rect 247862 274666 247868 274668
rect 247822 274606 247868 274666
rect 247932 274664 247979 274668
rect 247974 274608 247979 274664
rect 247862 274604 247868 274606
rect 247932 274604 247979 274608
rect 247913 274603 247979 274604
rect 253341 274666 253407 274669
rect 261437 274666 261503 274669
rect 253341 274664 261503 274666
rect 253341 274608 253346 274664
rect 253402 274608 261442 274664
rect 261498 274608 261503 274664
rect 253341 274606 261503 274608
rect 253341 274603 253407 274606
rect 261437 274603 261503 274606
rect 149054 274468 149060 274532
rect 149124 274530 149130 274532
rect 157753 274530 157819 274533
rect 149124 274528 157819 274530
rect 149124 274472 157758 274528
rect 157814 274472 157819 274528
rect 149124 274470 157819 274472
rect 149124 274468 149130 274470
rect 157753 274467 157819 274470
rect 158397 274530 158463 274533
rect 168558 274530 168564 274532
rect 158397 274528 168564 274530
rect 158397 274472 158402 274528
rect 158458 274472 168564 274528
rect 158397 274470 168564 274472
rect 158397 274467 158463 274470
rect 168558 274468 168564 274470
rect 168628 274468 168634 274532
rect 252053 274530 252119 274533
rect 262398 274530 262404 274532
rect 252053 274528 262404 274530
rect 252053 274472 252058 274528
rect 252114 274472 262404 274528
rect 252053 274470 262404 274472
rect 252053 274467 252119 274470
rect 262398 274468 262404 274470
rect 262468 274468 262474 274532
rect 157201 274394 157267 274397
rect 169110 274394 169116 274396
rect 157201 274392 169116 274394
rect 157201 274336 157206 274392
rect 157262 274336 169116 274392
rect 157201 274334 169116 274336
rect 157201 274331 157267 274334
rect 169110 274332 169116 274334
rect 169180 274332 169186 274396
rect 232733 274394 232799 274397
rect 247862 274394 247868 274396
rect 232733 274392 247868 274394
rect 232733 274336 232738 274392
rect 232794 274336 247868 274392
rect 232733 274334 247868 274336
rect 232733 274331 232799 274334
rect 247862 274332 247868 274334
rect 247932 274332 247938 274396
rect 250857 274394 250923 274397
rect 262950 274394 262956 274396
rect 250857 274392 262956 274394
rect 250857 274336 250862 274392
rect 250918 274336 262956 274392
rect 250857 274334 262956 274336
rect 250857 274331 250923 274334
rect 262950 274332 262956 274334
rect 263020 274332 263026 274396
rect 136910 273788 136916 273852
rect 136980 273850 136986 273852
rect 137513 273850 137579 273853
rect 136980 273848 137579 273850
rect 136980 273792 137518 273848
rect 137574 273792 137579 273848
rect 136980 273790 137579 273792
rect 136980 273788 136986 273790
rect 137513 273787 137579 273790
rect 242342 273788 242348 273852
rect 242412 273850 242418 273852
rect 250949 273850 251015 273853
rect 242412 273848 251015 273850
rect 242412 273792 250954 273848
rect 251010 273792 251015 273848
rect 242412 273790 251015 273792
rect 242412 273788 242418 273790
rect 250949 273787 251015 273790
rect 414249 273850 414315 273853
rect 415537 273850 415603 273853
rect 414249 273848 415603 273850
rect 414249 273792 414254 273848
rect 414310 273792 415542 273848
rect 415598 273792 415603 273848
rect 414249 273790 415603 273792
rect 414249 273787 414315 273790
rect 415537 273787 415603 273790
rect 241974 273652 241980 273716
rect 242044 273714 242050 273716
rect 246206 273714 246212 273716
rect 242044 273654 246212 273714
rect 242044 273652 242050 273654
rect 246206 273652 246212 273654
rect 246276 273714 246282 273716
rect 247269 273714 247335 273717
rect 246276 273712 247335 273714
rect 246276 273656 247274 273712
rect 247330 273656 247335 273712
rect 246276 273654 247335 273656
rect 246276 273652 246282 273654
rect 247269 273651 247335 273654
rect 138065 273442 138131 273445
rect 231629 273442 231695 273445
rect 325193 273442 325259 273445
rect 134740 273440 138131 273442
rect 134740 273384 138070 273440
rect 138126 273384 138131 273440
rect 134740 273382 138131 273384
rect 228764 273440 231695 273442
rect 228764 273384 231634 273440
rect 231690 273384 231695 273440
rect 228764 273382 231695 273384
rect 322788 273440 325259 273442
rect 322788 273384 325198 273440
rect 325254 273384 325259 273440
rect 322788 273382 325259 273384
rect 138065 273379 138131 273382
rect 231629 273379 231695 273382
rect 325193 273379 325259 273382
rect 9896 272898 10376 272928
rect 13037 272898 13103 272901
rect 9896 272896 13103 272898
rect 9896 272840 13042 272896
rect 13098 272840 13103 272896
rect 9896 272838 13103 272840
rect 9896 272808 10376 272838
rect 13037 272835 13103 272838
rect 54478 272292 54484 272356
rect 54548 272354 54554 272356
rect 55030 272354 55036 272356
rect 54548 272294 55036 272354
rect 54548 272292 54554 272294
rect 55030 272292 55036 272294
rect 55100 272292 55106 272356
rect 261437 272218 261503 272221
rect 261846 272218 261852 272220
rect 261437 272216 261852 272218
rect 261437 272160 261442 272216
rect 261498 272160 261852 272216
rect 261437 272158 261852 272160
rect 261437 272155 261503 272158
rect 261846 272156 261852 272158
rect 261916 272156 261922 272220
rect 138617 269772 138683 269773
rect 138566 269708 138572 269772
rect 138636 269770 138683 269772
rect 395113 269770 395179 269773
rect 395389 269770 395455 269773
rect 138636 269768 138728 269770
rect 138678 269712 138728 269768
rect 138636 269710 138728 269712
rect 395113 269768 395455 269770
rect 395113 269712 395118 269768
rect 395174 269712 395394 269768
rect 395450 269712 395455 269768
rect 395113 269710 395455 269712
rect 138636 269708 138683 269710
rect 138617 269707 138683 269708
rect 395113 269707 395179 269710
rect 395389 269707 395455 269710
rect 276433 269498 276499 269501
rect 276750 269498 276756 269500
rect 276433 269496 276756 269498
rect 276433 269440 276438 269496
rect 276494 269440 276756 269496
rect 276433 269438 276756 269440
rect 276433 269435 276499 269438
rect 276750 269436 276756 269438
rect 276820 269436 276826 269500
rect 429429 269498 429495 269501
rect 434416 269498 434896 269528
rect 429429 269496 434896 269498
rect 429429 269440 429434 269496
rect 429490 269440 434896 269496
rect 429429 269438 434896 269440
rect 429429 269435 429495 269438
rect 434416 269408 434896 269438
rect 218013 268410 218079 268413
rect 219710 268410 219716 268412
rect 218013 268408 219716 268410
rect 218013 268352 218018 268408
rect 218074 268352 219716 268408
rect 218013 268350 219716 268352
rect 218013 268347 218079 268350
rect 219710 268348 219716 268350
rect 219780 268348 219786 268412
rect 261846 268212 261852 268276
rect 261916 268274 261922 268276
rect 262214 268274 262220 268276
rect 261916 268214 262220 268274
rect 261916 268212 261922 268214
rect 262214 268212 262220 268214
rect 262284 268212 262290 268276
rect 52638 266716 52644 266780
rect 52708 266778 52714 266780
rect 53517 266778 53583 266781
rect 52708 266776 53583 266778
rect 52708 266720 53522 266776
rect 53578 266720 53583 266776
rect 52708 266718 53583 266720
rect 52708 266716 52714 266718
rect 53517 266715 53583 266718
rect 54529 266778 54595 266781
rect 54662 266778 54668 266780
rect 54529 266776 54668 266778
rect 54529 266720 54534 266776
rect 54590 266720 54668 266776
rect 54529 266718 54668 266720
rect 54529 266715 54595 266718
rect 54662 266716 54668 266718
rect 54732 266716 54738 266780
rect 55030 266716 55036 266780
rect 55100 266778 55106 266780
rect 55541 266778 55607 266781
rect 55100 266776 55607 266778
rect 55100 266720 55546 266776
rect 55602 266720 55607 266776
rect 55100 266718 55607 266720
rect 55100 266716 55106 266718
rect 55541 266715 55607 266718
rect 55950 266716 55956 266780
rect 56020 266778 56026 266780
rect 56553 266778 56619 266781
rect 56020 266776 56619 266778
rect 56020 266720 56558 266776
rect 56614 266720 56619 266776
rect 56020 266718 56619 266720
rect 56020 266716 56026 266718
rect 56553 266715 56619 266718
rect 351822 266716 351828 266780
rect 351892 266778 351898 266780
rect 352057 266778 352123 266781
rect 351892 266776 352123 266778
rect 351892 266720 352062 266776
rect 352118 266720 352123 266776
rect 351892 266718 352123 266720
rect 351892 266716 351898 266718
rect 352057 266715 352123 266718
rect 350953 266642 351019 266645
rect 352006 266642 352012 266644
rect 350953 266640 352012 266642
rect 350953 266584 350958 266640
rect 351014 266584 352012 266640
rect 350953 266582 352012 266584
rect 350953 266579 351019 266582
rect 352006 266580 352012 266582
rect 352076 266580 352082 266644
rect 74350 266036 74356 266100
rect 74420 266098 74426 266100
rect 75270 266098 75276 266100
rect 74420 266038 75276 266098
rect 74420 266036 74426 266038
rect 75270 266036 75276 266038
rect 75340 266036 75346 266100
rect 73430 265900 73436 265964
rect 73500 265962 73506 265964
rect 74350 265962 74356 265964
rect 73500 265902 74356 265962
rect 73500 265900 73506 265902
rect 74350 265900 74356 265902
rect 74420 265900 74426 265964
rect 156189 263922 156255 263925
rect 152006 263920 156255 263922
rect 152006 263864 156194 263920
rect 156250 263864 156255 263920
rect 152006 263862 156255 263864
rect 142389 263650 142455 263653
rect 152006 263650 152066 263862
rect 156189 263859 156255 263862
rect 142389 263648 152066 263650
rect 142389 263592 142394 263648
rect 142450 263592 152066 263648
rect 142389 263590 152066 263592
rect 327309 263650 327375 263653
rect 327309 263648 331098 263650
rect 327309 263592 327314 263648
rect 327370 263592 331098 263648
rect 327309 263590 331098 263592
rect 142389 263587 142455 263590
rect 327309 263587 327375 263590
rect 73849 263514 73915 263517
rect 73982 263514 73988 263516
rect 73849 263512 73988 263514
rect 73849 263456 73854 263512
rect 73910 263456 73988 263512
rect 73849 263454 73988 263456
rect 73849 263451 73915 263454
rect 73982 263452 73988 263454
rect 74052 263514 74058 263516
rect 74350 263514 74356 263516
rect 74052 263454 74356 263514
rect 74052 263452 74058 263454
rect 74350 263452 74356 263454
rect 74420 263452 74426 263516
rect 74534 263452 74540 263516
rect 74604 263514 74610 263516
rect 75638 263514 75644 263516
rect 74604 263454 75644 263514
rect 74604 263452 74610 263454
rect 75638 263452 75644 263454
rect 75708 263452 75714 263516
rect 237190 263452 237196 263516
rect 237260 263514 237266 263516
rect 242342 263514 242348 263516
rect 237260 263454 242348 263514
rect 237260 263452 237266 263454
rect 242342 263452 242348 263454
rect 242412 263452 242418 263516
rect 144086 263316 144092 263380
rect 144156 263378 144162 263380
rect 149054 263378 149060 263380
rect 144156 263318 149060 263378
rect 144156 263316 144162 263318
rect 149054 263316 149060 263318
rect 149124 263316 149130 263380
rect 237558 263316 237564 263380
rect 237628 263378 237634 263380
rect 241974 263378 241980 263380
rect 237628 263318 241980 263378
rect 237628 263316 237634 263318
rect 241974 263316 241980 263318
rect 242044 263316 242050 263380
rect 77253 263174 77319 263177
rect 76780 263172 77319 263174
rect 76780 263116 77258 263172
rect 77314 263116 77319 263172
rect 331038 263144 331098 263590
rect 76780 263114 77319 263116
rect 77253 263111 77319 263114
rect 139813 263106 139879 263109
rect 173393 263106 173459 263109
rect 139813 263104 143020 263106
rect 139813 263048 139818 263104
rect 139874 263048 143020 263104
rect 139813 263046 143020 263048
rect 170804 263104 173459 263106
rect 170804 263048 173398 263104
rect 173454 263048 173459 263104
rect 170804 263046 173459 263048
rect 139813 263043 139879 263046
rect 173393 263043 173459 263046
rect 233469 263106 233535 263109
rect 267509 263106 267575 263109
rect 233469 263104 237044 263106
rect 233469 263048 233474 263104
rect 233530 263048 237044 263104
rect 233469 263046 237044 263048
rect 264828 263104 267575 263106
rect 264828 263048 267514 263104
rect 267570 263048 267575 263104
rect 264828 263046 267575 263048
rect 233469 263043 233535 263046
rect 267509 263043 267575 263046
rect 138566 262772 138572 262836
rect 138636 262772 138642 262836
rect 49193 262562 49259 262565
rect 49150 262560 49259 262562
rect 49150 262504 49198 262560
rect 49254 262504 49259 262560
rect 49150 262499 49259 262504
rect 138574 262562 138634 262772
rect 138750 262562 138756 262564
rect 138574 262502 138756 262562
rect 138750 262500 138756 262502
rect 138820 262500 138826 262564
rect 49150 262260 49210 262499
rect 360797 262290 360863 262293
rect 358852 262288 360863 262290
rect 358852 262232 360802 262288
rect 360858 262232 360863 262288
rect 358852 262230 360863 262232
rect 360797 262227 360863 262230
rect 9896 262018 10376 262048
rect 13589 262018 13655 262021
rect 9896 262016 13655 262018
rect 9896 261960 13594 262016
rect 13650 261960 13655 262016
rect 9896 261958 13655 261960
rect 9896 261928 10376 261958
rect 13589 261955 13655 261958
rect 79737 261746 79803 261749
rect 76780 261744 79803 261746
rect 76780 261688 79742 261744
rect 79798 261688 79803 261744
rect 76780 261686 79803 261688
rect 79737 261683 79803 261686
rect 140365 261746 140431 261749
rect 173485 261746 173551 261749
rect 140365 261744 143020 261746
rect 140365 261688 140370 261744
rect 140426 261688 143020 261744
rect 140365 261686 143020 261688
rect 170804 261744 173551 261746
rect 170804 261688 173490 261744
rect 173546 261688 173551 261744
rect 170804 261686 173551 261688
rect 140365 261683 140431 261686
rect 173485 261683 173551 261686
rect 233469 261746 233535 261749
rect 267417 261746 267483 261749
rect 233469 261744 237044 261746
rect 233469 261688 233474 261744
rect 233530 261688 237044 261744
rect 233469 261686 237044 261688
rect 264828 261744 267483 261746
rect 264828 261688 267422 261744
rect 267478 261688 267483 261744
rect 264828 261686 267483 261688
rect 233469 261683 233535 261686
rect 267417 261683 267483 261686
rect 327217 261746 327283 261749
rect 327217 261744 331068 261746
rect 327217 261688 327222 261744
rect 327278 261688 331068 261744
rect 327217 261686 331068 261688
rect 327217 261683 327283 261686
rect 79737 260386 79803 260389
rect 76780 260384 79803 260386
rect 76780 260328 79742 260384
rect 79798 260328 79803 260384
rect 76780 260326 79803 260328
rect 79737 260323 79803 260326
rect 140365 260386 140431 260389
rect 173761 260386 173827 260389
rect 140365 260384 143020 260386
rect 140365 260328 140370 260384
rect 140426 260328 143020 260384
rect 140365 260326 143020 260328
rect 170804 260384 173827 260386
rect 170804 260328 173766 260384
rect 173822 260328 173827 260384
rect 170804 260326 173827 260328
rect 140365 260323 140431 260326
rect 173761 260323 173827 260326
rect 233469 260386 233535 260389
rect 267601 260386 267667 260389
rect 233469 260384 237044 260386
rect 233469 260328 233474 260384
rect 233530 260328 237044 260384
rect 233469 260326 237044 260328
rect 264828 260384 267667 260386
rect 264828 260328 267606 260384
rect 267662 260328 267667 260384
rect 264828 260326 267667 260328
rect 233469 260323 233535 260326
rect 267601 260323 267667 260326
rect 326757 260386 326823 260389
rect 326757 260384 331068 260386
rect 326757 260328 326762 260384
rect 326818 260328 331068 260384
rect 326757 260326 331068 260328
rect 326757 260323 326823 260326
rect 138801 259980 138867 259981
rect 138750 259978 138756 259980
rect 138710 259918 138756 259978
rect 138820 259976 138867 259980
rect 138862 259920 138867 259976
rect 138750 259916 138756 259918
rect 138820 259916 138867 259920
rect 138801 259915 138867 259916
rect 46709 259162 46775 259165
rect 360521 259162 360587 259165
rect 46709 259160 48996 259162
rect 46709 259104 46714 259160
rect 46770 259104 48996 259160
rect 46709 259102 48996 259104
rect 358852 259160 360587 259162
rect 358852 259104 360526 259160
rect 360582 259104 360587 259160
rect 358852 259102 360587 259104
rect 46709 259099 46775 259102
rect 360521 259099 360587 259102
rect 79737 258890 79803 258893
rect 76780 258888 79803 258890
rect 76780 258832 79742 258888
rect 79798 258832 79803 258888
rect 76780 258830 79803 258832
rect 79737 258827 79803 258830
rect 140549 258890 140615 258893
rect 173853 258890 173919 258893
rect 140549 258888 143020 258890
rect 140549 258832 140554 258888
rect 140610 258832 143020 258888
rect 140549 258830 143020 258832
rect 170804 258888 173919 258890
rect 170804 258832 173858 258888
rect 173914 258832 173919 258888
rect 170804 258830 173919 258832
rect 140549 258827 140615 258830
rect 173853 258827 173919 258830
rect 233469 258890 233535 258893
rect 267325 258890 267391 258893
rect 233469 258888 237044 258890
rect 233469 258832 233474 258888
rect 233530 258832 237044 258888
rect 233469 258830 237044 258832
rect 264828 258888 267391 258890
rect 264828 258832 267330 258888
rect 267386 258832 267391 258888
rect 264828 258830 267391 258832
rect 233469 258827 233535 258830
rect 267325 258827 267391 258830
rect 328413 258890 328479 258893
rect 328413 258888 331068 258890
rect 328413 258832 328418 258888
rect 328474 258832 331068 258888
rect 328413 258830 331068 258832
rect 328413 258827 328479 258830
rect 87189 258074 87255 258077
rect 87189 258072 90058 258074
rect 87189 258016 87194 258072
rect 87250 258016 90058 258072
rect 87189 258014 90058 258016
rect 87189 258011 87255 258014
rect 80289 257530 80355 257533
rect 76780 257528 80355 257530
rect 76780 257472 80294 257528
rect 80350 257472 80355 257528
rect 76780 257470 80355 257472
rect 80289 257467 80355 257470
rect 89998 257432 90058 258014
rect 140549 257530 140615 257533
rect 173945 257530 174011 257533
rect 140549 257528 143020 257530
rect 140549 257472 140554 257528
rect 140610 257472 143020 257528
rect 140549 257470 143020 257472
rect 170804 257528 174011 257530
rect 170804 257472 173950 257528
rect 174006 257472 174011 257528
rect 170804 257470 174011 257472
rect 140549 257467 140615 257470
rect 173945 257467 174011 257470
rect 233469 257530 233535 257533
rect 267785 257530 267851 257533
rect 233469 257528 237044 257530
rect 233469 257472 233474 257528
rect 233530 257472 237044 257528
rect 233469 257470 237044 257472
rect 264828 257528 267851 257530
rect 264828 257472 267790 257528
rect 267846 257472 267851 257528
rect 264828 257470 267851 257472
rect 233469 257467 233535 257470
rect 267785 257467 267851 257470
rect 327217 257530 327283 257533
rect 327217 257528 331068 257530
rect 327217 257472 327222 257528
rect 327278 257472 331068 257528
rect 327217 257470 331068 257472
rect 327217 257467 327283 257470
rect 131349 257394 131415 257397
rect 129772 257392 131415 257394
rect 129772 257336 131354 257392
rect 131410 257336 131415 257392
rect 129772 257334 131415 257336
rect 131349 257331 131415 257334
rect 182317 257394 182383 257397
rect 226385 257394 226451 257397
rect 182317 257392 184052 257394
rect 182317 257336 182322 257392
rect 182378 257336 184052 257392
rect 182317 257334 184052 257336
rect 223796 257392 226451 257394
rect 223796 257336 226390 257392
rect 226446 257336 226451 257392
rect 223796 257334 226451 257336
rect 182317 257331 182383 257334
rect 226385 257331 226451 257334
rect 274869 257394 274935 257397
rect 321237 257394 321303 257397
rect 274869 257392 278076 257394
rect 274869 257336 274874 257392
rect 274930 257336 278076 257392
rect 274869 257334 278076 257336
rect 317820 257392 321303 257394
rect 317820 257336 321242 257392
rect 321298 257336 321303 257392
rect 317820 257334 321303 257336
rect 274869 257331 274935 257334
rect 321237 257331 321303 257334
rect 428785 257394 428851 257397
rect 434416 257394 434896 257424
rect 428785 257392 434896 257394
rect 428785 257336 428790 257392
rect 428846 257336 434896 257392
rect 428785 257334 434896 257336
rect 428785 257331 428851 257334
rect 434416 257304 434896 257334
rect 87189 256850 87255 256853
rect 87189 256848 90058 256850
rect 87189 256792 87194 256848
rect 87250 256792 90058 256848
rect 87189 256790 90058 256792
rect 87189 256787 87255 256790
rect 89998 256480 90058 256790
rect 132361 256442 132427 256445
rect 129772 256440 132427 256442
rect 129772 256384 132366 256440
rect 132422 256384 132427 256440
rect 129772 256382 132427 256384
rect 132361 256379 132427 256382
rect 182317 256442 182383 256445
rect 226293 256442 226359 256445
rect 182317 256440 184052 256442
rect 182317 256384 182322 256440
rect 182378 256384 184052 256440
rect 182317 256382 184052 256384
rect 223796 256440 226359 256442
rect 223796 256384 226298 256440
rect 226354 256384 226359 256440
rect 223796 256382 226359 256384
rect 182317 256379 182383 256382
rect 226293 256379 226359 256382
rect 275053 256442 275119 256445
rect 321053 256442 321119 256445
rect 275053 256440 278076 256442
rect 275053 256384 275058 256440
rect 275114 256384 278076 256440
rect 275053 256382 278076 256384
rect 317820 256440 321119 256442
rect 317820 256384 321058 256440
rect 321114 256384 321119 256440
rect 317820 256382 321119 256384
rect 275053 256379 275119 256382
rect 321053 256379 321119 256382
rect 79737 256170 79803 256173
rect 76780 256168 79803 256170
rect 76780 256112 79742 256168
rect 79798 256112 79803 256168
rect 76780 256110 79803 256112
rect 79737 256107 79803 256110
rect 140549 256170 140615 256173
rect 174037 256170 174103 256173
rect 140549 256168 143020 256170
rect 140549 256112 140554 256168
rect 140610 256112 143020 256168
rect 140549 256110 143020 256112
rect 170804 256168 174103 256170
rect 170804 256112 174042 256168
rect 174098 256112 174103 256168
rect 170804 256110 174103 256112
rect 140549 256107 140615 256110
rect 174037 256107 174103 256110
rect 233469 256170 233535 256173
rect 266589 256170 266655 256173
rect 233469 256168 237044 256170
rect 233469 256112 233474 256168
rect 233530 256112 237044 256168
rect 233469 256110 237044 256112
rect 264828 256168 266655 256170
rect 264828 256112 266594 256168
rect 266650 256112 266655 256168
rect 264828 256110 266655 256112
rect 233469 256107 233535 256110
rect 266589 256107 266655 256110
rect 328045 256170 328111 256173
rect 328045 256168 331068 256170
rect 328045 256112 328050 256168
rect 328106 256112 331068 256168
rect 328045 256110 331068 256112
rect 328045 256107 328111 256110
rect 46617 256034 46683 256037
rect 48590 256034 48596 256036
rect 46617 256032 48596 256034
rect 46617 255976 46622 256032
rect 46678 255976 48596 256032
rect 46617 255974 48596 255976
rect 46617 255971 46683 255974
rect 48590 255972 48596 255974
rect 48660 256034 48666 256036
rect 360613 256034 360679 256037
rect 48660 255974 48996 256034
rect 358668 256032 360679 256034
rect 358668 256004 360618 256032
rect 358638 255976 360618 256004
rect 360674 255976 360679 256032
rect 358638 255974 360679 255976
rect 48660 255972 48666 255974
rect 358638 255900 358698 255974
rect 360613 255971 360679 255974
rect 358630 255836 358636 255900
rect 358700 255836 358706 255900
rect 87281 255626 87347 255629
rect 131441 255626 131507 255629
rect 87281 255624 90028 255626
rect 87281 255568 87286 255624
rect 87342 255568 90028 255624
rect 87281 255566 90028 255568
rect 129772 255624 131507 255626
rect 129772 255568 131446 255624
rect 131502 255568 131507 255624
rect 129772 255566 131507 255568
rect 87281 255563 87347 255566
rect 131441 255563 131507 255566
rect 181581 255626 181647 255629
rect 225557 255626 225623 255629
rect 181581 255624 184052 255626
rect 181581 255568 181586 255624
rect 181642 255568 184052 255624
rect 181581 255566 184052 255568
rect 223796 255624 225623 255626
rect 223796 255568 225562 255624
rect 225618 255568 225623 255624
rect 223796 255566 225623 255568
rect 181581 255563 181647 255566
rect 225557 255563 225623 255566
rect 275881 255626 275947 255629
rect 320869 255626 320935 255629
rect 275881 255624 278076 255626
rect 275881 255568 275886 255624
rect 275942 255568 278076 255624
rect 275881 255566 278076 255568
rect 317820 255624 320935 255626
rect 317820 255568 320874 255624
rect 320930 255568 320935 255624
rect 317820 255566 320935 255568
rect 275881 255563 275947 255566
rect 320869 255563 320935 255566
rect 87189 255354 87255 255357
rect 87189 255352 90058 255354
rect 87189 255296 87194 255352
rect 87250 255296 90058 255352
rect 87189 255294 90058 255296
rect 87189 255291 87255 255294
rect 89998 254712 90058 255294
rect 79829 254674 79895 254677
rect 131349 254674 131415 254677
rect 76780 254672 79895 254674
rect 76780 254616 79834 254672
rect 79890 254616 79895 254672
rect 76780 254614 79895 254616
rect 129772 254672 131415 254674
rect 129772 254616 131354 254672
rect 131410 254616 131415 254672
rect 129772 254614 131415 254616
rect 79829 254611 79895 254614
rect 131349 254611 131415 254614
rect 140549 254674 140615 254677
rect 173761 254674 173827 254677
rect 140549 254672 143020 254674
rect 140549 254616 140554 254672
rect 140610 254616 143020 254672
rect 140549 254614 143020 254616
rect 170804 254672 173827 254674
rect 170804 254616 173766 254672
rect 173822 254616 173827 254672
rect 170804 254614 173827 254616
rect 140549 254611 140615 254614
rect 173761 254611 173827 254614
rect 182317 254674 182383 254677
rect 226293 254674 226359 254677
rect 182317 254672 184052 254674
rect 182317 254616 182322 254672
rect 182378 254616 184052 254672
rect 182317 254614 184052 254616
rect 223796 254672 226359 254674
rect 223796 254616 226298 254672
rect 226354 254616 226359 254672
rect 223796 254614 226359 254616
rect 182317 254611 182383 254614
rect 226293 254611 226359 254614
rect 232733 254674 232799 254677
rect 266589 254674 266655 254677
rect 232733 254672 237044 254674
rect 232733 254616 232738 254672
rect 232794 254616 237044 254672
rect 232733 254614 237044 254616
rect 264828 254672 266655 254674
rect 264828 254616 266594 254672
rect 266650 254616 266655 254672
rect 264828 254614 266655 254616
rect 232733 254611 232799 254614
rect 266589 254611 266655 254614
rect 274409 254674 274475 254677
rect 320685 254674 320751 254677
rect 274409 254672 278076 254674
rect 274409 254616 274414 254672
rect 274470 254616 278076 254672
rect 274409 254614 278076 254616
rect 317820 254672 320751 254674
rect 317820 254616 320690 254672
rect 320746 254616 320751 254672
rect 317820 254614 320751 254616
rect 274409 254611 274475 254614
rect 320685 254611 320751 254614
rect 328413 254674 328479 254677
rect 328413 254672 331068 254674
rect 328413 254616 328418 254672
rect 328474 254616 331068 254672
rect 328413 254614 331068 254616
rect 328413 254611 328479 254614
rect 87373 254402 87439 254405
rect 87373 254400 90058 254402
rect 87373 254344 87378 254400
rect 87434 254344 90058 254400
rect 87373 254342 90058 254344
rect 87373 254339 87439 254342
rect 89998 253896 90058 254342
rect 236638 254068 236644 254132
rect 236708 254130 236714 254132
rect 237190 254130 237196 254132
rect 236708 254070 237196 254130
rect 236708 254068 236714 254070
rect 237190 254068 237196 254070
rect 237260 254068 237266 254132
rect 131349 253858 131415 253861
rect 129772 253856 131415 253858
rect 129772 253800 131354 253856
rect 131410 253800 131415 253856
rect 129772 253798 131415 253800
rect 131349 253795 131415 253798
rect 181765 253858 181831 253861
rect 225373 253858 225439 253861
rect 181765 253856 184052 253858
rect 181765 253800 181770 253856
rect 181826 253800 184052 253856
rect 181765 253798 184052 253800
rect 223796 253856 225439 253858
rect 223796 253800 225378 253856
rect 225434 253800 225439 253856
rect 223796 253798 225439 253800
rect 181765 253795 181831 253798
rect 225373 253795 225439 253798
rect 274869 253858 274935 253861
rect 321605 253858 321671 253861
rect 274869 253856 278076 253858
rect 274869 253800 274874 253856
rect 274930 253800 278076 253856
rect 274869 253798 278076 253800
rect 317820 253856 321671 253858
rect 317820 253800 321610 253856
rect 321666 253800 321671 253856
rect 317820 253798 321671 253800
rect 274869 253795 274935 253798
rect 321605 253795 321671 253798
rect 79737 253314 79803 253317
rect 76780 253312 79803 253314
rect 76780 253256 79742 253312
rect 79798 253256 79803 253312
rect 76780 253254 79803 253256
rect 79737 253251 79803 253254
rect 140457 253314 140523 253317
rect 172933 253314 172999 253317
rect 140457 253312 143020 253314
rect 140457 253256 140462 253312
rect 140518 253256 143020 253312
rect 140457 253254 143020 253256
rect 170804 253312 172999 253314
rect 170804 253256 172938 253312
rect 172994 253256 172999 253312
rect 170804 253254 172999 253256
rect 140457 253251 140523 253254
rect 172933 253251 172999 253254
rect 234205 253314 234271 253317
rect 266589 253314 266655 253317
rect 234205 253312 237044 253314
rect 234205 253256 234210 253312
rect 234266 253256 237044 253312
rect 234205 253254 237044 253256
rect 264828 253312 266655 253314
rect 264828 253256 266594 253312
rect 266650 253256 266655 253312
rect 264828 253254 266655 253256
rect 234205 253251 234271 253254
rect 266589 253251 266655 253254
rect 327217 253314 327283 253317
rect 327217 253312 331068 253314
rect 327217 253256 327222 253312
rect 327278 253256 331068 253312
rect 327217 253254 331068 253256
rect 327217 253251 327283 253254
rect 46525 252906 46591 252909
rect 87189 252906 87255 252909
rect 131349 252906 131415 252909
rect 46525 252904 49180 252906
rect 46525 252848 46530 252904
rect 46586 252876 49180 252904
rect 87189 252904 90028 252906
rect 46586 252848 49210 252876
rect 46525 252846 49210 252848
rect 46525 252843 46591 252846
rect 49150 252364 49210 252846
rect 87189 252848 87194 252904
rect 87250 252848 90028 252904
rect 87189 252846 90028 252848
rect 129772 252904 131415 252906
rect 129772 252848 131354 252904
rect 131410 252848 131415 252904
rect 129772 252846 131415 252848
rect 87189 252843 87255 252846
rect 131349 252843 131415 252846
rect 181581 252906 181647 252909
rect 225741 252906 225807 252909
rect 181581 252904 184052 252906
rect 181581 252848 181586 252904
rect 181642 252848 184052 252904
rect 181581 252846 184052 252848
rect 223796 252904 225807 252906
rect 223796 252848 225746 252904
rect 225802 252848 225807 252904
rect 223796 252846 225807 252848
rect 181581 252843 181647 252846
rect 225741 252843 225807 252846
rect 274317 252906 274383 252909
rect 321605 252906 321671 252909
rect 360470 252906 360476 252908
rect 274317 252904 278076 252906
rect 274317 252848 274322 252904
rect 274378 252848 278076 252904
rect 274317 252846 278076 252848
rect 317820 252904 321671 252906
rect 317820 252848 321610 252904
rect 321666 252848 321671 252904
rect 317820 252846 321671 252848
rect 358852 252846 360476 252906
rect 274317 252843 274383 252846
rect 321605 252843 321671 252846
rect 360470 252844 360476 252846
rect 360540 252906 360546 252908
rect 361165 252906 361231 252909
rect 360540 252904 361231 252906
rect 360540 252848 361170 252904
rect 361226 252848 361231 252904
rect 360540 252846 361231 252848
rect 360540 252844 360546 252846
rect 361165 252843 361231 252846
rect 87281 252770 87347 252773
rect 87281 252768 90058 252770
rect 87281 252712 87286 252768
rect 87342 252712 90058 252768
rect 87281 252710 90058 252712
rect 87281 252707 87347 252710
rect 49142 252300 49148 252364
rect 49212 252300 49218 252364
rect 89998 252128 90058 252710
rect 133373 252090 133439 252093
rect 129772 252088 133439 252090
rect 129772 252032 133378 252088
rect 133434 252032 133439 252088
rect 129772 252030 133439 252032
rect 133373 252027 133439 252030
rect 181765 252090 181831 252093
rect 227213 252090 227279 252093
rect 181765 252088 184052 252090
rect 181765 252032 181770 252088
rect 181826 252032 184052 252088
rect 181765 252030 184052 252032
rect 223796 252088 227279 252090
rect 223796 252032 227218 252088
rect 227274 252032 227279 252088
rect 223796 252030 227279 252032
rect 181765 252027 181831 252030
rect 227213 252027 227279 252030
rect 275605 252090 275671 252093
rect 321605 252090 321671 252093
rect 275605 252088 278076 252090
rect 275605 252032 275610 252088
rect 275666 252032 278076 252088
rect 275605 252030 278076 252032
rect 317820 252088 321671 252090
rect 317820 252032 321610 252088
rect 321666 252032 321671 252088
rect 317820 252030 321671 252032
rect 275605 252027 275671 252030
rect 321605 252027 321671 252030
rect 79737 251954 79803 251957
rect 76780 251952 79803 251954
rect 76780 251896 79742 251952
rect 79798 251896 79803 251952
rect 76780 251894 79803 251896
rect 79737 251891 79803 251894
rect 140733 251954 140799 251957
rect 173669 251954 173735 251957
rect 140733 251952 143020 251954
rect 140733 251896 140738 251952
rect 140794 251896 143020 251952
rect 140733 251894 143020 251896
rect 170804 251952 173735 251954
rect 170804 251896 173674 251952
rect 173730 251896 173735 251952
rect 170804 251894 173735 251896
rect 140733 251891 140799 251894
rect 173669 251891 173735 251894
rect 232825 251954 232891 251957
rect 266589 251954 266655 251957
rect 232825 251952 237044 251954
rect 232825 251896 232830 251952
rect 232886 251896 237044 251952
rect 232825 251894 237044 251896
rect 264828 251952 266655 251954
rect 264828 251896 266594 251952
rect 266650 251896 266655 251952
rect 264828 251894 266655 251896
rect 232825 251891 232891 251894
rect 266589 251891 266655 251894
rect 327125 251954 327191 251957
rect 327125 251952 331068 251954
rect 327125 251896 327130 251952
rect 327186 251896 331068 251952
rect 327125 251894 331068 251896
rect 327125 251891 327191 251894
rect 87189 251682 87255 251685
rect 87189 251680 90058 251682
rect 87189 251624 87194 251680
rect 87250 251624 90058 251680
rect 87189 251622 90058 251624
rect 87189 251619 87255 251622
rect 9896 251274 10376 251304
rect 13129 251274 13195 251277
rect 9896 251272 13195 251274
rect 9896 251216 13134 251272
rect 13190 251216 13195 251272
rect 9896 251214 13195 251216
rect 9896 251184 10376 251214
rect 13129 251211 13195 251214
rect 89998 251176 90058 251622
rect 132177 251138 132243 251141
rect 129772 251136 132243 251138
rect 129772 251080 132182 251136
rect 132238 251080 132243 251136
rect 129772 251078 132243 251080
rect 132177 251075 132243 251078
rect 182317 251138 182383 251141
rect 226017 251138 226083 251141
rect 182317 251136 184052 251138
rect 182317 251080 182322 251136
rect 182378 251080 184052 251136
rect 182317 251078 184052 251080
rect 223796 251136 226083 251138
rect 223796 251080 226022 251136
rect 226078 251080 226083 251136
rect 223796 251078 226083 251080
rect 182317 251075 182383 251078
rect 226017 251075 226083 251078
rect 275513 251138 275579 251141
rect 320593 251138 320659 251141
rect 275513 251136 278076 251138
rect 275513 251080 275518 251136
rect 275574 251080 278076 251136
rect 275513 251078 278076 251080
rect 317820 251136 320659 251138
rect 317820 251080 320598 251136
rect 320654 251080 320659 251136
rect 317820 251078 320659 251080
rect 275513 251075 275579 251078
rect 320593 251075 320659 251078
rect 233469 251002 233535 251005
rect 233469 251000 237074 251002
rect 233469 250944 233474 251000
rect 233530 250944 237074 251000
rect 233469 250942 237074 250944
rect 233469 250939 233535 250942
rect 237014 250632 237074 250942
rect 79737 250594 79803 250597
rect 76780 250592 79803 250594
rect 76780 250536 79742 250592
rect 79798 250536 79803 250592
rect 76780 250534 79803 250536
rect 79737 250531 79803 250534
rect 140365 250594 140431 250597
rect 173117 250594 173183 250597
rect 267325 250594 267391 250597
rect 140365 250592 143020 250594
rect 140365 250536 140370 250592
rect 140426 250536 143020 250592
rect 140365 250534 143020 250536
rect 170804 250592 173183 250594
rect 170804 250536 173122 250592
rect 173178 250536 173183 250592
rect 170804 250534 173183 250536
rect 264828 250592 267391 250594
rect 264828 250536 267330 250592
rect 267386 250536 267391 250592
rect 264828 250534 267391 250536
rect 140365 250531 140431 250534
rect 173117 250531 173183 250534
rect 267325 250531 267391 250534
rect 327217 250594 327283 250597
rect 327217 250592 331068 250594
rect 327217 250536 327222 250592
rect 327278 250536 331068 250592
rect 327217 250534 331068 250536
rect 327217 250531 327283 250534
rect 138801 250458 138867 250461
rect 138934 250458 138940 250460
rect 138801 250456 138940 250458
rect 138801 250400 138806 250456
rect 138862 250400 138940 250456
rect 138801 250398 138940 250400
rect 138801 250395 138867 250398
rect 138934 250396 138940 250398
rect 139004 250396 139010 250460
rect 87189 250322 87255 250325
rect 131993 250322 132059 250325
rect 87189 250320 90028 250322
rect 87189 250264 87194 250320
rect 87250 250264 90028 250320
rect 87189 250262 90028 250264
rect 129772 250320 132059 250322
rect 129772 250264 131998 250320
rect 132054 250264 132059 250320
rect 129772 250262 132059 250264
rect 87189 250259 87255 250262
rect 131993 250259 132059 250262
rect 182225 250322 182291 250325
rect 225373 250322 225439 250325
rect 182225 250320 184052 250322
rect 182225 250264 182230 250320
rect 182286 250264 184052 250320
rect 182225 250262 184052 250264
rect 223796 250320 225439 250322
rect 223796 250264 225378 250320
rect 225434 250264 225439 250320
rect 223796 250262 225439 250264
rect 182225 250259 182291 250262
rect 225373 250259 225439 250262
rect 274133 250322 274199 250325
rect 321053 250322 321119 250325
rect 274133 250320 278076 250322
rect 274133 250264 274138 250320
rect 274194 250264 278076 250320
rect 274133 250262 278076 250264
rect 317820 250320 321119 250322
rect 317820 250264 321058 250320
rect 321114 250264 321119 250320
rect 317820 250262 321119 250264
rect 274133 250259 274199 250262
rect 321053 250259 321119 250262
rect 324733 250322 324799 250325
rect 325142 250322 325148 250324
rect 324733 250320 325148 250322
rect 324733 250264 324738 250320
rect 324794 250264 325148 250320
rect 324733 250262 325148 250264
rect 324733 250259 324799 250262
rect 325142 250260 325148 250262
rect 325212 250260 325218 250324
rect 132085 250050 132151 250053
rect 129742 250048 132151 250050
rect 129742 249992 132090 250048
rect 132146 249992 132151 250048
rect 129742 249990 132151 249992
rect 46433 249778 46499 249781
rect 46433 249776 49180 249778
rect 46433 249720 46438 249776
rect 46494 249748 49180 249776
rect 46494 249720 49210 249748
rect 46433 249718 49210 249720
rect 46433 249715 46499 249718
rect 49150 249236 49210 249718
rect 129742 249408 129802 249990
rect 132085 249987 132151 249990
rect 274869 250050 274935 250053
rect 274869 250048 278106 250050
rect 274869 249992 274874 250048
rect 274930 249992 278106 250048
rect 274869 249990 278106 249992
rect 274869 249987 274935 249990
rect 181489 249778 181555 249781
rect 233469 249778 233535 249781
rect 181489 249776 184082 249778
rect 181489 249720 181494 249776
rect 181550 249720 184082 249776
rect 181489 249718 184082 249720
rect 181489 249715 181555 249718
rect 140549 249642 140615 249645
rect 140549 249640 143050 249642
rect 140549 249584 140554 249640
rect 140610 249584 143050 249640
rect 140549 249582 143050 249584
rect 140549 249579 140615 249582
rect 87189 249370 87255 249373
rect 87189 249368 90028 249370
rect 87189 249312 87194 249368
rect 87250 249312 90028 249368
rect 87189 249310 90028 249312
rect 87189 249307 87255 249310
rect 49142 249172 49148 249236
rect 49212 249172 49218 249236
rect 77253 249166 77319 249169
rect 76780 249164 77319 249166
rect 76780 249108 77258 249164
rect 77314 249108 77319 249164
rect 142990 249136 143050 249582
rect 184022 249408 184082 249718
rect 233469 249776 237074 249778
rect 233469 249720 233474 249776
rect 233530 249720 237074 249776
rect 233469 249718 237074 249720
rect 233469 249715 233535 249718
rect 225925 249370 225991 249373
rect 223796 249368 225991 249370
rect 223796 249312 225930 249368
rect 225986 249312 225991 249368
rect 223796 249310 225991 249312
rect 225925 249307 225991 249310
rect 237014 249136 237074 249718
rect 278046 249408 278106 249990
rect 361441 249778 361507 249781
rect 358668 249776 361507 249778
rect 358668 249748 361446 249776
rect 358638 249720 361446 249748
rect 361502 249720 361507 249776
rect 358638 249718 361507 249720
rect 321605 249370 321671 249373
rect 317820 249368 321671 249370
rect 317820 249312 321610 249368
rect 321666 249312 321671 249368
rect 317820 249310 321671 249312
rect 321605 249307 321671 249310
rect 358638 249236 358698 249718
rect 361441 249715 361507 249718
rect 358630 249172 358636 249236
rect 358700 249172 358706 249236
rect 76780 249106 77319 249108
rect 77253 249103 77319 249106
rect 173301 249098 173367 249101
rect 267141 249098 267207 249101
rect 170804 249096 173367 249098
rect 170804 249040 173306 249096
rect 173362 249040 173367 249096
rect 170804 249038 173367 249040
rect 264828 249096 267207 249098
rect 264828 249040 267146 249096
rect 267202 249040 267207 249096
rect 264828 249038 267207 249040
rect 173301 249035 173367 249038
rect 267141 249035 267207 249038
rect 328413 249098 328479 249101
rect 328413 249096 331068 249098
rect 328413 249040 328418 249096
rect 328474 249040 331068 249096
rect 328413 249038 331068 249040
rect 328413 249035 328479 249038
rect 131809 248962 131875 248965
rect 129742 248960 131875 248962
rect 129742 248904 131814 248960
rect 131870 248904 131875 248960
rect 129742 248902 131875 248904
rect 129742 248456 129802 248902
rect 131809 248899 131875 248902
rect 274869 248826 274935 248829
rect 274869 248824 278106 248826
rect 274869 248768 274874 248824
rect 274930 248768 278106 248824
rect 274869 248766 278106 248768
rect 274869 248763 274935 248766
rect 181949 248690 182015 248693
rect 181949 248688 184082 248690
rect 181949 248632 181954 248688
rect 182010 248632 184082 248688
rect 181949 248630 184082 248632
rect 181949 248627 182015 248630
rect 184022 248456 184082 248630
rect 278046 248456 278106 248766
rect 87189 248418 87255 248421
rect 139537 248418 139603 248421
rect 225833 248418 225899 248421
rect 87189 248416 90028 248418
rect 87189 248360 87194 248416
rect 87250 248360 90028 248416
rect 87189 248358 90028 248360
rect 139537 248416 143050 248418
rect 139537 248360 139542 248416
rect 139598 248360 143050 248416
rect 139537 248358 143050 248360
rect 223796 248416 225899 248418
rect 223796 248360 225838 248416
rect 225894 248360 225899 248416
rect 223796 248358 225899 248360
rect 87189 248355 87255 248358
rect 139537 248355 139603 248358
rect 131717 248282 131783 248285
rect 129742 248280 131783 248282
rect 129742 248224 131722 248280
rect 131778 248224 131783 248280
rect 129742 248222 131783 248224
rect 77253 247806 77319 247809
rect 76780 247804 77319 247806
rect 76780 247748 77258 247804
rect 77314 247748 77319 247804
rect 76780 247746 77319 247748
rect 77253 247743 77319 247746
rect 129742 247640 129802 248222
rect 131717 248219 131783 248222
rect 142990 247776 143050 248358
rect 225833 248355 225899 248358
rect 233561 248418 233627 248421
rect 321605 248418 321671 248421
rect 233561 248416 237074 248418
rect 233561 248360 233566 248416
rect 233622 248360 237074 248416
rect 233561 248358 237074 248360
rect 317820 248416 321671 248418
rect 317820 248360 321610 248416
rect 321666 248360 321671 248416
rect 317820 248358 321671 248360
rect 233561 248355 233627 248358
rect 181857 248282 181923 248285
rect 181857 248280 184082 248282
rect 181857 248224 181862 248280
rect 181918 248224 184082 248280
rect 181857 248222 184082 248224
rect 181857 248219 181923 248222
rect 173301 247738 173367 247741
rect 170804 247736 173367 247738
rect 170804 247680 173306 247736
rect 173362 247680 173367 247736
rect 170804 247678 173367 247680
rect 173301 247675 173367 247678
rect 184022 247640 184082 248222
rect 237014 247776 237074 248358
rect 321605 248355 321671 248358
rect 274961 248282 275027 248285
rect 274961 248280 278106 248282
rect 274961 248224 274966 248280
rect 275022 248224 278106 248280
rect 274961 248222 278106 248224
rect 274961 248219 275027 248222
rect 266589 247738 266655 247741
rect 264828 247736 266655 247738
rect 264828 247680 266594 247736
rect 266650 247680 266655 247736
rect 264828 247678 266655 247680
rect 266589 247675 266655 247678
rect 278046 247640 278106 248222
rect 328413 247738 328479 247741
rect 328413 247736 331068 247738
rect 328413 247680 328418 247736
rect 328474 247680 331068 247736
rect 328413 247678 331068 247680
rect 328413 247675 328479 247678
rect 88477 247602 88543 247605
rect 225649 247602 225715 247605
rect 321789 247602 321855 247605
rect 88477 247600 90028 247602
rect 88477 247544 88482 247600
rect 88538 247544 90028 247600
rect 88477 247542 90028 247544
rect 223796 247600 225715 247602
rect 223796 247544 225654 247600
rect 225710 247544 225715 247600
rect 223796 247542 225715 247544
rect 317820 247600 321855 247602
rect 317820 247544 321794 247600
rect 321850 247544 321855 247600
rect 317820 247542 321855 247544
rect 88477 247539 88543 247542
rect 225649 247539 225715 247542
rect 321789 247539 321855 247542
rect 182317 247330 182383 247333
rect 274869 247330 274935 247333
rect 182317 247328 184082 247330
rect 182317 247272 182322 247328
rect 182378 247272 184082 247328
rect 182317 247270 184082 247272
rect 182317 247267 182383 247270
rect 132453 247058 132519 247061
rect 129742 247056 132519 247058
rect 129742 247000 132458 247056
rect 132514 247000 132519 247056
rect 129742 246998 132519 247000
rect 129742 246688 129802 246998
rect 132453 246995 132519 246998
rect 140641 246922 140707 246925
rect 140641 246920 143050 246922
rect 140641 246864 140646 246920
rect 140702 246864 143050 246920
rect 140641 246862 143050 246864
rect 140641 246859 140707 246862
rect 48406 246588 48412 246652
rect 48476 246650 48482 246652
rect 87189 246650 87255 246653
rect 48476 246590 48996 246650
rect 87189 246648 90028 246650
rect 87189 246592 87194 246648
rect 87250 246592 90028 246648
rect 87189 246590 90028 246592
rect 48476 246588 48482 246590
rect 87189 246587 87255 246590
rect 77253 246446 77319 246449
rect 76780 246444 77319 246446
rect 76780 246388 77258 246444
rect 77314 246388 77319 246444
rect 142990 246416 143050 246862
rect 184022 246688 184082 247270
rect 274869 247328 278106 247330
rect 274869 247272 274874 247328
rect 274930 247272 278106 247328
rect 274869 247270 278106 247272
rect 274869 247267 274935 247270
rect 234297 246922 234363 246925
rect 234297 246920 237074 246922
rect 234297 246864 234302 246920
rect 234358 246864 237074 246920
rect 234297 246862 237074 246864
rect 234297 246859 234363 246862
rect 226201 246650 226267 246653
rect 223796 246648 226267 246650
rect 223796 246592 226206 246648
rect 226262 246592 226267 246648
rect 223796 246590 226267 246592
rect 226201 246587 226267 246590
rect 237014 246416 237074 246862
rect 278046 246688 278106 247270
rect 328413 246922 328479 246925
rect 328413 246920 331098 246922
rect 328413 246864 328418 246920
rect 328474 246864 331098 246920
rect 328413 246862 331098 246864
rect 328413 246859 328479 246862
rect 321237 246650 321303 246653
rect 317820 246648 321303 246650
rect 317820 246592 321242 246648
rect 321298 246592 321303 246648
rect 317820 246590 321303 246592
rect 321237 246587 321303 246590
rect 331038 246416 331098 246862
rect 360705 246650 360771 246653
rect 358852 246648 360771 246650
rect 358852 246592 360710 246648
rect 360766 246592 360771 246648
rect 358852 246590 360771 246592
rect 360705 246587 360771 246590
rect 76780 246386 77319 246388
rect 77253 246383 77319 246386
rect 173669 246378 173735 246381
rect 266589 246378 266655 246381
rect 170804 246376 173735 246378
rect 170804 246320 173674 246376
rect 173730 246320 173735 246376
rect 170804 246318 173735 246320
rect 264828 246376 266655 246378
rect 264828 246320 266594 246376
rect 266650 246320 266655 246376
rect 264828 246318 266655 246320
rect 173669 246315 173735 246318
rect 266589 246315 266655 246318
rect 132269 246106 132335 246109
rect 129742 246104 132335 246106
rect 129742 246048 132274 246104
rect 132330 246048 132335 246104
rect 129742 246046 132335 246048
rect 129742 245872 129802 246046
rect 132269 246043 132335 246046
rect 181673 246106 181739 246109
rect 274869 246106 274935 246109
rect 181673 246104 184082 246106
rect 181673 246048 181678 246104
rect 181734 246048 184082 246104
rect 181673 246046 184082 246048
rect 181673 246043 181739 246046
rect 184022 245872 184082 246046
rect 274869 246104 278106 246106
rect 274869 246048 274874 246104
rect 274930 246048 278106 246104
rect 274869 246046 278106 246048
rect 274869 246043 274935 246046
rect 278046 245872 278106 246046
rect 87281 245834 87347 245837
rect 226109 245834 226175 245837
rect 321605 245834 321671 245837
rect 87281 245832 90028 245834
rect 87281 245776 87286 245832
rect 87342 245776 90028 245832
rect 87281 245774 90028 245776
rect 223796 245832 226175 245834
rect 223796 245776 226114 245832
rect 226170 245776 226175 245832
rect 223796 245774 226175 245776
rect 317820 245832 321671 245834
rect 317820 245776 321610 245832
rect 321666 245776 321671 245832
rect 317820 245774 321671 245776
rect 87281 245771 87347 245774
rect 226109 245771 226175 245774
rect 321605 245771 321671 245774
rect 78909 245562 78975 245565
rect 131349 245562 131415 245565
rect 76750 245560 78975 245562
rect 76750 245504 78914 245560
rect 78970 245504 78975 245560
rect 76750 245502 78975 245504
rect 76750 244920 76810 245502
rect 78909 245499 78975 245502
rect 129742 245560 131415 245562
rect 129742 245504 131354 245560
rect 131410 245504 131415 245560
rect 129742 245502 131415 245504
rect 129742 244920 129802 245502
rect 131349 245499 131415 245502
rect 140549 245562 140615 245565
rect 181581 245562 181647 245565
rect 234205 245562 234271 245565
rect 275697 245562 275763 245565
rect 327861 245562 327927 245565
rect 140549 245560 143050 245562
rect 140549 245504 140554 245560
rect 140610 245504 143050 245560
rect 140549 245502 143050 245504
rect 140549 245499 140615 245502
rect 142990 244920 143050 245502
rect 181581 245560 184082 245562
rect 181581 245504 181586 245560
rect 181642 245504 184082 245560
rect 181581 245502 184082 245504
rect 181581 245499 181647 245502
rect 184022 244920 184082 245502
rect 234205 245560 237074 245562
rect 234205 245504 234210 245560
rect 234266 245504 237074 245560
rect 234205 245502 237074 245504
rect 234205 245499 234271 245502
rect 237014 244920 237074 245502
rect 275697 245560 278106 245562
rect 275697 245504 275702 245560
rect 275758 245504 278106 245560
rect 275697 245502 278106 245504
rect 275697 245499 275763 245502
rect 278046 244920 278106 245502
rect 327861 245560 331098 245562
rect 327861 245504 327866 245560
rect 327922 245504 331098 245560
rect 327861 245502 331098 245504
rect 327861 245499 327927 245502
rect 331038 244920 331098 245502
rect 429429 245154 429495 245157
rect 434416 245154 434896 245184
rect 429429 245152 434896 245154
rect 429429 245096 429434 245152
rect 429490 245096 434896 245152
rect 429429 245094 434896 245096
rect 429429 245091 429495 245094
rect 434416 245064 434896 245094
rect 87189 244882 87255 244885
rect 173301 244882 173367 244885
rect 225373 244882 225439 244885
rect 266589 244882 266655 244885
rect 321697 244882 321763 244885
rect 87189 244880 90028 244882
rect 87189 244824 87194 244880
rect 87250 244824 90028 244880
rect 87189 244822 90028 244824
rect 170804 244880 173367 244882
rect 170804 244824 173306 244880
rect 173362 244824 173367 244880
rect 170804 244822 173367 244824
rect 223796 244880 225439 244882
rect 223796 244824 225378 244880
rect 225434 244824 225439 244880
rect 223796 244822 225439 244824
rect 264828 244880 266655 244882
rect 264828 244824 266594 244880
rect 266650 244824 266655 244880
rect 264828 244822 266655 244824
rect 317820 244880 321763 244882
rect 317820 244824 321702 244880
rect 321758 244824 321763 244880
rect 317820 244822 321763 244824
rect 87189 244819 87255 244822
rect 173301 244819 173367 244822
rect 225373 244819 225439 244822
rect 266589 244819 266655 244822
rect 321697 244819 321763 244822
rect 274869 244746 274935 244749
rect 274869 244744 278106 244746
rect 274869 244688 274874 244744
rect 274930 244688 278106 244744
rect 274869 244686 278106 244688
rect 274869 244683 274935 244686
rect 182041 244610 182107 244613
rect 182041 244608 184082 244610
rect 182041 244552 182046 244608
rect 182102 244552 184082 244608
rect 182041 244550 184082 244552
rect 182041 244547 182107 244550
rect 131349 244474 131415 244477
rect 129742 244472 131415 244474
rect 129742 244416 131354 244472
rect 131410 244416 131415 244472
rect 129742 244414 131415 244416
rect 78909 244202 78975 244205
rect 76750 244200 78975 244202
rect 76750 244144 78914 244200
rect 78970 244144 78975 244200
rect 76750 244142 78975 244144
rect 76750 243560 76810 244142
rect 78909 244139 78975 244142
rect 129742 244104 129802 244414
rect 131349 244411 131415 244414
rect 138893 244202 138959 244205
rect 138893 244200 143050 244202
rect 138893 244144 138898 244200
rect 138954 244144 143050 244200
rect 138893 244142 143050 244144
rect 138893 244139 138959 244142
rect 87373 244066 87439 244069
rect 87373 244064 90028 244066
rect 87373 244008 87378 244064
rect 87434 244008 90028 244064
rect 87373 244006 90028 244008
rect 87373 244003 87439 244006
rect 138934 243658 138940 243660
rect 138758 243598 138940 243658
rect 49150 243388 49210 243492
rect 138758 243388 138818 243598
rect 138934 243596 138940 243598
rect 139004 243596 139010 243660
rect 142990 243560 143050 244142
rect 184022 244104 184082 244550
rect 233561 244202 233627 244205
rect 233561 244200 237074 244202
rect 233561 244144 233566 244200
rect 233622 244144 237074 244200
rect 233561 244142 237074 244144
rect 233561 244139 233627 244142
rect 225557 244066 225623 244069
rect 223796 244064 225623 244066
rect 223796 244008 225562 244064
rect 225618 244008 225623 244064
rect 223796 244006 225623 244008
rect 225557 244003 225623 244006
rect 237014 243560 237074 244142
rect 278046 244104 278106 244686
rect 321605 244066 321671 244069
rect 317820 244064 321671 244066
rect 317820 244008 321610 244064
rect 321666 244008 321671 244064
rect 317820 244006 321671 244008
rect 321605 244003 321671 244006
rect 327861 244066 327927 244069
rect 327861 244064 331098 244066
rect 327861 244008 327866 244064
rect 327922 244008 331098 244064
rect 327861 244006 331098 244008
rect 327861 244003 327927 244006
rect 331038 243560 331098 244006
rect 173301 243522 173367 243525
rect 267877 243522 267943 243525
rect 360613 243522 360679 243525
rect 170804 243520 173367 243522
rect 170804 243464 173306 243520
rect 173362 243464 173367 243520
rect 170804 243462 173367 243464
rect 264828 243520 267943 243522
rect 264828 243464 267882 243520
rect 267938 243464 267943 243520
rect 264828 243462 267943 243464
rect 358852 243520 360679 243522
rect 358852 243464 360618 243520
rect 360674 243464 360679 243520
rect 358852 243462 360679 243464
rect 173301 243459 173367 243462
rect 267877 243459 267943 243462
rect 360613 243459 360679 243462
rect 49142 243324 49148 243388
rect 49212 243324 49218 243388
rect 138750 243324 138756 243388
rect 138820 243324 138826 243388
rect 181029 243386 181095 243389
rect 181029 243384 184082 243386
rect 181029 243328 181034 243384
rect 181090 243328 184082 243384
rect 181029 243326 184082 243328
rect 181029 243323 181095 243326
rect 184022 243152 184082 243326
rect 87281 243114 87347 243117
rect 132637 243114 132703 243117
rect 226293 243114 226359 243117
rect 87281 243112 90028 243114
rect 87281 243056 87286 243112
rect 87342 243056 90028 243112
rect 87281 243054 90028 243056
rect 129772 243112 132703 243114
rect 129772 243056 132642 243112
rect 132698 243056 132703 243112
rect 129772 243054 132703 243056
rect 223796 243112 226359 243114
rect 223796 243056 226298 243112
rect 226354 243056 226359 243112
rect 223796 243054 226359 243056
rect 87281 243051 87347 243054
rect 132637 243051 132703 243054
rect 226293 243051 226359 243054
rect 274225 243114 274291 243117
rect 321605 243114 321671 243117
rect 274225 243112 278076 243114
rect 274225 243056 274230 243112
rect 274286 243056 278076 243112
rect 274225 243054 278076 243056
rect 317820 243112 321671 243114
rect 317820 243056 321610 243112
rect 321666 243056 321671 243112
rect 317820 243054 321671 243056
rect 274225 243051 274291 243054
rect 321605 243051 321671 243054
rect 275789 242978 275855 242981
rect 275789 242976 278106 242978
rect 275789 242920 275794 242976
rect 275850 242920 278106 242976
rect 275789 242918 278106 242920
rect 275789 242915 275855 242918
rect 80197 242842 80263 242845
rect 76750 242840 80263 242842
rect 76750 242784 80202 242840
rect 80258 242784 80263 242840
rect 76750 242782 80263 242784
rect 76750 242200 76810 242782
rect 80197 242779 80263 242782
rect 140641 242842 140707 242845
rect 180293 242842 180359 242845
rect 234113 242842 234179 242845
rect 140641 242840 143050 242842
rect 140641 242784 140646 242840
rect 140702 242784 143050 242840
rect 140641 242782 143050 242784
rect 140641 242779 140707 242782
rect 131901 242706 131967 242709
rect 129742 242704 131967 242706
rect 129742 242648 131906 242704
rect 131962 242648 131967 242704
rect 129742 242646 131967 242648
rect 129742 242336 129802 242646
rect 131901 242643 131967 242646
rect 87189 242298 87255 242301
rect 87189 242296 90028 242298
rect 87189 242240 87194 242296
rect 87250 242240 90028 242296
rect 87189 242238 90028 242240
rect 87189 242235 87255 242238
rect 142990 242200 143050 242782
rect 180293 242840 184082 242842
rect 180293 242784 180298 242840
rect 180354 242784 184082 242840
rect 180293 242782 184082 242784
rect 180293 242779 180359 242782
rect 184022 242336 184082 242782
rect 234113 242840 237074 242842
rect 234113 242784 234118 242840
rect 234174 242784 237074 242840
rect 234113 242782 237074 242784
rect 234113 242779 234179 242782
rect 226385 242298 226451 242301
rect 223796 242296 226451 242298
rect 223796 242240 226390 242296
rect 226446 242240 226451 242296
rect 223796 242238 226451 242240
rect 226385 242235 226451 242238
rect 237014 242200 237074 242782
rect 278046 242336 278106 242918
rect 327861 242706 327927 242709
rect 327861 242704 331098 242706
rect 327861 242648 327866 242704
rect 327922 242648 331098 242704
rect 327861 242646 331098 242648
rect 327861 242643 327927 242646
rect 320501 242298 320567 242301
rect 317820 242296 320567 242298
rect 317820 242240 320506 242296
rect 320562 242240 320567 242296
rect 317820 242238 320567 242240
rect 320501 242235 320567 242238
rect 331038 242200 331098 242646
rect 172933 242162 172999 242165
rect 267877 242162 267943 242165
rect 170804 242160 172999 242162
rect 170804 242104 172938 242160
rect 172994 242104 172999 242160
rect 170804 242102 172999 242104
rect 264828 242160 267943 242162
rect 264828 242104 267882 242160
rect 267938 242104 267943 242160
rect 264828 242102 267943 242104
rect 172933 242099 172999 242102
rect 267877 242099 267943 242102
rect 96062 241692 96068 241756
rect 96132 241754 96138 241756
rect 98919 241754 98985 241757
rect 104894 241754 104900 241756
rect 96132 241752 104900 241754
rect 96132 241696 98924 241752
rect 98980 241696 104900 241752
rect 96132 241694 104900 241696
rect 96132 241692 96138 241694
rect 98919 241691 98985 241694
rect 104894 241692 104900 241694
rect 104964 241692 104970 241756
rect 76558 241012 76564 241076
rect 76628 241074 76634 241076
rect 93854 241074 93860 241076
rect 76628 241014 93860 241074
rect 76628 241012 76634 241014
rect 93854 241012 93860 241014
rect 93924 241012 93930 241076
rect 78909 240666 78975 240669
rect 76780 240664 78975 240666
rect 76780 240608 78914 240664
rect 78970 240608 78975 240664
rect 76780 240606 78975 240608
rect 78909 240603 78975 240606
rect 140549 240666 140615 240669
rect 173577 240666 173643 240669
rect 140549 240664 143020 240666
rect 140549 240608 140554 240664
rect 140610 240608 143020 240664
rect 140549 240606 143020 240608
rect 170804 240664 173643 240666
rect 170804 240608 173582 240664
rect 173638 240608 173643 240664
rect 170804 240606 173643 240608
rect 140549 240603 140615 240606
rect 173577 240603 173643 240606
rect 222429 240666 222495 240669
rect 222797 240666 222863 240669
rect 222429 240664 222863 240666
rect 222429 240608 222434 240664
rect 222490 240608 222802 240664
rect 222858 240608 222863 240664
rect 222429 240606 222863 240608
rect 222429 240603 222495 240606
rect 222797 240603 222863 240606
rect 233469 240666 233535 240669
rect 267877 240666 267943 240669
rect 233469 240664 237044 240666
rect 233469 240608 233474 240664
rect 233530 240608 237044 240664
rect 233469 240606 237044 240608
rect 264828 240664 267943 240666
rect 264828 240608 267882 240664
rect 267938 240608 267943 240664
rect 264828 240606 267943 240608
rect 233469 240603 233535 240606
rect 267877 240603 267943 240606
rect 327033 240666 327099 240669
rect 327033 240664 331068 240666
rect 327033 240608 327038 240664
rect 327094 240608 331068 240664
rect 327033 240606 331068 240608
rect 327033 240603 327099 240606
rect 9896 240530 10376 240560
rect 13313 240530 13379 240533
rect 9896 240528 13379 240530
rect 9896 240472 13318 240528
rect 13374 240472 13379 240528
rect 9896 240470 13379 240472
rect 9896 240440 10376 240470
rect 13313 240467 13379 240470
rect 49150 239852 49210 240364
rect 106550 240332 106556 240396
rect 106620 240394 106626 240396
rect 118694 240394 118700 240396
rect 106620 240334 118700 240394
rect 106620 240332 106626 240334
rect 118694 240332 118700 240334
rect 118764 240332 118770 240396
rect 303798 240332 303804 240396
rect 303868 240394 303874 240396
rect 305137 240394 305203 240397
rect 360797 240394 360863 240397
rect 303868 240392 305203 240394
rect 303868 240336 305142 240392
rect 305198 240336 305203 240392
rect 303868 240334 305203 240336
rect 358852 240392 360863 240394
rect 358852 240336 360802 240392
rect 360858 240336 360863 240392
rect 358852 240334 360863 240336
rect 303868 240332 303874 240334
rect 305137 240331 305203 240334
rect 360797 240331 360863 240334
rect 125870 240196 125876 240260
rect 125940 240258 125946 240260
rect 128630 240258 128636 240260
rect 125940 240198 128636 240258
rect 125940 240196 125946 240198
rect 128630 240196 128636 240198
rect 128700 240196 128706 240260
rect 49142 239788 49148 239852
rect 49212 239788 49218 239852
rect 95193 239716 95259 239717
rect 95142 239652 95148 239716
rect 95212 239714 95259 239716
rect 95212 239712 95304 239714
rect 95254 239656 95304 239712
rect 95212 239654 95304 239656
rect 95212 239652 95259 239654
rect 187878 239652 187884 239716
rect 187948 239714 187954 239716
rect 189217 239714 189283 239717
rect 187948 239712 189283 239714
rect 187948 239656 189222 239712
rect 189278 239656 189283 239712
rect 187948 239654 189283 239656
rect 187948 239652 187954 239654
rect 95193 239651 95259 239652
rect 189217 239651 189283 239654
rect 211021 239714 211087 239717
rect 290509 239716 290575 239717
rect 211246 239714 211252 239716
rect 211021 239712 211252 239714
rect 211021 239656 211026 239712
rect 211082 239656 211252 239712
rect 211021 239654 211252 239656
rect 211021 239651 211087 239654
rect 211246 239652 211252 239654
rect 211316 239652 211322 239716
rect 290509 239714 290556 239716
rect 290464 239712 290556 239714
rect 290464 239656 290514 239712
rect 290464 239654 290556 239656
rect 290509 239652 290556 239654
rect 290620 239652 290626 239716
rect 290509 239651 290575 239652
rect 91697 239442 91763 239445
rect 92566 239442 92572 239444
rect 91697 239440 92572 239442
rect 91697 239384 91702 239440
rect 91758 239384 92572 239440
rect 91697 239382 92572 239384
rect 91697 239379 91763 239382
rect 92566 239380 92572 239382
rect 92636 239380 92642 239444
rect 283241 239442 283307 239445
rect 284294 239442 284300 239444
rect 283241 239440 284300 239442
rect 283241 239384 283246 239440
rect 283302 239384 284300 239440
rect 283241 239382 284300 239384
rect 283241 239379 283307 239382
rect 284294 239380 284300 239382
rect 284364 239380 284370 239444
rect 79001 239306 79067 239309
rect 76780 239304 79067 239306
rect 76780 239248 79006 239304
rect 79062 239248 79067 239304
rect 76780 239246 79067 239248
rect 79001 239243 79067 239246
rect 140549 239306 140615 239309
rect 173853 239306 173919 239309
rect 140549 239304 143020 239306
rect 140549 239248 140554 239304
rect 140610 239248 143020 239304
rect 140549 239246 143020 239248
rect 170804 239304 173919 239306
rect 170804 239248 173858 239304
rect 173914 239248 173919 239304
rect 170804 239246 173919 239248
rect 140549 239243 140615 239246
rect 173853 239243 173919 239246
rect 233469 239306 233535 239309
rect 267877 239306 267943 239309
rect 233469 239304 237044 239306
rect 233469 239248 233474 239304
rect 233530 239248 237044 239304
rect 233469 239246 237044 239248
rect 264828 239304 267943 239306
rect 264828 239248 267882 239304
rect 267938 239248 267943 239304
rect 264828 239246 267943 239248
rect 233469 239243 233535 239246
rect 267877 239243 267943 239246
rect 327217 239306 327283 239309
rect 327217 239304 331068 239306
rect 327217 239248 327222 239304
rect 327278 239248 331068 239304
rect 327217 239246 331068 239248
rect 327217 239243 327283 239246
rect 230985 239036 231051 239037
rect 230934 238972 230940 239036
rect 231004 239034 231051 239036
rect 325193 239034 325259 239037
rect 325326 239034 325332 239036
rect 231004 239032 231096 239034
rect 231046 238976 231096 239032
rect 231004 238974 231096 238976
rect 325193 239032 325332 239034
rect 325193 238976 325198 239032
rect 325254 238976 325332 239032
rect 325193 238974 325332 238976
rect 231004 238972 231051 238974
rect 230985 238971 231051 238972
rect 325193 238971 325259 238974
rect 325326 238972 325332 238974
rect 325396 238972 325402 239036
rect 79093 238626 79159 238629
rect 76750 238624 79159 238626
rect 76750 238568 79098 238624
rect 79154 238568 79159 238624
rect 76750 238566 79159 238568
rect 76750 237984 76810 238566
rect 79093 238563 79159 238566
rect 102318 238564 102324 238628
rect 102388 238626 102394 238628
rect 102553 238626 102619 238629
rect 136961 238626 137027 238629
rect 102388 238624 137027 238626
rect 102388 238568 102558 238624
rect 102614 238568 136966 238624
rect 137022 238568 137027 238624
rect 102388 238566 137027 238568
rect 102388 238564 102394 238566
rect 102553 238563 102619 238566
rect 136961 238563 137027 238566
rect 233561 238626 233627 238629
rect 327125 238626 327191 238629
rect 233561 238624 237074 238626
rect 233561 238568 233566 238624
rect 233622 238568 237074 238624
rect 233561 238566 237074 238568
rect 233561 238563 233627 238566
rect 140181 238490 140247 238493
rect 140181 238488 143050 238490
rect 140181 238432 140186 238488
rect 140242 238432 143050 238488
rect 140181 238430 143050 238432
rect 140181 238427 140247 238430
rect 142757 238356 142823 238357
rect 142757 238354 142804 238356
rect 142712 238352 142804 238354
rect 142712 238296 142762 238352
rect 142712 238294 142804 238296
rect 142757 238292 142804 238294
rect 142868 238292 142874 238356
rect 142757 238291 142823 238292
rect 142990 237984 143050 238430
rect 200022 238292 200028 238356
rect 200092 238354 200098 238356
rect 200165 238354 200231 238357
rect 200092 238352 200231 238354
rect 200092 238296 200170 238352
rect 200226 238296 200231 238352
rect 200092 238294 200231 238296
rect 200092 238292 200098 238294
rect 200165 238291 200231 238294
rect 230893 238354 230959 238357
rect 231854 238354 231860 238356
rect 230893 238352 231860 238354
rect 230893 238296 230898 238352
rect 230954 238296 231860 238352
rect 230893 238294 231860 238296
rect 230893 238291 230959 238294
rect 231854 238292 231860 238294
rect 231924 238292 231930 238356
rect 237014 237984 237074 238566
rect 327125 238624 331098 238626
rect 327125 238568 327130 238624
rect 327186 238568 331098 238624
rect 327125 238566 331098 238568
rect 327125 238563 327191 238566
rect 286921 238356 286987 238357
rect 286870 238292 286876 238356
rect 286940 238354 286987 238356
rect 286940 238352 287032 238354
rect 286982 238296 287032 238352
rect 286940 238294 287032 238296
rect 286940 238292 286987 238294
rect 286921 238291 286987 238292
rect 331038 237984 331098 238566
rect 174037 237946 174103 237949
rect 267509 237946 267575 237949
rect 170804 237944 174103 237946
rect 170804 237888 174042 237944
rect 174098 237888 174103 237944
rect 170804 237886 174103 237888
rect 264828 237944 267575 237946
rect 264828 237888 267514 237944
rect 267570 237888 267575 237944
rect 264828 237886 267575 237888
rect 174037 237883 174103 237886
rect 267509 237883 267575 237886
rect 219761 237812 219827 237813
rect 219710 237810 219716 237812
rect 219670 237750 219716 237810
rect 219780 237808 219827 237812
rect 219822 237752 219827 237808
rect 219710 237748 219716 237750
rect 219780 237748 219827 237752
rect 219761 237747 219827 237748
rect 47077 237402 47143 237405
rect 361165 237402 361231 237405
rect 47077 237400 48996 237402
rect 47077 237344 47082 237400
rect 47138 237344 48996 237400
rect 47077 237342 48996 237344
rect 358852 237400 361231 237402
rect 358852 237344 361170 237400
rect 361226 237344 361231 237400
rect 358852 237342 361231 237344
rect 47077 237339 47143 237342
rect 361165 237339 361231 237342
rect 140273 237266 140339 237269
rect 140273 237264 143050 237266
rect 140273 237208 140278 237264
rect 140334 237208 143050 237264
rect 140273 237206 143050 237208
rect 140273 237203 140339 237206
rect 142990 236624 143050 237206
rect 233469 237130 233535 237133
rect 233469 237128 237074 237130
rect 233469 237072 233474 237128
rect 233530 237072 237074 237128
rect 233469 237070 237074 237072
rect 233469 237067 233535 237070
rect 183830 236932 183836 236996
rect 183900 236994 183906 236996
rect 192897 236994 192963 236997
rect 183900 236992 192963 236994
rect 183900 236936 192902 236992
rect 192958 236936 192963 236992
rect 183900 236934 192963 236936
rect 183900 236932 183906 236934
rect 192897 236931 192963 236934
rect 237014 236624 237074 237070
rect 78909 236586 78975 236589
rect 172933 236586 172999 236589
rect 267233 236586 267299 236589
rect 76780 236584 78975 236586
rect 76780 236528 78914 236584
rect 78970 236528 78975 236584
rect 76780 236526 78975 236528
rect 170804 236584 172999 236586
rect 170804 236528 172938 236584
rect 172994 236528 172999 236584
rect 170804 236526 172999 236528
rect 264828 236584 267299 236586
rect 264828 236528 267238 236584
rect 267294 236528 267299 236584
rect 264828 236526 267299 236528
rect 78909 236523 78975 236526
rect 172933 236523 172999 236526
rect 267233 236523 267299 236526
rect 328413 236586 328479 236589
rect 369169 236586 369235 236589
rect 328413 236584 331068 236586
rect 328413 236528 328418 236584
rect 328474 236528 331068 236584
rect 328413 236526 331068 236528
rect 369169 236584 371916 236586
rect 369169 236528 369174 236584
rect 369230 236528 371916 236584
rect 369169 236526 371916 236528
rect 328413 236523 328479 236526
rect 369169 236523 369235 236526
rect 73982 236388 73988 236452
rect 74052 236450 74058 236452
rect 74166 236450 74172 236452
rect 74052 236390 74172 236450
rect 74052 236388 74058 236390
rect 74166 236388 74172 236390
rect 74236 236388 74242 236452
rect 74166 236252 74172 236316
rect 74236 236314 74242 236316
rect 75822 236314 75828 236316
rect 74236 236254 75828 236314
rect 74236 236252 74242 236254
rect 75822 236252 75828 236254
rect 75892 236252 75898 236316
rect 149238 236314 149244 236316
rect 147774 236254 149244 236314
rect 147449 236178 147515 236181
rect 147774 236178 147834 236254
rect 149238 236252 149244 236254
rect 149308 236252 149314 236316
rect 153470 236252 153476 236316
rect 153540 236314 153546 236316
rect 162854 236314 162860 236316
rect 153540 236254 162860 236314
rect 153540 236252 153546 236254
rect 162854 236252 162860 236254
rect 162924 236252 162930 236316
rect 147449 236176 147834 236178
rect 147449 236120 147454 236176
rect 147510 236120 147834 236176
rect 147449 236118 147834 236120
rect 148369 236178 148435 236181
rect 149606 236178 149612 236180
rect 148369 236176 149612 236178
rect 148369 236120 148374 236176
rect 148430 236120 149612 236176
rect 148369 236118 149612 236120
rect 147449 236115 147515 236118
rect 148369 236115 148435 236118
rect 149606 236116 149612 236118
rect 149676 236116 149682 236180
rect 238110 236116 238116 236180
rect 238180 236178 238186 236180
rect 243773 236178 243839 236181
rect 238180 236176 243839 236178
rect 238180 236120 243778 236176
rect 243834 236120 243839 236176
rect 238180 236118 243839 236120
rect 238180 236116 238186 236118
rect 243773 236115 243839 236118
rect 247269 236178 247335 236181
rect 248782 236178 248788 236180
rect 247269 236176 248788 236178
rect 247269 236120 247274 236176
rect 247330 236120 248788 236176
rect 247269 236118 248788 236120
rect 247269 236115 247335 236118
rect 248782 236116 248788 236118
rect 248852 236116 248858 236180
rect 369445 236178 369511 236181
rect 369445 236176 371916 236178
rect 369445 236120 369450 236176
rect 369506 236120 371916 236176
rect 369445 236118 371916 236120
rect 369445 236115 369511 236118
rect 148645 236044 148711 236045
rect 148645 236040 148692 236044
rect 148756 236042 148762 236044
rect 148645 235984 148650 236040
rect 148645 235980 148692 235984
rect 148756 235982 148802 236042
rect 148756 235980 148762 235982
rect 148645 235979 148711 235980
rect 147950 235844 147956 235908
rect 148020 235906 148026 235908
rect 148737 235906 148803 235909
rect 148020 235904 148803 235906
rect 148020 235848 148742 235904
rect 148798 235848 148803 235904
rect 148020 235846 148803 235848
rect 148020 235844 148026 235846
rect 148737 235843 148803 235846
rect 242485 235906 242551 235909
rect 262030 235906 262036 235908
rect 242485 235904 262036 235906
rect 242485 235848 242490 235904
rect 242546 235848 262036 235904
rect 242485 235846 262036 235848
rect 242485 235843 242551 235846
rect 262030 235844 262036 235846
rect 262100 235844 262106 235908
rect 109821 235770 109887 235773
rect 110414 235770 110420 235772
rect 109821 235768 110420 235770
rect 109821 235712 109826 235768
rect 109882 235712 110420 235768
rect 109821 235710 110420 235712
rect 109821 235707 109887 235710
rect 110414 235708 110420 235710
rect 110484 235770 110490 235772
rect 136961 235770 137027 235773
rect 110484 235768 137027 235770
rect 110484 235712 136966 235768
rect 137022 235712 137027 235768
rect 110484 235710 137027 235712
rect 110484 235708 110490 235710
rect 136961 235707 137027 235710
rect 262398 235708 262404 235772
rect 262468 235770 262474 235772
rect 262541 235770 262607 235773
rect 262468 235768 262607 235770
rect 262468 235712 262546 235768
rect 262602 235712 262607 235768
rect 262468 235710 262607 235712
rect 262468 235708 262474 235710
rect 262541 235707 262607 235710
rect 369629 235770 369695 235773
rect 369629 235768 371916 235770
rect 369629 235712 369634 235768
rect 369690 235712 371916 235768
rect 369629 235710 371916 235712
rect 369629 235707 369695 235710
rect 74677 235636 74743 235637
rect 74677 235634 74724 235636
rect 74596 235632 74724 235634
rect 74788 235634 74794 235636
rect 75822 235634 75828 235636
rect 74596 235576 74682 235632
rect 74596 235574 74724 235576
rect 74677 235572 74724 235574
rect 74788 235574 75828 235634
rect 74788 235572 74794 235574
rect 75822 235572 75828 235574
rect 75892 235572 75898 235636
rect 74677 235571 74743 235572
rect 369813 235362 369879 235365
rect 369813 235360 371916 235362
rect 369813 235304 369818 235360
rect 369874 235304 371916 235360
rect 369813 235302 371916 235304
rect 369813 235299 369879 235302
rect 74401 235090 74467 235093
rect 136961 235092 137027 235093
rect 74534 235090 74540 235092
rect 74401 235088 74540 235090
rect 74401 235032 74406 235088
rect 74462 235032 74540 235088
rect 74401 235030 74540 235032
rect 74401 235027 74467 235030
rect 74534 235028 74540 235030
rect 74604 235028 74610 235092
rect 136910 235090 136916 235092
rect 136870 235030 136916 235090
rect 136980 235090 137027 235092
rect 147817 235090 147883 235093
rect 136980 235088 147883 235090
rect 137022 235032 147822 235088
rect 147878 235032 147883 235088
rect 136910 235028 136916 235030
rect 136980 235030 147883 235032
rect 136980 235028 137027 235030
rect 136961 235027 137027 235028
rect 147817 235027 147883 235030
rect 74534 234892 74540 234956
rect 74604 234954 74610 234956
rect 74677 234954 74743 234957
rect 74604 234952 74743 234954
rect 74604 234896 74682 234952
rect 74738 234896 74743 234952
rect 74604 234894 74743 234896
rect 74604 234892 74610 234894
rect 74677 234891 74743 234894
rect 137697 234954 137763 234957
rect 137830 234954 137836 234956
rect 137697 234952 137836 234954
rect 137697 234896 137702 234952
rect 137758 234896 137836 234952
rect 137697 234894 137836 234896
rect 137697 234891 137763 234894
rect 137830 234892 137836 234894
rect 137900 234892 137906 234956
rect 139261 234954 139327 234957
rect 152049 234956 152115 234957
rect 207249 234956 207315 234957
rect 145006 234954 145012 234956
rect 139261 234952 145012 234954
rect 139261 234896 139266 234952
rect 139322 234896 145012 234952
rect 139261 234894 145012 234896
rect 139261 234891 139327 234894
rect 145006 234892 145012 234894
rect 145076 234892 145082 234956
rect 151998 234892 152004 234956
rect 152068 234954 152115 234956
rect 152068 234952 152160 234954
rect 152110 234896 152160 234952
rect 152068 234894 152160 234896
rect 152068 234892 152115 234894
rect 207198 234892 207204 234956
rect 207268 234954 207315 234956
rect 231813 234956 231879 234957
rect 231813 234954 231860 234956
rect 207268 234952 207360 234954
rect 207310 234896 207360 234952
rect 207268 234894 207360 234896
rect 231768 234952 231860 234954
rect 231768 234896 231818 234952
rect 231768 234894 231860 234896
rect 207268 234892 207315 234894
rect 152049 234891 152115 234892
rect 207249 234891 207315 234892
rect 231813 234892 231860 234894
rect 231924 234892 231930 234956
rect 234798 234892 234804 234956
rect 234868 234954 234874 234956
rect 237742 234954 237748 234956
rect 234868 234894 237748 234954
rect 234868 234892 234874 234894
rect 237742 234892 237748 234894
rect 237812 234954 237818 234956
rect 244366 234954 244372 234956
rect 237812 234894 244372 234954
rect 237812 234892 237818 234894
rect 244366 234892 244372 234894
rect 244436 234892 244442 234956
rect 301038 234892 301044 234956
rect 301108 234954 301114 234956
rect 301457 234954 301523 234957
rect 302009 234954 302075 234957
rect 301108 234952 302075 234954
rect 301108 234896 301462 234952
rect 301518 234896 302014 234952
rect 302070 234896 302075 234952
rect 301108 234894 302075 234896
rect 301108 234892 301114 234894
rect 231813 234891 231879 234892
rect 301457 234891 301523 234894
rect 302009 234891 302075 234894
rect 369997 234954 370063 234957
rect 369997 234952 371916 234954
rect 369997 234896 370002 234952
rect 370058 234896 371916 234952
rect 369997 234894 371916 234896
rect 369997 234891 370063 234894
rect 369905 234546 369971 234549
rect 369905 234544 371916 234546
rect 369905 234488 369910 234544
rect 369966 234488 371916 234544
rect 369905 234486 371916 234488
rect 369905 234483 369971 234486
rect 284294 234348 284300 234412
rect 284364 234410 284370 234412
rect 325653 234410 325719 234413
rect 284364 234408 325719 234410
rect 284364 234352 325658 234408
rect 325714 234352 325719 234408
rect 284364 234350 325719 234352
rect 284364 234348 284370 234350
rect 325653 234347 325719 234350
rect 245981 234276 246047 234277
rect 141142 234212 141148 234276
rect 141212 234274 141218 234276
rect 147766 234274 147772 234276
rect 141212 234214 147772 234274
rect 141212 234212 141218 234214
rect 147766 234212 147772 234214
rect 147836 234212 147842 234276
rect 147950 234212 147956 234276
rect 148020 234274 148026 234276
rect 153102 234274 153108 234276
rect 148020 234214 153108 234274
rect 148020 234212 148026 234214
rect 153102 234212 153108 234214
rect 153172 234212 153178 234276
rect 245981 234274 246028 234276
rect 245936 234272 246028 234274
rect 245936 234216 245986 234272
rect 245936 234214 246028 234216
rect 245981 234212 246028 234214
rect 246092 234212 246098 234276
rect 245981 234211 246047 234212
rect 368709 234138 368775 234141
rect 368709 234136 371916 234138
rect 368709 234080 368714 234136
rect 368770 234080 371916 234136
rect 368709 234078 371916 234080
rect 368709 234075 368775 234078
rect 73798 233940 73804 234004
rect 73868 234002 73874 234004
rect 75137 234002 75203 234005
rect 73868 234000 75203 234002
rect 73868 233944 75142 234000
rect 75198 233944 75203 234000
rect 73868 233942 75203 233944
rect 73868 233940 73874 233942
rect 75137 233939 75203 233942
rect 73430 233804 73436 233868
rect 73500 233866 73506 233868
rect 75454 233866 75460 233868
rect 73500 233806 75460 233866
rect 73500 233804 73506 233806
rect 75454 233804 75460 233806
rect 75524 233804 75530 233868
rect 73430 233668 73436 233732
rect 73500 233730 73506 233732
rect 73798 233730 73804 233732
rect 73500 233670 73804 233730
rect 73500 233668 73506 233670
rect 73798 233668 73804 233670
rect 73868 233668 73874 233732
rect 149289 233730 149355 233733
rect 150117 233730 150183 233733
rect 169110 233730 169116 233732
rect 149289 233728 169116 233730
rect 149289 233672 149294 233728
rect 149350 233672 150122 233728
rect 150178 233672 169116 233728
rect 149289 233670 169116 233672
rect 149289 233667 149355 233670
rect 150117 233667 150183 233670
rect 169110 233668 169116 233670
rect 169180 233668 169186 233732
rect 368709 233730 368775 233733
rect 368709 233728 371916 233730
rect 368709 233672 368714 233728
rect 368770 233672 371916 233728
rect 368709 233670 371916 233672
rect 368709 233667 368775 233670
rect 153102 233532 153108 233596
rect 153172 233594 153178 233596
rect 153245 233594 153311 233597
rect 167822 233594 167828 233596
rect 153172 233592 167828 233594
rect 153172 233536 153250 233592
rect 153306 233536 167828 233592
rect 153172 233534 167828 233536
rect 153172 233532 153178 233534
rect 153245 233531 153311 233534
rect 167822 233532 167828 233534
rect 167892 233532 167898 233596
rect 241473 233594 241539 233597
rect 249886 233594 249892 233596
rect 241473 233592 249892 233594
rect 241473 233536 241478 233592
rect 241534 233536 249892 233592
rect 241473 233534 249892 233536
rect 241473 233531 241539 233534
rect 249886 233532 249892 233534
rect 249956 233532 249962 233596
rect 289998 233532 290004 233596
rect 290068 233594 290074 233596
rect 297542 233594 297548 233596
rect 290068 233534 297548 233594
rect 290068 233532 290074 233534
rect 297542 233532 297548 233534
rect 297612 233532 297618 233596
rect 243037 233458 243103 233461
rect 262950 233458 262956 233460
rect 243037 233456 262956 233458
rect 243037 233400 243042 233456
rect 243098 233400 262956 233456
rect 243037 233398 262956 233400
rect 243037 233395 243103 233398
rect 262950 233396 262956 233398
rect 263020 233396 263026 233460
rect 368801 233458 368867 233461
rect 368801 233456 371916 233458
rect 368801 233400 368806 233456
rect 368862 233400 371916 233456
rect 368801 233398 371916 233400
rect 368801 233395 368867 233398
rect 137145 233050 137211 233053
rect 149289 233050 149355 233053
rect 137145 233048 149355 233050
rect 137145 232992 137150 233048
rect 137206 232992 149294 233048
rect 149350 232992 149355 233048
rect 137145 232990 149355 232992
rect 137145 232987 137211 232990
rect 149289 232987 149355 232990
rect 368893 233050 368959 233053
rect 429797 233050 429863 233053
rect 434416 233050 434896 233080
rect 368893 233048 371916 233050
rect 368893 232992 368898 233048
rect 368954 232992 371916 233048
rect 368893 232990 371916 232992
rect 429797 233048 434896 233050
rect 429797 232992 429802 233048
rect 429858 232992 434896 233048
rect 429797 232990 434896 232992
rect 368893 232987 368959 232990
rect 429797 232987 429863 232990
rect 434416 232960 434896 232990
rect 259638 232852 259644 232916
rect 259708 232914 259714 232916
rect 269206 232914 269212 232916
rect 259708 232854 269212 232914
rect 259708 232852 259714 232854
rect 269206 232852 269212 232854
rect 269276 232852 269282 232916
rect 282638 232852 282644 232916
rect 282708 232914 282714 232916
rect 285214 232914 285220 232916
rect 282708 232854 285220 232914
rect 282708 232852 282714 232854
rect 285214 232852 285220 232854
rect 285284 232852 285290 232916
rect 369721 232642 369787 232645
rect 369721 232640 371916 232642
rect 369721 232584 369726 232640
rect 369782 232584 371916 232640
rect 369721 232582 371916 232584
rect 369721 232579 369787 232582
rect 52638 232444 52644 232508
rect 52708 232506 52714 232508
rect 53517 232506 53583 232509
rect 52708 232504 53583 232506
rect 52708 232448 53522 232504
rect 53578 232448 53583 232504
rect 52708 232446 53583 232448
rect 52708 232444 52714 232446
rect 53517 232443 53583 232446
rect 54529 232506 54595 232509
rect 54662 232506 54668 232508
rect 54529 232504 54668 232506
rect 54529 232448 54534 232504
rect 54590 232448 54668 232504
rect 54529 232446 54668 232448
rect 54529 232443 54595 232446
rect 54662 232444 54668 232446
rect 54732 232444 54738 232508
rect 350953 232506 351019 232509
rect 351638 232506 351644 232508
rect 350953 232504 351644 232506
rect 350953 232448 350958 232504
rect 351014 232448 351644 232504
rect 350953 232446 351644 232448
rect 350953 232443 351019 232446
rect 351638 232444 351644 232446
rect 351708 232444 351714 232508
rect 351822 232444 351828 232508
rect 351892 232506 351898 232508
rect 352057 232506 352123 232509
rect 351892 232504 352123 232506
rect 351892 232448 352062 232504
rect 352118 232448 352123 232504
rect 351892 232446 352123 232448
rect 351892 232444 351898 232446
rect 352057 232443 352123 232446
rect 368709 232234 368775 232237
rect 368709 232232 371916 232234
rect 368709 232176 368714 232232
rect 368770 232176 371916 232232
rect 368709 232174 371916 232176
rect 368709 232171 368775 232174
rect 368801 231826 368867 231829
rect 368801 231824 371916 231826
rect 368801 231768 368806 231824
rect 368862 231768 371916 231824
rect 368801 231766 371916 231768
rect 368801 231763 368867 231766
rect 368893 231418 368959 231421
rect 368893 231416 371916 231418
rect 368893 231360 368898 231416
rect 368954 231360 371916 231416
rect 368893 231358 371916 231360
rect 368893 231355 368959 231358
rect 55398 230948 55404 231012
rect 55468 231010 55474 231012
rect 56553 231010 56619 231013
rect 74217 231012 74283 231013
rect 74166 231010 74172 231012
rect 55468 231008 56619 231010
rect 55468 230952 56558 231008
rect 56614 230952 56619 231008
rect 55468 230950 56619 230952
rect 74126 230950 74172 231010
rect 74236 231008 74283 231012
rect 74278 230952 74283 231008
rect 55468 230948 55474 230950
rect 56553 230947 56619 230950
rect 74166 230948 74172 230950
rect 74236 230948 74283 230952
rect 74217 230947 74283 230948
rect 368801 231010 368867 231013
rect 368801 231008 371916 231010
rect 368801 230952 368806 231008
rect 368862 230952 371916 231008
rect 368801 230950 371916 230952
rect 368801 230947 368867 230950
rect 368709 230602 368775 230605
rect 368709 230600 371916 230602
rect 368709 230544 368714 230600
rect 368770 230544 371916 230600
rect 368709 230542 371916 230544
rect 368709 230539 368775 230542
rect 368893 230194 368959 230197
rect 368893 230192 371916 230194
rect 368893 230136 368898 230192
rect 368954 230136 371916 230192
rect 368893 230134 371916 230136
rect 368893 230131 368959 230134
rect 369537 229922 369603 229925
rect 369537 229920 371916 229922
rect 369537 229864 369542 229920
rect 369598 229864 371916 229920
rect 369537 229862 371916 229864
rect 369537 229859 369603 229862
rect 9896 229786 10376 229816
rect 12853 229786 12919 229789
rect 9896 229784 12919 229786
rect 9896 229728 12858 229784
rect 12914 229728 12919 229784
rect 9896 229726 12919 229728
rect 9896 229696 10376 229726
rect 12853 229723 12919 229726
rect 55541 229652 55607 229653
rect 55541 229648 55588 229652
rect 55652 229650 55658 229652
rect 55541 229592 55546 229648
rect 55541 229588 55588 229592
rect 55652 229590 55698 229650
rect 55652 229588 55658 229590
rect 55541 229587 55607 229588
rect 368709 229514 368775 229517
rect 368709 229512 371916 229514
rect 368709 229456 368714 229512
rect 368770 229456 371916 229512
rect 368709 229454 371916 229456
rect 368709 229451 368775 229454
rect 73982 229044 73988 229108
rect 74052 229106 74058 229108
rect 74350 229106 74356 229108
rect 74052 229046 74356 229106
rect 74052 229044 74058 229046
rect 74350 229044 74356 229046
rect 74420 229044 74426 229108
rect 368801 229106 368867 229109
rect 368801 229104 371916 229106
rect 368801 229048 368806 229104
rect 368862 229048 371916 229104
rect 368801 229046 371916 229048
rect 368801 229043 368867 229046
rect 73982 228908 73988 228972
rect 74052 228970 74058 228972
rect 74534 228970 74540 228972
rect 74052 228910 74540 228970
rect 74052 228908 74058 228910
rect 74534 228908 74540 228910
rect 74604 228908 74610 228972
rect 368709 228698 368775 228701
rect 368709 228696 371916 228698
rect 368709 228640 368714 228696
rect 368770 228640 371916 228696
rect 368709 228638 371916 228640
rect 368709 228635 368775 228638
rect 324590 228228 324596 228292
rect 324660 228290 324666 228292
rect 325510 228290 325516 228292
rect 324660 228230 325516 228290
rect 324660 228228 324666 228230
rect 325510 228228 325516 228230
rect 325580 228228 325586 228292
rect 368709 228290 368775 228293
rect 368709 228288 371916 228290
rect 368709 228232 368714 228288
rect 368770 228232 371916 228288
rect 368709 228230 371916 228232
rect 368709 228227 368775 228230
rect 369537 227882 369603 227885
rect 369537 227880 371916 227882
rect 369537 227824 369542 227880
rect 369598 227824 371916 227880
rect 369537 227822 371916 227824
rect 369537 227819 369603 227822
rect 368801 227474 368867 227477
rect 368801 227472 371916 227474
rect 368801 227416 368806 227472
rect 368862 227416 371916 227472
rect 368801 227414 371916 227416
rect 368801 227411 368867 227414
rect 368709 227066 368775 227069
rect 368709 227064 371916 227066
rect 368709 227008 368714 227064
rect 368770 227008 371916 227064
rect 368709 227006 371916 227008
rect 368709 227003 368775 227006
rect 273949 226658 274015 226661
rect 276750 226658 276756 226660
rect 273949 226656 276756 226658
rect 273949 226600 273954 226656
rect 274010 226600 276756 226656
rect 273949 226598 276756 226600
rect 273949 226595 274015 226598
rect 276750 226596 276756 226598
rect 276820 226596 276826 226660
rect 369721 226658 369787 226661
rect 369721 226656 371916 226658
rect 369721 226600 369726 226656
rect 369782 226600 371916 226656
rect 369721 226598 371916 226600
rect 369721 226595 369787 226598
rect 92566 226460 92572 226524
rect 92636 226522 92642 226524
rect 368985 226522 369051 226525
rect 92636 226520 369051 226522
rect 92636 226464 368990 226520
rect 369046 226464 369051 226520
rect 92636 226462 369051 226464
rect 92636 226460 92642 226462
rect 368985 226459 369051 226462
rect 137697 226386 137763 226389
rect 230893 226386 230959 226389
rect 322985 226386 323051 226389
rect 134740 226384 137763 226386
rect 134740 226328 137702 226384
rect 137758 226328 137763 226384
rect 134740 226326 137763 226328
rect 228764 226384 230959 226386
rect 228764 226328 230898 226384
rect 230954 226328 230959 226384
rect 228764 226326 230959 226328
rect 322788 226384 323051 226386
rect 322788 226328 322990 226384
rect 323046 226328 323051 226384
rect 322788 226326 323051 226328
rect 137697 226323 137763 226326
rect 230893 226323 230959 226326
rect 322985 226323 323051 226326
rect 368893 226386 368959 226389
rect 368893 226384 371916 226386
rect 368893 226328 368898 226384
rect 368954 226328 371916 226384
rect 368893 226326 371916 226328
rect 368893 226323 368959 226326
rect 368801 225978 368867 225981
rect 368801 225976 371916 225978
rect 368801 225920 368806 225976
rect 368862 225920 371916 225976
rect 368801 225918 371916 225920
rect 368801 225915 368867 225918
rect 368709 225570 368775 225573
rect 368709 225568 371916 225570
rect 368709 225512 368714 225568
rect 368770 225512 371916 225568
rect 368709 225510 371916 225512
rect 368709 225507 368775 225510
rect 345709 225434 345775 225437
rect 355686 225434 355692 225436
rect 345709 225432 355692 225434
rect 345709 225376 345714 225432
rect 345770 225376 355692 225432
rect 345709 225374 355692 225376
rect 345709 225371 345775 225374
rect 355686 225372 355692 225374
rect 355756 225372 355762 225436
rect 368801 225162 368867 225165
rect 368801 225160 371916 225162
rect 368801 225104 368806 225160
rect 368862 225104 371916 225160
rect 368801 225102 371916 225104
rect 368801 225099 368867 225102
rect 341293 224890 341359 224893
rect 342673 224890 342739 224893
rect 341293 224888 342739 224890
rect 341293 224832 341298 224888
rect 341354 224832 342678 224888
rect 342734 224832 342739 224888
rect 341293 224830 342739 224832
rect 341293 224827 341359 224830
rect 342673 224827 342739 224830
rect 368709 224754 368775 224757
rect 368709 224752 371916 224754
rect 368709 224696 368714 224752
rect 368770 224696 371916 224752
rect 368709 224694 371916 224696
rect 368709 224691 368775 224694
rect 324958 224284 324964 224348
rect 325028 224346 325034 224348
rect 325377 224346 325443 224349
rect 325028 224344 325443 224346
rect 325028 224288 325382 224344
rect 325438 224288 325443 224344
rect 325028 224286 325443 224288
rect 325028 224284 325034 224286
rect 325377 224283 325443 224286
rect 369261 224346 369327 224349
rect 369261 224344 371916 224346
rect 369261 224288 369266 224344
rect 369322 224288 371916 224344
rect 369261 224286 371916 224288
rect 369261 224283 369327 224286
rect 368801 223938 368867 223941
rect 368801 223936 371916 223938
rect 368801 223880 368806 223936
rect 368862 223880 371916 223936
rect 368801 223878 371916 223880
rect 368801 223875 368867 223878
rect 368985 223530 369051 223533
rect 368985 223528 371916 223530
rect 368985 223472 368990 223528
rect 369046 223472 371916 223528
rect 368985 223470 371916 223472
rect 368985 223467 369051 223470
rect 137329 223258 137395 223261
rect 230985 223258 231051 223261
rect 324733 223258 324799 223261
rect 134740 223256 137395 223258
rect 134740 223200 137334 223256
rect 137390 223200 137395 223256
rect 134740 223198 137395 223200
rect 228764 223256 231051 223258
rect 228764 223200 230990 223256
rect 231046 223200 231051 223256
rect 228764 223198 231051 223200
rect 322788 223256 324799 223258
rect 322788 223200 324738 223256
rect 324794 223200 324799 223256
rect 322788 223198 324799 223200
rect 137329 223195 137395 223198
rect 230985 223195 231051 223198
rect 324733 223195 324799 223198
rect 368709 223258 368775 223261
rect 368709 223256 371916 223258
rect 368709 223200 368714 223256
rect 368770 223200 371916 223256
rect 368709 223198 371916 223200
rect 368709 223195 368775 223198
rect 368893 222850 368959 222853
rect 368893 222848 371916 222850
rect 368893 222792 368898 222848
rect 368954 222792 371916 222848
rect 368893 222790 371916 222792
rect 368893 222787 368959 222790
rect 368801 222442 368867 222445
rect 368801 222440 371916 222442
rect 368801 222384 368806 222440
rect 368862 222384 371916 222440
rect 368801 222382 371916 222384
rect 368801 222379 368867 222382
rect 55398 222034 55404 222036
rect 35718 221974 55404 222034
rect 35718 221528 35778 221974
rect 55398 221972 55404 221974
rect 55468 221972 55474 222036
rect 357669 222034 357735 222037
rect 358630 222034 358636 222036
rect 357669 222032 358636 222034
rect 357669 221976 357674 222032
rect 357730 221976 358636 222032
rect 357669 221974 358636 221976
rect 357669 221971 357735 221974
rect 358630 221972 358636 221974
rect 358700 221972 358706 222036
rect 368893 222034 368959 222037
rect 368893 222032 371916 222034
rect 368893 221976 368898 222032
rect 368954 221976 371916 222032
rect 368893 221974 371916 221976
rect 368893 221971 368959 221974
rect 405918 221972 405924 222036
rect 405988 222034 405994 222036
rect 405988 221974 408930 222034
rect 405988 221972 405994 221974
rect 368709 221626 368775 221629
rect 368709 221624 371916 221626
rect 368709 221568 368714 221624
rect 368770 221568 371916 221624
rect 368709 221566 371916 221568
rect 368709 221563 368775 221566
rect 74217 221490 74283 221493
rect 74350 221490 74356 221492
rect 74217 221488 74356 221490
rect 74217 221432 74222 221488
rect 74278 221432 74356 221488
rect 74217 221430 74356 221432
rect 74217 221427 74283 221430
rect 74350 221428 74356 221430
rect 74420 221428 74426 221492
rect 408870 221460 408930 221974
rect 53241 221354 53307 221357
rect 55582 221354 55588 221356
rect 53241 221352 55588 221354
rect 53241 221296 53246 221352
rect 53302 221296 55588 221352
rect 53241 221294 55588 221296
rect 53241 221291 53307 221294
rect 55582 221292 55588 221294
rect 55652 221354 55658 221356
rect 56318 221354 56324 221356
rect 55652 221294 56324 221354
rect 55652 221292 55658 221294
rect 56318 221292 56324 221294
rect 56388 221292 56394 221356
rect 368893 221218 368959 221221
rect 368893 221216 371916 221218
rect 368893 221160 368898 221216
rect 368954 221160 371916 221216
rect 368893 221158 371916 221160
rect 368893 221155 368959 221158
rect 428693 220946 428759 220949
rect 434416 220946 434896 220976
rect 428693 220944 434896 220946
rect 70678 220402 70738 220916
rect 428693 220888 428698 220944
rect 428754 220888 434896 220944
rect 428693 220886 434896 220888
rect 428693 220883 428759 220886
rect 434416 220856 434896 220886
rect 368801 220810 368867 220813
rect 368801 220808 371916 220810
rect 368801 220752 368806 220808
rect 368862 220752 371916 220808
rect 368801 220750 371916 220752
rect 368801 220747 368867 220750
rect 74309 220402 74375 220405
rect 70678 220400 74375 220402
rect 70678 220344 74314 220400
rect 74370 220344 74375 220400
rect 70678 220342 74375 220344
rect 74309 220339 74375 220342
rect 368709 220402 368775 220405
rect 368709 220400 371916 220402
rect 368709 220344 368714 220400
rect 368770 220344 371916 220400
rect 368709 220342 371916 220344
rect 368709 220339 368775 220342
rect 51861 220266 51927 220269
rect 355093 220266 355159 220269
rect 427405 220266 427471 220269
rect 51861 220264 55068 220266
rect 16165 219994 16231 219997
rect 20078 219994 20138 220236
rect 51861 220208 51866 220264
rect 51922 220208 55068 220264
rect 51861 220206 55068 220208
rect 352780 220264 355159 220266
rect 352780 220208 355098 220264
rect 355154 220208 355159 220264
rect 352780 220206 355159 220208
rect 424724 220264 427471 220266
rect 424724 220208 427410 220264
rect 427466 220208 427471 220264
rect 424724 220206 427471 220208
rect 51861 220203 51927 220206
rect 355093 220203 355159 220206
rect 427405 220203 427471 220206
rect 137237 220130 137303 220133
rect 230801 220130 230867 220133
rect 324549 220130 324615 220133
rect 134740 220128 137303 220130
rect 134740 220072 137242 220128
rect 137298 220072 137303 220128
rect 134740 220070 137303 220072
rect 228764 220128 230867 220130
rect 228764 220072 230806 220128
rect 230862 220072 230867 220128
rect 228764 220070 230867 220072
rect 322788 220128 324615 220130
rect 322788 220072 324554 220128
rect 324610 220072 324615 220128
rect 322788 220070 324615 220072
rect 137237 220067 137303 220070
rect 230801 220067 230867 220070
rect 324549 220067 324615 220070
rect 16165 219992 20138 219994
rect 16165 219936 16170 219992
rect 16226 219936 20138 219992
rect 16165 219934 20138 219936
rect 369813 219994 369879 219997
rect 369813 219992 371916 219994
rect 369813 219936 369818 219992
rect 369874 219936 371916 219992
rect 369813 219934 371916 219936
rect 16165 219931 16231 219934
rect 369813 219931 369879 219934
rect 368709 219722 368775 219725
rect 368709 219720 371916 219722
rect 368709 219664 368714 219720
rect 368770 219664 371916 219720
rect 368709 219662 371916 219664
rect 368709 219659 368775 219662
rect 81669 219586 81735 219589
rect 179281 219586 179347 219589
rect 272937 219586 273003 219589
rect 81669 219584 85060 219586
rect 81669 219528 81674 219584
rect 81730 219528 85060 219584
rect 81669 219526 85060 219528
rect 179268 219584 179347 219586
rect 179268 219528 179286 219584
rect 179342 219528 179347 219584
rect 179268 219526 179347 219528
rect 272924 219584 273003 219586
rect 272924 219528 272942 219584
rect 272998 219528 273003 219584
rect 272924 219526 273003 219528
rect 81669 219523 81735 219526
rect 179281 219523 179347 219526
rect 272937 219523 273003 219526
rect 38061 219450 38127 219453
rect 35718 219448 38127 219450
rect 35718 219392 38066 219448
rect 38122 219392 38127 219448
rect 35718 219390 38127 219392
rect 35718 219080 35778 219390
rect 38061 219387 38127 219390
rect 369077 219314 369143 219317
rect 369077 219312 371916 219314
rect 369077 219256 369082 219312
rect 369138 219256 371916 219312
rect 369077 219254 371916 219256
rect 369077 219251 369143 219254
rect 9896 218906 10376 218936
rect 13037 218906 13103 218909
rect 9896 218904 13103 218906
rect 9896 218848 13042 218904
rect 13098 218848 13103 218904
rect 9896 218846 13103 218848
rect 9896 218816 10376 218846
rect 13037 218843 13103 218846
rect 368801 218906 368867 218909
rect 368801 218904 371916 218906
rect 368801 218848 368806 218904
rect 368862 218848 371916 218904
rect 368801 218846 371916 218848
rect 368801 218843 368867 218846
rect 405969 218770 406035 218773
rect 409054 218770 409114 219012
rect 405969 218768 409114 218770
rect 405969 218712 405974 218768
rect 406030 218712 409114 218768
rect 405969 218710 409114 218712
rect 405969 218707 406035 218710
rect 369261 218498 369327 218501
rect 369261 218496 371916 218498
rect 369261 218440 369266 218496
rect 369322 218440 371916 218496
rect 369261 218438 371916 218440
rect 369261 218435 369327 218438
rect 368709 218090 368775 218093
rect 368709 218088 371916 218090
rect 368709 218032 368714 218088
rect 368770 218032 371916 218088
rect 368709 218030 371916 218032
rect 368709 218027 368775 218030
rect 368985 217682 369051 217685
rect 368985 217680 371916 217682
rect 368985 217624 368990 217680
rect 369046 217624 371916 217680
rect 368985 217622 371916 217624
rect 368985 217619 369051 217622
rect 75413 217410 75479 217413
rect 70862 217408 75479 217410
rect 70862 217352 75418 217408
rect 75474 217352 75479 217408
rect 70862 217350 75479 217352
rect 70862 217244 70922 217350
rect 75413 217347 75479 217350
rect 368801 217274 368867 217277
rect 368801 217272 371916 217274
rect 368801 217216 368806 217272
rect 368862 217216 371916 217272
rect 368801 217214 371916 217216
rect 368801 217211 368867 217214
rect 322934 217076 322940 217140
rect 323004 217138 323010 217140
rect 323004 217078 323554 217138
rect 323004 217076 323010 217078
rect 137145 217002 137211 217005
rect 230709 217002 230775 217005
rect 134740 217000 137211 217002
rect 134740 216944 137150 217000
rect 137206 216944 137211 217000
rect 134740 216942 137211 216944
rect 228764 217000 230775 217002
rect 228764 216944 230714 217000
rect 230770 216944 230775 217000
rect 228764 216942 230775 216944
rect 137145 216939 137211 216942
rect 230709 216939 230775 216942
rect 231537 217002 231603 217005
rect 242710 217002 242716 217004
rect 231537 217000 242716 217002
rect 231537 216944 231542 217000
rect 231598 216944 242716 217000
rect 231537 216942 242716 216944
rect 231537 216939 231603 216942
rect 242710 216940 242716 216942
rect 242780 216940 242786 217004
rect 258718 216940 258724 217004
rect 258788 217002 258794 217004
rect 272702 217002 272708 217004
rect 258788 216942 272708 217002
rect 258788 216940 258794 216942
rect 272702 216940 272708 216942
rect 272772 216940 272778 217004
rect 323494 217002 323554 217078
rect 336918 217002 336924 217004
rect 38521 216866 38587 216869
rect 35718 216864 38587 216866
rect 35718 216808 38526 216864
rect 38582 216808 38587 216864
rect 35718 216806 38587 216808
rect 35718 216496 35778 216806
rect 38521 216803 38587 216806
rect 322758 216730 322818 216972
rect 323494 216942 336924 217002
rect 336918 216940 336924 216942
rect 336988 216940 336994 217004
rect 352742 216940 352748 217004
rect 352812 217002 352818 217004
rect 369077 217002 369143 217005
rect 352812 217000 369143 217002
rect 352812 216944 369082 217000
rect 369138 216944 369143 217000
rect 352812 216942 369143 216944
rect 352812 216940 352818 216942
rect 369077 216939 369143 216942
rect 369077 216866 369143 216869
rect 369077 216864 371916 216866
rect 369077 216808 369082 216864
rect 369138 216808 371916 216864
rect 369077 216806 371916 216808
rect 369077 216803 369143 216806
rect 325837 216730 325903 216733
rect 322758 216728 325903 216730
rect 322758 216672 325842 216728
rect 325898 216672 325903 216728
rect 322758 216670 325903 216672
rect 325837 216667 325903 216670
rect 137697 216594 137763 216597
rect 148686 216594 148692 216596
rect 137697 216592 148692 216594
rect 137697 216536 137702 216592
rect 137758 216536 148692 216592
rect 137697 216534 148692 216536
rect 137697 216531 137763 216534
rect 148686 216532 148692 216534
rect 148756 216532 148762 216596
rect 164878 216532 164884 216596
rect 164948 216594 164954 216596
rect 177574 216594 177580 216596
rect 164948 216534 177580 216594
rect 164948 216532 164954 216534
rect 177574 216532 177580 216534
rect 177644 216532 177650 216596
rect 228910 216532 228916 216596
rect 228980 216594 228986 216596
rect 242710 216594 242716 216596
rect 228980 216534 242716 216594
rect 228980 216532 228986 216534
rect 242710 216532 242716 216534
rect 242780 216532 242786 216596
rect 258718 216532 258724 216596
rect 258788 216594 258794 216596
rect 272702 216594 272708 216596
rect 258788 216534 272708 216594
rect 258788 216532 258794 216534
rect 272702 216532 272708 216534
rect 272772 216532 272778 216596
rect 322934 216532 322940 216596
rect 323004 216594 323010 216596
rect 336734 216594 336740 216596
rect 323004 216534 336740 216594
rect 323004 216532 323010 216534
rect 336734 216532 336740 216534
rect 336804 216532 336810 216596
rect 352742 216532 352748 216596
rect 352812 216594 352818 216596
rect 368985 216594 369051 216597
rect 352812 216592 369051 216594
rect 352812 216536 368990 216592
rect 369046 216536 369051 216592
rect 352812 216534 369051 216536
rect 352812 216532 352818 216534
rect 368985 216531 369051 216534
rect 368709 216458 368775 216461
rect 368709 216456 371916 216458
rect 368709 216400 368714 216456
rect 368770 216400 371916 216456
rect 368709 216398 371916 216400
rect 368709 216395 368775 216398
rect 148326 216194 148908 216254
rect 242350 216194 242932 216254
rect 145149 216186 145215 216189
rect 148326 216186 148386 216194
rect 145149 216184 148386 216186
rect 145149 216128 145154 216184
rect 145210 216128 148386 216184
rect 145149 216126 148386 216128
rect 240921 216186 240987 216189
rect 242350 216186 242410 216194
rect 240921 216184 242410 216186
rect 240921 216128 240926 216184
rect 240982 216128 242410 216184
rect 240921 216126 242410 216128
rect 334209 216186 334275 216189
rect 368801 216186 368867 216189
rect 334209 216184 336956 216186
rect 334209 216128 334214 216184
rect 334270 216128 336956 216184
rect 334209 216126 336956 216128
rect 368801 216184 371916 216186
rect 368801 216128 368806 216184
rect 368862 216128 371916 216184
rect 368801 216126 371916 216128
rect 145149 216123 145215 216126
rect 240921 216123 240987 216126
rect 334209 216123 334275 216126
rect 368801 216123 368867 216126
rect 356289 215914 356355 215917
rect 357526 215914 357532 215916
rect 356289 215912 357532 215914
rect 356289 215856 356294 215912
rect 356350 215856 357532 215912
rect 356289 215854 357532 215856
rect 356289 215851 356355 215854
rect 357526 215852 357532 215854
rect 357596 215852 357602 215916
rect 405918 215852 405924 215916
rect 405988 215914 405994 215916
rect 409054 215914 409114 216428
rect 405988 215854 409114 215914
rect 405988 215852 405994 215854
rect 368709 215778 368775 215781
rect 368709 215776 371916 215778
rect 368709 215720 368714 215776
rect 368770 215720 371916 215776
rect 368709 215718 371916 215720
rect 368709 215715 368775 215718
rect 369077 215370 369143 215373
rect 369077 215368 371916 215370
rect 369077 215312 369082 215368
rect 369138 215312 371916 215368
rect 369077 215310 371916 215312
rect 369077 215307 369143 215310
rect 51677 215234 51743 215237
rect 356197 215234 356263 215237
rect 428693 215234 428759 215237
rect 51677 215232 55068 215234
rect 16349 214554 16415 214557
rect 20078 214554 20138 215204
rect 51677 215176 51682 215232
rect 51738 215176 55068 215232
rect 51677 215174 55068 215176
rect 352780 215232 356263 215234
rect 352780 215176 356202 215232
rect 356258 215176 356263 215232
rect 352780 215174 356263 215176
rect 424724 215232 428759 215234
rect 424724 215176 428698 215232
rect 428754 215176 428759 215232
rect 424724 215174 428759 215176
rect 51677 215171 51743 215174
rect 356197 215171 356263 215174
rect 428693 215171 428759 215174
rect 368801 214962 368867 214965
rect 368801 214960 371916 214962
rect 368801 214904 368806 214960
rect 368862 214904 371916 214960
rect 368801 214902 371916 214904
rect 368801 214899 368867 214902
rect 16349 214552 20138 214554
rect 16349 214496 16354 214552
rect 16410 214496 20138 214552
rect 16349 214494 20138 214496
rect 16349 214491 16415 214494
rect 73430 214492 73436 214556
rect 73500 214554 73506 214556
rect 73798 214554 73804 214556
rect 73500 214494 73804 214554
rect 73500 214492 73506 214494
rect 73798 214492 73804 214494
rect 73868 214492 73874 214556
rect 368985 214554 369051 214557
rect 368985 214552 371916 214554
rect 368985 214496 368990 214552
rect 369046 214496 371916 214552
rect 368985 214494 371916 214496
rect 368985 214491 369051 214494
rect 38521 214282 38587 214285
rect 35718 214280 38587 214282
rect 35718 214224 38526 214280
rect 38582 214224 38587 214280
rect 35718 214222 38587 214224
rect 35718 214048 35778 214222
rect 38521 214219 38587 214222
rect 368893 214146 368959 214149
rect 405969 214146 406035 214149
rect 368893 214144 371916 214146
rect 368893 214088 368898 214144
rect 368954 214088 371916 214144
rect 368893 214086 371916 214088
rect 405969 214144 408930 214146
rect 405969 214088 405974 214144
rect 406030 214088 408930 214144
rect 405969 214086 408930 214088
rect 368893 214083 368959 214086
rect 405969 214083 406035 214086
rect 408870 213980 408930 214086
rect 137053 213874 137119 213877
rect 231721 213874 231787 213877
rect 325745 213874 325811 213877
rect 134740 213872 137119 213874
rect 134740 213816 137058 213872
rect 137114 213816 137119 213872
rect 134740 213814 137119 213816
rect 228764 213872 231787 213874
rect 228764 213816 231726 213872
rect 231782 213816 231787 213872
rect 228764 213814 231787 213816
rect 322788 213872 325811 213874
rect 322788 213816 325750 213872
rect 325806 213816 325811 213872
rect 322788 213814 325811 213816
rect 137053 213811 137119 213814
rect 231721 213811 231787 213814
rect 325745 213811 325811 213814
rect 368709 213738 368775 213741
rect 368709 213736 371916 213738
rect 368709 213680 368714 213736
rect 368770 213680 371916 213736
rect 368709 213678 371916 213680
rect 368709 213675 368775 213678
rect 70678 213194 70738 213572
rect 368893 213330 368959 213333
rect 368893 213328 371916 213330
rect 368893 213272 368898 213328
rect 368954 213272 371916 213328
rect 368893 213270 371916 213272
rect 368893 213267 368959 213270
rect 74217 213196 74283 213197
rect 74166 213194 74172 213196
rect 70678 213134 74172 213194
rect 74236 213194 74283 213196
rect 74236 213192 74328 213194
rect 74278 213136 74328 213192
rect 74166 213132 74172 213134
rect 74236 213134 74328 213136
rect 74236 213132 74283 213134
rect 74217 213131 74283 213132
rect 368709 213058 368775 213061
rect 368709 213056 371916 213058
rect 368709 213000 368714 213056
rect 368770 213000 371916 213056
rect 368709 212998 371916 213000
rect 368709 212995 368775 212998
rect 167965 212786 168031 212789
rect 262357 212786 262423 212789
rect 164732 212784 168031 212786
rect 164732 212728 167970 212784
rect 168026 212728 168031 212784
rect 164732 212726 168031 212728
rect 258756 212784 262423 212786
rect 258756 212728 262362 212784
rect 262418 212728 262423 212784
rect 258756 212726 262423 212728
rect 167965 212723 168031 212726
rect 262357 212723 262423 212726
rect 74401 211700 74467 211701
rect 74350 211636 74356 211700
rect 74420 211698 74467 211700
rect 74420 211696 74512 211698
rect 74462 211640 74512 211696
rect 74420 211638 74512 211640
rect 74420 211636 74467 211638
rect 74401 211635 74467 211636
rect 38705 211562 38771 211565
rect 35748 211560 38771 211562
rect 35748 211504 38710 211560
rect 38766 211504 38771 211560
rect 35748 211502 38771 211504
rect 38705 211499 38771 211502
rect 54069 211018 54135 211021
rect 54662 211018 54668 211020
rect 54069 211016 54668 211018
rect 54069 210960 54074 211016
rect 54130 210960 54668 211016
rect 54069 210958 54668 210960
rect 54069 210955 54135 210958
rect 54662 210956 54668 210958
rect 54732 210956 54738 211020
rect 405969 211018 406035 211021
rect 409054 211018 409114 211532
rect 405969 211016 409114 211018
rect 405969 210960 405974 211016
rect 406030 210960 409114 211016
rect 405969 210958 409114 210960
rect 405969 210955 406035 210958
rect 136961 210746 137027 210749
rect 231629 210746 231695 210749
rect 325561 210746 325627 210749
rect 134740 210744 137027 210746
rect 134740 210688 136966 210744
rect 137022 210688 137027 210744
rect 134740 210686 137027 210688
rect 228764 210744 231695 210746
rect 228764 210688 231634 210744
rect 231690 210688 231695 210744
rect 228764 210686 231695 210688
rect 322788 210744 325627 210746
rect 322788 210688 325566 210744
rect 325622 210688 325627 210744
rect 322788 210686 325627 210688
rect 136961 210683 137027 210686
rect 231629 210683 231695 210686
rect 325561 210683 325627 210686
rect 51401 210202 51467 210205
rect 72653 210202 72719 210205
rect 73481 210202 73547 210205
rect 356013 210202 356079 210205
rect 427497 210202 427563 210205
rect 51401 210200 55068 210202
rect 17545 209658 17611 209661
rect 20078 209658 20138 210172
rect 51401 210144 51406 210200
rect 51462 210144 55068 210200
rect 51401 210142 55068 210144
rect 70862 210200 73547 210202
rect 70862 210144 72658 210200
rect 72714 210144 73486 210200
rect 73542 210144 73547 210200
rect 70862 210142 73547 210144
rect 352780 210200 356079 210202
rect 352780 210144 356018 210200
rect 356074 210144 356079 210200
rect 352780 210142 356079 210144
rect 424724 210200 427563 210202
rect 424724 210144 427502 210200
rect 427558 210144 427563 210200
rect 424724 210142 427563 210144
rect 51401 210139 51467 210142
rect 70862 210036 70922 210142
rect 72653 210139 72719 210142
rect 73481 210139 73547 210142
rect 356013 210139 356079 210142
rect 427497 210139 427563 210142
rect 17545 209656 20138 209658
rect 17545 209600 17550 209656
rect 17606 209600 20138 209656
rect 17545 209598 20138 209600
rect 17545 209595 17611 209598
rect 405969 209522 406035 209525
rect 405969 209520 408930 209522
rect 405969 209464 405974 209520
rect 406030 209464 408930 209520
rect 405969 209462 408930 209464
rect 405969 209459 406035 209462
rect 38521 209250 38587 209253
rect 35718 209248 38587 209250
rect 35718 209192 38526 209248
rect 38582 209192 38587 209248
rect 35718 209190 38587 209192
rect 35718 209016 35778 209190
rect 38521 209187 38587 209190
rect 16533 208978 16599 208981
rect 17545 208978 17611 208981
rect 16533 208976 17611 208978
rect 16533 208920 16538 208976
rect 16594 208920 17550 208976
rect 17606 208920 17611 208976
rect 408870 208948 408930 209462
rect 16533 208918 17611 208920
rect 16533 208915 16599 208918
rect 17545 208915 17611 208918
rect 429613 208842 429679 208845
rect 434416 208842 434896 208872
rect 429613 208840 434896 208842
rect 429613 208784 429618 208840
rect 429674 208784 434896 208840
rect 429613 208782 434896 208784
rect 429613 208779 429679 208782
rect 434416 208752 434896 208782
rect 138157 208298 138223 208301
rect 147030 208298 147036 208300
rect 138157 208296 147036 208298
rect 138157 208240 138162 208296
rect 138218 208240 147036 208296
rect 138157 208238 147036 208240
rect 138157 208235 138223 208238
rect 147030 208236 147036 208238
rect 147100 208236 147106 208300
rect 9896 208162 10376 208192
rect 13037 208162 13103 208165
rect 9896 208160 13103 208162
rect 9896 208104 13042 208160
rect 13098 208104 13103 208160
rect 9896 208102 13103 208104
rect 9896 208072 10376 208102
rect 13037 208099 13103 208102
rect 231445 207754 231511 207757
rect 231854 207754 231860 207756
rect 228734 207752 231860 207754
rect 228734 207696 231450 207752
rect 231506 207696 231860 207752
rect 228734 207694 231860 207696
rect 138157 207618 138223 207621
rect 134740 207616 138223 207618
rect 134740 207560 138162 207616
rect 138218 207560 138223 207616
rect 228734 207588 228794 207694
rect 231445 207691 231511 207694
rect 231854 207692 231860 207694
rect 231924 207692 231930 207756
rect 325653 207618 325719 207621
rect 322788 207616 325719 207618
rect 134740 207558 138223 207560
rect 322788 207560 325658 207616
rect 325714 207560 325719 207616
rect 322788 207558 325719 207560
rect 138157 207555 138223 207558
rect 325653 207555 325719 207558
rect 51401 206802 51467 206805
rect 52638 206802 52644 206804
rect 51401 206800 52644 206802
rect 51401 206744 51406 206800
rect 51462 206744 52644 206800
rect 51401 206742 52644 206744
rect 51401 206739 51467 206742
rect 52638 206740 52644 206742
rect 52708 206740 52714 206804
rect 405969 206802 406035 206805
rect 405969 206800 408930 206802
rect 405969 206744 405974 206800
rect 406030 206744 408930 206800
rect 405969 206742 408930 206744
rect 405969 206739 406035 206742
rect 38521 206666 38587 206669
rect 73757 206666 73823 206669
rect 73982 206666 73988 206668
rect 35718 206664 38587 206666
rect 35718 206608 38526 206664
rect 38582 206608 38587 206664
rect 35718 206606 38587 206608
rect 35718 206568 35778 206606
rect 38521 206603 38587 206606
rect 70862 206664 73988 206666
rect 70862 206608 73762 206664
rect 73818 206608 73988 206664
rect 70862 206606 73988 206608
rect 70862 206364 70922 206606
rect 73757 206603 73823 206606
rect 73982 206604 73988 206606
rect 74052 206604 74058 206668
rect 408870 206500 408930 206742
rect 74401 205444 74467 205445
rect 74350 205442 74356 205444
rect 74310 205382 74356 205442
rect 74420 205440 74467 205444
rect 74462 205384 74467 205440
rect 74350 205380 74356 205382
rect 74420 205380 74467 205384
rect 74401 205379 74467 205380
rect 51401 205306 51467 205309
rect 356197 205306 356263 205309
rect 427313 205306 427379 205309
rect 51401 205304 55068 205306
rect 16441 204898 16507 204901
rect 20078 204898 20138 205276
rect 51401 205248 51406 205304
rect 51462 205248 55068 205304
rect 51401 205246 55068 205248
rect 352780 205304 356263 205306
rect 352780 205248 356202 205304
rect 356258 205248 356263 205304
rect 352780 205246 356263 205248
rect 424724 205304 427379 205306
rect 424724 205248 427318 205304
rect 427374 205248 427379 205304
rect 424724 205246 427379 205248
rect 51401 205243 51467 205246
rect 356197 205243 356263 205246
rect 427313 205243 427379 205246
rect 73430 204972 73436 205036
rect 73500 205034 73506 205036
rect 73941 205034 74007 205037
rect 73500 205032 74007 205034
rect 73500 204976 73946 205032
rect 74002 204976 74007 205032
rect 73500 204974 74007 204976
rect 73500 204972 73506 204974
rect 73941 204971 74007 204974
rect 134702 204972 134708 205036
rect 134772 204972 134778 205036
rect 16441 204896 20138 204898
rect 16441 204840 16446 204896
rect 16502 204840 20138 204896
rect 16441 204838 20138 204840
rect 16441 204835 16507 204838
rect 73430 204836 73436 204900
rect 73500 204898 73506 204900
rect 73982 204898 73988 204900
rect 73500 204838 73988 204898
rect 73500 204836 73506 204838
rect 73982 204836 73988 204838
rect 74052 204836 74058 204900
rect 38521 204490 38587 204493
rect 35718 204488 38587 204490
rect 35718 204432 38526 204488
rect 38582 204432 38587 204488
rect 35718 204430 38587 204432
rect 35718 204120 35778 204430
rect 38521 204427 38587 204430
rect 73614 204428 73620 204492
rect 73684 204490 73690 204492
rect 74217 204490 74283 204493
rect 84654 204490 84660 204492
rect 73684 204488 84660 204490
rect 73684 204432 74222 204488
rect 74278 204432 84660 204488
rect 73684 204430 84660 204432
rect 73684 204428 73690 204430
rect 74217 204427 74283 204430
rect 84654 204428 84660 204430
rect 84724 204428 84730 204492
rect 134710 204490 134770 204972
rect 406061 204626 406127 204629
rect 406061 204624 408930 204626
rect 406061 204568 406066 204624
rect 406122 204568 408930 204624
rect 406061 204566 408930 204568
rect 406061 204563 406127 204566
rect 136869 204490 136935 204493
rect 231997 204490 232063 204493
rect 325469 204490 325535 204493
rect 134710 204488 136935 204490
rect 134710 204460 136874 204488
rect 134740 204432 136874 204460
rect 136930 204432 136935 204488
rect 134740 204430 136935 204432
rect 228764 204488 232063 204490
rect 228764 204432 232002 204488
rect 232058 204432 232063 204488
rect 228764 204430 232063 204432
rect 322788 204488 325535 204490
rect 322788 204432 325474 204488
rect 325530 204432 325535 204488
rect 322788 204430 325535 204432
rect 136869 204427 136935 204430
rect 231997 204427 232063 204430
rect 325469 204427 325535 204430
rect 408870 204052 408930 204566
rect 73614 203266 73620 203268
rect 70862 203206 73620 203266
rect 70862 202692 70922 203206
rect 73614 203204 73620 203206
rect 73684 203266 73690 203268
rect 74125 203266 74191 203269
rect 73684 203264 74191 203266
rect 73684 203208 74130 203264
rect 74186 203208 74191 203264
rect 73684 203206 74191 203208
rect 73684 203204 73690 203206
rect 74125 203203 74191 203206
rect 148326 202866 148908 202926
rect 242350 202866 242932 202926
rect 81669 202858 81735 202861
rect 145425 202858 145491 202861
rect 148326 202858 148386 202866
rect 178913 202858 178979 202861
rect 81669 202856 85060 202858
rect 81669 202800 81674 202856
rect 81730 202800 85060 202856
rect 81669 202798 85060 202800
rect 145425 202856 148386 202858
rect 145425 202800 145430 202856
rect 145486 202800 148386 202856
rect 145425 202798 148386 202800
rect 178900 202856 178979 202858
rect 178900 202800 178918 202856
rect 178974 202800 178979 202856
rect 178900 202798 178979 202800
rect 81669 202795 81735 202798
rect 145425 202795 145491 202798
rect 178913 202795 178979 202798
rect 240645 202858 240711 202861
rect 242350 202858 242410 202866
rect 272937 202858 273003 202861
rect 240645 202856 242410 202858
rect 240645 202800 240650 202856
rect 240706 202800 242410 202856
rect 240645 202798 242410 202800
rect 272924 202856 273003 202858
rect 272924 202800 272942 202856
rect 272998 202800 273003 202856
rect 272924 202798 273003 202800
rect 240645 202795 240711 202798
rect 272937 202795 273003 202798
rect 334209 202858 334275 202861
rect 334209 202856 336956 202858
rect 334209 202800 334214 202856
rect 334270 202800 336956 202856
rect 334209 202798 336956 202800
rect 334209 202795 334275 202798
rect 38521 201498 38587 201501
rect 35748 201496 38587 201498
rect 35748 201440 38526 201496
rect 38582 201440 38587 201496
rect 35748 201438 38587 201440
rect 38521 201435 38587 201438
rect 405969 201362 406035 201365
rect 409054 201362 409114 201468
rect 405969 201360 409114 201362
rect 134710 200954 134770 201264
rect 136869 200954 136935 200957
rect 137830 200954 137836 200956
rect 134710 200952 137836 200954
rect 134710 200896 136874 200952
rect 136930 200896 137836 200952
rect 134710 200894 137836 200896
rect 136869 200891 136935 200894
rect 137830 200892 137836 200894
rect 137900 200892 137906 200956
rect 228734 200682 228794 201264
rect 322758 200956 322818 201332
rect 405969 201304 405974 201360
rect 406030 201304 409114 201360
rect 405969 201302 409114 201304
rect 405969 201299 406035 201302
rect 322750 200892 322756 200956
rect 322820 200892 322826 200956
rect 230750 200682 230756 200684
rect 228734 200622 230756 200682
rect 230750 200620 230756 200622
rect 230820 200682 230826 200684
rect 230893 200682 230959 200685
rect 230820 200680 230959 200682
rect 230820 200624 230898 200680
rect 230954 200624 230959 200680
rect 230820 200622 230959 200624
rect 230820 200620 230826 200622
rect 230893 200619 230959 200622
rect 74309 200548 74375 200549
rect 74309 200546 74356 200548
rect 74264 200544 74356 200546
rect 74264 200488 74314 200544
rect 74264 200486 74356 200488
rect 74309 200484 74356 200486
rect 74420 200484 74426 200548
rect 74309 200483 74375 200484
rect 51769 200274 51835 200277
rect 355921 200274 355987 200277
rect 427129 200274 427195 200277
rect 51769 200272 55068 200274
rect 17637 199730 17703 199733
rect 20078 199730 20138 200244
rect 51769 200216 51774 200272
rect 51830 200216 55068 200272
rect 51769 200214 55068 200216
rect 352780 200272 355987 200274
rect 352780 200216 355926 200272
rect 355982 200216 355987 200272
rect 352780 200214 355987 200216
rect 424724 200272 427195 200274
rect 424724 200216 427134 200272
rect 427190 200216 427195 200272
rect 424724 200214 427195 200216
rect 51769 200211 51835 200214
rect 355921 200211 355987 200214
rect 427129 200211 427195 200214
rect 17637 199728 20138 199730
rect 17637 199672 17642 199728
rect 17698 199672 20138 199728
rect 17637 199670 20138 199672
rect 17637 199667 17703 199670
rect 73757 199324 73823 199325
rect 73757 199322 73804 199324
rect 73712 199320 73804 199322
rect 73712 199264 73762 199320
rect 73712 199262 73804 199264
rect 73757 199260 73804 199262
rect 73868 199260 73874 199324
rect 73941 199322 74007 199325
rect 74166 199322 74172 199324
rect 73941 199320 74172 199322
rect 73941 199264 73946 199320
rect 74002 199264 74172 199320
rect 73941 199262 74172 199264
rect 73757 199259 73823 199260
rect 73941 199259 74007 199262
rect 74166 199260 74172 199262
rect 74236 199260 74242 199324
rect 38521 199186 38587 199189
rect 74534 199186 74540 199188
rect 35718 199184 38587 199186
rect 35718 199128 38526 199184
rect 38582 199128 38587 199184
rect 35718 199126 38587 199128
rect 35718 199088 35778 199126
rect 38521 199123 38587 199126
rect 70862 199126 74540 199186
rect 70862 199020 70922 199126
rect 74534 199124 74540 199126
rect 74604 199124 74610 199188
rect 405969 199186 406035 199189
rect 405969 199184 408930 199186
rect 405969 199128 405974 199184
rect 406030 199128 408930 199184
rect 405969 199126 408930 199128
rect 405969 199123 406035 199126
rect 408870 199020 408930 199126
rect 322750 198716 322756 198780
rect 322820 198778 322826 198780
rect 324825 198778 324891 198781
rect 322820 198776 324891 198778
rect 322820 198720 324830 198776
rect 324886 198720 324891 198776
rect 322820 198718 324891 198720
rect 322820 198716 322826 198718
rect 230709 198236 230775 198237
rect 138014 198234 138020 198236
rect 134740 198174 138020 198234
rect 138014 198172 138020 198174
rect 138084 198172 138090 198236
rect 230709 198234 230756 198236
rect 228764 198232 230756 198234
rect 228764 198176 230714 198232
rect 228764 198174 230756 198176
rect 230709 198172 230756 198174
rect 230820 198172 230826 198236
rect 322758 198204 322818 198716
rect 324825 198715 324891 198718
rect 230709 198171 230775 198172
rect 73982 197900 73988 197964
rect 74052 197962 74058 197964
rect 74534 197962 74540 197964
rect 74052 197902 74540 197962
rect 74052 197900 74058 197902
rect 74534 197900 74540 197902
rect 74604 197900 74610 197964
rect 9896 197418 10376 197448
rect 13037 197418 13103 197421
rect 9896 197416 13103 197418
rect 9896 197360 13042 197416
rect 13098 197360 13103 197416
rect 9896 197358 13103 197360
rect 9896 197328 10376 197358
rect 13037 197355 13103 197358
rect 429521 196738 429587 196741
rect 434416 196738 434896 196768
rect 429521 196736 434896 196738
rect 429521 196680 429526 196736
rect 429582 196680 434896 196736
rect 429521 196678 434896 196680
rect 429521 196675 429587 196678
rect 434416 196648 434896 196678
rect 38521 196466 38587 196469
rect 35748 196464 38587 196466
rect 35748 196408 38526 196464
rect 38582 196408 38587 196464
rect 35748 196406 38587 196408
rect 38521 196403 38587 196406
rect 405969 195922 406035 195925
rect 409054 195922 409114 196436
rect 405969 195920 409114 195922
rect 405969 195864 405974 195920
rect 406030 195864 409114 195920
rect 405969 195862 409114 195864
rect 405969 195859 406035 195862
rect 16257 195378 16323 195381
rect 16257 195376 19954 195378
rect 16257 195320 16262 195376
rect 16318 195320 19954 195376
rect 16257 195318 19954 195320
rect 16257 195315 16323 195318
rect 19894 195212 19954 195318
rect 51309 195242 51375 195245
rect 70678 195242 70738 195484
rect 74166 195242 74172 195244
rect 51309 195240 55068 195242
rect 51309 195184 51314 195240
rect 51370 195184 55068 195240
rect 51309 195182 55068 195184
rect 70678 195182 74172 195242
rect 51309 195179 51375 195182
rect 74166 195180 74172 195182
rect 74236 195242 74242 195244
rect 74534 195242 74540 195244
rect 74236 195182 74540 195242
rect 74236 195180 74242 195182
rect 74534 195180 74540 195182
rect 74604 195180 74610 195244
rect 356197 195242 356263 195245
rect 427589 195242 427655 195245
rect 352780 195240 356263 195242
rect 352780 195184 356202 195240
rect 356258 195184 356263 195240
rect 352780 195182 356263 195184
rect 424724 195240 427655 195242
rect 424724 195184 427594 195240
rect 427650 195184 427655 195240
rect 424724 195182 427655 195184
rect 356197 195179 356263 195182
rect 427589 195179 427655 195182
rect 134710 194698 134770 195008
rect 138014 194698 138020 194700
rect 134710 194638 138020 194698
rect 138014 194636 138020 194638
rect 138084 194636 138090 194700
rect 38797 194562 38863 194565
rect 35718 194560 38863 194562
rect 35718 194504 38802 194560
rect 38858 194504 38863 194560
rect 35718 194502 38863 194504
rect 35718 194056 35778 194502
rect 38797 194499 38863 194502
rect 228734 194428 228794 195008
rect 322758 194836 322818 195076
rect 322750 194772 322756 194836
rect 322820 194772 322826 194836
rect 235309 194562 235375 194565
rect 236086 194562 236092 194564
rect 235309 194560 236092 194562
rect 235309 194504 235314 194560
rect 235370 194504 236092 194560
rect 235309 194502 236092 194504
rect 235309 194499 235375 194502
rect 236086 194500 236092 194502
rect 236156 194500 236162 194564
rect 406061 194562 406127 194565
rect 406061 194560 408930 194562
rect 406061 194504 406066 194560
rect 406122 194504 408930 194560
rect 406061 194502 408930 194504
rect 406061 194499 406127 194502
rect 228726 194364 228732 194428
rect 228796 194426 228802 194428
rect 230801 194426 230867 194429
rect 228796 194424 230867 194426
rect 228796 194368 230806 194424
rect 230862 194368 230867 194424
rect 228796 194366 230867 194368
rect 228796 194364 228802 194366
rect 230801 194363 230867 194366
rect 408870 193988 408930 194502
rect 169253 192794 169319 192797
rect 263093 192794 263159 192797
rect 164732 192792 169319 192794
rect 164732 192736 169258 192792
rect 169314 192736 169319 192792
rect 164732 192734 169319 192736
rect 258756 192792 263159 192794
rect 258756 192736 263098 192792
rect 263154 192736 263159 192792
rect 258756 192734 263159 192736
rect 169253 192731 169319 192734
rect 263093 192731 263159 192734
rect 74309 191978 74375 191981
rect 137697 191978 137763 191981
rect 231537 191978 231603 191981
rect 325377 191978 325443 191981
rect 70862 191976 74375 191978
rect 70862 191920 74314 191976
rect 74370 191920 74375 191976
rect 70862 191918 74375 191920
rect 134740 191976 137763 191978
rect 134740 191920 137702 191976
rect 137758 191920 137763 191976
rect 134740 191918 137763 191920
rect 228764 191976 231603 191978
rect 228764 191920 231542 191976
rect 231598 191920 231603 191976
rect 228764 191918 231603 191920
rect 322788 191976 325443 191978
rect 322788 191920 325382 191976
rect 325438 191920 325443 191976
rect 322788 191918 325443 191920
rect 70862 191812 70922 191918
rect 74309 191915 74375 191918
rect 137697 191915 137763 191918
rect 231537 191915 231603 191918
rect 325377 191915 325443 191918
rect 405969 191706 406035 191709
rect 405969 191704 408930 191706
rect 405969 191648 405974 191704
rect 406030 191648 408930 191704
rect 405969 191646 408930 191648
rect 405969 191643 406035 191646
rect 38797 191570 38863 191573
rect 35748 191568 38863 191570
rect 35748 191512 38802 191568
rect 38858 191512 38863 191568
rect 408870 191540 408930 191646
rect 35748 191510 38863 191512
rect 38797 191507 38863 191510
rect 352742 191372 352748 191436
rect 352812 191434 352818 191436
rect 352885 191434 352951 191437
rect 352812 191432 352951 191434
rect 352812 191376 352890 191432
rect 352946 191376 352951 191432
rect 352812 191374 352951 191376
rect 352812 191372 352818 191374
rect 352885 191371 352951 191374
rect 74309 191028 74375 191029
rect 74309 191024 74356 191028
rect 74420 191026 74426 191028
rect 74309 190968 74314 191024
rect 74309 190964 74356 190968
rect 74420 190966 74466 191026
rect 74420 190964 74426 190966
rect 74309 190963 74375 190964
rect 51769 190210 51835 190213
rect 355185 190210 355251 190213
rect 426853 190210 426919 190213
rect 51769 190208 55068 190210
rect 17085 189802 17151 189805
rect 20078 189802 20138 190180
rect 51769 190152 51774 190208
rect 51830 190152 55068 190208
rect 51769 190150 55068 190152
rect 352780 190208 355251 190210
rect 352780 190152 355190 190208
rect 355246 190152 355251 190208
rect 352780 190150 355251 190152
rect 424724 190208 426919 190210
rect 424724 190152 426858 190208
rect 426914 190152 426919 190208
rect 424724 190150 426919 190152
rect 51769 190147 51835 190150
rect 355185 190147 355251 190150
rect 426853 190147 426919 190150
rect 17085 189800 20138 189802
rect 17085 189744 17090 189800
rect 17146 189744 20138 189800
rect 17085 189742 20138 189744
rect 17085 189739 17151 189742
rect 148326 189538 148908 189598
rect 242350 189538 242932 189598
rect 73757 189532 73823 189533
rect 73757 189530 73804 189532
rect 73712 189528 73804 189530
rect 73712 189472 73762 189528
rect 73712 189470 73804 189472
rect 73757 189468 73804 189470
rect 73868 189468 73874 189532
rect 145609 189530 145675 189533
rect 148326 189530 148386 189538
rect 145609 189528 148386 189530
rect 145609 189472 145614 189528
rect 145670 189472 148386 189528
rect 145609 189470 148386 189472
rect 240921 189530 240987 189533
rect 242350 189530 242410 189538
rect 240921 189528 242410 189530
rect 240921 189472 240926 189528
rect 240982 189472 242410 189528
rect 240921 189470 242410 189472
rect 334209 189530 334275 189533
rect 405969 189530 406035 189533
rect 334209 189528 336956 189530
rect 334209 189472 334214 189528
rect 334270 189472 336956 189528
rect 334209 189470 336956 189472
rect 405969 189528 408930 189530
rect 405969 189472 405974 189528
rect 406030 189472 408930 189528
rect 405969 189470 408930 189472
rect 73757 189467 73823 189468
rect 145609 189467 145675 189470
rect 240921 189467 240987 189470
rect 334209 189467 334275 189470
rect 405969 189467 406035 189470
rect 38061 189258 38127 189261
rect 35718 189256 38127 189258
rect 35718 189200 38066 189256
rect 38122 189200 38127 189256
rect 35718 189198 38127 189200
rect 35718 189024 35778 189198
rect 38061 189195 38127 189198
rect 408870 188956 408930 189470
rect 231997 188850 232063 188853
rect 324549 188850 324615 188853
rect 228764 188848 232063 188850
rect 228764 188792 232002 188848
rect 232058 188792 232063 188848
rect 228764 188790 232063 188792
rect 322788 188848 324615 188850
rect 322788 188792 324554 188848
rect 324610 188792 324615 188848
rect 322788 188790 324615 188792
rect 231997 188787 232063 188790
rect 324549 188787 324615 188790
rect 134710 188578 134770 188752
rect 137789 188578 137855 188581
rect 134710 188576 137855 188578
rect 134710 188520 137794 188576
rect 137850 188520 137855 188576
rect 134710 188518 137855 188520
rect 137789 188515 137855 188518
rect 70678 188034 70738 188140
rect 74217 188034 74283 188037
rect 70678 188032 74283 188034
rect 70678 187976 74222 188032
rect 74278 187976 74283 188032
rect 70678 187974 74283 187976
rect 74217 187971 74283 187974
rect 74493 187084 74559 187085
rect 74493 187082 74540 187084
rect 74448 187080 74540 187082
rect 74448 187024 74498 187080
rect 74448 187022 74540 187024
rect 74493 187020 74540 187022
rect 74604 187020 74610 187084
rect 74493 187019 74559 187020
rect 74217 186946 74283 186949
rect 74534 186946 74540 186948
rect 74217 186944 74540 186946
rect 74217 186888 74222 186944
rect 74278 186888 74540 186944
rect 74217 186886 74540 186888
rect 74217 186883 74283 186886
rect 74534 186884 74540 186886
rect 74604 186884 74610 186948
rect 9896 186674 10376 186704
rect 13037 186674 13103 186677
rect 9896 186672 13103 186674
rect 9896 186616 13042 186672
rect 13098 186616 13103 186672
rect 9896 186614 13103 186616
rect 9896 186584 10376 186614
rect 13037 186611 13103 186614
rect 38061 186538 38127 186541
rect 35748 186536 38127 186538
rect 35748 186480 38066 186536
rect 38122 186480 38127 186536
rect 35748 186478 38127 186480
rect 38061 186475 38127 186478
rect 81669 186266 81735 186269
rect 178913 186266 178979 186269
rect 272937 186266 273003 186269
rect 81669 186264 85060 186266
rect 81669 186208 81674 186264
rect 81730 186208 85060 186264
rect 81669 186206 85060 186208
rect 178900 186264 178979 186266
rect 178900 186208 178918 186264
rect 178974 186208 178979 186264
rect 178900 186206 178979 186208
rect 272924 186264 273003 186266
rect 272924 186208 272942 186264
rect 272998 186208 273003 186264
rect 272924 186206 273003 186208
rect 81669 186203 81735 186206
rect 178913 186203 178979 186206
rect 272937 186203 273003 186206
rect 405969 186266 406035 186269
rect 409054 186266 409114 186508
rect 405969 186264 409114 186266
rect 405969 186208 405974 186264
rect 406030 186208 409114 186264
rect 405969 186206 409114 186208
rect 405969 186203 406035 186206
rect 137605 185722 137671 185725
rect 231353 185722 231419 185725
rect 325285 185722 325351 185725
rect 134740 185720 137671 185722
rect 134740 185664 137610 185720
rect 137666 185664 137671 185720
rect 134740 185662 137671 185664
rect 228764 185720 231419 185722
rect 228764 185664 231358 185720
rect 231414 185664 231419 185720
rect 228764 185662 231419 185664
rect 322788 185720 325351 185722
rect 322788 185664 325290 185720
rect 325346 185664 325351 185720
rect 322788 185662 325351 185664
rect 137605 185659 137671 185662
rect 231353 185659 231419 185662
rect 325285 185659 325351 185662
rect 427681 185450 427747 185453
rect 424694 185448 427747 185450
rect 424694 185392 427686 185448
rect 427742 185392 427747 185448
rect 424694 185390 427747 185392
rect 424694 185352 424754 185390
rect 427681 185387 427747 185390
rect 51401 185314 51467 185317
rect 356197 185314 356263 185317
rect 51401 185312 55068 185314
rect 16073 184226 16139 184229
rect 20078 184226 20138 185284
rect 51401 185256 51406 185312
rect 51462 185256 55068 185312
rect 51401 185254 55068 185256
rect 352780 185312 356263 185314
rect 352780 185256 356202 185312
rect 356258 185256 356263 185312
rect 352780 185254 356263 185256
rect 51401 185251 51467 185254
rect 356197 185251 356263 185254
rect 74033 185178 74099 185181
rect 70862 185176 74099 185178
rect 70862 185120 74038 185176
rect 74094 185120 74099 185176
rect 70862 185118 74099 185120
rect 70862 184604 70922 185118
rect 74033 185115 74099 185118
rect 429337 184634 429403 184637
rect 434416 184634 434896 184664
rect 429337 184632 434896 184634
rect 429337 184576 429342 184632
rect 429398 184576 434896 184632
rect 429337 184574 434896 184576
rect 429337 184571 429403 184574
rect 434416 184544 434896 184574
rect 16073 184224 20138 184226
rect 16073 184168 16078 184224
rect 16134 184168 20138 184224
rect 16073 184166 20138 184168
rect 16073 184163 16139 184166
rect 38797 184090 38863 184093
rect 35748 184088 38863 184090
rect 35748 184032 38802 184088
rect 38858 184032 38863 184088
rect 35748 184030 38863 184032
rect 38797 184027 38863 184030
rect 351638 184028 351644 184092
rect 351708 184090 351714 184092
rect 352793 184090 352859 184093
rect 351708 184088 352859 184090
rect 351708 184032 352798 184088
rect 352854 184032 352859 184088
rect 351708 184030 352859 184032
rect 351708 184028 351714 184030
rect 352793 184027 352859 184030
rect 405969 183954 406035 183957
rect 409054 183954 409114 184060
rect 405969 183952 409114 183954
rect 405969 183896 405974 183952
rect 406030 183896 409114 183952
rect 405969 183894 409114 183896
rect 405969 183891 406035 183894
rect 242526 183076 242532 183140
rect 242596 183138 242602 183140
rect 248925 183138 248991 183141
rect 242596 183136 248991 183138
rect 242596 183080 248930 183136
rect 248986 183080 248991 183136
rect 242596 183078 248991 183080
rect 242596 183076 242602 183078
rect 248925 183075 248991 183078
rect 137881 182594 137947 182597
rect 231445 182594 231511 182597
rect 325469 182594 325535 182597
rect 134740 182592 137947 182594
rect 134740 182536 137886 182592
rect 137942 182536 137947 182592
rect 134740 182534 137947 182536
rect 228764 182592 231511 182594
rect 228764 182536 231450 182592
rect 231506 182536 231511 182592
rect 228764 182534 231511 182536
rect 322788 182592 325535 182594
rect 322788 182536 325474 182592
rect 325530 182536 325535 182592
rect 322788 182534 325535 182536
rect 137881 182531 137947 182534
rect 231445 182531 231511 182534
rect 325469 182531 325535 182534
rect 249017 182186 249083 182189
rect 271414 182186 271420 182188
rect 249017 182184 271420 182186
rect 249017 182128 249022 182184
rect 249078 182128 271420 182184
rect 249017 182126 271420 182128
rect 249017 182123 249083 182126
rect 271414 182124 271420 182126
rect 271484 182124 271490 182188
rect 323118 182124 323124 182188
rect 323188 182186 323194 182188
rect 352885 182186 352951 182189
rect 323188 182184 352951 182186
rect 323188 182128 352890 182184
rect 352946 182128 352951 182184
rect 323188 182126 352951 182128
rect 323188 182124 323194 182126
rect 352885 182123 352951 182126
rect 154717 182050 154783 182053
rect 174814 182050 174820 182052
rect 154717 182048 174820 182050
rect 154717 181992 154722 182048
rect 154778 181992 174820 182048
rect 154717 181990 174820 181992
rect 154717 181987 154783 181990
rect 174814 181988 174820 181990
rect 174884 181988 174890 182052
rect 228726 181988 228732 182052
rect 228796 182050 228802 182052
rect 261069 182050 261135 182053
rect 228796 182048 261135 182050
rect 228796 181992 261074 182048
rect 261130 181992 261135 182048
rect 228796 181990 261135 181992
rect 228796 181988 228802 181990
rect 261069 181987 261135 181990
rect 323486 181988 323492 182052
rect 323556 182050 323562 182052
rect 352977 182050 353043 182053
rect 323556 182048 353043 182050
rect 323556 181992 352982 182048
rect 353038 181992 353043 182048
rect 323556 181990 353043 181992
rect 323556 181988 323562 181990
rect 352977 181987 353043 181990
rect 74401 181236 74467 181237
rect 74350 181172 74356 181236
rect 74420 181234 74467 181236
rect 74420 181232 74512 181234
rect 74462 181176 74512 181232
rect 74420 181174 74512 181176
rect 74420 181172 74467 181174
rect 147030 181172 147036 181236
rect 147100 181234 147106 181236
rect 155269 181234 155335 181237
rect 267509 181236 267575 181237
rect 267509 181234 267556 181236
rect 147100 181232 155335 181234
rect 147100 181176 155274 181232
rect 155330 181176 155335 181232
rect 147100 181174 155335 181176
rect 267464 181232 267556 181234
rect 267464 181176 267514 181232
rect 267464 181174 267556 181176
rect 147100 181172 147106 181174
rect 74401 181171 74467 181172
rect 155269 181171 155335 181174
rect 267509 181172 267556 181174
rect 267620 181172 267626 181236
rect 267509 181171 267575 181172
rect 158397 181098 158463 181101
rect 168558 181098 168564 181100
rect 158397 181096 168564 181098
rect 158397 181040 158402 181096
rect 158458 181040 168564 181096
rect 158397 181038 168564 181040
rect 158397 181035 158463 181038
rect 168558 181036 168564 181038
rect 168628 181036 168634 181100
rect 157201 180962 157267 180965
rect 167822 180962 167828 180964
rect 157201 180960 167828 180962
rect 157201 180904 157206 180960
rect 157262 180904 167828 180960
rect 157201 180902 167828 180904
rect 157201 180899 157267 180902
rect 167822 180900 167828 180902
rect 167892 180900 167898 180964
rect 157753 180826 157819 180829
rect 169294 180826 169300 180828
rect 157753 180824 169300 180826
rect 157753 180768 157758 180824
rect 157814 180768 169300 180824
rect 157753 180766 169300 180768
rect 157753 180763 157819 180766
rect 169294 180764 169300 180766
rect 169364 180764 169370 180828
rect 253341 180826 253407 180829
rect 261662 180826 261668 180828
rect 253341 180824 261668 180826
rect 253341 180768 253346 180824
rect 253402 180768 261668 180824
rect 253341 180766 261668 180768
rect 253341 180763 253407 180766
rect 261662 180764 261668 180766
rect 261732 180764 261738 180828
rect 156557 180690 156623 180693
rect 167638 180690 167644 180692
rect 156557 180688 167644 180690
rect 156557 180632 156562 180688
rect 156618 180632 167644 180688
rect 156557 180630 167644 180632
rect 156557 180627 156623 180630
rect 167638 180628 167644 180630
rect 167708 180628 167714 180692
rect 252697 180690 252763 180693
rect 262398 180690 262404 180692
rect 252697 180688 262404 180690
rect 252697 180632 252702 180688
rect 252758 180632 262404 180688
rect 252697 180630 262404 180632
rect 252697 180627 252763 180630
rect 262398 180628 262404 180630
rect 262468 180628 262474 180692
rect 141510 180492 141516 180556
rect 141580 180554 141586 180556
rect 159041 180554 159107 180557
rect 141580 180552 159107 180554
rect 141580 180496 159046 180552
rect 159102 180496 159107 180552
rect 141580 180494 159107 180496
rect 141580 180492 141586 180494
rect 159041 180491 159107 180494
rect 252053 180554 252119 180557
rect 262950 180554 262956 180556
rect 252053 180552 262956 180554
rect 252053 180496 252058 180552
rect 252114 180496 262956 180552
rect 252053 180494 262956 180496
rect 252053 180491 252119 180494
rect 262950 180492 262956 180494
rect 263020 180492 263026 180556
rect 242342 180220 242348 180284
rect 242412 180282 242418 180284
rect 250857 180282 250923 180285
rect 242412 180280 250923 180282
rect 242412 180224 250862 180280
rect 250918 180224 250923 180280
rect 242412 180222 250923 180224
rect 242412 180220 242418 180222
rect 250857 180219 250923 180222
rect 241790 180084 241796 180148
rect 241860 180146 241866 180148
rect 250213 180146 250279 180149
rect 241860 180144 250279 180146
rect 241860 180088 250218 180144
rect 250274 180088 250279 180144
rect 241860 180086 250279 180088
rect 241860 180084 241866 180086
rect 250213 180083 250279 180086
rect 73757 180012 73823 180013
rect 73757 180008 73804 180012
rect 73868 180010 73874 180012
rect 73757 179952 73762 180008
rect 73757 179948 73804 179952
rect 73868 179950 73914 180010
rect 73868 179948 73874 179950
rect 74166 179948 74172 180012
rect 74236 180010 74242 180012
rect 74493 180010 74559 180013
rect 74236 180008 74559 180010
rect 74236 179952 74498 180008
rect 74554 179952 74559 180008
rect 74236 179950 74559 179952
rect 74236 179948 74242 179950
rect 73757 179947 73823 179948
rect 74493 179947 74559 179950
rect 148737 180010 148803 180013
rect 155913 180010 155979 180013
rect 148737 180008 155979 180010
rect 148737 179952 148742 180008
rect 148798 179952 155918 180008
rect 155974 179952 155979 180008
rect 148737 179950 155979 179952
rect 148737 179947 148803 179950
rect 155913 179947 155979 179950
rect 242526 179948 242532 180012
rect 242596 180010 242602 180012
rect 249569 180010 249635 180013
rect 242596 180008 249635 180010
rect 242596 179952 249574 180008
rect 249630 179952 249635 180008
rect 242596 179950 249635 179952
rect 242596 179948 242602 179950
rect 249569 179947 249635 179950
rect 138893 179466 138959 179469
rect 230985 179466 231051 179469
rect 324549 179466 324615 179469
rect 134740 179464 138959 179466
rect 134740 179408 138898 179464
rect 138954 179408 138959 179464
rect 134740 179406 138959 179408
rect 228764 179464 231051 179466
rect 228764 179408 230990 179464
rect 231046 179408 231051 179464
rect 228764 179406 231051 179408
rect 322788 179464 324615 179466
rect 322788 179408 324554 179464
rect 324610 179408 324615 179464
rect 322788 179406 324615 179408
rect 138893 179403 138959 179406
rect 230985 179403 231051 179406
rect 324549 179403 324615 179406
rect 309870 179268 309876 179332
rect 309940 179330 309946 179332
rect 312630 179330 312636 179332
rect 309940 179270 312636 179330
rect 309940 179268 309946 179270
rect 312630 179268 312636 179270
rect 312700 179268 312706 179332
rect 311158 179132 311164 179196
rect 311228 179194 311234 179196
rect 313734 179194 313740 179196
rect 311228 179134 313740 179194
rect 311228 179132 311234 179134
rect 313734 179132 313740 179134
rect 313804 179132 313810 179196
rect 9896 175794 10376 175824
rect 13037 175794 13103 175797
rect 9896 175792 13103 175794
rect 9896 175736 13042 175792
rect 13098 175736 13103 175792
rect 9896 175734 13103 175736
rect 9896 175704 10376 175734
rect 13037 175731 13103 175734
rect 74534 175732 74540 175796
rect 74604 175794 74610 175796
rect 75086 175794 75092 175796
rect 74604 175734 75092 175794
rect 74604 175732 74610 175734
rect 75086 175732 75092 175734
rect 75156 175732 75162 175796
rect 218013 175522 218079 175525
rect 219710 175522 219716 175524
rect 218013 175520 219716 175522
rect 218013 175464 218018 175520
rect 218074 175464 219716 175520
rect 218013 175462 219716 175464
rect 218013 175459 218079 175462
rect 219710 175460 219716 175462
rect 219780 175460 219786 175524
rect 182961 174980 183027 174981
rect 182910 174978 182916 174980
rect 182870 174918 182916 174978
rect 182980 174976 183027 174980
rect 183022 174920 183027 174976
rect 182910 174916 182916 174918
rect 182980 174916 183027 174920
rect 182961 174915 183027 174916
rect 241790 173964 241796 174028
rect 241860 174026 241866 174028
rect 242526 174026 242532 174028
rect 241860 173966 242532 174026
rect 241860 173964 241866 173966
rect 242526 173964 242532 173966
rect 242596 173964 242602 174028
rect 148737 173076 148803 173077
rect 148686 173074 148692 173076
rect 148646 173014 148692 173074
rect 148756 173072 148803 173076
rect 148798 173016 148803 173072
rect 148686 173012 148692 173014
rect 148756 173012 148803 173016
rect 148737 173011 148803 173012
rect 55541 172940 55607 172941
rect 55541 172938 55588 172940
rect 55496 172936 55588 172938
rect 55496 172880 55546 172936
rect 55496 172878 55588 172880
rect 55541 172876 55588 172878
rect 55652 172876 55658 172940
rect 169294 172876 169300 172940
rect 169364 172876 169370 172940
rect 350953 172938 351019 172941
rect 351638 172938 351644 172940
rect 350953 172936 351644 172938
rect 350953 172880 350958 172936
rect 351014 172880 351644 172936
rect 350953 172878 351644 172880
rect 55541 172875 55607 172876
rect 55398 172740 55404 172804
rect 55468 172802 55474 172804
rect 56553 172802 56619 172805
rect 55468 172800 56619 172802
rect 55468 172744 56558 172800
rect 56614 172744 56619 172800
rect 55468 172742 56619 172744
rect 55468 172740 55474 172742
rect 56553 172739 56619 172742
rect 168742 172740 168748 172804
rect 168812 172802 168818 172804
rect 169302 172802 169362 172876
rect 350953 172875 351019 172878
rect 351638 172876 351644 172878
rect 351708 172876 351714 172940
rect 351822 172876 351828 172940
rect 351892 172938 351898 172940
rect 352057 172938 352123 172941
rect 351892 172936 352123 172938
rect 351892 172880 352062 172936
rect 352118 172880 352123 172936
rect 351892 172878 352123 172880
rect 351892 172876 351898 172878
rect 352057 172875 352123 172878
rect 168812 172742 169362 172802
rect 168812 172740 168818 172742
rect 429889 172530 429955 172533
rect 434416 172530 434896 172560
rect 429889 172528 434896 172530
rect 429889 172472 429894 172528
rect 429950 172472 434896 172528
rect 429889 172470 434896 172472
rect 429889 172467 429955 172470
rect 434416 172440 434896 172470
rect 52638 171652 52644 171716
rect 52708 171714 52714 171716
rect 53517 171714 53583 171717
rect 52708 171712 53583 171714
rect 52708 171656 53522 171712
rect 53578 171656 53583 171712
rect 52708 171654 53583 171656
rect 52708 171652 52714 171654
rect 53517 171651 53583 171654
rect 54529 171714 54595 171717
rect 74401 171716 74467 171717
rect 54662 171714 54668 171716
rect 54529 171712 54668 171714
rect 54529 171656 54534 171712
rect 54590 171656 54668 171712
rect 54529 171654 54668 171656
rect 54529 171651 54595 171654
rect 54662 171652 54668 171654
rect 54732 171652 54738 171716
rect 74350 171714 74356 171716
rect 74310 171654 74356 171714
rect 74420 171712 74467 171716
rect 74462 171656 74467 171712
rect 74350 171652 74356 171654
rect 74420 171652 74467 171656
rect 74401 171651 74467 171652
rect 72653 169810 72719 169813
rect 75638 169810 75644 169812
rect 72653 169808 75644 169810
rect 72653 169752 72658 169808
rect 72714 169752 75644 169808
rect 72653 169750 75644 169752
rect 72653 169747 72719 169750
rect 75638 169748 75644 169750
rect 75708 169748 75714 169812
rect 73982 169612 73988 169676
rect 74052 169674 74058 169676
rect 75454 169674 75460 169676
rect 74052 169614 75460 169674
rect 74052 169612 74058 169614
rect 75454 169612 75460 169614
rect 75524 169612 75530 169676
rect 73481 169540 73547 169541
rect 73430 169476 73436 169540
rect 73500 169538 73547 169540
rect 76006 169538 76012 169540
rect 73500 169536 76012 169538
rect 73542 169480 76012 169536
rect 73500 169478 76012 169480
rect 73500 169476 73547 169478
rect 76006 169476 76012 169478
rect 76076 169476 76082 169540
rect 237374 169476 237380 169540
rect 237444 169538 237450 169540
rect 243446 169538 243452 169540
rect 237444 169478 243452 169538
rect 237444 169476 237450 169478
rect 243446 169476 243452 169478
rect 243516 169476 243522 169540
rect 73481 169475 73547 169476
rect 73798 169204 73804 169268
rect 73868 169266 73874 169268
rect 74718 169266 74724 169268
rect 73868 169206 74724 169266
rect 73868 169204 73874 169206
rect 74718 169204 74724 169206
rect 74788 169204 74794 169268
rect 144086 169204 144092 169268
rect 144156 169266 144162 169268
rect 148686 169266 148692 169268
rect 144156 169206 148692 169266
rect 144156 169204 144162 169206
rect 148686 169204 148692 169206
rect 148756 169204 148762 169268
rect 238110 169204 238116 169268
rect 238180 169266 238186 169268
rect 242342 169266 242348 169268
rect 238180 169206 242348 169266
rect 238180 169204 238186 169206
rect 242342 169204 242348 169206
rect 242412 169204 242418 169268
rect 242526 169204 242532 169268
rect 242596 169266 242602 169268
rect 247126 169266 247132 169268
rect 242596 169206 247132 169266
rect 242596 169204 242602 169206
rect 247126 169204 247132 169206
rect 247196 169204 247202 169268
rect 79185 169130 79251 169133
rect 76780 169128 79251 169130
rect 76780 169072 79190 169128
rect 79246 169072 79251 169128
rect 76780 169070 79251 169072
rect 79185 169067 79251 169070
rect 140549 169130 140615 169133
rect 173577 169130 173643 169133
rect 140549 169128 143020 169130
rect 140549 169072 140554 169128
rect 140610 169072 143020 169128
rect 140549 169070 143020 169072
rect 170804 169128 173643 169130
rect 170804 169072 173582 169128
rect 173638 169072 173643 169128
rect 170804 169070 173643 169072
rect 140549 169067 140615 169070
rect 173577 169067 173643 169070
rect 233469 169130 233535 169133
rect 267417 169130 267483 169133
rect 233469 169128 237044 169130
rect 233469 169072 233474 169128
rect 233530 169072 237044 169128
rect 233469 169070 237044 169072
rect 264828 169128 267483 169130
rect 264828 169072 267422 169128
rect 267478 169072 267483 169128
rect 264828 169070 267483 169072
rect 233469 169067 233535 169070
rect 267417 169067 267483 169070
rect 328413 169130 328479 169133
rect 328413 169128 331068 169130
rect 328413 169072 328418 169128
rect 328474 169072 331068 169128
rect 328413 169070 331068 169072
rect 328413 169067 328479 169070
rect 49193 168858 49259 168861
rect 49150 168856 49259 168858
rect 49150 168800 49198 168856
rect 49254 168800 49259 168856
rect 49150 168795 49259 168800
rect 49150 168284 49210 168795
rect 360429 168314 360495 168317
rect 361165 168314 361231 168317
rect 358852 168312 361231 168314
rect 358852 168256 360434 168312
rect 360490 168256 361170 168312
rect 361226 168256 361231 168312
rect 358852 168254 361231 168256
rect 360429 168251 360495 168254
rect 361165 168251 361231 168254
rect 140549 167770 140615 167773
rect 173485 167770 173551 167773
rect 140549 167768 143020 167770
rect 140549 167712 140554 167768
rect 140610 167712 143020 167768
rect 140549 167710 143020 167712
rect 170804 167768 173551 167770
rect 170804 167712 173490 167768
rect 173546 167712 173551 167768
rect 170804 167710 173551 167712
rect 140549 167707 140615 167710
rect 173485 167707 173551 167710
rect 233469 167770 233535 167773
rect 267601 167770 267667 167773
rect 233469 167768 237044 167770
rect 233469 167712 233474 167768
rect 233530 167712 237044 167768
rect 233469 167710 237044 167712
rect 264828 167768 267667 167770
rect 264828 167712 267606 167768
rect 267662 167712 267667 167768
rect 264828 167710 267667 167712
rect 233469 167707 233535 167710
rect 267601 167707 267667 167710
rect 327217 167770 327283 167773
rect 327217 167768 331068 167770
rect 327217 167712 327222 167768
rect 327278 167712 331068 167768
rect 327217 167710 331068 167712
rect 327217 167707 327283 167710
rect 77253 167702 77319 167705
rect 76780 167700 77319 167702
rect 76780 167644 77258 167700
rect 77314 167644 77319 167700
rect 76780 167642 77319 167644
rect 77253 167639 77319 167642
rect 140549 166410 140615 166413
rect 173393 166410 173459 166413
rect 140549 166408 143020 166410
rect 140549 166352 140554 166408
rect 140610 166352 143020 166408
rect 140549 166350 143020 166352
rect 170804 166408 173459 166410
rect 170804 166352 173398 166408
rect 173454 166352 173459 166408
rect 170804 166350 173459 166352
rect 140549 166347 140615 166350
rect 173393 166347 173459 166350
rect 233469 166410 233535 166413
rect 267509 166410 267575 166413
rect 233469 166408 237044 166410
rect 233469 166352 233474 166408
rect 233530 166352 237044 166408
rect 233469 166350 237044 166352
rect 264828 166408 267575 166410
rect 264828 166352 267514 166408
rect 267570 166352 267575 166408
rect 264828 166350 267575 166352
rect 233469 166347 233535 166350
rect 267509 166347 267575 166350
rect 327493 166410 327559 166413
rect 327493 166408 331068 166410
rect 327493 166352 327498 166408
rect 327554 166352 331068 166408
rect 327493 166350 331068 166352
rect 327493 166347 327559 166350
rect 77253 166342 77319 166345
rect 76780 166340 77319 166342
rect 76780 166284 77258 166340
rect 77314 166284 77319 166340
rect 76780 166282 77319 166284
rect 77253 166279 77319 166282
rect 46893 165186 46959 165189
rect 360521 165186 360587 165189
rect 361717 165186 361783 165189
rect 46893 165184 48996 165186
rect 46893 165128 46898 165184
rect 46954 165128 48996 165184
rect 46893 165126 48996 165128
rect 358852 165184 361783 165186
rect 358852 165128 360526 165184
rect 360582 165128 361722 165184
rect 361778 165128 361783 165184
rect 358852 165126 361783 165128
rect 46893 165123 46959 165126
rect 360521 165123 360587 165126
rect 361717 165123 361783 165126
rect 9896 165050 10376 165080
rect 13405 165050 13471 165053
rect 9896 165048 13471 165050
rect 9896 164992 13410 165048
rect 13466 164992 13471 165048
rect 9896 164990 13471 164992
rect 9896 164960 10376 164990
rect 13405 164987 13471 164990
rect 139629 164914 139695 164917
rect 172933 164914 172999 164917
rect 139629 164912 143020 164914
rect 139629 164856 139634 164912
rect 139690 164856 143020 164912
rect 139629 164854 143020 164856
rect 170804 164912 172999 164914
rect 170804 164856 172938 164912
rect 172994 164856 172999 164912
rect 170804 164854 172999 164856
rect 139629 164851 139695 164854
rect 172933 164851 172999 164854
rect 233469 164914 233535 164917
rect 267141 164914 267207 164917
rect 233469 164912 237044 164914
rect 233469 164856 233474 164912
rect 233530 164856 237044 164912
rect 233469 164854 237044 164856
rect 264828 164912 267207 164914
rect 264828 164856 267146 164912
rect 267202 164856 267207 164912
rect 264828 164854 267207 164856
rect 233469 164851 233535 164854
rect 267141 164851 267207 164854
rect 328413 164914 328479 164917
rect 328413 164912 331068 164914
rect 328413 164856 328418 164912
rect 328474 164856 331068 164912
rect 328413 164854 331068 164856
rect 328413 164851 328479 164854
rect 77253 164846 77319 164849
rect 76780 164844 77319 164846
rect 76780 164788 77258 164844
rect 77314 164788 77319 164844
rect 76780 164786 77319 164788
rect 77253 164783 77319 164786
rect 87189 164098 87255 164101
rect 87189 164096 90058 164098
rect 87189 164040 87194 164096
rect 87250 164040 90058 164096
rect 87189 164038 90058 164040
rect 87189 164035 87255 164038
rect 77253 163486 77319 163489
rect 76780 163484 77319 163486
rect 76780 163428 77258 163484
rect 77314 163428 77319 163484
rect 89998 163456 90058 164038
rect 139629 163554 139695 163557
rect 173117 163554 173183 163557
rect 139629 163552 143020 163554
rect 139629 163496 139634 163552
rect 139690 163496 143020 163552
rect 139629 163494 143020 163496
rect 170804 163552 173183 163554
rect 170804 163496 173122 163552
rect 173178 163496 173183 163552
rect 170804 163494 173183 163496
rect 139629 163491 139695 163494
rect 173117 163491 173183 163494
rect 233469 163554 233535 163557
rect 267877 163554 267943 163557
rect 233469 163552 237044 163554
rect 233469 163496 233474 163552
rect 233530 163496 237044 163552
rect 233469 163494 237044 163496
rect 264828 163552 267943 163554
rect 264828 163496 267882 163552
rect 267938 163496 267943 163552
rect 264828 163494 267943 163496
rect 233469 163491 233535 163494
rect 267877 163491 267943 163494
rect 76780 163426 77319 163428
rect 77253 163423 77319 163426
rect 330486 163426 331068 163486
rect 131349 163418 131415 163421
rect 129772 163416 131415 163418
rect 129772 163360 131354 163416
rect 131410 163360 131415 163416
rect 129772 163358 131415 163360
rect 131349 163355 131415 163358
rect 181765 163418 181831 163421
rect 226293 163418 226359 163421
rect 181765 163416 184052 163418
rect 181765 163360 181770 163416
rect 181826 163360 184052 163416
rect 181765 163358 184052 163360
rect 223796 163416 226359 163418
rect 223796 163360 226298 163416
rect 226354 163360 226359 163416
rect 223796 163358 226359 163360
rect 181765 163355 181831 163358
rect 226293 163355 226359 163358
rect 274869 163418 274935 163421
rect 321605 163418 321671 163421
rect 274869 163416 278076 163418
rect 274869 163360 274874 163416
rect 274930 163360 278076 163416
rect 274869 163358 278076 163360
rect 317820 163416 321671 163418
rect 317820 163360 321610 163416
rect 321666 163360 321671 163416
rect 317820 163358 321671 163360
rect 274869 163355 274935 163358
rect 321605 163355 321671 163358
rect 327217 163418 327283 163421
rect 330486 163418 330546 163426
rect 327217 163416 330546 163418
rect 327217 163360 327222 163416
rect 327278 163360 330546 163416
rect 327217 163358 330546 163360
rect 327217 163355 327283 163358
rect 87097 163146 87163 163149
rect 87097 163144 90058 163146
rect 87097 163088 87102 163144
rect 87158 163088 90058 163144
rect 87097 163086 90058 163088
rect 87097 163083 87163 163086
rect 46617 162602 46683 162605
rect 46617 162600 49210 162602
rect 46617 162544 46622 162600
rect 46678 162544 49210 162600
rect 46617 162542 49210 162544
rect 46617 162539 46683 162542
rect 49150 162332 49210 162542
rect 89998 162504 90058 163086
rect 131993 162466 132059 162469
rect 129772 162464 132059 162466
rect 129772 162408 131998 162464
rect 132054 162408 132059 162464
rect 129772 162406 132059 162408
rect 131993 162403 132059 162406
rect 181305 162466 181371 162469
rect 226201 162466 226267 162469
rect 181305 162464 184052 162466
rect 181305 162408 181310 162464
rect 181366 162408 184052 162464
rect 181305 162406 184052 162408
rect 223796 162464 226267 162466
rect 223796 162408 226206 162464
rect 226262 162408 226267 162464
rect 223796 162406 226267 162408
rect 181305 162403 181371 162406
rect 226201 162403 226267 162406
rect 275053 162466 275119 162469
rect 321605 162466 321671 162469
rect 275053 162464 278076 162466
rect 275053 162408 275058 162464
rect 275114 162408 278076 162464
rect 275053 162406 278076 162408
rect 317820 162464 321671 162466
rect 317820 162408 321610 162464
rect 321666 162408 321671 162464
rect 317820 162406 321671 162408
rect 275053 162403 275119 162406
rect 321605 162403 321671 162406
rect 49142 162330 49148 162332
rect 49020 162270 49148 162330
rect 49142 162268 49148 162270
rect 49212 162268 49218 162332
rect 49150 162028 49210 162268
rect 139629 162194 139695 162197
rect 173761 162194 173827 162197
rect 139629 162192 143020 162194
rect 139629 162136 139634 162192
rect 139690 162136 143020 162192
rect 139629 162134 143020 162136
rect 170804 162192 173827 162194
rect 170804 162136 173766 162192
rect 173822 162136 173827 162192
rect 170804 162134 173827 162136
rect 139629 162131 139695 162134
rect 173761 162131 173827 162134
rect 233469 162194 233535 162197
rect 267049 162194 267115 162197
rect 233469 162192 237044 162194
rect 233469 162136 233474 162192
rect 233530 162136 237044 162192
rect 233469 162134 237044 162136
rect 264828 162192 267115 162194
rect 264828 162136 267054 162192
rect 267110 162136 267115 162192
rect 264828 162134 267115 162136
rect 233469 162131 233535 162134
rect 267049 162131 267115 162134
rect 327309 162194 327375 162197
rect 327309 162192 331068 162194
rect 327309 162136 327314 162192
rect 327370 162136 331068 162192
rect 327309 162134 331068 162136
rect 327309 162131 327375 162134
rect 77253 162126 77319 162129
rect 76780 162124 77319 162126
rect 76780 162068 77258 162124
rect 77314 162068 77319 162124
rect 76780 162066 77319 162068
rect 77253 162063 77319 162066
rect 360613 162058 360679 162061
rect 361717 162058 361783 162061
rect 358852 162056 361783 162058
rect 358852 162000 360618 162056
rect 360674 162000 361722 162056
rect 361778 162000 361783 162056
rect 358852 161998 361783 162000
rect 360613 161995 360679 161998
rect 361717 161995 361783 161998
rect 87281 161922 87347 161925
rect 87281 161920 90058 161922
rect 87281 161864 87286 161920
rect 87342 161864 90058 161920
rect 87281 161862 90058 161864
rect 87281 161859 87347 161862
rect 89998 161688 90058 161862
rect 131441 161650 131507 161653
rect 226293 161650 226359 161653
rect 129772 161648 131507 161650
rect 129772 161592 131446 161648
rect 131502 161592 131507 161648
rect 223796 161648 226359 161650
rect 129772 161590 131507 161592
rect 131441 161587 131507 161590
rect 87189 161378 87255 161381
rect 87189 161376 90058 161378
rect 87189 161320 87194 161376
rect 87250 161320 90058 161376
rect 87189 161318 90058 161320
rect 87189 161315 87255 161318
rect 89998 160736 90058 161318
rect 180293 160970 180359 160973
rect 184022 160970 184082 161620
rect 223796 161592 226298 161648
rect 226354 161592 226359 161648
rect 223796 161590 226359 161592
rect 226293 161587 226359 161590
rect 275145 161650 275211 161653
rect 321605 161650 321671 161653
rect 275145 161648 278076 161650
rect 275145 161592 275150 161648
rect 275206 161592 278076 161648
rect 275145 161590 278076 161592
rect 317820 161648 321671 161650
rect 317820 161592 321610 161648
rect 321666 161592 321671 161648
rect 317820 161590 321671 161592
rect 275145 161587 275211 161590
rect 321605 161587 321671 161590
rect 180293 160968 184082 160970
rect 180293 160912 180298 160968
rect 180354 160912 184082 160968
rect 180293 160910 184082 160912
rect 180293 160907 180359 160910
rect 131349 160698 131415 160701
rect 129772 160696 131415 160698
rect 129772 160640 131354 160696
rect 131410 160640 131415 160696
rect 129772 160638 131415 160640
rect 131349 160635 131415 160638
rect 140641 160698 140707 160701
rect 174037 160698 174103 160701
rect 140641 160696 143020 160698
rect 140641 160640 140646 160696
rect 140702 160640 143020 160696
rect 140641 160638 143020 160640
rect 170804 160696 174103 160698
rect 170804 160640 174042 160696
rect 174098 160640 174103 160696
rect 170804 160638 174103 160640
rect 140641 160635 140707 160638
rect 174037 160635 174103 160638
rect 182317 160698 182383 160701
rect 225741 160698 225807 160701
rect 182317 160696 184052 160698
rect 182317 160640 182322 160696
rect 182378 160640 184052 160696
rect 182317 160638 184052 160640
rect 223796 160696 225807 160698
rect 223796 160640 225746 160696
rect 225802 160640 225807 160696
rect 223796 160638 225807 160640
rect 182317 160635 182383 160638
rect 225741 160635 225807 160638
rect 232733 160698 232799 160701
rect 266589 160698 266655 160701
rect 232733 160696 237044 160698
rect 232733 160640 232738 160696
rect 232794 160640 237044 160696
rect 232733 160638 237044 160640
rect 264828 160696 266655 160698
rect 264828 160640 266594 160696
rect 266650 160640 266655 160696
rect 264828 160638 266655 160640
rect 232733 160635 232799 160638
rect 266589 160635 266655 160638
rect 275789 160698 275855 160701
rect 321053 160698 321119 160701
rect 275789 160696 278076 160698
rect 275789 160640 275794 160696
rect 275850 160640 278076 160696
rect 275789 160638 278076 160640
rect 317820 160696 321119 160698
rect 317820 160640 321058 160696
rect 321114 160640 321119 160696
rect 317820 160638 321119 160640
rect 275789 160635 275855 160638
rect 321053 160635 321119 160638
rect 327401 160698 327467 160701
rect 327401 160696 331068 160698
rect 327401 160640 327406 160696
rect 327462 160640 331068 160696
rect 327401 160638 331068 160640
rect 327401 160635 327467 160638
rect 76750 160018 76810 160600
rect 87189 160426 87255 160429
rect 87189 160424 90058 160426
rect 87189 160368 87194 160424
rect 87250 160368 90058 160424
rect 87189 160366 90058 160368
rect 87189 160363 87255 160366
rect 81761 160018 81827 160021
rect 76750 160016 81827 160018
rect 76750 159960 81766 160016
rect 81822 159960 81827 160016
rect 76750 159958 81827 159960
rect 81761 159955 81827 159958
rect 89998 159920 90058 160366
rect 428785 160290 428851 160293
rect 434416 160290 434896 160320
rect 428785 160288 434896 160290
rect 428785 160232 428790 160288
rect 428846 160232 434896 160288
rect 428785 160230 434896 160232
rect 428785 160227 428851 160230
rect 434416 160200 434896 160230
rect 131349 159882 131415 159885
rect 129772 159880 131415 159882
rect 129772 159824 131354 159880
rect 131410 159824 131415 159880
rect 129772 159822 131415 159824
rect 131349 159819 131415 159822
rect 181673 159882 181739 159885
rect 226109 159882 226175 159885
rect 181673 159880 184052 159882
rect 181673 159824 181678 159880
rect 181734 159824 184052 159880
rect 181673 159822 184052 159824
rect 223796 159880 226175 159882
rect 223796 159824 226114 159880
rect 226170 159824 226175 159880
rect 223796 159822 226175 159824
rect 181673 159819 181739 159822
rect 226109 159819 226175 159822
rect 275145 159882 275211 159885
rect 320593 159882 320659 159885
rect 275145 159880 278076 159882
rect 275145 159824 275150 159880
rect 275206 159824 278076 159880
rect 275145 159822 278076 159824
rect 317820 159880 320659 159882
rect 317820 159824 320598 159880
rect 320654 159824 320659 159880
rect 317820 159822 320659 159824
rect 275145 159819 275211 159822
rect 320593 159819 320659 159822
rect 79277 159338 79343 159341
rect 76780 159336 79343 159338
rect 76780 159280 79282 159336
rect 79338 159280 79343 159336
rect 76780 159278 79343 159280
rect 79277 159275 79343 159278
rect 139629 159338 139695 159341
rect 173669 159338 173735 159341
rect 139629 159336 143020 159338
rect 139629 159280 139634 159336
rect 139690 159280 143020 159336
rect 139629 159278 143020 159280
rect 170804 159336 173735 159338
rect 170804 159280 173674 159336
rect 173730 159280 173735 159336
rect 170804 159278 173735 159280
rect 139629 159275 139695 159278
rect 173669 159275 173735 159278
rect 233469 159338 233535 159341
rect 266589 159338 266655 159341
rect 233469 159336 237044 159338
rect 233469 159280 233474 159336
rect 233530 159280 237044 159336
rect 233469 159278 237044 159280
rect 264828 159336 266655 159338
rect 264828 159280 266594 159336
rect 266650 159280 266655 159336
rect 264828 159278 266655 159280
rect 233469 159275 233535 159278
rect 266589 159275 266655 159278
rect 327217 159338 327283 159341
rect 327217 159336 331068 159338
rect 327217 159280 327222 159336
rect 327278 159280 331068 159336
rect 327217 159278 331068 159280
rect 327217 159275 327283 159278
rect 46525 158930 46591 158933
rect 87189 158930 87255 158933
rect 132177 158930 132243 158933
rect 46525 158928 49180 158930
rect 46525 158872 46530 158928
rect 46586 158900 49180 158928
rect 87189 158928 90028 158930
rect 46586 158872 49210 158900
rect 46525 158870 49210 158872
rect 46525 158867 46591 158870
rect 49150 158388 49210 158870
rect 87189 158872 87194 158928
rect 87250 158872 90028 158928
rect 87189 158870 90028 158872
rect 129772 158928 132243 158930
rect 129772 158872 132182 158928
rect 132238 158872 132243 158928
rect 129772 158870 132243 158872
rect 87189 158867 87255 158870
rect 132177 158867 132243 158870
rect 181397 158930 181463 158933
rect 227213 158930 227279 158933
rect 181397 158928 184052 158930
rect 181397 158872 181402 158928
rect 181458 158872 184052 158928
rect 181397 158870 184052 158872
rect 223796 158928 227279 158930
rect 223796 158872 227218 158928
rect 227274 158872 227279 158928
rect 223796 158870 227279 158872
rect 181397 158867 181463 158870
rect 227213 158867 227279 158870
rect 274869 158930 274935 158933
rect 321053 158930 321119 158933
rect 360705 158930 360771 158933
rect 361717 158930 361783 158933
rect 274869 158928 278076 158930
rect 274869 158872 274874 158928
rect 274930 158872 278076 158928
rect 274869 158870 278076 158872
rect 317820 158928 321119 158930
rect 317820 158872 321058 158928
rect 321114 158872 321119 158928
rect 317820 158870 321119 158872
rect 358852 158928 361783 158930
rect 358852 158872 360710 158928
rect 360766 158872 361722 158928
rect 361778 158872 361783 158928
rect 358852 158870 361783 158872
rect 274869 158867 274935 158870
rect 321053 158867 321119 158870
rect 360705 158867 360771 158870
rect 361717 158867 361783 158870
rect 87281 158658 87347 158661
rect 87281 158656 90058 158658
rect 87281 158600 87286 158656
rect 87342 158600 90058 158656
rect 87281 158598 90058 158600
rect 87281 158595 87347 158598
rect 49142 158324 49148 158388
rect 49212 158324 49218 158388
rect 89998 158152 90058 158598
rect 132545 158114 132611 158117
rect 129772 158112 132611 158114
rect 129772 158056 132550 158112
rect 132606 158056 132611 158112
rect 129772 158054 132611 158056
rect 132545 158051 132611 158054
rect 182317 158114 182383 158117
rect 226293 158114 226359 158117
rect 182317 158112 184052 158114
rect 182317 158056 182322 158112
rect 182378 158056 184052 158112
rect 182317 158054 184052 158056
rect 223796 158112 226359 158114
rect 223796 158056 226298 158112
rect 226354 158056 226359 158112
rect 223796 158054 226359 158056
rect 182317 158051 182383 158054
rect 226293 158051 226359 158054
rect 275513 158114 275579 158117
rect 321605 158114 321671 158117
rect 275513 158112 278076 158114
rect 275513 158056 275518 158112
rect 275574 158056 278076 158112
rect 275513 158054 278076 158056
rect 317820 158112 321671 158114
rect 317820 158056 321610 158112
rect 321666 158056 321671 158112
rect 317820 158054 321671 158056
rect 275513 158051 275579 158054
rect 321605 158051 321671 158054
rect 79737 157978 79803 157981
rect 76780 157976 79803 157978
rect 76780 157920 79742 157976
rect 79798 157920 79803 157976
rect 76780 157918 79803 157920
rect 79737 157915 79803 157918
rect 140733 157978 140799 157981
rect 173669 157978 173735 157981
rect 140733 157976 143020 157978
rect 140733 157920 140738 157976
rect 140794 157920 143020 157976
rect 140733 157918 143020 157920
rect 170804 157976 173735 157978
rect 170804 157920 173674 157976
rect 173730 157920 173735 157976
rect 170804 157918 173735 157920
rect 140733 157915 140799 157918
rect 173669 157915 173735 157918
rect 234113 157978 234179 157981
rect 266589 157978 266655 157981
rect 234113 157976 237044 157978
rect 234113 157920 234118 157976
rect 234174 157920 237044 157976
rect 234113 157918 237044 157920
rect 264828 157976 266655 157978
rect 264828 157920 266594 157976
rect 266650 157920 266655 157976
rect 264828 157918 266655 157920
rect 234113 157915 234179 157918
rect 266589 157915 266655 157918
rect 327217 157978 327283 157981
rect 327217 157976 331068 157978
rect 327217 157920 327222 157976
rect 327278 157920 331068 157976
rect 327217 157918 331068 157920
rect 327217 157915 327283 157918
rect 87189 157706 87255 157709
rect 87189 157704 90058 157706
rect 87189 157648 87194 157704
rect 87250 157648 90058 157704
rect 87189 157646 90058 157648
rect 87189 157643 87255 157646
rect 89998 157200 90058 157646
rect 132269 157162 132335 157165
rect 129772 157160 132335 157162
rect 129772 157104 132274 157160
rect 132330 157104 132335 157160
rect 129772 157102 132335 157104
rect 132269 157099 132335 157102
rect 182317 157162 182383 157165
rect 226109 157162 226175 157165
rect 182317 157160 184052 157162
rect 182317 157104 182322 157160
rect 182378 157104 184052 157160
rect 182317 157102 184052 157104
rect 223796 157160 226175 157162
rect 223796 157104 226114 157160
rect 226170 157104 226175 157160
rect 223796 157102 226175 157104
rect 182317 157099 182383 157102
rect 226109 157099 226175 157102
rect 275605 157162 275671 157165
rect 321605 157162 321671 157165
rect 275605 157160 278076 157162
rect 275605 157104 275610 157160
rect 275666 157104 278076 157160
rect 275605 157102 278076 157104
rect 317820 157160 321671 157162
rect 317820 157104 321610 157160
rect 321666 157104 321671 157160
rect 317820 157102 321671 157104
rect 275605 157099 275671 157102
rect 321605 157099 321671 157102
rect 140365 156618 140431 156621
rect 173301 156618 173367 156621
rect 140365 156616 143020 156618
rect 140365 156560 140370 156616
rect 140426 156560 143020 156616
rect 140365 156558 143020 156560
rect 170804 156616 173367 156618
rect 170804 156560 173306 156616
rect 173362 156560 173367 156616
rect 170804 156558 173367 156560
rect 140365 156555 140431 156558
rect 173301 156555 173367 156558
rect 233469 156618 233535 156621
rect 267325 156618 267391 156621
rect 233469 156616 237044 156618
rect 233469 156560 233474 156616
rect 233530 156560 237044 156616
rect 233469 156558 237044 156560
rect 264828 156616 267391 156618
rect 264828 156560 267330 156616
rect 267386 156560 267391 156616
rect 264828 156558 267391 156560
rect 233469 156555 233535 156558
rect 267325 156555 267391 156558
rect 327217 156618 327283 156621
rect 327217 156616 331068 156618
rect 327217 156560 327222 156616
rect 327278 156560 331068 156616
rect 327217 156558 331068 156560
rect 327217 156555 327283 156558
rect 77253 156550 77319 156553
rect 76780 156548 77319 156550
rect 76780 156492 77258 156548
rect 77314 156492 77319 156548
rect 76780 156490 77319 156492
rect 77253 156487 77319 156490
rect 87189 156346 87255 156349
rect 132361 156346 132427 156349
rect 87189 156344 90028 156346
rect 87189 156288 87194 156344
rect 87250 156288 90028 156344
rect 87189 156286 90028 156288
rect 129772 156344 132427 156346
rect 129772 156288 132366 156344
rect 132422 156288 132427 156344
rect 129772 156286 132427 156288
rect 87189 156283 87255 156286
rect 132361 156283 132427 156286
rect 182317 156346 182383 156349
rect 226385 156346 226451 156349
rect 182317 156344 184052 156346
rect 182317 156288 182322 156344
rect 182378 156288 184052 156344
rect 182317 156286 184052 156288
rect 223796 156344 226451 156346
rect 223796 156288 226390 156344
rect 226446 156288 226451 156344
rect 223796 156286 226451 156288
rect 182317 156283 182383 156286
rect 226385 156283 226451 156286
rect 274961 156346 275027 156349
rect 321053 156346 321119 156349
rect 274961 156344 278076 156346
rect 274961 156288 274966 156344
rect 275022 156288 278076 156344
rect 274961 156286 278076 156288
rect 317820 156344 321119 156346
rect 317820 156288 321058 156344
rect 321114 156288 321119 156344
rect 317820 156286 321119 156288
rect 274961 156283 275027 156286
rect 321053 156283 321119 156286
rect 132085 156074 132151 156077
rect 129742 156072 132151 156074
rect 129742 156016 132090 156072
rect 132146 156016 132151 156072
rect 129742 156014 132151 156016
rect 46433 155802 46499 155805
rect 46433 155800 49180 155802
rect 46433 155744 46438 155800
rect 46494 155772 49180 155800
rect 46494 155744 49210 155772
rect 46433 155742 49210 155744
rect 46433 155739 46499 155742
rect 49150 155396 49210 155742
rect 129742 155432 129802 156014
rect 132085 156011 132151 156014
rect 182133 156074 182199 156077
rect 274869 156074 274935 156077
rect 182133 156072 184082 156074
rect 182133 156016 182138 156072
rect 182194 156016 184082 156072
rect 182133 156014 184082 156016
rect 182133 156011 182199 156014
rect 184022 155432 184082 156014
rect 274869 156072 278106 156074
rect 274869 156016 274874 156072
rect 274930 156016 278106 156072
rect 274869 156014 278106 156016
rect 274869 156011 274935 156014
rect 278046 155432 278106 156014
rect 360889 155802 360955 155805
rect 361717 155802 361783 155805
rect 358852 155800 361783 155802
rect 358852 155744 360894 155800
rect 360950 155744 361722 155800
rect 361778 155744 361783 155800
rect 358852 155742 361783 155744
rect 360889 155739 360955 155742
rect 361717 155739 361783 155742
rect 49142 155332 49148 155396
rect 49212 155332 49218 155396
rect 87189 155394 87255 155397
rect 226017 155394 226083 155397
rect 321605 155394 321671 155397
rect 87189 155392 90028 155394
rect 87189 155336 87194 155392
rect 87250 155336 90028 155392
rect 87189 155334 90028 155336
rect 223796 155392 226083 155394
rect 223796 155336 226022 155392
rect 226078 155336 226083 155392
rect 223796 155334 226083 155336
rect 317820 155392 321671 155394
rect 317820 155336 321610 155392
rect 321666 155336 321671 155392
rect 317820 155334 321671 155336
rect 87189 155331 87255 155334
rect 226017 155331 226083 155334
rect 321605 155331 321671 155334
rect 79737 155122 79803 155125
rect 131993 155122 132059 155125
rect 76780 155120 79803 155122
rect 76780 155064 79742 155120
rect 79798 155064 79803 155120
rect 76780 155062 79803 155064
rect 79737 155059 79803 155062
rect 129742 155120 132059 155122
rect 129742 155064 131998 155120
rect 132054 155064 132059 155120
rect 129742 155062 132059 155064
rect 129742 154480 129802 155062
rect 131993 155059 132059 155062
rect 139629 155122 139695 155125
rect 173577 155122 173643 155125
rect 139629 155120 143020 155122
rect 139629 155064 139634 155120
rect 139690 155064 143020 155120
rect 139629 155062 143020 155064
rect 170804 155120 173643 155122
rect 170804 155064 173582 155120
rect 173638 155064 173643 155120
rect 170804 155062 173643 155064
rect 139629 155059 139695 155062
rect 173577 155059 173643 155062
rect 233469 155122 233535 155125
rect 266589 155122 266655 155125
rect 233469 155120 237044 155122
rect 233469 155064 233474 155120
rect 233530 155064 237044 155120
rect 233469 155062 237044 155064
rect 264828 155120 266655 155122
rect 264828 155064 266594 155120
rect 266650 155064 266655 155120
rect 264828 155062 266655 155064
rect 233469 155059 233535 155062
rect 266589 155059 266655 155062
rect 328413 155122 328479 155125
rect 328413 155120 331068 155122
rect 328413 155064 328418 155120
rect 328474 155064 331068 155120
rect 328413 155062 331068 155064
rect 328413 155059 328479 155062
rect 182317 154986 182383 154989
rect 274869 154986 274935 154989
rect 182317 154984 184082 154986
rect 182317 154928 182322 154984
rect 182378 154928 184082 154984
rect 182317 154926 184082 154928
rect 182317 154923 182383 154926
rect 184022 154480 184082 154926
rect 274869 154984 278106 154986
rect 274869 154928 274874 154984
rect 274930 154928 278106 154984
rect 274869 154926 278106 154928
rect 274869 154923 274935 154926
rect 278046 154480 278106 154926
rect 87189 154442 87255 154445
rect 225925 154442 225991 154445
rect 320869 154442 320935 154445
rect 87189 154440 90028 154442
rect 87189 154384 87194 154440
rect 87250 154384 90028 154440
rect 87189 154382 90028 154384
rect 223796 154440 225991 154442
rect 223796 154384 225930 154440
rect 225986 154384 225991 154440
rect 223796 154382 225991 154384
rect 317820 154440 320935 154442
rect 317820 154384 320874 154440
rect 320930 154384 320935 154440
rect 317820 154382 320935 154384
rect 87189 154379 87255 154382
rect 225925 154379 225991 154382
rect 320869 154379 320935 154382
rect 9896 154306 10376 154336
rect 12669 154306 12735 154309
rect 9896 154304 12735 154306
rect 9896 154248 12674 154304
rect 12730 154248 12735 154304
rect 9896 154246 12735 154248
rect 9896 154216 10376 154246
rect 12669 154243 12735 154246
rect 81761 153762 81827 153765
rect 76780 153760 81827 153762
rect 76780 153704 81766 153760
rect 81822 153704 81827 153760
rect 76780 153702 81827 153704
rect 81761 153699 81827 153702
rect 139537 153762 139603 153765
rect 173393 153762 173459 153765
rect 139537 153760 143020 153762
rect 139537 153704 139542 153760
rect 139598 153704 143020 153760
rect 139537 153702 143020 153704
rect 170804 153760 173459 153762
rect 170804 153704 173398 153760
rect 173454 153704 173459 153760
rect 170804 153702 173459 153704
rect 139537 153699 139603 153702
rect 173393 153699 173459 153702
rect 234573 153762 234639 153765
rect 266681 153762 266747 153765
rect 234573 153760 237044 153762
rect 234573 153704 234578 153760
rect 234634 153704 237044 153760
rect 234573 153702 237044 153704
rect 264828 153760 266747 153762
rect 264828 153704 266686 153760
rect 266742 153704 266747 153760
rect 264828 153702 266747 153704
rect 234573 153699 234639 153702
rect 266681 153699 266747 153702
rect 328413 153762 328479 153765
rect 328413 153760 331068 153762
rect 328413 153704 328418 153760
rect 328474 153704 331068 153760
rect 328413 153702 331068 153704
rect 328413 153699 328479 153702
rect 87189 153626 87255 153629
rect 131901 153626 131967 153629
rect 87189 153624 90028 153626
rect 87189 153568 87194 153624
rect 87250 153568 90028 153624
rect 87189 153566 90028 153568
rect 129772 153624 131967 153626
rect 129772 153568 131906 153624
rect 131962 153568 131967 153624
rect 129772 153566 131967 153568
rect 87189 153563 87255 153566
rect 131901 153563 131967 153566
rect 182317 153626 182383 153629
rect 225833 153626 225899 153629
rect 182317 153624 184052 153626
rect 182317 153568 182322 153624
rect 182378 153568 184052 153624
rect 182317 153566 184052 153568
rect 223796 153624 225899 153626
rect 223796 153568 225838 153624
rect 225894 153568 225899 153624
rect 223796 153566 225899 153568
rect 182317 153563 182383 153566
rect 225833 153563 225899 153566
rect 274869 153626 274935 153629
rect 321605 153626 321671 153629
rect 274869 153624 278076 153626
rect 274869 153568 274874 153624
rect 274930 153568 278076 153624
rect 274869 153566 278076 153568
rect 317820 153624 321671 153626
rect 317820 153568 321610 153624
rect 321666 153568 321671 153624
rect 317820 153566 321671 153568
rect 274869 153563 274935 153566
rect 321605 153563 321671 153566
rect 132637 153354 132703 153357
rect 129742 153352 132703 153354
rect 129742 153296 132642 153352
rect 132698 153296 132703 153352
rect 129742 153294 132703 153296
rect 49142 152884 49148 152948
rect 49212 152884 49218 152948
rect 49150 152644 49210 152884
rect 129742 152712 129802 153294
rect 132637 153291 132703 153294
rect 274961 153354 275027 153357
rect 274961 153352 278106 153354
rect 274961 153296 274966 153352
rect 275022 153296 278106 153352
rect 274961 153294 278106 153296
rect 274961 153291 275027 153294
rect 181397 153218 181463 153221
rect 181397 153216 184082 153218
rect 181397 153160 181402 153216
rect 181458 153160 184082 153216
rect 181397 153158 184082 153160
rect 181397 153155 181463 153158
rect 184022 152712 184082 153158
rect 278046 152712 278106 153294
rect 87189 152674 87255 152677
rect 225649 152674 225715 152677
rect 320501 152674 320567 152677
rect 360797 152674 360863 152677
rect 87189 152672 90028 152674
rect 87189 152616 87194 152672
rect 87250 152616 90028 152672
rect 87189 152614 90028 152616
rect 223796 152672 225715 152674
rect 223796 152616 225654 152672
rect 225710 152616 225715 152672
rect 223796 152614 225715 152616
rect 317820 152672 320567 152674
rect 317820 152616 320506 152672
rect 320562 152616 320567 152672
rect 317820 152614 320567 152616
rect 358852 152672 360863 152674
rect 358852 152616 360802 152672
rect 360858 152616 360863 152672
rect 358852 152614 360863 152616
rect 87189 152611 87255 152614
rect 225649 152611 225715 152614
rect 320501 152611 320567 152614
rect 360797 152611 360863 152614
rect 81761 152402 81827 152405
rect 76780 152400 81827 152402
rect 76780 152344 81766 152400
rect 81822 152344 81827 152400
rect 76780 152342 81827 152344
rect 81761 152339 81827 152342
rect 140825 152402 140891 152405
rect 173577 152402 173643 152405
rect 140825 152400 143020 152402
rect 140825 152344 140830 152400
rect 140886 152344 143020 152400
rect 140825 152342 143020 152344
rect 170804 152400 173643 152402
rect 170804 152344 173582 152400
rect 173638 152344 173643 152400
rect 170804 152342 173643 152344
rect 140825 152339 140891 152342
rect 173577 152339 173643 152342
rect 234297 152402 234363 152405
rect 266589 152402 266655 152405
rect 234297 152400 237044 152402
rect 234297 152344 234302 152400
rect 234358 152344 237044 152400
rect 234297 152342 237044 152344
rect 264828 152400 266655 152402
rect 264828 152344 266594 152400
rect 266650 152344 266655 152400
rect 264828 152342 266655 152344
rect 234297 152339 234363 152342
rect 266589 152339 266655 152342
rect 328229 152402 328295 152405
rect 328229 152400 331068 152402
rect 328229 152344 328234 152400
rect 328290 152344 331068 152400
rect 328229 152342 331068 152344
rect 328229 152339 328295 152342
rect 131625 152266 131691 152269
rect 129742 152264 131691 152266
rect 129742 152208 131630 152264
rect 131686 152208 131691 152264
rect 129742 152206 131691 152208
rect 129742 151896 129802 152206
rect 131625 152203 131691 152206
rect 182317 152130 182383 152133
rect 274869 152130 274935 152133
rect 182317 152128 184082 152130
rect 182317 152072 182322 152128
rect 182378 152072 184082 152128
rect 182317 152070 184082 152072
rect 182317 152067 182383 152070
rect 184022 151896 184082 152070
rect 274869 152128 278106 152130
rect 274869 152072 274874 152128
rect 274930 152072 278106 152128
rect 274869 152070 278106 152072
rect 274869 152067 274935 152070
rect 278046 151896 278106 152070
rect 88109 151858 88175 151861
rect 226201 151858 226267 151861
rect 320777 151858 320843 151861
rect 88109 151856 90028 151858
rect 88109 151800 88114 151856
rect 88170 151800 90028 151856
rect 88109 151798 90028 151800
rect 223796 151856 226267 151858
rect 223796 151800 226206 151856
rect 226262 151800 226267 151856
rect 223796 151798 226267 151800
rect 317820 151856 320843 151858
rect 317820 151800 320782 151856
rect 320838 151800 320843 151856
rect 317820 151798 320843 151800
rect 88109 151795 88175 151798
rect 226201 151795 226267 151798
rect 320777 151795 320843 151798
rect 79737 150906 79803 150909
rect 76780 150904 79803 150906
rect 76780 150848 79742 150904
rect 79798 150848 79803 150904
rect 76780 150846 79803 150848
rect 79737 150843 79803 150846
rect 87097 150906 87163 150909
rect 132453 150906 132519 150909
rect 87097 150904 90028 150906
rect 87097 150848 87102 150904
rect 87158 150848 90028 150904
rect 87097 150846 90028 150848
rect 129772 150904 132519 150906
rect 129772 150848 132458 150904
rect 132514 150848 132519 150904
rect 129772 150846 132519 150848
rect 87097 150843 87163 150846
rect 132453 150843 132519 150846
rect 140457 150906 140523 150909
rect 173577 150906 173643 150909
rect 140457 150904 143020 150906
rect 140457 150848 140462 150904
rect 140518 150848 143020 150904
rect 140457 150846 143020 150848
rect 170804 150904 173643 150906
rect 170804 150848 173582 150904
rect 173638 150848 173643 150904
rect 170804 150846 173643 150848
rect 140457 150843 140523 150846
rect 173577 150843 173643 150846
rect 182317 150906 182383 150909
rect 226477 150906 226543 150909
rect 182317 150904 184052 150906
rect 182317 150848 182322 150904
rect 182378 150848 184052 150904
rect 182317 150846 184052 150848
rect 223796 150904 226543 150906
rect 223796 150848 226482 150904
rect 226538 150848 226543 150904
rect 223796 150846 226543 150848
rect 182317 150843 182383 150846
rect 226477 150843 226543 150846
rect 233469 150906 233535 150909
rect 266589 150906 266655 150909
rect 233469 150904 237044 150906
rect 233469 150848 233474 150904
rect 233530 150848 237044 150904
rect 233469 150846 237044 150848
rect 264828 150904 266655 150906
rect 264828 150848 266594 150904
rect 266650 150848 266655 150904
rect 264828 150846 266655 150848
rect 233469 150843 233535 150846
rect 266589 150843 266655 150846
rect 274869 150906 274935 150909
rect 321697 150906 321763 150909
rect 274869 150904 278076 150906
rect 274869 150848 274874 150904
rect 274930 150848 278076 150904
rect 274869 150846 278076 150848
rect 317820 150904 321763 150906
rect 317820 150848 321702 150904
rect 321758 150848 321763 150904
rect 317820 150846 321763 150848
rect 274869 150843 274935 150846
rect 321697 150843 321763 150846
rect 328413 150906 328479 150909
rect 328413 150904 331068 150906
rect 328413 150848 328418 150904
rect 328474 150848 331068 150904
rect 328413 150846 331068 150848
rect 328413 150843 328479 150846
rect 182225 150634 182291 150637
rect 274961 150634 275027 150637
rect 182225 150632 184082 150634
rect 182225 150576 182230 150632
rect 182286 150576 184082 150632
rect 182225 150574 184082 150576
rect 182225 150571 182291 150574
rect 131349 150498 131415 150501
rect 129742 150496 131415 150498
rect 129742 150440 131354 150496
rect 131410 150440 131415 150496
rect 129742 150438 131415 150440
rect 129742 150128 129802 150438
rect 131349 150435 131415 150438
rect 184022 150128 184082 150574
rect 274961 150632 278106 150634
rect 274961 150576 274966 150632
rect 275022 150576 278106 150632
rect 274961 150574 278106 150576
rect 274961 150571 275027 150574
rect 278046 150128 278106 150574
rect 87189 150090 87255 150093
rect 225557 150090 225623 150093
rect 321605 150090 321671 150093
rect 87189 150088 90028 150090
rect 87189 150032 87194 150088
rect 87250 150032 90028 150088
rect 87189 150030 90028 150032
rect 223796 150088 225623 150090
rect 223796 150032 225562 150088
rect 225618 150032 225623 150088
rect 223796 150030 225623 150032
rect 317820 150088 321671 150090
rect 317820 150032 321610 150088
rect 321666 150032 321671 150088
rect 317820 150030 321671 150032
rect 87189 150027 87255 150030
rect 225557 150027 225623 150030
rect 321605 150027 321671 150030
rect 81761 149546 81827 149549
rect 131809 149546 131875 149549
rect 76780 149544 81827 149546
rect 49150 149004 49210 149516
rect 76780 149488 81766 149544
rect 81822 149488 81827 149544
rect 76780 149486 81827 149488
rect 81761 149483 81827 149486
rect 129742 149544 131875 149546
rect 129742 149488 131814 149544
rect 131870 149488 131875 149544
rect 129742 149486 131875 149488
rect 129742 149176 129802 149486
rect 131809 149483 131875 149486
rect 140549 149546 140615 149549
rect 172749 149546 172815 149549
rect 140549 149544 143020 149546
rect 140549 149488 140554 149544
rect 140610 149488 143020 149544
rect 140549 149486 143020 149488
rect 170804 149544 172815 149546
rect 170804 149488 172754 149544
rect 172810 149488 172815 149544
rect 170804 149486 172815 149488
rect 140549 149483 140615 149486
rect 172749 149483 172815 149486
rect 181673 149546 181739 149549
rect 233469 149546 233535 149549
rect 266589 149546 266655 149549
rect 181673 149544 184082 149546
rect 181673 149488 181678 149544
rect 181734 149488 184082 149544
rect 181673 149486 184082 149488
rect 181673 149483 181739 149486
rect 184022 149176 184082 149486
rect 233469 149544 237044 149546
rect 233469 149488 233474 149544
rect 233530 149488 237044 149544
rect 233469 149486 237044 149488
rect 264828 149544 266655 149546
rect 264828 149488 266594 149544
rect 266650 149488 266655 149544
rect 264828 149486 266655 149488
rect 233469 149483 233535 149486
rect 266589 149483 266655 149486
rect 275697 149546 275763 149549
rect 328413 149546 328479 149549
rect 360981 149546 361047 149549
rect 275697 149544 278106 149546
rect 275697 149488 275702 149544
rect 275758 149488 278106 149544
rect 275697 149486 278106 149488
rect 275697 149483 275763 149486
rect 278046 149176 278106 149486
rect 328413 149544 331068 149546
rect 328413 149488 328418 149544
rect 328474 149488 331068 149544
rect 328413 149486 331068 149488
rect 358852 149544 361047 149546
rect 358852 149488 360986 149544
rect 361042 149488 361047 149544
rect 358852 149486 361047 149488
rect 328413 149483 328479 149486
rect 360981 149483 361047 149486
rect 87189 149138 87255 149141
rect 226293 149138 226359 149141
rect 321053 149138 321119 149141
rect 87189 149136 90028 149138
rect 87189 149080 87194 149136
rect 87250 149080 90028 149136
rect 87189 149078 90028 149080
rect 223796 149136 226359 149138
rect 223796 149080 226298 149136
rect 226354 149080 226359 149136
rect 223796 149078 226359 149080
rect 317820 149136 321119 149138
rect 317820 149080 321058 149136
rect 321114 149080 321119 149136
rect 317820 149078 321119 149080
rect 87189 149075 87255 149078
rect 226293 149075 226359 149078
rect 321053 149075 321119 149078
rect 49142 148940 49148 149004
rect 49212 148940 49218 149004
rect 131349 148866 131415 148869
rect 129742 148864 131415 148866
rect 129742 148808 131354 148864
rect 131410 148808 131415 148864
rect 129742 148806 131415 148808
rect 129742 148360 129802 148806
rect 131349 148803 131415 148806
rect 181857 148866 181923 148869
rect 274869 148866 274935 148869
rect 181857 148864 184082 148866
rect 181857 148808 181862 148864
rect 181918 148808 184082 148864
rect 181857 148806 184082 148808
rect 181857 148803 181923 148806
rect 184022 148360 184082 148806
rect 274869 148864 278106 148866
rect 274869 148808 274874 148864
rect 274930 148808 278106 148864
rect 274869 148806 278106 148808
rect 274869 148803 274935 148806
rect 278046 148360 278106 148806
rect 87281 148322 87347 148325
rect 225925 148322 225991 148325
rect 321605 148322 321671 148325
rect 87281 148320 90028 148322
rect 87281 148264 87286 148320
rect 87342 148264 90028 148320
rect 87281 148262 90028 148264
rect 223796 148320 225991 148322
rect 223796 148264 225930 148320
rect 225986 148264 225991 148320
rect 223796 148262 225991 148264
rect 317820 148320 321671 148322
rect 317820 148264 321610 148320
rect 321666 148264 321671 148320
rect 317820 148262 321671 148264
rect 87281 148259 87347 148262
rect 225925 148259 225991 148262
rect 321605 148259 321671 148262
rect 79737 148186 79803 148189
rect 76780 148184 79803 148186
rect 76780 148128 79742 148184
rect 79798 148128 79803 148184
rect 76780 148126 79803 148128
rect 79737 148123 79803 148126
rect 138893 148186 138959 148189
rect 173577 148186 173643 148189
rect 138893 148184 143020 148186
rect 138893 148128 138898 148184
rect 138954 148128 143020 148184
rect 138893 148126 143020 148128
rect 170804 148184 173643 148186
rect 170804 148128 173582 148184
rect 173638 148128 173643 148184
rect 170804 148126 173643 148128
rect 138893 148123 138959 148126
rect 173577 148123 173643 148126
rect 233469 148186 233535 148189
rect 266957 148186 267023 148189
rect 233469 148184 237044 148186
rect 233469 148128 233474 148184
rect 233530 148128 237044 148184
rect 233469 148126 237044 148128
rect 264828 148184 267023 148186
rect 264828 148128 266962 148184
rect 267018 148128 267023 148184
rect 264828 148126 267023 148128
rect 233469 148123 233535 148126
rect 266957 148123 267023 148126
rect 328413 148186 328479 148189
rect 429429 148186 429495 148189
rect 434416 148186 434896 148216
rect 328413 148184 331068 148186
rect 328413 148128 328418 148184
rect 328474 148128 331068 148184
rect 328413 148126 331068 148128
rect 429429 148184 434896 148186
rect 429429 148128 429434 148184
rect 429490 148128 434896 148184
rect 429429 148126 434896 148128
rect 328413 148123 328479 148126
rect 429429 148123 429495 148126
rect 434416 148096 434896 148126
rect 80105 146690 80171 146693
rect 76780 146688 80171 146690
rect 76780 146632 80110 146688
rect 80166 146632 80171 146688
rect 76780 146630 80171 146632
rect 80105 146627 80171 146630
rect 139629 146690 139695 146693
rect 173853 146690 173919 146693
rect 139629 146688 143020 146690
rect 139629 146632 139634 146688
rect 139690 146632 143020 146688
rect 139629 146630 143020 146632
rect 170804 146688 173919 146690
rect 170804 146632 173858 146688
rect 173914 146632 173919 146688
rect 170804 146630 173919 146632
rect 139629 146627 139695 146630
rect 173853 146627 173919 146630
rect 233469 146690 233535 146693
rect 267877 146690 267943 146693
rect 233469 146688 237044 146690
rect 233469 146632 233474 146688
rect 233530 146632 237044 146688
rect 233469 146630 237044 146632
rect 264828 146688 267943 146690
rect 264828 146632 267882 146688
rect 267938 146632 267943 146688
rect 264828 146630 267943 146632
rect 233469 146627 233535 146630
rect 267877 146627 267943 146630
rect 327217 146690 327283 146693
rect 327217 146688 331068 146690
rect 327217 146632 327222 146688
rect 327278 146632 331068 146688
rect 327217 146630 331068 146632
rect 327217 146627 327283 146630
rect 361165 146418 361231 146421
rect 358852 146416 361231 146418
rect 49150 146148 49210 146388
rect 358852 146360 361170 146416
rect 361226 146360 361231 146416
rect 358852 146358 361231 146360
rect 361165 146355 361231 146358
rect 49142 146084 49148 146148
rect 49212 146084 49218 146148
rect 79737 145330 79803 145333
rect 76780 145328 79803 145330
rect 76780 145272 79742 145328
rect 79798 145272 79803 145328
rect 76780 145270 79803 145272
rect 79737 145267 79803 145270
rect 139629 145330 139695 145333
rect 173945 145330 174011 145333
rect 139629 145328 143020 145330
rect 139629 145272 139634 145328
rect 139690 145272 143020 145328
rect 139629 145270 143020 145272
rect 170804 145328 174011 145330
rect 170804 145272 173950 145328
rect 174006 145272 174011 145328
rect 170804 145270 174011 145272
rect 139629 145267 139695 145270
rect 173945 145267 174011 145270
rect 233469 145330 233535 145333
rect 266773 145330 266839 145333
rect 233469 145328 237044 145330
rect 233469 145272 233474 145328
rect 233530 145272 237044 145328
rect 233469 145270 237044 145272
rect 264828 145328 266839 145330
rect 264828 145272 266778 145328
rect 266834 145272 266839 145328
rect 264828 145270 266839 145272
rect 233469 145267 233535 145270
rect 266773 145267 266839 145270
rect 328505 145330 328571 145333
rect 328505 145328 331068 145330
rect 328505 145272 328510 145328
rect 328566 145272 331068 145328
rect 328505 145270 331068 145272
rect 328505 145267 328571 145270
rect 98873 145196 98939 145197
rect 98822 145132 98828 145196
rect 98892 145194 98939 145196
rect 98892 145192 98984 145194
rect 98934 145136 98984 145192
rect 98892 145134 98984 145136
rect 98892 145132 98939 145134
rect 98873 145131 98939 145132
rect 192897 144650 192963 144653
rect 197630 144650 197636 144652
rect 192897 144648 197636 144650
rect 192897 144592 192902 144648
rect 192958 144592 197636 144648
rect 192897 144590 197636 144592
rect 192897 144587 192963 144590
rect 197630 144588 197636 144590
rect 197700 144588 197706 144652
rect 292574 144588 292580 144652
rect 292644 144650 292650 144652
rect 294189 144650 294255 144653
rect 292644 144648 294255 144650
rect 292644 144592 294194 144648
rect 294250 144592 294255 144648
rect 292644 144590 294255 144592
rect 292644 144588 292650 144590
rect 294189 144587 294255 144590
rect 95193 144516 95259 144517
rect 95142 144452 95148 144516
rect 95212 144514 95259 144516
rect 95212 144512 95304 144514
rect 95254 144456 95304 144512
rect 95212 144454 95304 144456
rect 95212 144452 95259 144454
rect 187878 144452 187884 144516
rect 187948 144514 187954 144516
rect 189217 144514 189283 144517
rect 187948 144512 189283 144514
rect 187948 144456 189222 144512
rect 189278 144456 189283 144512
rect 187948 144454 189283 144456
rect 187948 144452 187954 144454
rect 95193 144451 95259 144452
rect 189217 144451 189283 144454
rect 79737 143970 79803 143973
rect 76780 143968 79803 143970
rect 76780 143912 79742 143968
rect 79798 143912 79803 143968
rect 76780 143910 79803 143912
rect 79737 143907 79803 143910
rect 139629 143970 139695 143973
rect 174037 143970 174103 143973
rect 139629 143968 143020 143970
rect 139629 143912 139634 143968
rect 139690 143912 143020 143968
rect 139629 143910 143020 143912
rect 170804 143968 174103 143970
rect 170804 143912 174042 143968
rect 174098 143912 174103 143968
rect 170804 143910 174103 143912
rect 139629 143907 139695 143910
rect 174037 143907 174103 143910
rect 233469 143970 233535 143973
rect 267785 143970 267851 143973
rect 233469 143968 237044 143970
rect 233469 143912 233474 143968
rect 233530 143912 237044 143968
rect 233469 143910 237044 143912
rect 264828 143968 267851 143970
rect 264828 143912 267790 143968
rect 267846 143912 267851 143968
rect 264828 143910 267851 143912
rect 233469 143907 233535 143910
rect 267785 143907 267851 143910
rect 328321 143970 328387 143973
rect 328321 143968 331068 143970
rect 328321 143912 328326 143968
rect 328382 143912 331068 143968
rect 328321 143910 331068 143912
rect 328321 143907 328387 143910
rect 282454 143772 282460 143836
rect 282524 143834 282530 143836
rect 283742 143834 283748 143836
rect 282524 143774 283748 143834
rect 282524 143772 282530 143774
rect 283742 143772 283748 143774
rect 283812 143772 283818 143836
rect 302326 143772 302332 143836
rect 302396 143834 302402 143836
rect 303849 143834 303915 143837
rect 302396 143832 303915 143834
rect 302396 143776 303854 143832
rect 303910 143776 303915 143832
rect 302396 143774 303915 143776
rect 302396 143772 302402 143774
rect 303849 143771 303915 143774
rect 9896 143562 10376 143592
rect 13313 143562 13379 143565
rect 9896 143560 13379 143562
rect 9896 143504 13318 143560
rect 13374 143504 13379 143560
rect 9896 143502 13379 143504
rect 9896 143472 10376 143502
rect 13313 143499 13379 143502
rect 47077 143426 47143 143429
rect 361073 143426 361139 143429
rect 47077 143424 48996 143426
rect 47077 143368 47082 143424
rect 47138 143368 48996 143424
rect 47077 143366 48996 143368
rect 358852 143424 361139 143426
rect 358852 143368 361078 143424
rect 361134 143368 361139 143424
rect 358852 143366 361139 143368
rect 47077 143363 47143 143366
rect 361073 143363 361139 143366
rect 203150 143228 203156 143292
rect 203220 143290 203226 143292
rect 203753 143290 203819 143293
rect 231670 143290 231676 143292
rect 203220 143288 231676 143290
rect 203220 143232 203758 143288
rect 203814 143232 231676 143288
rect 203220 143230 231676 143232
rect 203220 143228 203226 143230
rect 203753 143227 203819 143230
rect 231670 143228 231676 143230
rect 231740 143228 231746 143292
rect 109729 143156 109795 143157
rect 109678 143092 109684 143156
rect 109748 143154 109795 143156
rect 230985 143154 231051 143157
rect 297777 143156 297843 143157
rect 231118 143154 231124 143156
rect 109748 143152 109840 143154
rect 109790 143096 109840 143152
rect 109748 143094 109840 143096
rect 230985 143152 231124 143154
rect 230985 143096 230990 143152
rect 231046 143096 231124 143152
rect 230985 143094 231124 143096
rect 109748 143092 109795 143094
rect 109729 143091 109795 143092
rect 230985 143091 231051 143094
rect 231118 143092 231124 143094
rect 231188 143092 231194 143156
rect 297726 143092 297732 143156
rect 297796 143154 297843 143156
rect 297796 143152 297888 143154
rect 297838 143096 297888 143152
rect 297796 143094 297888 143096
rect 297796 143092 297843 143094
rect 297777 143091 297843 143092
rect 105998 142548 106004 142612
rect 106068 142610 106074 142612
rect 106141 142610 106207 142613
rect 106068 142608 106207 142610
rect 106068 142552 106146 142608
rect 106202 142552 106207 142608
rect 106068 142550 106207 142552
rect 106068 142548 106074 142550
rect 106141 142547 106207 142550
rect 140273 142610 140339 142613
rect 173577 142610 173643 142613
rect 267233 142610 267299 142613
rect 140273 142608 143020 142610
rect 140273 142552 140278 142608
rect 140334 142552 143020 142608
rect 140273 142550 143020 142552
rect 170804 142608 173643 142610
rect 170804 142552 173582 142608
rect 173638 142552 173643 142608
rect 170804 142550 173643 142552
rect 264828 142608 267299 142610
rect 264828 142552 267238 142608
rect 267294 142552 267299 142608
rect 264828 142550 267299 142552
rect 140273 142547 140339 142550
rect 173577 142547 173643 142550
rect 267233 142547 267299 142550
rect 77253 142542 77319 142545
rect 76780 142540 77319 142542
rect 76780 142484 77258 142540
rect 77314 142484 77319 142540
rect 76780 142482 77319 142484
rect 77253 142479 77319 142482
rect 73982 142412 73988 142476
rect 74052 142474 74058 142476
rect 74902 142474 74908 142476
rect 74052 142414 74908 142474
rect 74052 142412 74058 142414
rect 74902 142412 74908 142414
rect 74972 142412 74978 142476
rect 147030 142412 147036 142476
rect 147100 142474 147106 142476
rect 150342 142474 150348 142476
rect 147100 142414 150348 142474
rect 147100 142412 147106 142414
rect 150342 142412 150348 142414
rect 150412 142412 150418 142476
rect 74166 142276 74172 142340
rect 74236 142338 74242 142340
rect 77110 142338 77116 142340
rect 74236 142278 77116 142338
rect 74236 142276 74242 142278
rect 77110 142276 77116 142278
rect 77180 142276 77186 142340
rect 144086 142140 144092 142204
rect 144156 142202 144162 142204
rect 147909 142202 147975 142205
rect 144156 142200 147975 142202
rect 144156 142144 147914 142200
rect 147970 142144 147975 142200
rect 144156 142142 147975 142144
rect 150350 142202 150410 142412
rect 150669 142202 150735 142205
rect 150350 142200 150735 142202
rect 150350 142144 150674 142200
rect 150730 142144 150735 142200
rect 150350 142142 150735 142144
rect 144156 142140 144162 142142
rect 147909 142139 147975 142142
rect 150669 142139 150735 142142
rect 167781 142204 167847 142205
rect 167781 142200 167828 142204
rect 167892 142202 167898 142204
rect 167781 142144 167786 142200
rect 167781 142140 167828 142144
rect 167892 142142 167938 142202
rect 167892 142140 167898 142142
rect 167781 142139 167847 142140
rect 76374 142004 76380 142068
rect 76444 142066 76450 142068
rect 77662 142066 77668 142068
rect 76444 142006 77668 142066
rect 76444 142004 76450 142006
rect 77662 142004 77668 142006
rect 77732 142004 77738 142068
rect 147449 142066 147515 142069
rect 219669 142068 219735 142069
rect 147766 142066 147772 142068
rect 147449 142064 147772 142066
rect 147449 142008 147454 142064
rect 147510 142008 147772 142064
rect 147449 142006 147772 142008
rect 147449 142003 147515 142006
rect 147766 142004 147772 142006
rect 147836 142066 147842 142068
rect 148318 142066 148324 142068
rect 147836 142006 148324 142066
rect 147836 142004 147842 142006
rect 148318 142004 148324 142006
rect 148388 142004 148394 142068
rect 219669 142064 219716 142068
rect 219780 142066 219786 142068
rect 233469 142066 233535 142069
rect 237014 142066 237074 142512
rect 242894 142412 242900 142476
rect 242964 142474 242970 142476
rect 247310 142474 247316 142476
rect 242964 142414 247316 142474
rect 242964 142412 242970 142414
rect 246766 142205 246826 142414
rect 247310 142412 247316 142414
rect 247380 142412 247386 142476
rect 249886 142412 249892 142476
rect 249956 142412 249962 142476
rect 250438 142412 250444 142476
rect 250508 142474 250514 142476
rect 255222 142474 255228 142476
rect 250508 142414 255228 142474
rect 250508 142412 250514 142414
rect 255222 142412 255228 142414
rect 255292 142412 255298 142476
rect 289998 142412 290004 142476
rect 290068 142474 290074 142476
rect 290509 142474 290575 142477
rect 290969 142474 291035 142477
rect 290068 142472 291035 142474
rect 290068 142416 290514 142472
rect 290570 142416 290974 142472
rect 291030 142416 291035 142472
rect 290068 142414 291035 142416
rect 290068 142412 290074 142414
rect 242485 142204 242551 142205
rect 242485 142202 242532 142204
rect 242440 142200 242532 142202
rect 242440 142144 242490 142200
rect 242440 142142 242532 142144
rect 242485 142140 242532 142142
rect 242596 142140 242602 142204
rect 246766 142200 246875 142205
rect 246766 142144 246814 142200
rect 246870 142144 246875 142200
rect 246766 142142 246875 142144
rect 242485 142139 242551 142140
rect 246809 142139 246875 142142
rect 219669 142008 219674 142064
rect 219669 142004 219716 142008
rect 219780 142006 219826 142066
rect 233469 142064 237074 142066
rect 233469 142008 233474 142064
rect 233530 142008 237074 142064
rect 233469 142006 237074 142008
rect 243405 142066 243471 142069
rect 246390 142066 246396 142068
rect 243405 142064 246396 142066
rect 243405 142008 243410 142064
rect 243466 142008 246396 142064
rect 243405 142006 246396 142008
rect 219780 142004 219786 142006
rect 219669 142003 219735 142004
rect 233469 142003 233535 142006
rect 243405 142003 243471 142006
rect 246390 142004 246396 142006
rect 246460 142066 246466 142068
rect 249894 142066 249954 142412
rect 290509 142411 290575 142414
rect 290969 142411 291035 142414
rect 246460 142006 249954 142066
rect 328413 142066 328479 142069
rect 331038 142066 331098 142512
rect 328413 142064 331098 142066
rect 328413 142008 328418 142064
rect 328474 142008 331098 142064
rect 328413 142006 331098 142008
rect 246460 142004 246466 142006
rect 328413 142003 328479 142006
rect 105998 141868 106004 141932
rect 106068 141930 106074 141932
rect 136961 141930 137027 141933
rect 106068 141928 137027 141930
rect 106068 141872 136966 141928
rect 137022 141872 137027 141928
rect 106068 141870 137027 141872
rect 106068 141868 106074 141870
rect 136961 141867 137027 141870
rect 74309 141796 74375 141797
rect 74309 141794 74356 141796
rect 74264 141792 74356 141794
rect 74264 141736 74314 141792
rect 74264 141734 74356 141736
rect 74309 141732 74356 141734
rect 74420 141732 74426 141796
rect 74309 141731 74375 141732
rect 74033 141658 74099 141661
rect 75638 141658 75644 141660
rect 74033 141656 75644 141658
rect 74033 141600 74038 141656
rect 74094 141600 75644 141656
rect 74033 141598 75644 141600
rect 74033 141595 74099 141598
rect 75638 141596 75644 141598
rect 75708 141658 75714 141660
rect 82313 141658 82379 141661
rect 75708 141656 82379 141658
rect 75708 141600 82318 141656
rect 82374 141600 82379 141656
rect 75708 141598 82379 141600
rect 75708 141596 75714 141598
rect 82313 141595 82379 141598
rect 74125 141522 74191 141525
rect 76006 141522 76012 141524
rect 74125 141520 76012 141522
rect 74125 141464 74130 141520
rect 74186 141464 76012 141520
rect 74125 141462 76012 141464
rect 74125 141459 74191 141462
rect 76006 141460 76012 141462
rect 76076 141522 76082 141524
rect 77713 141522 77779 141525
rect 76076 141520 77779 141522
rect 76076 141464 77718 141520
rect 77774 141464 77779 141520
rect 76076 141462 77779 141464
rect 76076 141460 76082 141462
rect 77713 141459 77779 141462
rect 73798 141324 73804 141388
rect 73868 141386 73874 141388
rect 74718 141386 74724 141388
rect 73868 141326 74724 141386
rect 73868 141324 73874 141326
rect 74718 141324 74724 141326
rect 74788 141324 74794 141388
rect 74534 141188 74540 141252
rect 74604 141250 74610 141252
rect 76374 141250 76380 141252
rect 74604 141190 76380 141250
rect 74604 141188 74610 141190
rect 76374 141188 76380 141190
rect 76444 141188 76450 141252
rect 137329 141114 137395 141117
rect 149105 141116 149171 141117
rect 152049 141116 152115 141117
rect 137462 141114 137468 141116
rect 137329 141112 137468 141114
rect 137329 141056 137334 141112
rect 137390 141056 137468 141112
rect 137329 141054 137468 141056
rect 137329 141051 137395 141054
rect 137462 141052 137468 141054
rect 137532 141052 137538 141116
rect 146478 141052 146484 141116
rect 146548 141114 146554 141116
rect 149054 141114 149060 141116
rect 146548 141054 149060 141114
rect 149124 141114 149171 141116
rect 149124 141112 149252 141114
rect 149166 141056 149252 141112
rect 146548 141052 146554 141054
rect 149054 141052 149060 141054
rect 149124 141054 149252 141056
rect 149124 141052 149171 141054
rect 151998 141052 152004 141116
rect 152068 141114 152115 141116
rect 207249 141114 207315 141117
rect 207566 141114 207572 141116
rect 152068 141112 152160 141114
rect 152110 141056 152160 141112
rect 152068 141054 152160 141056
rect 207249 141112 207572 141114
rect 207249 141056 207254 141112
rect 207310 141056 207572 141112
rect 207249 141054 207572 141056
rect 152068 141052 152115 141054
rect 149105 141051 149171 141052
rect 152049 141051 152115 141052
rect 207249 141051 207315 141054
rect 207566 141052 207572 141054
rect 207636 141114 207642 141116
rect 207893 141114 207959 141117
rect 207636 141112 207959 141114
rect 207636 141056 207898 141112
rect 207954 141056 207959 141112
rect 207636 141054 207959 141056
rect 207636 141052 207642 141054
rect 207893 141051 207959 141054
rect 301089 141114 301155 141117
rect 302009 141116 302075 141117
rect 301958 141114 301964 141116
rect 301089 141112 301964 141114
rect 302028 141114 302075 141116
rect 302028 141112 302120 141114
rect 301089 141056 301094 141112
rect 301150 141056 301964 141112
rect 302070 141056 302120 141112
rect 301089 141054 301964 141056
rect 301089 141051 301155 141054
rect 301958 141052 301964 141054
rect 302028 141054 302120 141056
rect 302028 141052 302075 141054
rect 302009 141051 302075 141052
rect 196209 140570 196275 140573
rect 197262 140570 197268 140572
rect 196209 140568 197268 140570
rect 196209 140512 196214 140568
rect 196270 140512 197268 140568
rect 196209 140510 197268 140512
rect 196209 140507 196275 140510
rect 197262 140508 197268 140510
rect 197332 140570 197338 140572
rect 231445 140570 231511 140573
rect 243037 140570 243103 140573
rect 197332 140568 243103 140570
rect 197332 140512 231450 140568
rect 231506 140512 243042 140568
rect 243098 140512 243103 140568
rect 197332 140510 243103 140512
rect 197332 140508 197338 140510
rect 231445 140507 231511 140510
rect 243037 140507 243103 140510
rect 137605 140436 137671 140437
rect 137605 140434 137652 140436
rect 137560 140432 137652 140434
rect 137560 140376 137610 140432
rect 137560 140374 137652 140376
rect 137605 140372 137652 140374
rect 137716 140372 137722 140436
rect 137605 140371 137671 140372
rect 231077 140026 231143 140029
rect 231670 140026 231676 140028
rect 231077 140024 231676 140026
rect 231077 139968 231082 140024
rect 231138 139968 231676 140024
rect 231077 139966 231676 139968
rect 231077 139963 231143 139966
rect 231670 139964 231676 139966
rect 231740 139964 231746 140028
rect 136869 139890 136935 139893
rect 141510 139890 141516 139892
rect 136869 139888 141516 139890
rect 136869 139832 136874 139888
rect 136930 139832 141516 139888
rect 136869 139830 141516 139832
rect 136869 139827 136935 139830
rect 141510 139828 141516 139830
rect 141580 139890 141586 139892
rect 141837 139890 141903 139893
rect 141580 139888 141903 139890
rect 141580 139832 141842 139888
rect 141898 139832 141903 139888
rect 141580 139830 141903 139832
rect 141580 139828 141586 139830
rect 141837 139827 141903 139830
rect 148185 139890 148251 139893
rect 148502 139890 148508 139892
rect 148185 139888 148508 139890
rect 148185 139832 148190 139888
rect 148246 139832 148508 139888
rect 148185 139830 148508 139832
rect 148185 139827 148251 139830
rect 148502 139828 148508 139830
rect 148572 139828 148578 139892
rect 246165 139890 246231 139893
rect 246441 139890 246507 139893
rect 251358 139890 251364 139892
rect 246165 139888 251364 139890
rect 246165 139832 246170 139888
rect 246226 139832 246446 139888
rect 246502 139832 251364 139888
rect 246165 139830 251364 139832
rect 246165 139827 246231 139830
rect 246441 139827 246507 139830
rect 251358 139828 251364 139830
rect 251428 139828 251434 139892
rect 231353 139754 231419 139757
rect 238110 139754 238116 139756
rect 231353 139752 238116 139754
rect 231353 139696 231358 139752
rect 231414 139696 238116 139752
rect 231353 139694 238116 139696
rect 231353 139691 231419 139694
rect 238110 139692 238116 139694
rect 238180 139754 238186 139756
rect 243773 139754 243839 139757
rect 238180 139752 243839 139754
rect 238180 139696 243778 139752
rect 243834 139696 243839 139752
rect 238180 139694 243839 139696
rect 238180 139692 238186 139694
rect 243773 139691 243839 139694
rect 52638 139556 52644 139620
rect 52708 139618 52714 139620
rect 53517 139618 53583 139621
rect 52708 139616 53583 139618
rect 52708 139560 53522 139616
rect 53578 139560 53583 139616
rect 52708 139558 53583 139560
rect 52708 139556 52714 139558
rect 53517 139555 53583 139558
rect 54529 139618 54595 139621
rect 245337 139620 245403 139621
rect 54662 139618 54668 139620
rect 54529 139616 54668 139618
rect 54529 139560 54534 139616
rect 54590 139560 54668 139616
rect 54529 139558 54668 139560
rect 54529 139555 54595 139558
rect 54662 139556 54668 139558
rect 54732 139556 54738 139620
rect 73798 139556 73804 139620
rect 73868 139618 73874 139620
rect 74534 139618 74540 139620
rect 73868 139558 74540 139618
rect 73868 139556 73874 139558
rect 74534 139556 74540 139558
rect 74604 139556 74610 139620
rect 245286 139618 245292 139620
rect 245210 139558 245292 139618
rect 245356 139618 245403 139620
rect 262950 139618 262956 139620
rect 245356 139616 262956 139618
rect 245398 139560 262956 139616
rect 245286 139556 245292 139558
rect 245356 139558 262956 139560
rect 245356 139556 245403 139558
rect 262950 139556 262956 139558
rect 263020 139556 263026 139620
rect 350953 139618 351019 139621
rect 351638 139618 351644 139620
rect 350953 139616 351644 139618
rect 350953 139560 350958 139616
rect 351014 139560 351644 139616
rect 350953 139558 351644 139560
rect 245337 139555 245403 139556
rect 350953 139555 351019 139558
rect 351638 139556 351644 139558
rect 351708 139556 351714 139620
rect 351822 139556 351828 139620
rect 351892 139618 351898 139620
rect 352057 139618 352123 139621
rect 351892 139616 352123 139618
rect 351892 139560 352062 139616
rect 352118 139560 352123 139616
rect 351892 139558 352123 139560
rect 351892 139556 351898 139558
rect 352057 139555 352123 139558
rect 73982 138876 73988 138940
rect 74052 138938 74058 138940
rect 74718 138938 74724 138940
rect 74052 138878 74724 138938
rect 74052 138876 74058 138878
rect 74718 138876 74724 138878
rect 74788 138876 74794 138940
rect 231353 138666 231419 138669
rect 231997 138666 232063 138669
rect 231353 138664 232063 138666
rect 231353 138608 231358 138664
rect 231414 138608 232002 138664
rect 232058 138608 232063 138664
rect 231353 138606 232063 138608
rect 231353 138603 231419 138606
rect 231997 138603 232063 138606
rect 249109 138530 249175 138533
rect 285909 138530 285975 138533
rect 287197 138530 287263 138533
rect 249109 138528 287263 138530
rect 249109 138472 249114 138528
rect 249170 138472 285914 138528
rect 285970 138472 287202 138528
rect 287258 138472 287263 138528
rect 249109 138470 287263 138472
rect 249109 138467 249175 138470
rect 285909 138467 285975 138470
rect 287197 138467 287263 138470
rect 249109 137308 249175 137309
rect 249109 137304 249156 137308
rect 249220 137306 249226 137308
rect 249109 137248 249114 137304
rect 249109 137244 249156 137248
rect 249220 137246 249266 137306
rect 249220 137244 249226 137246
rect 249109 137243 249175 137244
rect 429429 136082 429495 136085
rect 434416 136082 434896 136112
rect 429429 136080 434896 136082
rect 429429 136024 429434 136080
rect 429490 136024 434896 136080
rect 429429 136022 434896 136024
rect 429429 136019 429495 136022
rect 434416 135992 434896 136022
rect 137094 134388 137100 134452
rect 137164 134450 137170 134452
rect 137237 134450 137303 134453
rect 137164 134448 137303 134450
rect 137164 134392 137242 134448
rect 137298 134392 137303 134448
rect 137164 134390 137303 134392
rect 137164 134388 137170 134390
rect 137237 134387 137303 134390
rect 249661 134314 249727 134317
rect 283149 134314 283215 134317
rect 249661 134312 283215 134314
rect 249661 134256 249666 134312
rect 249722 134256 283154 134312
rect 283210 134256 283215 134312
rect 249661 134254 283215 134256
rect 249661 134251 249727 134254
rect 283149 134251 283215 134254
rect 249661 133092 249727 133093
rect 249661 133090 249708 133092
rect 249616 133088 249708 133090
rect 249616 133032 249666 133088
rect 249616 133030 249708 133032
rect 249661 133028 249708 133030
rect 249772 133028 249778 133092
rect 249661 133027 249727 133028
rect 136869 132954 136935 132957
rect 230985 132954 231051 132957
rect 134710 132952 136935 132954
rect 134710 132896 136874 132952
rect 136930 132896 136935 132952
rect 134710 132894 136935 132896
rect 9896 132682 10376 132712
rect 13037 132682 13103 132685
rect 9896 132680 13103 132682
rect 9896 132624 13042 132680
rect 13098 132624 13103 132680
rect 9896 132622 13103 132624
rect 9896 132592 10376 132622
rect 13037 132619 13103 132622
rect 55398 132348 55404 132412
rect 55468 132410 55474 132412
rect 55633 132410 55699 132413
rect 55468 132408 55699 132410
rect 55468 132352 55638 132408
rect 55694 132352 55699 132408
rect 55468 132350 55699 132352
rect 55468 132348 55474 132350
rect 55633 132347 55699 132350
rect 134710 132312 134770 132894
rect 136869 132891 136935 132894
rect 228734 132952 231051 132954
rect 228734 132896 230990 132952
rect 231046 132896 231051 132952
rect 228734 132894 231051 132896
rect 197630 132484 197636 132548
rect 197700 132546 197706 132548
rect 198550 132546 198556 132548
rect 197700 132486 198556 132546
rect 197700 132484 197706 132486
rect 198550 132484 198556 132486
rect 198620 132484 198626 132548
rect 228734 132312 228794 132894
rect 230985 132891 231051 132894
rect 324641 132410 324707 132413
rect 322758 132408 324707 132410
rect 322758 132352 324646 132408
rect 324702 132352 324707 132408
rect 322758 132350 324707 132352
rect 322758 132312 322818 132350
rect 324641 132347 324707 132350
rect 54110 131532 54116 131596
rect 54180 131594 54186 131596
rect 55449 131594 55515 131597
rect 54180 131592 55515 131594
rect 54180 131536 55454 131592
rect 55510 131536 55515 131592
rect 54180 131534 55515 131536
rect 54180 131532 54186 131534
rect 55449 131531 55515 131534
rect 246206 130172 246212 130236
rect 246276 130234 246282 130236
rect 246441 130234 246507 130237
rect 246276 130232 246507 130234
rect 246276 130176 246446 130232
rect 246502 130176 246507 130232
rect 246276 130174 246507 130176
rect 246276 130172 246282 130174
rect 246441 130171 246507 130174
rect 137605 129826 137671 129829
rect 231261 129826 231327 129829
rect 325469 129826 325535 129829
rect 134710 129824 137671 129826
rect 134710 129768 137610 129824
rect 137666 129768 137671 129824
rect 134710 129766 137671 129768
rect 134710 129184 134770 129766
rect 137605 129763 137671 129766
rect 228734 129824 231327 129826
rect 228734 129768 231266 129824
rect 231322 129768 231327 129824
rect 228734 129766 231327 129768
rect 228734 129184 228794 129766
rect 231261 129763 231327 129766
rect 322758 129824 325535 129826
rect 322758 129768 325474 129824
rect 325530 129768 325535 129824
rect 322758 129766 325535 129768
rect 322758 129184 322818 129766
rect 325469 129763 325535 129766
rect 38797 127514 38863 127517
rect 35748 127512 38863 127514
rect 35748 127456 38802 127512
rect 38858 127456 38863 127512
rect 35748 127454 38863 127456
rect 38797 127451 38863 127454
rect 54069 127242 54135 127245
rect 55398 127242 55404 127244
rect 54069 127240 55404 127242
rect 54069 127184 54074 127240
rect 54130 127184 55404 127240
rect 54069 127182 55404 127184
rect 54069 127179 54135 127182
rect 55398 127180 55404 127182
rect 55468 127180 55474 127244
rect 405969 126970 406035 126973
rect 409054 126970 409114 127484
rect 405969 126968 409114 126970
rect 70678 126426 70738 126940
rect 405969 126912 405974 126968
rect 406030 126912 409114 126968
rect 405969 126910 409114 126912
rect 405969 126907 406035 126910
rect 248598 126772 248604 126836
rect 248668 126834 248674 126836
rect 249702 126834 249708 126836
rect 248668 126774 249708 126834
rect 248668 126772 248674 126774
rect 249702 126772 249708 126774
rect 249772 126772 249778 126836
rect 74401 126426 74467 126429
rect 70678 126424 74467 126426
rect 70678 126368 74406 126424
rect 74462 126368 74467 126424
rect 70678 126366 74467 126368
rect 74401 126363 74467 126366
rect 51217 126290 51283 126293
rect 356197 126290 356263 126293
rect 427313 126290 427379 126293
rect 51217 126288 55068 126290
rect 16073 126154 16139 126157
rect 19894 126154 19954 126260
rect 51217 126232 51222 126288
rect 51278 126232 55068 126288
rect 51217 126230 55068 126232
rect 352780 126288 356263 126290
rect 352780 126232 356202 126288
rect 356258 126232 356263 126288
rect 352780 126230 356263 126232
rect 424724 126288 427379 126290
rect 424724 126232 427318 126288
rect 427374 126232 427379 126288
rect 424724 126230 427379 126232
rect 51217 126227 51283 126230
rect 356197 126227 356263 126230
rect 427313 126227 427379 126230
rect 16073 126152 19954 126154
rect 16073 126096 16078 126152
rect 16134 126096 19954 126152
rect 16073 126094 19954 126096
rect 16073 126091 16139 126094
rect 134710 126018 134770 126052
rect 137053 126018 137119 126021
rect 134710 126016 137119 126018
rect 134710 125960 137058 126016
rect 137114 125960 137119 126016
rect 134710 125958 137119 125960
rect 228734 126018 228794 126052
rect 231077 126018 231143 126021
rect 228734 126016 231143 126018
rect 228734 125960 231082 126016
rect 231138 125960 231143 126016
rect 228734 125958 231143 125960
rect 322758 126018 322818 126056
rect 325377 126018 325443 126021
rect 322758 126016 325443 126018
rect 322758 125960 325382 126016
rect 325438 125960 325443 126016
rect 322758 125958 325443 125960
rect 137053 125955 137119 125958
rect 231077 125955 231143 125958
rect 325377 125955 325443 125958
rect 38245 125610 38311 125613
rect 35718 125608 38311 125610
rect 35718 125552 38250 125608
rect 38306 125552 38311 125608
rect 35718 125550 38311 125552
rect 35718 125104 35778 125550
rect 38245 125547 38311 125550
rect 405969 125610 406035 125613
rect 405969 125608 408930 125610
rect 405969 125552 405974 125608
rect 406030 125552 408930 125608
rect 405969 125550 408930 125552
rect 405969 125547 406035 125550
rect 84662 125482 85060 125542
rect 178318 125482 178900 125542
rect 272342 125482 272924 125542
rect 81669 125474 81735 125477
rect 84662 125474 84722 125482
rect 81669 125472 84722 125474
rect 81669 125416 81674 125472
rect 81730 125416 84722 125472
rect 81669 125414 84722 125416
rect 175509 125474 175575 125477
rect 178318 125474 178378 125482
rect 175509 125472 178378 125474
rect 175509 125416 175514 125472
rect 175570 125416 178378 125472
rect 175509 125414 178378 125416
rect 270361 125474 270427 125477
rect 272342 125474 272402 125482
rect 270361 125472 272402 125474
rect 270361 125416 270366 125472
rect 270422 125416 272402 125472
rect 270361 125414 272402 125416
rect 81669 125411 81735 125414
rect 175509 125411 175575 125414
rect 270361 125411 270427 125414
rect 408870 125036 408930 125550
rect 322750 124052 322756 124116
rect 322820 124114 322826 124116
rect 323169 124114 323235 124117
rect 322820 124112 323235 124114
rect 322820 124056 323174 124112
rect 323230 124056 323235 124112
rect 322820 124054 323235 124056
rect 322820 124052 322826 124054
rect 323169 124051 323235 124054
rect 428693 123978 428759 123981
rect 434416 123978 434896 124008
rect 428693 123976 434896 123978
rect 428693 123920 428698 123976
rect 428754 123920 434896 123976
rect 428693 123918 434896 123920
rect 428693 123915 428759 123918
rect 434416 123888 434896 123918
rect 136961 123298 137027 123301
rect 134710 123296 137027 123298
rect 38797 122754 38863 122757
rect 35534 122752 38863 122754
rect 35534 122696 38802 122752
rect 38858 122696 38863 122752
rect 35534 122694 38863 122696
rect 35534 122520 35594 122694
rect 38797 122691 38863 122694
rect 53149 122754 53215 122757
rect 54110 122754 54116 122756
rect 53149 122752 54116 122754
rect 53149 122696 53154 122752
rect 53210 122696 54116 122752
rect 53149 122694 54116 122696
rect 53149 122691 53215 122694
rect 54110 122692 54116 122694
rect 54180 122692 54186 122756
rect 70678 122754 70738 123268
rect 134710 123240 136966 123296
rect 137022 123240 137027 123296
rect 134710 123238 137027 123240
rect 134710 122928 134770 123238
rect 136961 123235 137027 123238
rect 323169 122958 323235 122961
rect 322788 122956 323235 122958
rect 74125 122754 74191 122757
rect 70678 122752 74191 122754
rect 70678 122696 74130 122752
rect 74186 122696 74191 122752
rect 70678 122694 74191 122696
rect 74125 122691 74191 122694
rect 228734 122618 228794 122924
rect 322788 122900 323174 122956
rect 323230 122900 323235 122956
rect 322788 122898 323235 122900
rect 323169 122895 323235 122898
rect 231997 122618 232063 122621
rect 242710 122618 242716 122620
rect 228734 122616 242716 122618
rect 228734 122560 232002 122616
rect 232058 122560 242716 122616
rect 228734 122558 242716 122560
rect 231997 122555 232063 122558
rect 242710 122556 242716 122558
rect 242780 122556 242786 122620
rect 258718 122556 258724 122620
rect 258788 122618 258794 122620
rect 260333 122618 260399 122621
rect 272702 122618 272708 122620
rect 258788 122616 272708 122618
rect 258788 122560 260338 122616
rect 260394 122560 272708 122616
rect 258788 122558 272708 122560
rect 258788 122556 258794 122558
rect 260333 122555 260399 122558
rect 272702 122556 272708 122558
rect 272772 122556 272778 122620
rect 405969 122618 406035 122621
rect 405969 122616 408930 122618
rect 405969 122560 405974 122616
rect 406030 122560 408930 122616
rect 405969 122558 408930 122560
rect 405969 122555 406035 122558
rect 408870 122452 408930 122558
rect 144229 122346 144295 122349
rect 148686 122346 148692 122348
rect 144229 122344 148692 122346
rect 144229 122288 144234 122344
rect 144290 122288 148692 122344
rect 144229 122286 148692 122288
rect 144229 122283 144295 122286
rect 148686 122284 148692 122286
rect 148756 122284 148762 122348
rect 148870 122148 148876 122212
rect 148940 122148 148946 122212
rect 240369 122210 240435 122213
rect 334209 122210 334275 122213
rect 240369 122208 242932 122210
rect 240369 122152 240374 122208
rect 240430 122152 242932 122208
rect 240369 122150 242932 122152
rect 334209 122208 336956 122210
rect 334209 122152 334214 122208
rect 334270 122152 336956 122208
rect 334209 122150 336956 122152
rect 240369 122147 240435 122150
rect 334209 122147 334275 122150
rect 9896 121938 10376 121968
rect 13221 121938 13287 121941
rect 9896 121936 13287 121938
rect 9896 121880 13226 121936
rect 13282 121880 13287 121936
rect 9896 121878 13287 121880
rect 9896 121848 10376 121878
rect 13221 121875 13287 121878
rect 52597 121258 52663 121261
rect 356197 121258 356263 121261
rect 427497 121258 427563 121261
rect 52597 121256 55068 121258
rect 16257 120714 16323 120717
rect 19894 120714 19954 121228
rect 52597 121200 52602 121256
rect 52658 121200 55068 121256
rect 52597 121198 55068 121200
rect 352780 121256 356263 121258
rect 352780 121200 356202 121256
rect 356258 121200 356263 121256
rect 352780 121198 356263 121200
rect 424724 121256 427563 121258
rect 424724 121200 427502 121256
rect 427558 121200 427563 121256
rect 424724 121198 427563 121200
rect 52597 121195 52663 121198
rect 356197 121195 356263 121198
rect 427497 121195 427563 121198
rect 16257 120712 19954 120714
rect 16257 120656 16262 120712
rect 16318 120656 19954 120712
rect 16257 120654 19954 120656
rect 16257 120651 16323 120654
rect 73389 120578 73455 120581
rect 74309 120578 74375 120581
rect 73389 120576 74375 120578
rect 73389 120520 73394 120576
rect 73450 120520 74314 120576
rect 74370 120520 74375 120576
rect 73389 120518 74375 120520
rect 73389 120515 73455 120518
rect 74309 120515 74375 120518
rect 405969 120578 406035 120581
rect 405969 120576 408930 120578
rect 405969 120520 405974 120576
rect 406030 120520 408930 120576
rect 405969 120518 408930 120520
rect 405969 120515 406035 120518
rect 136869 120442 136935 120445
rect 230985 120442 231051 120445
rect 134710 120440 136935 120442
rect 134710 120384 136874 120440
rect 136930 120384 136935 120440
rect 134710 120382 136935 120384
rect 38797 120306 38863 120309
rect 35718 120304 38863 120306
rect 35718 120248 38802 120304
rect 38858 120248 38863 120304
rect 35718 120246 38863 120248
rect 35718 120072 35778 120246
rect 38797 120243 38863 120246
rect 134710 119800 134770 120382
rect 136869 120379 136935 120382
rect 228734 120440 231051 120442
rect 228734 120384 230990 120440
rect 231046 120384 231051 120440
rect 228734 120382 231051 120384
rect 228734 119800 228794 120382
rect 230985 120379 231051 120382
rect 408870 120004 408930 120518
rect 324549 119898 324615 119901
rect 322758 119896 324615 119898
rect 322758 119840 324554 119896
rect 324610 119840 324615 119896
rect 322758 119838 324615 119840
rect 322758 119800 322818 119838
rect 324549 119835 324615 119838
rect 73389 119762 73455 119765
rect 70862 119760 73455 119762
rect 70862 119704 73394 119760
rect 73450 119704 73455 119760
rect 70862 119702 73455 119704
rect 70862 119596 70922 119702
rect 73389 119699 73455 119702
rect 167873 118810 167939 118813
rect 261161 118810 261227 118813
rect 164732 118808 167939 118810
rect 164732 118752 167878 118808
rect 167934 118752 167939 118808
rect 164732 118750 167939 118752
rect 258756 118808 261227 118810
rect 258756 118752 261166 118808
rect 261222 118752 261227 118808
rect 258756 118750 261227 118752
rect 167873 118747 167939 118750
rect 261161 118747 261227 118750
rect 177574 117796 177580 117860
rect 177644 117858 177650 117860
rect 178678 117858 178684 117860
rect 177644 117798 178684 117858
rect 177644 117796 177650 117798
rect 178678 117796 178684 117798
rect 178748 117796 178754 117860
rect 38245 117586 38311 117589
rect 35748 117584 38311 117586
rect 35748 117528 38250 117584
rect 38306 117528 38311 117584
rect 35748 117526 38311 117528
rect 38245 117523 38311 117526
rect 405969 117450 406035 117453
rect 409054 117450 409114 117556
rect 405969 117448 409114 117450
rect 405969 117392 405974 117448
rect 406030 117392 409114 117448
rect 405969 117390 409114 117392
rect 405969 117387 406035 117390
rect 325469 117314 325535 117317
rect 322758 117312 325535 117314
rect 322758 117256 325474 117312
rect 325530 117256 325535 117312
rect 322758 117254 325535 117256
rect 54069 117178 54135 117181
rect 54662 117178 54668 117180
rect 54069 117176 54668 117178
rect 54069 117120 54074 117176
rect 54130 117120 54668 117176
rect 54069 117118 54668 117120
rect 54069 117115 54135 117118
rect 54662 117116 54668 117118
rect 54732 117116 54738 117180
rect 322758 116672 322818 117254
rect 325469 117251 325535 117254
rect 134710 116634 134770 116668
rect 136910 116634 136916 116636
rect 134710 116574 136916 116634
rect 136910 116572 136916 116574
rect 136980 116572 136986 116636
rect 138198 116572 138204 116636
rect 138268 116634 138274 116636
rect 145006 116634 145012 116636
rect 138268 116574 145012 116634
rect 138268 116572 138274 116574
rect 145006 116572 145012 116574
rect 145076 116572 145082 116636
rect 228734 116500 228794 116668
rect 228726 116436 228732 116500
rect 228796 116436 228802 116500
rect 51217 116226 51283 116229
rect 73481 116226 73547 116229
rect 356197 116226 356263 116229
rect 428693 116226 428759 116229
rect 51217 116224 55068 116226
rect 16441 115138 16507 115141
rect 19894 115138 19954 116196
rect 51217 116168 51222 116224
rect 51278 116168 55068 116224
rect 51217 116166 55068 116168
rect 70862 116224 73547 116226
rect 70862 116168 73486 116224
rect 73542 116168 73547 116224
rect 70862 116166 73547 116168
rect 352780 116224 356263 116226
rect 352780 116168 356202 116224
rect 356258 116168 356263 116224
rect 352780 116166 356263 116168
rect 424724 116224 428759 116226
rect 424724 116168 428698 116224
rect 428754 116168 428759 116224
rect 424724 116166 428759 116168
rect 51217 116163 51283 116166
rect 70862 116060 70922 116166
rect 73481 116163 73547 116166
rect 356197 116163 356263 116166
rect 428693 116163 428759 116166
rect 369813 115274 369879 115277
rect 369813 115272 369922 115274
rect 369813 115216 369818 115272
rect 369874 115216 369922 115272
rect 369813 115211 369922 115216
rect 16441 115136 19954 115138
rect 16441 115080 16446 115136
rect 16502 115080 19954 115136
rect 16441 115078 19954 115080
rect 369862 115141 369922 115211
rect 369862 115136 369971 115141
rect 369862 115080 369910 115136
rect 369966 115080 369971 115136
rect 369862 115078 369971 115080
rect 16441 115075 16507 115078
rect 369905 115075 369971 115078
rect 38797 115002 38863 115005
rect 35748 115000 38863 115002
rect 35748 114944 38802 115000
rect 38858 114944 38863 115000
rect 35748 114942 38863 114944
rect 38797 114939 38863 114942
rect 177574 114940 177580 115004
rect 177644 114940 177650 115004
rect 177582 114869 177642 114940
rect 177582 114864 177691 114869
rect 177582 114808 177630 114864
rect 177686 114808 177691 114864
rect 177582 114806 177691 114808
rect 177625 114803 177691 114806
rect 405969 114866 406035 114869
rect 409054 114866 409114 114972
rect 405969 114864 409114 114866
rect 405969 114808 405974 114864
rect 406030 114808 409114 114864
rect 405969 114806 409114 114808
rect 405969 114803 406035 114806
rect 147357 113642 147423 113645
rect 147766 113642 147772 113644
rect 147357 113640 147772 113642
rect 147357 113584 147362 113640
rect 147418 113584 147772 113640
rect 147357 113582 147772 113584
rect 147357 113579 147423 113582
rect 147766 113580 147772 113582
rect 147836 113580 147842 113644
rect 324549 113642 324615 113645
rect 322758 113640 324615 113642
rect 322758 113584 324554 113640
rect 324610 113584 324615 113640
rect 322758 113582 324615 113584
rect 322758 113544 322818 113582
rect 324549 113579 324615 113582
rect 134710 113234 134770 113540
rect 136869 113234 136935 113237
rect 134710 113232 136935 113234
rect 134710 113176 136874 113232
rect 136930 113176 136935 113232
rect 134710 113174 136935 113176
rect 136869 113171 136935 113174
rect 52137 113098 52203 113101
rect 52638 113098 52644 113100
rect 52137 113096 52644 113098
rect 52137 113040 52142 113096
rect 52198 113040 52644 113096
rect 52137 113038 52644 113040
rect 52137 113035 52203 113038
rect 52638 113036 52644 113038
rect 52708 113036 52714 113100
rect 228734 112962 228794 113540
rect 230750 112962 230756 112964
rect 228734 112902 230756 112962
rect 230750 112900 230756 112902
rect 230820 112900 230826 112964
rect 38797 112826 38863 112829
rect 73430 112826 73436 112828
rect 35534 112824 38863 112826
rect 35534 112768 38802 112824
rect 38858 112768 38863 112824
rect 35534 112766 38863 112768
rect 35534 112592 35594 112766
rect 38797 112763 38863 112766
rect 70862 112766 73436 112826
rect 70862 112388 70922 112766
rect 73430 112764 73436 112766
rect 73500 112826 73506 112828
rect 73573 112826 73639 112829
rect 73500 112824 73639 112826
rect 73500 112768 73578 112824
rect 73634 112768 73639 112824
rect 73500 112766 73639 112768
rect 73500 112764 73506 112766
rect 73573 112763 73639 112766
rect 405969 112690 406035 112693
rect 405969 112688 408930 112690
rect 405969 112632 405974 112688
rect 406030 112632 408930 112688
rect 405969 112630 408930 112632
rect 405969 112627 406035 112630
rect 147357 112554 147423 112557
rect 147766 112554 147772 112556
rect 147357 112552 147772 112554
rect 147357 112496 147362 112552
rect 147418 112496 147772 112552
rect 147357 112494 147772 112496
rect 147357 112491 147423 112494
rect 147766 112492 147772 112494
rect 147836 112492 147842 112556
rect 408870 112524 408930 112630
rect 429429 111874 429495 111877
rect 434416 111874 434896 111904
rect 429429 111872 434896 111874
rect 429429 111816 429434 111872
rect 429490 111816 434896 111872
rect 429429 111814 434896 111816
rect 429429 111811 429495 111814
rect 434416 111784 434896 111814
rect 52597 111330 52663 111333
rect 356197 111330 356263 111333
rect 427589 111330 427655 111333
rect 52597 111328 55068 111330
rect 9896 111194 10376 111224
rect 12853 111194 12919 111197
rect 9896 111192 12919 111194
rect 9896 111136 12858 111192
rect 12914 111136 12919 111192
rect 9896 111134 12919 111136
rect 9896 111104 10376 111134
rect 12853 111131 12919 111134
rect 16533 111058 16599 111061
rect 19894 111058 19954 111300
rect 52597 111272 52602 111328
rect 52658 111272 55068 111328
rect 52597 111270 55068 111272
rect 352780 111328 356263 111330
rect 352780 111272 356202 111328
rect 356258 111272 356263 111328
rect 352780 111270 356263 111272
rect 424724 111328 427655 111330
rect 424724 111272 427594 111328
rect 427650 111272 427655 111328
rect 424724 111270 427655 111272
rect 52597 111267 52663 111270
rect 356197 111267 356263 111270
rect 427589 111267 427655 111270
rect 16533 111056 19954 111058
rect 16533 111000 16538 111056
rect 16594 111000 19954 111056
rect 16533 110998 19954 111000
rect 16533 110995 16599 110998
rect 78030 110860 78036 110924
rect 78100 110922 78106 110924
rect 78173 110922 78239 110925
rect 231629 110922 231695 110925
rect 325285 110922 325351 110925
rect 78100 110920 78239 110922
rect 78100 110864 78178 110920
rect 78234 110864 78239 110920
rect 78100 110862 78239 110864
rect 78100 110860 78106 110862
rect 78173 110859 78239 110862
rect 228734 110920 231695 110922
rect 228734 110864 231634 110920
rect 231690 110864 231695 110920
rect 228734 110862 231695 110864
rect 136869 110786 136935 110789
rect 134710 110784 136935 110786
rect 134710 110728 136874 110784
rect 136930 110728 136935 110784
rect 134710 110726 136935 110728
rect 38245 110514 38311 110517
rect 35718 110512 38311 110514
rect 35718 110456 38250 110512
rect 38306 110456 38311 110512
rect 35718 110454 38311 110456
rect 35718 110144 35778 110454
rect 38245 110451 38311 110454
rect 134710 109836 134770 110726
rect 136869 110723 136935 110726
rect 228734 110416 228794 110862
rect 231629 110859 231695 110862
rect 322758 110920 325351 110922
rect 322758 110864 325290 110920
rect 325346 110864 325351 110920
rect 322758 110862 325351 110864
rect 240093 109836 240159 109837
rect 322758 109836 322818 110862
rect 325285 110859 325351 110862
rect 406061 110650 406127 110653
rect 406061 110648 408930 110650
rect 406061 110592 406066 110648
rect 406122 110592 408930 110648
rect 406061 110590 408930 110592
rect 406061 110587 406127 110590
rect 408870 110076 408930 110590
rect 134702 109772 134708 109836
rect 134772 109772 134778 109836
rect 240093 109834 240140 109836
rect 240048 109832 240140 109834
rect 240048 109776 240098 109832
rect 240048 109774 240140 109776
rect 240093 109772 240140 109774
rect 240204 109772 240210 109836
rect 322750 109772 322756 109836
rect 322820 109772 322826 109836
rect 240093 109771 240159 109772
rect 78173 109698 78239 109701
rect 84654 109698 84660 109700
rect 78173 109696 84660 109698
rect 78173 109640 78178 109696
rect 78234 109640 84660 109696
rect 78173 109638 84660 109640
rect 78173 109635 78239 109638
rect 84654 109636 84660 109638
rect 84724 109636 84730 109700
rect 73665 109562 73731 109565
rect 74534 109562 74540 109564
rect 73665 109560 74540 109562
rect 73665 109504 73670 109560
rect 73726 109504 74540 109560
rect 73665 109502 74540 109504
rect 73665 109499 73731 109502
rect 74534 109500 74540 109502
rect 74604 109500 74610 109564
rect 73665 108882 73731 108885
rect 70862 108880 73731 108882
rect 70862 108824 73670 108880
rect 73726 108824 73731 108880
rect 70862 108822 73731 108824
rect 70862 108716 70922 108822
rect 73665 108819 73731 108822
rect 81669 108882 81735 108885
rect 143953 108882 144019 108885
rect 148686 108882 148692 108884
rect 81669 108880 84722 108882
rect 81669 108824 81674 108880
rect 81730 108824 84722 108880
rect 81669 108822 84722 108824
rect 81669 108819 81735 108822
rect 84662 108810 84722 108822
rect 143953 108880 148692 108882
rect 143953 108824 143958 108880
rect 144014 108824 148692 108880
rect 143953 108822 148692 108824
rect 143953 108819 144019 108822
rect 148686 108820 148692 108822
rect 148756 108820 148762 108884
rect 148870 108820 148876 108884
rect 148940 108820 148946 108884
rect 174865 108882 174931 108885
rect 240369 108882 240435 108885
rect 268613 108882 268679 108885
rect 334209 108882 334275 108885
rect 174865 108880 178378 108882
rect 174865 108824 174870 108880
rect 174926 108824 178378 108880
rect 174865 108822 178378 108824
rect 174865 108819 174931 108822
rect 178318 108814 178378 108822
rect 240369 108880 242932 108882
rect 240369 108824 240374 108880
rect 240430 108824 242932 108880
rect 240369 108822 242932 108824
rect 268613 108880 272402 108882
rect 268613 108824 268618 108880
rect 268674 108824 272402 108880
rect 268613 108822 272402 108824
rect 240369 108819 240435 108822
rect 268613 108819 268679 108822
rect 272342 108814 272402 108822
rect 334209 108880 336956 108882
rect 334209 108824 334214 108880
rect 334270 108824 336956 108880
rect 334209 108822 336956 108824
rect 334209 108819 334275 108822
rect 84662 108750 85060 108810
rect 178318 108754 178900 108814
rect 272342 108754 272924 108814
rect 405969 107658 406035 107661
rect 405969 107656 408930 107658
rect 405969 107600 405974 107656
rect 406030 107600 408930 107656
rect 405969 107598 408930 107600
rect 405969 107595 406035 107598
rect 38797 107522 38863 107525
rect 35748 107520 38863 107522
rect 35748 107464 38802 107520
rect 38858 107464 38863 107520
rect 408870 107492 408930 107598
rect 35748 107462 38863 107464
rect 38797 107459 38863 107462
rect 230893 107388 230959 107389
rect 230893 107386 230940 107388
rect 228734 107384 230940 107386
rect 231004 107386 231010 107388
rect 228734 107328 230898 107384
rect 228734 107326 230940 107328
rect 134710 107114 134770 107284
rect 136910 107114 136916 107116
rect 134710 107054 136916 107114
rect 136910 107052 136916 107054
rect 136980 107052 136986 107116
rect 228734 106844 228794 107326
rect 230893 107324 230940 107326
rect 231004 107326 231086 107386
rect 231004 107324 231010 107326
rect 230893 107323 230959 107324
rect 228726 106780 228732 106844
rect 228796 106780 228802 106844
rect 322758 106842 322818 107288
rect 324641 106842 324707 106845
rect 322758 106840 324707 106842
rect 322758 106784 324646 106840
rect 324702 106784 324707 106840
rect 322758 106782 324707 106784
rect 324641 106779 324707 106782
rect 18097 106298 18163 106301
rect 52597 106298 52663 106301
rect 356197 106298 356263 106301
rect 427681 106298 427747 106301
rect 18097 106296 19924 106298
rect 18097 106240 18102 106296
rect 18158 106240 19924 106296
rect 18097 106238 19924 106240
rect 52597 106296 55068 106298
rect 52597 106240 52602 106296
rect 52658 106240 55068 106296
rect 52597 106238 55068 106240
rect 352780 106296 356263 106298
rect 352780 106240 356202 106296
rect 356258 106240 356263 106296
rect 352780 106238 356263 106240
rect 424724 106296 427747 106298
rect 424724 106240 427686 106296
rect 427742 106240 427747 106296
rect 424724 106238 427747 106240
rect 18097 106235 18163 106238
rect 52597 106235 52663 106238
rect 356197 106235 356263 106238
rect 427681 106235 427747 106238
rect 369905 105618 369971 105621
rect 369862 105616 369971 105618
rect 369862 105560 369910 105616
rect 369966 105560 369971 105616
rect 369862 105555 369971 105560
rect 369862 105485 369922 105555
rect 74217 105482 74283 105485
rect 74036 105480 74283 105482
rect 74036 105424 74222 105480
rect 74278 105424 74283 105480
rect 74036 105422 74283 105424
rect 38797 105346 38863 105349
rect 74036 105346 74096 105422
rect 74217 105419 74283 105422
rect 177625 105482 177691 105485
rect 177758 105482 177764 105484
rect 177625 105480 177764 105482
rect 177625 105424 177630 105480
rect 177686 105424 177764 105480
rect 177625 105422 177764 105424
rect 177625 105419 177691 105422
rect 177758 105420 177764 105422
rect 177828 105420 177834 105484
rect 242158 105420 242164 105484
rect 242228 105482 242234 105484
rect 242526 105482 242532 105484
rect 242228 105422 242532 105482
rect 242228 105420 242234 105422
rect 242526 105420 242532 105422
rect 242596 105420 242602 105484
rect 369813 105480 369922 105485
rect 369813 105424 369818 105480
rect 369874 105424 369922 105480
rect 369813 105422 369922 105424
rect 369813 105419 369879 105422
rect 74217 105346 74283 105349
rect 35534 105344 38863 105346
rect 35534 105288 38802 105344
rect 38858 105288 38863 105344
rect 35534 105286 38863 105288
rect 35534 105112 35594 105286
rect 38797 105283 38863 105286
rect 70862 105344 74283 105346
rect 70862 105288 74222 105344
rect 74278 105288 74283 105344
rect 70862 105286 74283 105288
rect 70862 105044 70922 105286
rect 74217 105283 74283 105286
rect 405969 105346 406035 105349
rect 405969 105344 408930 105346
rect 405969 105288 405974 105344
rect 406030 105288 408930 105344
rect 405969 105286 408930 105288
rect 405969 105283 406035 105286
rect 352793 105212 352859 105213
rect 352742 105148 352748 105212
rect 352812 105210 352859 105212
rect 352812 105208 352904 105210
rect 352854 105152 352904 105208
rect 352812 105150 352904 105152
rect 352812 105148 352859 105150
rect 352793 105147 352859 105148
rect 408870 105044 408930 105286
rect 134710 104122 134770 104156
rect 137789 104122 137855 104125
rect 134710 104120 137855 104122
rect 134710 104064 137794 104120
rect 137850 104064 137855 104120
rect 134710 104062 137855 104064
rect 228734 104122 228794 104156
rect 230709 104122 230775 104125
rect 228734 104120 230775 104122
rect 228734 104064 230714 104120
rect 230770 104064 230775 104120
rect 228734 104062 230775 104064
rect 322758 104122 322818 104160
rect 324549 104122 324615 104125
rect 322758 104120 324615 104122
rect 322758 104064 324554 104120
rect 324610 104064 324615 104120
rect 322758 104062 324615 104064
rect 137789 104059 137855 104062
rect 230709 104059 230775 104062
rect 324549 104059 324615 104062
rect 38613 102490 38679 102493
rect 35748 102488 38679 102490
rect 35748 102432 38618 102488
rect 38674 102432 38679 102488
rect 35748 102430 38679 102432
rect 38613 102427 38679 102430
rect 405969 102218 406035 102221
rect 409054 102218 409114 102460
rect 405969 102216 409114 102218
rect 405969 102160 405974 102216
rect 406030 102160 409114 102216
rect 405969 102158 409114 102160
rect 405969 102155 406035 102158
rect 74166 102082 74172 102084
rect 70862 102022 74172 102082
rect 70862 101508 70922 102022
rect 74166 102020 74172 102022
rect 74236 102020 74242 102084
rect 230801 101674 230867 101677
rect 228734 101672 230867 101674
rect 228734 101616 230806 101672
rect 230862 101616 230867 101672
rect 228734 101614 230867 101616
rect 17453 101266 17519 101269
rect 52597 101266 52663 101269
rect 17453 101264 19924 101266
rect 17453 101208 17458 101264
rect 17514 101208 19924 101264
rect 17453 101206 19924 101208
rect 52597 101264 55068 101266
rect 52597 101208 52602 101264
rect 52658 101208 55068 101264
rect 52597 101206 55068 101208
rect 17453 101203 17519 101206
rect 52597 101203 52663 101206
rect 134710 100994 134770 101028
rect 136910 100994 136916 100996
rect 134710 100934 136916 100994
rect 136910 100932 136916 100934
rect 136980 100932 136986 100996
rect 228734 100860 228794 101614
rect 230801 101611 230867 101614
rect 356197 101266 356263 101269
rect 427405 101266 427471 101269
rect 352780 101264 356263 101266
rect 352780 101208 356202 101264
rect 356258 101208 356263 101264
rect 352780 101206 356263 101208
rect 424724 101264 427471 101266
rect 424724 101208 427410 101264
rect 427466 101208 427471 101264
rect 424724 101206 427471 101208
rect 356197 101203 356263 101206
rect 427405 101203 427471 101206
rect 228726 100796 228732 100860
rect 228796 100796 228802 100860
rect 164878 100660 164884 100724
rect 164948 100722 164954 100724
rect 178126 100722 178132 100724
rect 164948 100662 178132 100722
rect 164948 100660 164954 100662
rect 178126 100660 178132 100662
rect 178196 100660 178202 100724
rect 258902 100660 258908 100724
rect 258972 100722 258978 100724
rect 272702 100722 272708 100724
rect 258972 100662 272708 100722
rect 258972 100660 258978 100662
rect 272702 100660 272708 100662
rect 272772 100660 272778 100724
rect 9896 100450 10376 100480
rect 12853 100450 12919 100453
rect 322758 100452 322818 101032
rect 323118 100932 323124 100996
rect 323188 100994 323194 100996
rect 324641 100994 324707 100997
rect 323188 100992 324707 100994
rect 323188 100936 324646 100992
rect 324702 100936 324707 100992
rect 323188 100934 324707 100936
rect 323188 100932 323194 100934
rect 324641 100931 324707 100934
rect 405969 100586 406035 100589
rect 405969 100584 408930 100586
rect 405969 100528 405974 100584
rect 406030 100528 408930 100584
rect 405969 100526 408930 100528
rect 405969 100523 406035 100526
rect 322750 100450 322756 100452
rect 9896 100448 12919 100450
rect 9896 100392 12858 100448
rect 12914 100392 12919 100448
rect 9896 100390 12919 100392
rect 322628 100390 322756 100450
rect 9896 100360 10376 100390
rect 12853 100387 12919 100390
rect 322750 100388 322756 100390
rect 322820 100450 322826 100452
rect 325285 100450 325351 100453
rect 322820 100448 325351 100450
rect 322820 100392 325290 100448
rect 325346 100392 325351 100448
rect 322820 100390 325351 100392
rect 322820 100388 322826 100390
rect 325285 100387 325351 100390
rect 38797 100314 38863 100317
rect 35718 100312 38863 100314
rect 35718 100256 38802 100312
rect 38858 100256 38863 100312
rect 35718 100254 38863 100256
rect 35718 100080 35778 100254
rect 38797 100251 38863 100254
rect 176102 100252 176108 100316
rect 176172 100314 176178 100316
rect 177022 100314 177028 100316
rect 176172 100254 177028 100314
rect 176172 100252 176178 100254
rect 177022 100252 177028 100254
rect 177092 100252 177098 100316
rect 263134 100252 263140 100316
rect 263204 100314 263210 100316
rect 264422 100314 264428 100316
rect 263204 100254 264428 100314
rect 263204 100252 263210 100254
rect 264422 100252 264428 100254
rect 264492 100252 264498 100316
rect 408870 100012 408930 100526
rect 429429 99770 429495 99773
rect 434416 99770 434896 99800
rect 429429 99768 434896 99770
rect 429429 99712 429434 99768
rect 429490 99712 434896 99768
rect 429429 99710 434896 99712
rect 429429 99707 429495 99710
rect 434416 99680 434896 99710
rect 168241 98818 168307 98821
rect 263093 98818 263159 98821
rect 164732 98816 168307 98818
rect 164732 98760 168246 98816
rect 168302 98760 168307 98816
rect 164732 98758 168307 98760
rect 258756 98816 263159 98818
rect 258756 98760 263098 98816
rect 263154 98760 263159 98816
rect 258756 98758 263159 98760
rect 168241 98755 168307 98758
rect 263093 98755 263159 98758
rect 137513 98546 137579 98549
rect 134710 98544 137579 98546
rect 134710 98488 137518 98544
rect 137574 98488 137579 98544
rect 134710 98486 137579 98488
rect 73614 98274 73620 98276
rect 70862 98214 73620 98274
rect 38797 97866 38863 97869
rect 35534 97864 38863 97866
rect 35534 97808 38802 97864
rect 38858 97808 38863 97864
rect 70862 97836 70922 98214
rect 73614 98212 73620 98214
rect 73684 98212 73690 98276
rect 134710 97904 134770 98486
rect 137513 98483 137579 98486
rect 231353 98274 231419 98277
rect 325193 98274 325259 98277
rect 228734 98272 231419 98274
rect 228734 98216 231358 98272
rect 231414 98216 231419 98272
rect 228734 98214 231419 98216
rect 228734 97904 228794 98214
rect 231353 98211 231419 98214
rect 322758 98272 325259 98274
rect 322758 98216 325198 98272
rect 325254 98216 325259 98272
rect 322758 98214 325259 98216
rect 322758 97904 322818 98214
rect 325193 98211 325259 98214
rect 35534 97806 38863 97808
rect 35534 97632 35594 97806
rect 38797 97803 38863 97806
rect 405969 97730 406035 97733
rect 405969 97728 408930 97730
rect 405969 97672 405974 97728
rect 406030 97672 408930 97728
rect 405969 97670 408930 97672
rect 405969 97667 406035 97670
rect 352793 97596 352859 97597
rect 352742 97594 352748 97596
rect 352702 97534 352748 97594
rect 352812 97592 352859 97596
rect 352854 97536 352859 97592
rect 408870 97564 408930 97670
rect 352742 97532 352748 97534
rect 352812 97532 352859 97536
rect 352793 97531 352859 97532
rect 18097 96234 18163 96237
rect 52597 96234 52663 96237
rect 356197 96234 356263 96237
rect 427221 96234 427287 96237
rect 18097 96232 19924 96234
rect 18097 96176 18102 96232
rect 18158 96176 19924 96232
rect 18097 96174 19924 96176
rect 52597 96232 55068 96234
rect 52597 96176 52602 96232
rect 52658 96176 55068 96232
rect 52597 96174 55068 96176
rect 352780 96232 356263 96234
rect 352780 96176 356202 96232
rect 356258 96176 356263 96232
rect 352780 96174 356263 96176
rect 424724 96232 427287 96234
rect 424724 96176 427226 96232
rect 427282 96176 427287 96232
rect 424724 96174 427287 96176
rect 18097 96171 18163 96174
rect 52597 96171 52663 96174
rect 356197 96171 356263 96174
rect 427221 96171 427287 96174
rect 144413 95554 144479 95557
rect 148686 95554 148692 95556
rect 144413 95552 148692 95554
rect 144413 95496 144418 95552
rect 144474 95496 148692 95552
rect 144413 95494 148692 95496
rect 144413 95491 144479 95494
rect 148686 95492 148692 95494
rect 148756 95492 148762 95556
rect 148870 95492 148876 95556
rect 148940 95492 148946 95556
rect 240369 95554 240435 95557
rect 334209 95554 334275 95557
rect 405969 95554 406035 95557
rect 240369 95552 242932 95554
rect 240369 95496 240374 95552
rect 240430 95496 242932 95552
rect 240369 95494 242932 95496
rect 334209 95552 336956 95554
rect 334209 95496 334214 95552
rect 334270 95496 336956 95552
rect 334209 95494 336956 95496
rect 405969 95552 408930 95554
rect 405969 95496 405974 95552
rect 406030 95496 408930 95552
rect 405969 95494 408930 95496
rect 240369 95491 240435 95494
rect 334209 95491 334275 95494
rect 405969 95491 406035 95494
rect 38061 95418 38127 95421
rect 35718 95416 38127 95418
rect 35718 95360 38066 95416
rect 38122 95360 38127 95416
rect 35718 95358 38127 95360
rect 35718 95048 35778 95358
rect 38061 95355 38127 95358
rect 230709 95418 230775 95421
rect 242526 95418 242532 95420
rect 230709 95416 242532 95418
rect 230709 95360 230714 95416
rect 230770 95360 242532 95416
rect 230709 95358 242532 95360
rect 230709 95355 230775 95358
rect 242526 95356 242532 95358
rect 242596 95356 242602 95420
rect 137789 95282 137855 95285
rect 148502 95282 148508 95284
rect 137789 95280 148508 95282
rect 137789 95224 137794 95280
rect 137850 95224 148508 95280
rect 137789 95222 148508 95224
rect 137789 95219 137855 95222
rect 148502 95220 148508 95222
rect 148572 95220 148578 95284
rect 164878 95220 164884 95284
rect 164948 95282 164954 95284
rect 178678 95282 178684 95284
rect 164948 95222 178684 95282
rect 164948 95220 164954 95222
rect 178678 95220 178684 95222
rect 178748 95220 178754 95284
rect 258718 95220 258724 95284
rect 258788 95282 258794 95284
rect 272702 95282 272708 95284
rect 258788 95222 272708 95282
rect 258788 95220 258794 95222
rect 272702 95220 272708 95222
rect 272772 95220 272778 95284
rect 231813 95010 231879 95013
rect 228734 95008 231879 95010
rect 228734 94952 231818 95008
rect 231874 94952 231879 95008
rect 408870 94980 408930 95494
rect 228734 94950 231879 94952
rect 228734 94776 228794 94950
rect 231813 94947 231879 94950
rect 229094 94812 229100 94876
rect 229164 94874 229170 94876
rect 230709 94874 230775 94877
rect 229164 94872 230775 94874
rect 229164 94816 230714 94872
rect 230770 94816 230775 94872
rect 229164 94814 230775 94816
rect 229164 94812 229170 94814
rect 230709 94811 230775 94814
rect 134710 94602 134770 94772
rect 322758 94738 322818 94776
rect 325837 94738 325903 94741
rect 322758 94736 325903 94738
rect 322758 94680 325842 94736
rect 325898 94680 325903 94736
rect 322758 94678 325903 94680
rect 325837 94675 325903 94678
rect 138157 94602 138223 94605
rect 134710 94600 138223 94602
rect 134710 94544 138162 94600
rect 138218 94544 138223 94600
rect 134710 94542 138223 94544
rect 138157 94539 138223 94542
rect 322750 94404 322756 94468
rect 322820 94466 322826 94468
rect 324549 94466 324615 94469
rect 322820 94464 324615 94466
rect 322820 94408 324554 94464
rect 324610 94408 324615 94464
rect 322820 94406 324615 94408
rect 322820 94404 322826 94406
rect 324549 94403 324615 94406
rect 74677 94330 74743 94333
rect 70862 94328 74743 94330
rect 70862 94272 74682 94328
rect 74738 94272 74743 94328
rect 70862 94270 74743 94272
rect 70862 94164 70922 94270
rect 74677 94267 74743 94270
rect 37601 92562 37667 92565
rect 35748 92560 37667 92562
rect 35748 92504 37606 92560
rect 37662 92504 37667 92560
rect 35748 92502 37667 92504
rect 37601 92499 37667 92502
rect 405969 92426 406035 92429
rect 409054 92426 409114 92532
rect 405969 92424 409114 92426
rect 405969 92368 405974 92424
rect 406030 92368 409114 92424
rect 405969 92366 409114 92368
rect 405969 92363 406035 92366
rect 81669 92290 81735 92293
rect 137605 92290 137671 92293
rect 81669 92288 84722 92290
rect 81669 92232 81674 92288
rect 81730 92232 84722 92288
rect 81669 92230 84722 92232
rect 81669 92227 81735 92230
rect 84662 92218 84722 92230
rect 134710 92288 137671 92290
rect 134710 92232 137610 92288
rect 137666 92232 137671 92288
rect 134710 92230 137671 92232
rect 84662 92158 85060 92218
rect 134710 91648 134770 92230
rect 137605 92227 137671 92230
rect 175509 92290 175575 92293
rect 231445 92290 231511 92293
rect 175509 92288 178378 92290
rect 175509 92232 175514 92288
rect 175570 92232 178378 92288
rect 175509 92230 178378 92232
rect 175509 92227 175575 92230
rect 178318 92222 178378 92230
rect 228734 92288 231511 92290
rect 228734 92232 231450 92288
rect 231506 92232 231511 92288
rect 228734 92230 231511 92232
rect 178318 92162 178900 92222
rect 228734 91648 228794 92230
rect 231445 92227 231511 92230
rect 270361 92290 270427 92293
rect 325377 92290 325443 92293
rect 270361 92288 272402 92290
rect 270361 92232 270366 92288
rect 270422 92232 272402 92288
rect 270361 92230 272402 92232
rect 270361 92227 270427 92230
rect 272342 92222 272402 92230
rect 322758 92288 325443 92290
rect 322758 92232 325382 92288
rect 325438 92232 325443 92288
rect 322758 92230 325443 92232
rect 272342 92162 272924 92222
rect 322758 91648 322818 92230
rect 325377 92227 325443 92230
rect 427681 91610 427747 91613
rect 424694 91608 427747 91610
rect 424694 91552 427686 91608
rect 427742 91552 427747 91608
rect 424694 91550 427747 91552
rect 424694 91376 424754 91550
rect 427681 91547 427747 91550
rect 17269 91338 17335 91341
rect 52597 91338 52663 91341
rect 356197 91338 356263 91341
rect 17269 91336 19924 91338
rect 17269 91280 17274 91336
rect 17330 91280 19924 91336
rect 17269 91278 19924 91280
rect 52597 91336 55068 91338
rect 52597 91280 52602 91336
rect 52658 91280 55068 91336
rect 52597 91278 55068 91280
rect 352780 91336 356263 91338
rect 352780 91280 356202 91336
rect 356258 91280 356263 91336
rect 352780 91278 356263 91280
rect 17269 91275 17335 91278
rect 52597 91275 52663 91278
rect 356197 91275 356263 91278
rect 73849 91202 73915 91205
rect 70862 91200 73915 91202
rect 70862 91144 73854 91200
rect 73910 91144 73915 91200
rect 70862 91142 73915 91144
rect 70862 90628 70922 91142
rect 73849 91139 73915 91142
rect 405969 90250 406035 90253
rect 405969 90248 408930 90250
rect 405969 90192 405974 90248
rect 406030 90192 408930 90248
rect 405969 90190 408930 90192
rect 405969 90187 406035 90190
rect 38797 90114 38863 90117
rect 35748 90112 38863 90114
rect 35748 90056 38802 90112
rect 38858 90056 38863 90112
rect 35748 90054 38863 90056
rect 38797 90051 38863 90054
rect 152182 90052 152188 90116
rect 152252 90114 152258 90116
rect 155310 90114 155316 90116
rect 152252 90054 155316 90114
rect 152252 90052 152258 90054
rect 155310 90052 155316 90054
rect 155380 90052 155386 90116
rect 246206 90052 246212 90116
rect 246276 90114 246282 90116
rect 249150 90114 249156 90116
rect 246276 90054 249156 90114
rect 246276 90052 246282 90054
rect 249150 90052 249156 90054
rect 249220 90052 249226 90116
rect 351638 90052 351644 90116
rect 351708 90114 351714 90116
rect 352793 90114 352859 90117
rect 351708 90112 352859 90114
rect 351708 90056 352798 90112
rect 352854 90056 352859 90112
rect 408870 90084 408930 90190
rect 351708 90054 352859 90056
rect 351708 90052 351714 90054
rect 352793 90051 352859 90054
rect 9896 89570 10376 89600
rect 13221 89570 13287 89573
rect 9896 89568 13287 89570
rect 9896 89512 13226 89568
rect 13282 89512 13287 89568
rect 9896 89510 13287 89512
rect 9896 89480 10376 89510
rect 13221 89507 13287 89510
rect 155361 89164 155427 89165
rect 155310 89100 155316 89164
rect 155380 89162 155427 89164
rect 155380 89160 155472 89162
rect 155422 89104 155472 89160
rect 155380 89102 155472 89104
rect 155380 89100 155427 89102
rect 245838 89100 245844 89164
rect 245908 89162 245914 89164
rect 248925 89162 248991 89165
rect 245908 89160 248991 89162
rect 245908 89104 248930 89160
rect 248986 89104 248991 89160
rect 245908 89102 248991 89104
rect 245908 89100 245914 89102
rect 155361 89099 155427 89100
rect 248925 89099 248991 89102
rect 137697 88890 137763 88893
rect 231537 88890 231603 88893
rect 134710 88888 137763 88890
rect 134710 88832 137702 88888
rect 137758 88832 137763 88888
rect 134710 88830 137763 88832
rect 134710 88520 134770 88830
rect 137697 88827 137763 88830
rect 228734 88888 231603 88890
rect 228734 88832 231542 88888
rect 231598 88832 231603 88888
rect 228734 88830 231603 88832
rect 228734 88520 228794 88830
rect 231537 88827 231603 88830
rect 249150 88828 249156 88892
rect 249220 88890 249226 88892
rect 249569 88890 249635 88893
rect 325561 88890 325627 88893
rect 249220 88888 249635 88890
rect 249220 88832 249574 88888
rect 249630 88832 249635 88888
rect 249220 88830 249635 88832
rect 249220 88828 249226 88830
rect 249569 88827 249635 88830
rect 322758 88888 325627 88890
rect 322758 88832 325566 88888
rect 325622 88832 325627 88888
rect 322758 88830 325627 88832
rect 322758 88520 322818 88830
rect 325561 88827 325627 88830
rect 249109 88484 249175 88485
rect 249109 88480 249156 88484
rect 249220 88482 249226 88484
rect 249109 88424 249114 88480
rect 249109 88420 249156 88424
rect 249220 88422 249266 88482
rect 249220 88420 249226 88422
rect 249109 88419 249175 88420
rect 72561 88348 72627 88349
rect 72510 88346 72516 88348
rect 72470 88286 72516 88346
rect 72580 88344 72627 88348
rect 72622 88288 72627 88344
rect 72510 88284 72516 88286
rect 72580 88284 72627 88288
rect 72561 88283 72627 88284
rect 252145 88076 252211 88077
rect 252094 88074 252100 88076
rect 252054 88014 252100 88074
rect 252164 88072 252211 88076
rect 252206 88016 252211 88072
rect 252094 88012 252100 88014
rect 252164 88012 252211 88016
rect 252145 88011 252211 88012
rect 260057 87530 260123 87533
rect 260333 87530 260399 87533
rect 261662 87530 261668 87532
rect 260057 87528 261668 87530
rect 260057 87472 260062 87528
rect 260118 87472 260338 87528
rect 260394 87472 261668 87528
rect 260057 87470 261668 87472
rect 260057 87467 260123 87470
rect 260333 87467 260399 87470
rect 261662 87468 261668 87470
rect 261732 87468 261738 87532
rect 430165 87530 430231 87533
rect 434416 87530 434896 87560
rect 430165 87528 434896 87530
rect 430165 87472 430170 87528
rect 430226 87472 434896 87528
rect 430165 87470 434896 87472
rect 430165 87467 430231 87470
rect 434416 87440 434896 87470
rect 155913 87394 155979 87397
rect 163774 87394 163780 87396
rect 155913 87392 163780 87394
rect 155913 87336 155918 87392
rect 155974 87336 163780 87392
rect 155913 87334 163780 87336
rect 155913 87331 155979 87334
rect 163774 87332 163780 87334
rect 163844 87394 163850 87396
rect 167638 87394 167644 87396
rect 163844 87334 167644 87394
rect 163844 87332 163850 87334
rect 167638 87332 167644 87334
rect 167708 87332 167714 87396
rect 356790 87332 356796 87396
rect 356860 87394 356866 87396
rect 360429 87394 360495 87397
rect 415537 87394 415603 87397
rect 356860 87392 415603 87394
rect 356860 87336 360434 87392
rect 360490 87336 415542 87392
rect 415598 87336 415603 87392
rect 356860 87334 415603 87336
rect 356860 87332 356866 87334
rect 360429 87331 360495 87334
rect 415537 87331 415603 87334
rect 148502 87060 148508 87124
rect 148572 87122 148578 87124
rect 157753 87122 157819 87125
rect 148572 87120 157819 87122
rect 148572 87064 157758 87120
rect 157814 87064 157819 87120
rect 148572 87062 157819 87064
rect 148572 87060 148578 87062
rect 157753 87059 157819 87062
rect 159041 87122 159107 87125
rect 168742 87122 168748 87124
rect 159041 87120 168748 87122
rect 159041 87064 159046 87120
rect 159102 87064 168748 87120
rect 159041 87062 168748 87064
rect 159041 87059 159107 87062
rect 168742 87060 168748 87062
rect 168812 87060 168818 87124
rect 158397 86986 158463 86989
rect 169294 86986 169300 86988
rect 158397 86984 169300 86986
rect 158397 86928 158402 86984
rect 158458 86928 169300 86984
rect 158397 86926 169300 86928
rect 158397 86923 158463 86926
rect 169294 86924 169300 86926
rect 169364 86924 169370 86988
rect 253065 86986 253131 86989
rect 262766 86986 262772 86988
rect 253065 86984 262772 86986
rect 253065 86928 253070 86984
rect 253126 86928 262772 86984
rect 253065 86926 262772 86928
rect 253065 86923 253131 86926
rect 262766 86924 262772 86926
rect 262836 86924 262842 86988
rect 156557 86850 156623 86853
rect 168006 86850 168012 86852
rect 156557 86848 168012 86850
rect 156557 86792 156562 86848
rect 156618 86792 168012 86848
rect 156557 86790 168012 86792
rect 156557 86787 156623 86790
rect 168006 86788 168012 86790
rect 168076 86788 168082 86852
rect 252053 86850 252119 86853
rect 263502 86850 263508 86852
rect 252053 86848 263508 86850
rect 252053 86792 252058 86848
rect 252114 86792 263508 86848
rect 252053 86790 263508 86792
rect 252053 86787 252119 86790
rect 263502 86788 263508 86790
rect 263572 86788 263578 86852
rect 157201 86714 157267 86717
rect 169110 86714 169116 86716
rect 157201 86712 169116 86714
rect 157201 86656 157206 86712
rect 157262 86656 169116 86712
rect 157201 86654 169116 86656
rect 157201 86651 157267 86654
rect 169110 86652 169116 86654
rect 169180 86652 169186 86716
rect 250857 86714 250923 86717
rect 263134 86714 263140 86716
rect 250857 86712 263140 86714
rect 250857 86656 250862 86712
rect 250918 86656 263140 86712
rect 250857 86654 263140 86656
rect 250857 86651 250923 86654
rect 263134 86652 263140 86654
rect 263204 86652 263210 86716
rect 73573 86442 73639 86445
rect 73982 86442 73988 86444
rect 73573 86440 73988 86442
rect 73573 86384 73578 86440
rect 73634 86384 73988 86440
rect 73573 86382 73988 86384
rect 73573 86379 73639 86382
rect 73982 86380 73988 86382
rect 74052 86380 74058 86444
rect 73246 86244 73252 86308
rect 73316 86306 73322 86308
rect 73665 86306 73731 86309
rect 73316 86304 73731 86306
rect 73316 86248 73670 86304
rect 73726 86248 73731 86304
rect 73316 86246 73731 86248
rect 73316 86244 73322 86246
rect 73665 86243 73731 86246
rect 72694 86108 72700 86172
rect 72764 86170 72770 86172
rect 73481 86170 73547 86173
rect 72764 86168 73547 86170
rect 72764 86112 73486 86168
rect 73542 86112 73547 86168
rect 72764 86110 73547 86112
rect 72764 86108 72770 86110
rect 73481 86107 73547 86110
rect 73757 86170 73823 86173
rect 74350 86170 74356 86172
rect 73757 86168 74356 86170
rect 73757 86112 73762 86168
rect 73818 86112 74356 86168
rect 73757 86110 74356 86112
rect 73757 86107 73823 86110
rect 74350 86108 74356 86110
rect 74420 86108 74426 86172
rect 252145 86170 252211 86173
rect 252646 86170 252652 86172
rect 252145 86168 252652 86170
rect 252145 86112 252150 86168
rect 252206 86112 252652 86168
rect 252145 86110 252652 86112
rect 252145 86107 252211 86110
rect 252646 86108 252652 86110
rect 252716 86108 252722 86172
rect 242526 85972 242532 86036
rect 242596 85972 242602 86036
rect 242534 85901 242594 85972
rect 72694 85836 72700 85900
rect 72764 85898 72770 85900
rect 72837 85898 72903 85901
rect 72764 85896 72903 85898
rect 72764 85840 72842 85896
rect 72898 85840 72903 85896
rect 72764 85838 72903 85840
rect 242534 85896 242643 85901
rect 242534 85840 242582 85896
rect 242638 85840 242643 85896
rect 242534 85838 242643 85840
rect 72764 85836 72770 85838
rect 72837 85835 72903 85838
rect 242577 85835 242643 85838
rect 230985 85762 231051 85765
rect 228734 85760 231051 85762
rect 228734 85704 230990 85760
rect 231046 85704 231051 85760
rect 228734 85702 231051 85704
rect 138157 85490 138223 85493
rect 134710 85488 138223 85490
rect 134710 85432 138162 85488
rect 138218 85432 138223 85488
rect 134710 85430 138223 85432
rect 134710 85392 134770 85430
rect 138157 85427 138223 85430
rect 228734 85392 228794 85702
rect 230985 85699 231051 85702
rect 324549 85626 324615 85629
rect 322758 85624 324615 85626
rect 322758 85568 324554 85624
rect 324610 85568 324615 85624
rect 322758 85566 324615 85568
rect 322758 85392 322818 85566
rect 324549 85563 324615 85566
rect 182501 83724 182567 83725
rect 182501 83722 182548 83724
rect 182456 83720 182548 83722
rect 182456 83664 182506 83720
rect 182456 83662 182548 83664
rect 182501 83660 182548 83662
rect 182612 83660 182618 83724
rect 182501 83659 182567 83660
rect 52638 79036 52644 79100
rect 52708 79098 52714 79100
rect 53057 79098 53123 79101
rect 52708 79096 53123 79098
rect 52708 79040 53062 79096
rect 53118 79040 53123 79096
rect 52708 79038 53123 79040
rect 52708 79036 52714 79038
rect 53057 79035 53123 79038
rect 54069 79098 54135 79101
rect 54662 79098 54668 79100
rect 54069 79096 54668 79098
rect 54069 79040 54074 79096
rect 54130 79040 54668 79096
rect 54069 79038 54668 79040
rect 54069 79035 54135 79038
rect 54662 79036 54668 79038
rect 54732 79036 54738 79100
rect 55398 79036 55404 79100
rect 55468 79098 55474 79100
rect 56093 79098 56159 79101
rect 55468 79096 56159 79098
rect 55468 79040 56098 79096
rect 56154 79040 56159 79096
rect 55468 79038 56159 79040
rect 55468 79036 55474 79038
rect 56093 79035 56159 79038
rect 54110 78900 54116 78964
rect 54180 78962 54186 78964
rect 55081 78962 55147 78965
rect 54180 78960 55147 78962
rect 54180 78904 55086 78960
rect 55142 78904 55147 78960
rect 54180 78902 55147 78904
rect 54180 78900 54186 78902
rect 55081 78899 55147 78902
rect 9896 78826 10376 78856
rect 13497 78826 13563 78829
rect 9896 78824 13563 78826
rect 9896 78768 13502 78824
rect 13558 78768 13563 78824
rect 9896 78766 13563 78768
rect 9896 78736 10376 78766
rect 13497 78763 13563 78766
rect 350953 77874 351019 77877
rect 351638 77874 351644 77876
rect 350953 77872 351644 77874
rect 350953 77816 350958 77872
rect 351014 77816 351644 77872
rect 350953 77814 351644 77816
rect 350953 77811 351019 77814
rect 351638 77812 351644 77814
rect 351708 77812 351714 77876
rect 351822 77812 351828 77876
rect 351892 77874 351898 77876
rect 352057 77874 352123 77877
rect 351892 77872 352123 77874
rect 351892 77816 352062 77872
rect 352118 77816 352123 77872
rect 351892 77814 352123 77816
rect 351892 77812 351898 77814
rect 352057 77811 352123 77814
rect 72837 76514 72903 76517
rect 73062 76514 73068 76516
rect 72837 76512 73068 76514
rect 72837 76456 72842 76512
rect 72898 76456 73068 76512
rect 72837 76454 73068 76456
rect 72837 76451 72903 76454
rect 73062 76452 73068 76454
rect 73132 76452 73138 76516
rect 242577 76514 242643 76517
rect 242710 76514 242716 76516
rect 242577 76512 242716 76514
rect 242577 76456 242582 76512
rect 242638 76456 242716 76512
rect 242577 76454 242716 76456
rect 242577 76451 242643 76454
rect 242710 76452 242716 76454
rect 242780 76452 242786 76516
rect 73062 76316 73068 76380
rect 73132 76316 73138 76380
rect 73070 76108 73130 76316
rect 73062 76044 73068 76108
rect 73132 76044 73138 76108
rect 78909 75834 78975 75837
rect 76198 75832 78975 75834
rect 76198 75776 78914 75832
rect 78970 75776 78975 75832
rect 76198 75774 78975 75776
rect 73246 75364 73252 75428
rect 73316 75426 73322 75428
rect 73798 75426 73804 75428
rect 73316 75366 73804 75426
rect 73316 75364 73322 75366
rect 73798 75364 73804 75366
rect 73868 75364 73874 75428
rect 76198 75260 76258 75774
rect 78909 75771 78975 75774
rect 155361 75564 155427 75565
rect 249201 75564 249267 75565
rect 155310 75562 155316 75564
rect 155270 75502 155316 75562
rect 155380 75560 155427 75564
rect 249150 75562 249156 75564
rect 155422 75504 155427 75560
rect 155310 75500 155316 75502
rect 155380 75500 155427 75504
rect 249110 75502 249156 75562
rect 249220 75560 249267 75564
rect 249262 75504 249267 75560
rect 249150 75500 249156 75502
rect 249220 75500 249267 75504
rect 155361 75499 155427 75500
rect 249201 75499 249267 75500
rect 252646 75364 252652 75428
rect 252716 75426 252722 75428
rect 261846 75426 261852 75428
rect 252716 75366 261852 75426
rect 252716 75364 252722 75366
rect 261846 75364 261852 75366
rect 261916 75364 261922 75428
rect 429429 75426 429495 75429
rect 434416 75426 434896 75456
rect 429429 75424 434896 75426
rect 429429 75368 429434 75424
rect 429490 75368 434896 75424
rect 429429 75366 434896 75368
rect 429429 75363 429495 75366
rect 434416 75336 434896 75366
rect 139629 75290 139695 75293
rect 173853 75290 173919 75293
rect 139629 75288 143020 75290
rect 139629 75232 139634 75288
rect 139690 75232 143020 75288
rect 139629 75230 143020 75232
rect 170804 75288 173919 75290
rect 170804 75232 173858 75288
rect 173914 75232 173919 75288
rect 170804 75230 173919 75232
rect 139629 75227 139695 75230
rect 173853 75227 173919 75230
rect 233469 75290 233535 75293
rect 266589 75290 266655 75293
rect 233469 75288 237044 75290
rect 233469 75232 233474 75288
rect 233530 75232 237044 75288
rect 233469 75230 237044 75232
rect 264828 75288 266655 75290
rect 264828 75232 266594 75288
rect 266650 75232 266655 75288
rect 264828 75230 266655 75232
rect 233469 75227 233535 75230
rect 266589 75227 266655 75230
rect 328413 75290 328479 75293
rect 328413 75288 331068 75290
rect 328413 75232 328418 75288
rect 328474 75232 331068 75288
rect 328413 75230 331068 75232
rect 328413 75227 328479 75230
rect 172933 74202 172999 74205
rect 267417 74202 267483 74205
rect 170804 74200 172999 74202
rect 76382 73930 76442 74172
rect 170804 74144 172938 74200
rect 172994 74144 172999 74200
rect 170804 74142 172999 74144
rect 264828 74200 267483 74202
rect 264828 74144 267422 74200
rect 267478 74144 267483 74200
rect 264828 74142 267483 74144
rect 172933 74139 172999 74142
rect 267417 74139 267483 74142
rect 78909 73930 78975 73933
rect 76382 73928 78975 73930
rect 76382 73872 78914 73928
rect 78970 73872 78975 73928
rect 76382 73870 78975 73872
rect 78909 73867 78975 73870
rect 139813 73794 139879 73797
rect 142990 73794 143050 74104
rect 233929 73930 233995 73933
rect 237014 73930 237074 74104
rect 233929 73928 237074 73930
rect 233929 73872 233934 73928
rect 233990 73872 237074 73928
rect 233929 73870 237074 73872
rect 327033 73930 327099 73933
rect 331038 73930 331098 74104
rect 327033 73928 331098 73930
rect 327033 73872 327038 73928
rect 327094 73872 331098 73928
rect 327033 73870 331098 73872
rect 233929 73867 233995 73870
rect 327033 73867 327099 73870
rect 139813 73792 143050 73794
rect 139813 73736 139818 73792
rect 139874 73736 143050 73792
rect 139813 73734 143050 73736
rect 139813 73731 139879 73734
rect 173485 73250 173551 73253
rect 266589 73250 266655 73253
rect 170804 73248 173551 73250
rect 76382 72842 76442 73220
rect 170804 73192 173490 73248
rect 173546 73192 173551 73248
rect 170804 73190 173551 73192
rect 264828 73248 266655 73250
rect 264828 73192 266594 73248
rect 266650 73192 266655 73248
rect 264828 73190 266655 73192
rect 173485 73187 173551 73190
rect 266589 73187 266655 73190
rect 78909 72842 78975 72845
rect 76382 72840 78975 72842
rect 76382 72784 78914 72840
rect 78970 72784 78975 72840
rect 76382 72782 78975 72784
rect 78909 72779 78975 72782
rect 139629 72570 139695 72573
rect 142990 72570 143050 73152
rect 139629 72568 143050 72570
rect 139629 72512 139634 72568
rect 139690 72512 143050 72568
rect 139629 72510 143050 72512
rect 233469 72570 233535 72573
rect 237014 72570 237074 73152
rect 233469 72568 237074 72570
rect 233469 72512 233474 72568
rect 233530 72512 237074 72568
rect 233469 72510 237074 72512
rect 327861 72570 327927 72573
rect 331038 72570 331098 73152
rect 327861 72568 331098 72570
rect 327861 72512 327866 72568
rect 327922 72512 331098 72568
rect 327861 72510 331098 72512
rect 139629 72507 139695 72510
rect 233469 72507 233535 72510
rect 327861 72507 327927 72510
rect 173485 72162 173551 72165
rect 266681 72162 266747 72165
rect 170804 72160 173551 72162
rect 76382 71618 76442 72132
rect 170804 72104 173490 72160
rect 173546 72104 173551 72160
rect 170804 72102 173551 72104
rect 264828 72160 266747 72162
rect 264828 72104 266686 72160
rect 266742 72104 266747 72160
rect 264828 72102 266747 72104
rect 173485 72099 173551 72102
rect 266681 72099 266747 72102
rect 78909 71618 78975 71621
rect 76382 71616 78975 71618
rect 76382 71560 78914 71616
rect 78970 71560 78975 71616
rect 76382 71558 78975 71560
rect 78909 71555 78975 71558
rect 139721 71482 139787 71485
rect 142990 71482 143050 72064
rect 139721 71480 143050 71482
rect 139721 71424 139726 71480
rect 139782 71424 143050 71480
rect 139721 71422 143050 71424
rect 233469 71482 233535 71485
rect 237014 71482 237074 72064
rect 233469 71480 237074 71482
rect 233469 71424 233474 71480
rect 233530 71424 237074 71480
rect 233469 71422 237074 71424
rect 327125 71482 327191 71485
rect 331038 71482 331098 72064
rect 327125 71480 331098 71482
rect 327125 71424 327130 71480
rect 327186 71424 331098 71480
rect 327125 71422 331098 71424
rect 139721 71419 139787 71422
rect 233469 71419 233535 71422
rect 327125 71419 327191 71422
rect 80197 71210 80263 71213
rect 76198 71208 80263 71210
rect 76198 71152 80202 71208
rect 80258 71152 80263 71208
rect 76198 71150 80263 71152
rect 76198 71044 76258 71150
rect 80197 71147 80263 71150
rect 139997 71074 140063 71077
rect 173301 71074 173367 71077
rect 139997 71072 143020 71074
rect 139997 71016 140002 71072
rect 140058 71016 143020 71072
rect 139997 71014 143020 71016
rect 170804 71072 173367 71074
rect 170804 71016 173306 71072
rect 173362 71016 173367 71072
rect 170804 71014 173367 71016
rect 139997 71011 140063 71014
rect 173301 71011 173367 71014
rect 233745 71074 233811 71077
rect 266589 71074 266655 71077
rect 233745 71072 237044 71074
rect 233745 71016 233750 71072
rect 233806 71016 237044 71072
rect 233745 71014 237044 71016
rect 264828 71072 266655 71074
rect 264828 71016 266594 71072
rect 266650 71016 266655 71072
rect 264828 71014 266655 71016
rect 233745 71011 233811 71014
rect 266589 71011 266655 71014
rect 326849 71074 326915 71077
rect 326849 71072 331068 71074
rect 326849 71016 326854 71072
rect 326910 71016 331068 71072
rect 326849 71014 331068 71016
rect 326849 71011 326915 71014
rect 173301 70122 173367 70125
rect 266589 70122 266655 70125
rect 170804 70120 173367 70122
rect 76382 69850 76442 70092
rect 170804 70064 173306 70120
rect 173362 70064 173367 70120
rect 170804 70062 173367 70064
rect 264828 70120 266655 70122
rect 264828 70064 266594 70120
rect 266650 70064 266655 70120
rect 264828 70062 266655 70064
rect 173301 70059 173367 70062
rect 266589 70059 266655 70062
rect 78909 69850 78975 69853
rect 76382 69848 78975 69850
rect 76382 69792 78914 69848
rect 78970 69792 78975 69848
rect 76382 69790 78975 69792
rect 78909 69787 78975 69790
rect 139905 69578 139971 69581
rect 142990 69578 143050 70024
rect 233561 69714 233627 69717
rect 237014 69714 237074 70024
rect 233561 69712 237074 69714
rect 233561 69656 233566 69712
rect 233622 69656 237074 69712
rect 233561 69654 237074 69656
rect 233561 69651 233627 69654
rect 139905 69576 143050 69578
rect 139905 69520 139910 69576
rect 139966 69520 143050 69576
rect 139905 69518 143050 69520
rect 326941 69578 327007 69581
rect 331038 69578 331098 70024
rect 326941 69576 331098 69578
rect 326941 69520 326946 69576
rect 327002 69520 331098 69576
rect 326941 69518 331098 69520
rect 139905 69515 139971 69518
rect 326941 69515 327007 69518
rect 87373 69442 87439 69445
rect 131349 69442 131415 69445
rect 87373 69440 90028 69442
rect 87373 69384 87378 69440
rect 87434 69384 90028 69440
rect 87373 69382 90028 69384
rect 129772 69440 131415 69442
rect 129772 69384 131354 69440
rect 131410 69384 131415 69440
rect 129772 69382 131415 69384
rect 87373 69379 87439 69382
rect 131349 69379 131415 69382
rect 182317 69442 182383 69445
rect 226293 69442 226359 69445
rect 182317 69440 184052 69442
rect 182317 69384 182322 69440
rect 182378 69384 184052 69440
rect 182317 69382 184052 69384
rect 223796 69440 226359 69442
rect 223796 69384 226298 69440
rect 226354 69384 226359 69440
rect 223796 69382 226359 69384
rect 182317 69379 182383 69382
rect 226293 69379 226359 69382
rect 274869 69442 274935 69445
rect 321605 69442 321671 69445
rect 274869 69440 278076 69442
rect 274869 69384 274874 69440
rect 274930 69384 278076 69440
rect 274869 69382 278076 69384
rect 317820 69440 321671 69442
rect 317820 69384 321610 69440
rect 321666 69384 321671 69440
rect 317820 69382 321671 69384
rect 274869 69379 274935 69382
rect 321605 69379 321671 69382
rect 173117 69034 173183 69037
rect 266589 69034 266655 69037
rect 170804 69032 173183 69034
rect 76382 68626 76442 69004
rect 170804 68976 173122 69032
rect 173178 68976 173183 69032
rect 170804 68974 173183 68976
rect 264828 69032 266655 69034
rect 264828 68976 266594 69032
rect 266650 68976 266655 69032
rect 264828 68974 266655 68976
rect 173117 68971 173183 68974
rect 266589 68971 266655 68974
rect 78909 68626 78975 68629
rect 76382 68624 78975 68626
rect 76382 68568 78914 68624
rect 78970 68568 78975 68624
rect 76382 68566 78975 68568
rect 78909 68563 78975 68566
rect 87189 68490 87255 68493
rect 131441 68490 131507 68493
rect 87189 68488 90028 68490
rect 87189 68432 87194 68488
rect 87250 68432 90028 68488
rect 87189 68430 90028 68432
rect 129772 68488 131507 68490
rect 129772 68432 131446 68488
rect 131502 68432 131507 68488
rect 129772 68430 131507 68432
rect 87189 68427 87255 68430
rect 131441 68427 131507 68430
rect 139629 68354 139695 68357
rect 142990 68354 143050 68936
rect 181673 68490 181739 68493
rect 226385 68490 226451 68493
rect 181673 68488 184052 68490
rect 181673 68432 181678 68488
rect 181734 68432 184052 68488
rect 181673 68430 184052 68432
rect 223796 68488 226451 68490
rect 223796 68432 226390 68488
rect 226446 68432 226451 68488
rect 223796 68430 226451 68432
rect 181673 68427 181739 68430
rect 226385 68427 226451 68430
rect 139629 68352 143050 68354
rect 139629 68296 139634 68352
rect 139690 68296 143050 68352
rect 139629 68294 143050 68296
rect 233653 68354 233719 68357
rect 237014 68354 237074 68936
rect 274961 68490 275027 68493
rect 321605 68490 321671 68493
rect 274961 68488 278076 68490
rect 274961 68432 274966 68488
rect 275022 68432 278076 68488
rect 274961 68430 278076 68432
rect 317820 68488 321671 68490
rect 317820 68432 321610 68488
rect 321666 68432 321671 68488
rect 317820 68430 321671 68432
rect 274961 68427 275027 68430
rect 321605 68427 321671 68430
rect 233653 68352 237074 68354
rect 233653 68296 233658 68352
rect 233714 68296 237074 68352
rect 233653 68294 237074 68296
rect 327033 68354 327099 68357
rect 331038 68354 331098 68936
rect 327033 68352 331098 68354
rect 327033 68296 327038 68352
rect 327094 68296 331098 68352
rect 327033 68294 331098 68296
rect 139629 68291 139695 68294
rect 233653 68291 233719 68294
rect 327033 68291 327099 68294
rect 9896 68082 10376 68112
rect 13405 68082 13471 68085
rect 9896 68080 13471 68082
rect 9896 68024 13410 68080
rect 13466 68024 13471 68080
rect 9896 68022 13471 68024
rect 9896 67992 10376 68022
rect 13405 68019 13471 68022
rect 173669 67946 173735 67949
rect 266681 67946 266747 67949
rect 170804 67944 173735 67946
rect 76382 67538 76442 67916
rect 170804 67888 173674 67944
rect 173730 67888 173735 67944
rect 170804 67886 173735 67888
rect 264828 67944 266747 67946
rect 264828 67888 266686 67944
rect 266742 67888 266747 67944
rect 264828 67886 266747 67888
rect 173669 67883 173735 67886
rect 266681 67883 266747 67886
rect 87189 67674 87255 67677
rect 132361 67674 132427 67677
rect 87189 67672 90028 67674
rect 87189 67616 87194 67672
rect 87250 67616 90028 67672
rect 87189 67614 90028 67616
rect 129772 67672 132427 67674
rect 129772 67616 132366 67672
rect 132422 67616 132427 67672
rect 129772 67614 132427 67616
rect 87189 67611 87255 67614
rect 132361 67611 132427 67614
rect 78909 67538 78975 67541
rect 76382 67536 78975 67538
rect 76382 67480 78914 67536
rect 78970 67480 78975 67536
rect 76382 67478 78975 67480
rect 78909 67475 78975 67478
rect 139721 67402 139787 67405
rect 142990 67402 143050 67848
rect 181397 67674 181463 67677
rect 226293 67674 226359 67677
rect 181397 67672 184052 67674
rect 181397 67616 181402 67672
rect 181458 67616 184052 67672
rect 181397 67614 184052 67616
rect 223796 67672 226359 67674
rect 223796 67616 226298 67672
rect 226354 67616 226359 67672
rect 223796 67614 226359 67616
rect 181397 67611 181463 67614
rect 226293 67611 226359 67614
rect 139721 67400 143050 67402
rect 139721 67344 139726 67400
rect 139782 67344 143050 67400
rect 139721 67342 143050 67344
rect 139721 67339 139787 67342
rect 233561 67266 233627 67269
rect 237014 67266 237074 67848
rect 274777 67674 274843 67677
rect 320501 67674 320567 67677
rect 274777 67672 278076 67674
rect 274777 67616 274782 67672
rect 274838 67616 278076 67672
rect 274777 67614 278076 67616
rect 317820 67672 320567 67674
rect 317820 67616 320506 67672
rect 320562 67616 320567 67672
rect 317820 67614 320567 67616
rect 274777 67611 274843 67614
rect 320501 67611 320567 67614
rect 233561 67264 237074 67266
rect 233561 67208 233566 67264
rect 233622 67208 237074 67264
rect 233561 67206 237074 67208
rect 327677 67266 327743 67269
rect 331038 67266 331098 67848
rect 327677 67264 331098 67266
rect 327677 67208 327682 67264
rect 327738 67208 331098 67264
rect 327677 67206 331098 67208
rect 233561 67203 233627 67206
rect 327677 67203 327743 67206
rect 139629 67130 139695 67133
rect 139629 67128 142314 67130
rect 139629 67072 139634 67128
rect 139690 67072 142314 67128
rect 139629 67070 142314 67072
rect 139629 67067 139695 67070
rect 76382 66858 76442 66964
rect 142254 66926 142314 67070
rect 174037 66994 174103 66997
rect 170804 66992 174103 66994
rect 170804 66936 174042 66992
rect 174098 66936 174103 66992
rect 170804 66934 174103 66936
rect 174037 66931 174103 66934
rect 233469 66994 233535 66997
rect 266589 66994 266655 66997
rect 233469 66992 237044 66994
rect 233469 66936 233474 66992
rect 233530 66936 237044 66992
rect 233469 66934 237044 66936
rect 264828 66992 266655 66994
rect 264828 66936 266594 66992
rect 266650 66936 266655 66992
rect 264828 66934 266655 66936
rect 233469 66931 233535 66934
rect 266589 66931 266655 66934
rect 328413 66994 328479 66997
rect 328413 66992 331068 66994
rect 328413 66936 328418 66992
rect 328474 66936 331068 66992
rect 328413 66934 331068 66936
rect 328413 66931 328479 66934
rect 142254 66866 143020 66926
rect 78909 66858 78975 66861
rect 76382 66856 78975 66858
rect 76382 66800 78914 66856
rect 78970 66800 78975 66856
rect 76382 66798 78975 66800
rect 78909 66795 78975 66798
rect 87189 66722 87255 66725
rect 131349 66722 131415 66725
rect 226293 66722 226359 66725
rect 87189 66720 90028 66722
rect 87189 66664 87194 66720
rect 87250 66664 90028 66720
rect 87189 66662 90028 66664
rect 129772 66720 131415 66722
rect 129772 66664 131354 66720
rect 131410 66664 131415 66720
rect 129772 66662 131415 66664
rect 223796 66720 226359 66722
rect 223796 66664 226298 66720
rect 226354 66664 226359 66720
rect 223796 66662 226359 66664
rect 87189 66659 87255 66662
rect 131349 66659 131415 66662
rect 226293 66659 226359 66662
rect 274685 66722 274751 66725
rect 321421 66722 321487 66725
rect 274685 66720 278076 66722
rect 274685 66664 274690 66720
rect 274746 66664 278076 66720
rect 274685 66662 278076 66664
rect 317820 66720 321487 66722
rect 317820 66664 321426 66720
rect 321482 66664 321487 66720
rect 317820 66662 321487 66664
rect 274685 66659 274751 66662
rect 321421 66659 321487 66662
rect 181029 66178 181095 66181
rect 184022 66178 184082 66624
rect 181029 66176 184082 66178
rect 181029 66120 181034 66176
rect 181090 66120 184082 66176
rect 181029 66118 184082 66120
rect 181029 66115 181095 66118
rect 87281 65906 87347 65909
rect 132361 65906 132427 65909
rect 174037 65906 174103 65909
rect 87281 65904 90028 65906
rect 76382 65634 76442 65876
rect 87281 65848 87286 65904
rect 87342 65848 90028 65904
rect 87281 65846 90028 65848
rect 129772 65904 132427 65906
rect 129772 65848 132366 65904
rect 132422 65848 132427 65904
rect 129772 65846 132427 65848
rect 170804 65904 174103 65906
rect 170804 65848 174042 65904
rect 174098 65848 174103 65904
rect 170804 65846 174103 65848
rect 87281 65843 87347 65846
rect 132361 65843 132427 65846
rect 174037 65843 174103 65846
rect 181765 65906 181831 65909
rect 226293 65906 226359 65909
rect 266589 65906 266655 65909
rect 181765 65904 184052 65906
rect 181765 65848 181770 65904
rect 181826 65848 184052 65904
rect 181765 65846 184052 65848
rect 223796 65904 226359 65906
rect 223796 65848 226298 65904
rect 226354 65848 226359 65904
rect 223796 65846 226359 65848
rect 264828 65904 266655 65906
rect 264828 65848 266594 65904
rect 266650 65848 266655 65904
rect 264828 65846 266655 65848
rect 181765 65843 181831 65846
rect 226293 65843 226359 65846
rect 266589 65843 266655 65846
rect 274869 65906 274935 65909
rect 321605 65906 321671 65909
rect 274869 65904 278076 65906
rect 274869 65848 274874 65904
rect 274930 65848 278076 65904
rect 274869 65846 278076 65848
rect 317820 65904 321671 65906
rect 317820 65848 321610 65904
rect 321666 65848 321671 65904
rect 317820 65846 321671 65848
rect 274869 65843 274935 65846
rect 321605 65843 321671 65846
rect 328413 65906 328479 65909
rect 328413 65904 331068 65906
rect 328413 65848 328418 65904
rect 328474 65848 331068 65904
rect 328413 65846 331068 65848
rect 328413 65843 328479 65846
rect 78909 65634 78975 65637
rect 76382 65632 78975 65634
rect 76382 65576 78914 65632
rect 78970 65576 78975 65632
rect 76382 65574 78975 65576
rect 78909 65571 78975 65574
rect 139905 65498 139971 65501
rect 142990 65498 143050 65808
rect 139905 65496 143050 65498
rect 139905 65440 139910 65496
rect 139966 65440 143050 65496
rect 139905 65438 143050 65440
rect 180845 65498 180911 65501
rect 181029 65498 181095 65501
rect 180845 65496 181095 65498
rect 180845 65440 180850 65496
rect 180906 65440 181034 65496
rect 181090 65440 181095 65496
rect 180845 65438 181095 65440
rect 139905 65435 139971 65438
rect 180845 65435 180911 65438
rect 181029 65435 181095 65438
rect 233469 65498 233535 65501
rect 237014 65498 237074 65808
rect 233469 65496 237074 65498
rect 233469 65440 233474 65496
rect 233530 65440 237074 65496
rect 233469 65438 237074 65440
rect 233469 65435 233535 65438
rect 87281 64954 87347 64957
rect 131349 64954 131415 64957
rect 173117 64954 173183 64957
rect 87281 64952 90028 64954
rect 76382 64682 76442 64924
rect 87281 64896 87286 64952
rect 87342 64896 90028 64952
rect 87281 64894 90028 64896
rect 129772 64952 131415 64954
rect 129772 64896 131354 64952
rect 131410 64896 131415 64952
rect 129772 64894 131415 64896
rect 170804 64952 173183 64954
rect 170804 64896 173122 64952
rect 173178 64896 173183 64952
rect 170804 64894 173183 64896
rect 87281 64891 87347 64894
rect 131349 64891 131415 64894
rect 173117 64891 173183 64894
rect 182317 64954 182383 64957
rect 226201 64954 226267 64957
rect 266589 64954 266655 64957
rect 182317 64952 184052 64954
rect 182317 64896 182322 64952
rect 182378 64896 184052 64952
rect 182317 64894 184052 64896
rect 223796 64952 226267 64954
rect 223796 64896 226206 64952
rect 226262 64896 226267 64952
rect 223796 64894 226267 64896
rect 264828 64952 266655 64954
rect 264828 64896 266594 64952
rect 266650 64896 266655 64952
rect 264828 64894 266655 64896
rect 182317 64891 182383 64894
rect 226201 64891 226267 64894
rect 266589 64891 266655 64894
rect 275053 64954 275119 64957
rect 321605 64954 321671 64957
rect 275053 64952 278076 64954
rect 275053 64896 275058 64952
rect 275114 64896 278076 64952
rect 275053 64894 278076 64896
rect 317820 64952 321671 64954
rect 317820 64896 321610 64952
rect 321666 64896 321671 64952
rect 317820 64894 321671 64896
rect 275053 64891 275119 64894
rect 321605 64891 321671 64894
rect 78909 64682 78975 64685
rect 76382 64680 78975 64682
rect 76382 64624 78914 64680
rect 78970 64624 78975 64680
rect 76382 64622 78975 64624
rect 78909 64619 78975 64622
rect 139629 64274 139695 64277
rect 142990 64274 143050 64856
rect 234573 64546 234639 64549
rect 237014 64546 237074 64856
rect 234573 64544 237074 64546
rect 234573 64488 234578 64544
rect 234634 64488 237074 64544
rect 234573 64486 237074 64488
rect 327309 64546 327375 64549
rect 331038 64546 331098 64856
rect 327309 64544 331098 64546
rect 327309 64488 327314 64544
rect 327370 64488 331098 64544
rect 327309 64486 331098 64488
rect 234573 64483 234639 64486
rect 327309 64483 327375 64486
rect 139629 64272 143050 64274
rect 139629 64216 139634 64272
rect 139690 64216 143050 64272
rect 139629 64214 143050 64216
rect 139629 64211 139695 64214
rect 87189 64138 87255 64141
rect 131441 64138 131507 64141
rect 87189 64136 90028 64138
rect 87189 64080 87194 64136
rect 87250 64080 90028 64136
rect 87189 64078 90028 64080
rect 129772 64136 131507 64138
rect 129772 64080 131446 64136
rect 131502 64080 131507 64136
rect 129772 64078 131507 64080
rect 87189 64075 87255 64078
rect 131441 64075 131507 64078
rect 181581 64138 181647 64141
rect 225925 64138 225991 64141
rect 181581 64136 184052 64138
rect 181581 64080 181586 64136
rect 181642 64080 184052 64136
rect 181581 64078 184052 64080
rect 223796 64136 225991 64138
rect 223796 64080 225930 64136
rect 225986 64080 225991 64136
rect 223796 64078 225991 64080
rect 181581 64075 181647 64078
rect 225925 64075 225991 64078
rect 274869 64138 274935 64141
rect 321421 64138 321487 64141
rect 274869 64136 278076 64138
rect 274869 64080 274874 64136
rect 274930 64080 278076 64136
rect 274869 64078 278076 64080
rect 317820 64136 321487 64138
rect 317820 64080 321426 64136
rect 321482 64080 321487 64136
rect 317820 64078 321487 64080
rect 274869 64075 274935 64078
rect 321421 64075 321487 64078
rect 173485 63866 173551 63869
rect 266681 63866 266747 63869
rect 170804 63864 173551 63866
rect 76382 63458 76442 63836
rect 170804 63808 173490 63864
rect 173546 63808 173551 63864
rect 170804 63806 173551 63808
rect 264828 63864 266747 63866
rect 264828 63808 266686 63864
rect 266742 63808 266747 63864
rect 264828 63806 266747 63808
rect 173485 63803 173551 63806
rect 266681 63803 266747 63806
rect 78909 63458 78975 63461
rect 76382 63456 78975 63458
rect 76382 63400 78914 63456
rect 78970 63400 78975 63456
rect 76382 63398 78975 63400
rect 78909 63395 78975 63398
rect 87189 63186 87255 63189
rect 132361 63186 132427 63189
rect 87189 63184 90028 63186
rect 87189 63128 87194 63184
rect 87250 63128 90028 63184
rect 87189 63126 90028 63128
rect 129772 63184 132427 63186
rect 129772 63128 132366 63184
rect 132422 63128 132427 63184
rect 129772 63126 132427 63128
rect 87189 63123 87255 63126
rect 132361 63123 132427 63126
rect 139721 63186 139787 63189
rect 142990 63186 143050 63768
rect 139721 63184 143050 63186
rect 139721 63128 139726 63184
rect 139782 63128 143050 63184
rect 139721 63126 143050 63128
rect 182317 63186 182383 63189
rect 225741 63186 225807 63189
rect 182317 63184 184052 63186
rect 182317 63128 182322 63184
rect 182378 63128 184052 63184
rect 182317 63126 184052 63128
rect 223796 63184 225807 63186
rect 223796 63128 225746 63184
rect 225802 63128 225807 63184
rect 223796 63126 225807 63128
rect 139721 63123 139787 63126
rect 182317 63123 182383 63126
rect 225741 63123 225807 63126
rect 233469 63186 233535 63189
rect 237014 63186 237074 63768
rect 233469 63184 237074 63186
rect 233469 63128 233474 63184
rect 233530 63128 237074 63184
rect 233469 63126 237074 63128
rect 274869 63186 274935 63189
rect 321053 63186 321119 63189
rect 274869 63184 278076 63186
rect 274869 63128 274874 63184
rect 274930 63128 278076 63184
rect 274869 63126 278076 63128
rect 317820 63184 321119 63186
rect 317820 63128 321058 63184
rect 321114 63128 321119 63184
rect 317820 63126 321119 63128
rect 233469 63123 233535 63126
rect 274869 63123 274935 63126
rect 321053 63123 321119 63126
rect 328045 63186 328111 63189
rect 331038 63186 331098 63768
rect 430073 63322 430139 63325
rect 434416 63322 434896 63352
rect 430073 63320 434896 63322
rect 430073 63264 430078 63320
rect 430134 63264 434896 63320
rect 430073 63262 434896 63264
rect 430073 63259 430139 63262
rect 434416 63232 434896 63262
rect 328045 63184 331098 63186
rect 328045 63128 328050 63184
rect 328106 63128 331098 63184
rect 328045 63126 331098 63128
rect 328045 63123 328111 63126
rect 78909 62914 78975 62917
rect 76198 62912 78975 62914
rect 76198 62856 78914 62912
rect 78970 62856 78975 62912
rect 76198 62854 78975 62856
rect 76198 62748 76258 62854
rect 78909 62851 78975 62854
rect 139813 62778 139879 62781
rect 174037 62778 174103 62781
rect 139813 62776 143020 62778
rect 139813 62720 139818 62776
rect 139874 62720 143020 62776
rect 139813 62718 143020 62720
rect 170804 62776 174103 62778
rect 170804 62720 174042 62776
rect 174098 62720 174103 62776
rect 170804 62718 174103 62720
rect 139813 62715 139879 62718
rect 174037 62715 174103 62718
rect 233561 62778 233627 62781
rect 266589 62778 266655 62781
rect 233561 62776 237044 62778
rect 233561 62720 233566 62776
rect 233622 62720 237044 62776
rect 233561 62718 237044 62720
rect 264828 62776 266655 62778
rect 264828 62720 266594 62776
rect 266650 62720 266655 62776
rect 264828 62718 266655 62720
rect 233561 62715 233627 62718
rect 266589 62715 266655 62718
rect 328321 62778 328387 62781
rect 328321 62776 331068 62778
rect 328321 62720 328326 62776
rect 328382 62720 331068 62776
rect 328321 62718 331068 62720
rect 328321 62715 328387 62718
rect 87281 62370 87347 62373
rect 131349 62370 131415 62373
rect 87281 62368 90028 62370
rect 87281 62312 87286 62368
rect 87342 62312 90028 62368
rect 87281 62310 90028 62312
rect 129772 62368 131415 62370
rect 129772 62312 131354 62368
rect 131410 62312 131415 62368
rect 129772 62310 131415 62312
rect 87281 62307 87347 62310
rect 131349 62307 131415 62310
rect 182317 62370 182383 62373
rect 226293 62370 226359 62373
rect 182317 62368 184052 62370
rect 182317 62312 182322 62368
rect 182378 62312 184052 62368
rect 182317 62310 184052 62312
rect 223796 62368 226359 62370
rect 223796 62312 226298 62368
rect 226354 62312 226359 62368
rect 223796 62310 226359 62312
rect 182317 62307 182383 62310
rect 226293 62307 226359 62310
rect 274961 62370 275027 62373
rect 321697 62370 321763 62373
rect 274961 62368 278076 62370
rect 274961 62312 274966 62368
rect 275022 62312 278076 62368
rect 274961 62310 278076 62312
rect 317820 62368 321763 62370
rect 317820 62312 321702 62368
rect 321758 62312 321763 62368
rect 317820 62310 321763 62312
rect 274961 62307 275027 62310
rect 321697 62307 321763 62310
rect 173117 61826 173183 61829
rect 266589 61826 266655 61829
rect 170804 61824 173183 61826
rect 76382 61554 76442 61796
rect 170804 61768 173122 61824
rect 173178 61768 173183 61824
rect 170804 61766 173183 61768
rect 264828 61824 266655 61826
rect 264828 61768 266594 61824
rect 266650 61768 266655 61824
rect 264828 61766 266655 61768
rect 173117 61763 173183 61766
rect 266589 61763 266655 61766
rect 78909 61554 78975 61557
rect 76382 61552 78975 61554
rect 76382 61496 78914 61552
rect 78970 61496 78975 61552
rect 76382 61494 78975 61496
rect 78909 61491 78975 61494
rect 87189 61418 87255 61421
rect 131717 61418 131783 61421
rect 87189 61416 90028 61418
rect 87189 61360 87194 61416
rect 87250 61360 90028 61416
rect 87189 61358 90028 61360
rect 129772 61416 131783 61418
rect 129772 61360 131722 61416
rect 131778 61360 131783 61416
rect 129772 61358 131783 61360
rect 87189 61355 87255 61358
rect 131717 61355 131783 61358
rect 139629 61418 139695 61421
rect 142990 61418 143050 61728
rect 139629 61416 143050 61418
rect 139629 61360 139634 61416
rect 139690 61360 143050 61416
rect 139629 61358 143050 61360
rect 181581 61418 181647 61421
rect 225925 61418 225991 61421
rect 181581 61416 184052 61418
rect 181581 61360 181586 61416
rect 181642 61360 184052 61416
rect 181581 61358 184052 61360
rect 223796 61416 225991 61418
rect 223796 61360 225930 61416
rect 225986 61360 225991 61416
rect 223796 61358 225991 61360
rect 139629 61355 139695 61358
rect 181581 61355 181647 61358
rect 225925 61355 225991 61358
rect 233469 61418 233535 61421
rect 237014 61418 237074 61728
rect 328505 61554 328571 61557
rect 331038 61554 331098 61728
rect 328505 61552 331098 61554
rect 328505 61496 328510 61552
rect 328566 61496 331098 61552
rect 328505 61494 331098 61496
rect 328505 61491 328571 61494
rect 233469 61416 237074 61418
rect 233469 61360 233474 61416
rect 233530 61360 237074 61416
rect 233469 61358 237074 61360
rect 274869 61418 274935 61421
rect 321237 61418 321303 61421
rect 274869 61416 278076 61418
rect 274869 61360 274874 61416
rect 274930 61360 278076 61416
rect 274869 61358 278076 61360
rect 317820 61416 321303 61418
rect 317820 61360 321242 61416
rect 321298 61360 321303 61416
rect 317820 61358 321303 61360
rect 233469 61355 233535 61358
rect 274869 61355 274935 61358
rect 321237 61355 321303 61358
rect 173485 60738 173551 60741
rect 266589 60738 266655 60741
rect 170804 60736 173551 60738
rect 76382 60330 76442 60708
rect 170804 60680 173490 60736
rect 173546 60680 173551 60736
rect 170804 60678 173551 60680
rect 264828 60736 266655 60738
rect 264828 60680 266594 60736
rect 266650 60680 266655 60736
rect 264828 60678 266655 60680
rect 173485 60675 173551 60678
rect 266589 60675 266655 60678
rect 87189 60466 87255 60469
rect 131349 60466 131415 60469
rect 87189 60464 90028 60466
rect 87189 60408 87194 60464
rect 87250 60408 90028 60464
rect 87189 60406 90028 60408
rect 129772 60464 131415 60466
rect 129772 60408 131354 60464
rect 131410 60408 131415 60464
rect 129772 60406 131415 60408
rect 87189 60403 87255 60406
rect 131349 60403 131415 60406
rect 78909 60330 78975 60333
rect 76382 60328 78975 60330
rect 76382 60272 78914 60328
rect 78970 60272 78975 60328
rect 76382 60270 78975 60272
rect 78909 60267 78975 60270
rect 139721 60058 139787 60061
rect 142990 60058 143050 60640
rect 181213 60466 181279 60469
rect 226293 60466 226359 60469
rect 181213 60464 184052 60466
rect 181213 60408 181218 60464
rect 181274 60408 184052 60464
rect 181213 60406 184052 60408
rect 223796 60464 226359 60466
rect 223796 60408 226298 60464
rect 226354 60408 226359 60464
rect 223796 60406 226359 60408
rect 181213 60403 181279 60406
rect 226293 60403 226359 60406
rect 139721 60056 143050 60058
rect 139721 60000 139726 60056
rect 139782 60000 143050 60056
rect 139721 59998 143050 60000
rect 233653 60058 233719 60061
rect 237014 60058 237074 60640
rect 274869 60466 274935 60469
rect 320869 60466 320935 60469
rect 274869 60464 278076 60466
rect 274869 60408 274874 60464
rect 274930 60408 278076 60464
rect 274869 60406 278076 60408
rect 317820 60464 320935 60466
rect 317820 60408 320874 60464
rect 320930 60408 320935 60464
rect 317820 60406 320935 60408
rect 274869 60403 274935 60406
rect 320869 60403 320935 60406
rect 233653 60056 237074 60058
rect 233653 60000 233658 60056
rect 233714 60000 237074 60056
rect 233653 59998 237074 60000
rect 328413 60058 328479 60061
rect 331038 60058 331098 60640
rect 328413 60056 331098 60058
rect 328413 60000 328418 60056
rect 328474 60000 331098 60056
rect 328413 59998 331098 60000
rect 139721 59995 139787 59998
rect 233653 59995 233719 59998
rect 328413 59995 328479 59998
rect 87373 59650 87439 59653
rect 132637 59650 132703 59653
rect 174037 59650 174103 59653
rect 87373 59648 90028 59650
rect 76382 59106 76442 59620
rect 87373 59592 87378 59648
rect 87434 59592 90028 59648
rect 87373 59590 90028 59592
rect 129772 59648 132703 59650
rect 129772 59592 132642 59648
rect 132698 59592 132703 59648
rect 129772 59590 132703 59592
rect 170804 59648 174103 59650
rect 170804 59592 174042 59648
rect 174098 59592 174103 59648
rect 170804 59590 174103 59592
rect 87373 59587 87439 59590
rect 132637 59587 132703 59590
rect 174037 59587 174103 59590
rect 182317 59650 182383 59653
rect 226109 59650 226175 59653
rect 266681 59650 266747 59653
rect 182317 59648 184052 59650
rect 182317 59592 182322 59648
rect 182378 59592 184052 59648
rect 182317 59590 184052 59592
rect 223796 59648 226175 59650
rect 223796 59592 226114 59648
rect 226170 59592 226175 59648
rect 223796 59590 226175 59592
rect 264828 59648 266747 59650
rect 264828 59592 266686 59648
rect 266742 59592 266747 59648
rect 264828 59590 266747 59592
rect 182317 59587 182383 59590
rect 226109 59587 226175 59590
rect 266681 59587 266747 59590
rect 275053 59650 275119 59653
rect 321605 59650 321671 59653
rect 275053 59648 278076 59650
rect 275053 59592 275058 59648
rect 275114 59592 278076 59648
rect 275053 59590 278076 59592
rect 317820 59648 321671 59650
rect 317820 59592 321610 59648
rect 321666 59592 321671 59648
rect 317820 59590 321671 59592
rect 275053 59587 275119 59590
rect 321605 59587 321671 59590
rect 80197 59106 80263 59109
rect 76382 59104 80263 59106
rect 76382 59048 80202 59104
rect 80258 59048 80263 59104
rect 76382 59046 80263 59048
rect 80197 59043 80263 59046
rect 139721 58970 139787 58973
rect 142990 58970 143050 59552
rect 139721 58968 143050 58970
rect 139721 58912 139726 58968
rect 139782 58912 143050 58968
rect 139721 58910 143050 58912
rect 233561 58970 233627 58973
rect 237014 58970 237074 59552
rect 233561 58968 237074 58970
rect 233561 58912 233566 58968
rect 233622 58912 237074 58968
rect 233561 58910 237074 58912
rect 328505 58970 328571 58973
rect 331038 58970 331098 59552
rect 328505 58968 331098 58970
rect 328505 58912 328510 58968
rect 328566 58912 331098 58968
rect 328505 58910 331098 58912
rect 139721 58907 139787 58910
rect 233561 58907 233627 58910
rect 328505 58907 328571 58910
rect 87189 58698 87255 58701
rect 132545 58698 132611 58701
rect 87189 58696 90028 58698
rect 76382 58562 76442 58668
rect 87189 58640 87194 58696
rect 87250 58640 90028 58696
rect 87189 58638 90028 58640
rect 129772 58696 132611 58698
rect 129772 58640 132550 58696
rect 132606 58640 132611 58696
rect 129772 58638 132611 58640
rect 87189 58635 87255 58638
rect 132545 58635 132611 58638
rect 139629 58698 139695 58701
rect 174037 58698 174103 58701
rect 139629 58696 143020 58698
rect 139629 58640 139634 58696
rect 139690 58640 143020 58696
rect 139629 58638 143020 58640
rect 170804 58696 174103 58698
rect 170804 58640 174042 58696
rect 174098 58640 174103 58696
rect 170804 58638 174103 58640
rect 139629 58635 139695 58638
rect 174037 58635 174103 58638
rect 181581 58698 181647 58701
rect 226293 58698 226359 58701
rect 181581 58696 184052 58698
rect 181581 58640 181586 58696
rect 181642 58640 184052 58696
rect 181581 58638 184052 58640
rect 223796 58696 226359 58698
rect 223796 58640 226298 58696
rect 226354 58640 226359 58696
rect 223796 58638 226359 58640
rect 181581 58635 181647 58638
rect 226293 58635 226359 58638
rect 233469 58698 233535 58701
rect 266589 58698 266655 58701
rect 233469 58696 237044 58698
rect 233469 58640 233474 58696
rect 233530 58640 237044 58696
rect 233469 58638 237044 58640
rect 264828 58696 266655 58698
rect 264828 58640 266594 58696
rect 266650 58640 266655 58696
rect 264828 58638 266655 58640
rect 233469 58635 233535 58638
rect 266589 58635 266655 58638
rect 274869 58698 274935 58701
rect 321053 58698 321119 58701
rect 274869 58696 278076 58698
rect 274869 58640 274874 58696
rect 274930 58640 278076 58696
rect 274869 58638 278076 58640
rect 317820 58696 321119 58698
rect 317820 58640 321058 58696
rect 321114 58640 321119 58696
rect 317820 58638 321119 58640
rect 274869 58635 274935 58638
rect 321053 58635 321119 58638
rect 327677 58698 327743 58701
rect 327677 58696 331068 58698
rect 327677 58640 327682 58696
rect 327738 58640 331068 58696
rect 327677 58638 331068 58640
rect 327677 58635 327743 58638
rect 80197 58562 80263 58565
rect 76382 58560 80263 58562
rect 76382 58504 80202 58560
rect 80258 58504 80263 58560
rect 76382 58502 80263 58504
rect 80197 58499 80263 58502
rect 87189 57882 87255 57885
rect 132637 57882 132703 57885
rect 87189 57880 90028 57882
rect 87189 57824 87194 57880
rect 87250 57824 90028 57880
rect 87189 57822 90028 57824
rect 129772 57880 132703 57882
rect 129772 57824 132642 57880
rect 132698 57824 132703 57880
rect 129772 57822 132703 57824
rect 87189 57819 87255 57822
rect 132637 57819 132703 57822
rect 182317 57882 182383 57885
rect 226293 57882 226359 57885
rect 182317 57880 184052 57882
rect 182317 57824 182322 57880
rect 182378 57824 184052 57880
rect 182317 57822 184052 57824
rect 223796 57880 226359 57882
rect 223796 57824 226298 57880
rect 226354 57824 226359 57880
rect 223796 57822 226359 57824
rect 182317 57819 182383 57822
rect 226293 57819 226359 57822
rect 274961 57882 275027 57885
rect 320869 57882 320935 57885
rect 274961 57880 278076 57882
rect 274961 57824 274966 57880
rect 275022 57824 278076 57880
rect 274961 57822 278076 57824
rect 317820 57880 320935 57882
rect 317820 57824 320874 57880
rect 320930 57824 320935 57880
rect 317820 57822 320935 57824
rect 274961 57819 275027 57822
rect 320869 57819 320935 57822
rect 173485 57610 173551 57613
rect 266589 57610 266655 57613
rect 170804 57608 173551 57610
rect 9896 57338 10376 57368
rect 13313 57338 13379 57341
rect 9896 57336 13379 57338
rect 9896 57280 13318 57336
rect 13374 57280 13379 57336
rect 9896 57278 13379 57280
rect 76382 57338 76442 57580
rect 170804 57552 173490 57608
rect 173546 57552 173551 57608
rect 170804 57550 173551 57552
rect 264828 57608 266655 57610
rect 264828 57552 266594 57608
rect 266650 57552 266655 57608
rect 264828 57550 266655 57552
rect 173485 57547 173551 57550
rect 266589 57547 266655 57550
rect 78909 57338 78975 57341
rect 76382 57336 78975 57338
rect 76382 57280 78914 57336
rect 78970 57280 78975 57336
rect 76382 57278 78975 57280
rect 9896 57248 10376 57278
rect 13313 57275 13379 57278
rect 78909 57275 78975 57278
rect 139629 57338 139695 57341
rect 142990 57338 143050 57512
rect 139629 57336 143050 57338
rect 139629 57280 139634 57336
rect 139690 57280 143050 57336
rect 139629 57278 143050 57280
rect 139629 57275 139695 57278
rect 233469 57202 233535 57205
rect 237014 57202 237074 57512
rect 233469 57200 237074 57202
rect 233469 57144 233474 57200
rect 233530 57144 237074 57200
rect 233469 57142 237074 57144
rect 328321 57202 328387 57205
rect 331038 57202 331098 57512
rect 328321 57200 331098 57202
rect 328321 57144 328326 57200
rect 328382 57144 331098 57200
rect 328321 57142 331098 57144
rect 233469 57139 233535 57142
rect 328321 57139 328387 57142
rect 87189 56930 87255 56933
rect 132637 56930 132703 56933
rect 226293 56930 226359 56933
rect 87189 56928 90028 56930
rect 87189 56872 87194 56928
rect 87250 56872 90028 56928
rect 87189 56870 90028 56872
rect 129772 56928 132703 56930
rect 129772 56872 132642 56928
rect 132698 56872 132703 56928
rect 129772 56870 132703 56872
rect 223796 56928 226359 56930
rect 223796 56872 226298 56928
rect 226354 56872 226359 56928
rect 223796 56870 226359 56872
rect 87189 56867 87255 56870
rect 132637 56867 132703 56870
rect 226293 56867 226359 56870
rect 274869 56930 274935 56933
rect 321053 56930 321119 56933
rect 274869 56928 278076 56930
rect 274869 56872 274874 56928
rect 274930 56872 278076 56928
rect 274869 56870 278076 56872
rect 317820 56928 321119 56930
rect 317820 56872 321058 56928
rect 321114 56872 321119 56928
rect 317820 56870 321119 56872
rect 274869 56867 274935 56870
rect 321053 56867 321119 56870
rect 172749 56658 172815 56661
rect 170804 56656 172815 56658
rect 76382 56250 76442 56628
rect 170804 56600 172754 56656
rect 172810 56600 172815 56656
rect 170804 56598 172815 56600
rect 172749 56595 172815 56598
rect 78909 56250 78975 56253
rect 76382 56248 78975 56250
rect 76382 56192 78914 56248
rect 78970 56192 78975 56248
rect 76382 56190 78975 56192
rect 78909 56187 78975 56190
rect 87281 56114 87347 56117
rect 132545 56114 132611 56117
rect 87281 56112 90028 56114
rect 87281 56056 87286 56112
rect 87342 56056 90028 56112
rect 87281 56054 90028 56056
rect 129772 56112 132611 56114
rect 129772 56056 132550 56112
rect 132606 56056 132611 56112
rect 129772 56054 132611 56056
rect 87281 56051 87347 56054
rect 132545 56051 132611 56054
rect 139537 55978 139603 55981
rect 142990 55978 143050 56560
rect 182317 56522 182383 56525
rect 184022 56522 184082 56832
rect 266589 56658 266655 56661
rect 264828 56656 266655 56658
rect 264828 56600 266594 56656
rect 266650 56600 266655 56656
rect 264828 56598 266655 56600
rect 266589 56595 266655 56598
rect 182317 56520 184082 56522
rect 182317 56464 182322 56520
rect 182378 56464 184082 56520
rect 182317 56462 184082 56464
rect 182317 56459 182383 56462
rect 181765 56114 181831 56117
rect 225373 56114 225439 56117
rect 181765 56112 184052 56114
rect 181765 56056 181770 56112
rect 181826 56056 184052 56112
rect 181765 56054 184052 56056
rect 223796 56112 225439 56114
rect 223796 56056 225378 56112
rect 225434 56056 225439 56112
rect 223796 56054 225439 56056
rect 181765 56051 181831 56054
rect 225373 56051 225439 56054
rect 139537 55976 143050 55978
rect 139537 55920 139542 55976
rect 139598 55920 143050 55976
rect 139537 55918 143050 55920
rect 234389 55978 234455 55981
rect 237014 55978 237074 56560
rect 327493 56250 327559 56253
rect 331038 56250 331098 56560
rect 327493 56248 331098 56250
rect 327493 56192 327498 56248
rect 327554 56192 331098 56248
rect 327493 56190 331098 56192
rect 327493 56187 327559 56190
rect 275053 56114 275119 56117
rect 321605 56114 321671 56117
rect 275053 56112 278076 56114
rect 275053 56056 275058 56112
rect 275114 56056 278076 56112
rect 275053 56054 278076 56056
rect 317820 56112 321671 56114
rect 317820 56056 321610 56112
rect 321666 56056 321671 56112
rect 317820 56054 321671 56056
rect 275053 56051 275119 56054
rect 321605 56051 321671 56054
rect 234389 55976 237074 55978
rect 234389 55920 234394 55976
rect 234450 55920 237074 55976
rect 234389 55918 237074 55920
rect 139537 55915 139603 55918
rect 234389 55915 234455 55918
rect 79553 55706 79619 55709
rect 76198 55704 79619 55706
rect 76198 55648 79558 55704
rect 79614 55648 79619 55704
rect 76198 55646 79619 55648
rect 76198 55540 76258 55646
rect 79553 55643 79619 55646
rect 173393 55570 173459 55573
rect 267233 55570 267299 55573
rect 170804 55568 173459 55570
rect 170804 55512 173398 55568
rect 173454 55512 173459 55568
rect 170804 55510 173459 55512
rect 264828 55568 267299 55570
rect 264828 55512 267238 55568
rect 267294 55512 267299 55568
rect 264828 55510 267299 55512
rect 173393 55507 173459 55510
rect 267233 55507 267299 55510
rect 87373 55162 87439 55165
rect 132637 55162 132703 55165
rect 87373 55160 90028 55162
rect 87373 55104 87378 55160
rect 87434 55104 90028 55160
rect 87373 55102 90028 55104
rect 129772 55160 132703 55162
rect 129772 55104 132642 55160
rect 132698 55104 132703 55160
rect 129772 55102 132703 55104
rect 87373 55099 87439 55102
rect 132637 55099 132703 55102
rect 134201 55162 134267 55165
rect 142990 55162 143050 55472
rect 233469 55298 233535 55301
rect 237014 55298 237074 55472
rect 233469 55296 237074 55298
rect 233469 55240 233474 55296
rect 233530 55240 237074 55296
rect 233469 55238 237074 55240
rect 328505 55298 328571 55301
rect 331038 55298 331098 55472
rect 328505 55296 331098 55298
rect 328505 55240 328510 55296
rect 328566 55240 331098 55296
rect 328505 55238 331098 55240
rect 233469 55235 233535 55238
rect 328505 55235 328571 55238
rect 134201 55160 143050 55162
rect 134201 55104 134206 55160
rect 134262 55104 143050 55160
rect 134201 55102 143050 55104
rect 181673 55162 181739 55165
rect 225373 55162 225439 55165
rect 181673 55160 184052 55162
rect 181673 55104 181678 55160
rect 181734 55104 184052 55160
rect 181673 55102 184052 55104
rect 223796 55160 225439 55162
rect 223796 55104 225378 55160
rect 225434 55104 225439 55160
rect 223796 55102 225439 55104
rect 134201 55099 134267 55102
rect 181673 55099 181739 55102
rect 225373 55099 225439 55102
rect 274961 55162 275027 55165
rect 321605 55162 321671 55165
rect 274961 55160 278076 55162
rect 274961 55104 274966 55160
rect 275022 55104 278076 55160
rect 274961 55102 278076 55104
rect 317820 55160 321671 55162
rect 317820 55104 321610 55160
rect 321666 55104 321671 55160
rect 317820 55102 321671 55104
rect 274961 55099 275027 55102
rect 321605 55099 321671 55102
rect 78909 54618 78975 54621
rect 76198 54616 78975 54618
rect 76198 54560 78914 54616
rect 78970 54560 78975 54616
rect 76198 54558 78975 54560
rect 76198 54452 76258 54558
rect 78909 54555 78975 54558
rect 139629 54482 139695 54485
rect 174037 54482 174103 54485
rect 139629 54480 143020 54482
rect 139629 54424 139634 54480
rect 139690 54424 143020 54480
rect 139629 54422 143020 54424
rect 170804 54480 174103 54482
rect 170804 54424 174042 54480
rect 174098 54424 174103 54480
rect 170804 54422 174103 54424
rect 139629 54419 139695 54422
rect 174037 54419 174103 54422
rect 233469 54482 233535 54485
rect 266589 54482 266655 54485
rect 233469 54480 237044 54482
rect 233469 54424 233474 54480
rect 233530 54424 237044 54480
rect 233469 54422 237044 54424
rect 264828 54480 266655 54482
rect 264828 54424 266594 54480
rect 266650 54424 266655 54480
rect 264828 54422 266655 54424
rect 233469 54419 233535 54422
rect 266589 54419 266655 54422
rect 328413 54482 328479 54485
rect 328413 54480 331068 54482
rect 328413 54424 328418 54480
rect 328474 54424 331068 54480
rect 328413 54422 331068 54424
rect 328413 54419 328479 54422
rect 87189 54346 87255 54349
rect 132637 54346 132703 54349
rect 87189 54344 90028 54346
rect 87189 54288 87194 54344
rect 87250 54288 90028 54344
rect 87189 54286 90028 54288
rect 129772 54344 132703 54346
rect 129772 54288 132642 54344
rect 132698 54288 132703 54344
rect 129772 54286 132703 54288
rect 87189 54283 87255 54286
rect 132637 54283 132703 54286
rect 182317 54346 182383 54349
rect 226293 54346 226359 54349
rect 182317 54344 184052 54346
rect 182317 54288 182322 54344
rect 182378 54288 184052 54344
rect 182317 54286 184052 54288
rect 223796 54344 226359 54346
rect 223796 54288 226298 54344
rect 226354 54288 226359 54344
rect 223796 54286 226359 54288
rect 182317 54283 182383 54286
rect 226293 54283 226359 54286
rect 274869 54346 274935 54349
rect 320961 54346 321027 54349
rect 274869 54344 278076 54346
rect 274869 54288 274874 54344
rect 274930 54288 278076 54344
rect 274869 54286 278076 54288
rect 317820 54344 321027 54346
rect 317820 54288 320966 54344
rect 321022 54288 321027 54344
rect 317820 54286 321027 54288
rect 274869 54283 274935 54286
rect 320961 54283 321027 54286
rect 78909 53666 78975 53669
rect 76198 53664 78975 53666
rect 76198 53608 78914 53664
rect 78970 53608 78975 53664
rect 76198 53606 78975 53608
rect 76198 53500 76258 53606
rect 78909 53603 78975 53606
rect 139629 53530 139695 53533
rect 174037 53530 174103 53533
rect 139629 53528 143020 53530
rect 139629 53472 139634 53528
rect 139690 53472 143020 53528
rect 139629 53470 143020 53472
rect 170804 53528 174103 53530
rect 170804 53472 174042 53528
rect 174098 53472 174103 53528
rect 170804 53470 174103 53472
rect 139629 53467 139695 53470
rect 174037 53467 174103 53470
rect 233469 53530 233535 53533
rect 266589 53530 266655 53533
rect 233469 53528 237044 53530
rect 233469 53472 233474 53528
rect 233530 53472 237044 53528
rect 233469 53470 237044 53472
rect 264828 53528 266655 53530
rect 264828 53472 266594 53528
rect 266650 53472 266655 53528
rect 264828 53470 266655 53472
rect 233469 53467 233535 53470
rect 266589 53467 266655 53470
rect 328413 53530 328479 53533
rect 328413 53528 331068 53530
rect 328413 53472 328418 53528
rect 328474 53472 331068 53528
rect 328413 53470 331068 53472
rect 328413 53467 328479 53470
rect 306977 53394 307043 53397
rect 307110 53394 307116 53396
rect 306977 53392 307116 53394
rect 306977 53336 306982 53392
rect 307038 53336 307116 53392
rect 306977 53334 307116 53336
rect 306977 53331 307043 53334
rect 307110 53332 307116 53334
rect 307180 53332 307186 53396
rect 118193 53124 118259 53125
rect 212033 53124 212099 53125
rect 118142 53122 118148 53124
rect 118102 53062 118148 53122
rect 118212 53120 118259 53124
rect 211982 53122 211988 53124
rect 118254 53064 118259 53120
rect 118142 53060 118148 53062
rect 118212 53060 118259 53064
rect 211942 53062 211988 53122
rect 212052 53120 212099 53124
rect 212094 53064 212099 53120
rect 211982 53060 211988 53062
rect 212052 53060 212099 53064
rect 118193 53059 118259 53060
rect 212033 53059 212099 53060
rect 78950 52850 78956 52852
rect 76198 52790 78956 52850
rect 76198 52412 76258 52790
rect 78950 52788 78956 52790
rect 79020 52788 79026 52852
rect 173894 52442 173900 52444
rect 170804 52382 173900 52442
rect 173894 52380 173900 52382
rect 173964 52380 173970 52444
rect 266630 52442 266636 52444
rect 264828 52382 266636 52442
rect 266630 52380 266636 52382
rect 266700 52380 266706 52444
rect 134150 51700 134156 51764
rect 134220 51762 134226 51764
rect 142990 51762 143050 52344
rect 134220 51702 143050 51762
rect 134220 51700 134226 51702
rect 227990 51700 227996 51764
rect 228060 51762 228066 51764
rect 237014 51762 237074 52344
rect 228060 51702 237074 51762
rect 228060 51700 228066 51702
rect 321830 51700 321836 51764
rect 321900 51762 321906 51764
rect 331038 51762 331098 52344
rect 321900 51702 331098 51762
rect 321900 51700 321906 51702
rect 102369 51354 102435 51357
rect 102502 51354 102508 51356
rect 102369 51352 102508 51354
rect 76382 50810 76442 51324
rect 102369 51296 102374 51352
rect 102430 51296 102508 51352
rect 102369 51294 102508 51296
rect 102369 51291 102435 51294
rect 102502 51292 102508 51294
rect 102572 51292 102578 51356
rect 173945 51354 174011 51357
rect 266681 51354 266747 51357
rect 170804 51352 174011 51354
rect 170804 51296 173950 51352
rect 174006 51296 174011 51352
rect 170804 51294 174011 51296
rect 264828 51352 266747 51354
rect 264828 51296 266686 51352
rect 266742 51296 266747 51352
rect 264828 51294 266747 51296
rect 173945 51291 174011 51294
rect 266681 51291 266747 51294
rect 142849 51084 142915 51085
rect 142798 51082 142804 51084
rect 142758 51022 142804 51082
rect 142868 51080 142915 51084
rect 142910 51024 142915 51080
rect 142798 51020 142804 51022
rect 142868 51020 142915 51024
rect 142849 51019 142915 51020
rect 79001 50810 79067 50813
rect 76382 50808 79067 50810
rect 76382 50752 79006 50808
rect 79062 50752 79067 50808
rect 76382 50750 79067 50752
rect 79001 50747 79067 50750
rect 93629 50676 93695 50677
rect 93629 50674 93676 50676
rect 93584 50672 93676 50674
rect 93584 50616 93634 50672
rect 93584 50614 93676 50616
rect 93629 50612 93676 50614
rect 93740 50612 93746 50676
rect 139721 50674 139787 50677
rect 142990 50674 143050 51256
rect 233561 50810 233627 50813
rect 237014 50810 237074 51256
rect 327677 50946 327743 50949
rect 331038 50946 331098 51256
rect 429797 51218 429863 51221
rect 434416 51218 434896 51248
rect 429797 51216 434896 51218
rect 429797 51160 429802 51216
rect 429858 51160 434896 51216
rect 429797 51158 434896 51160
rect 429797 51155 429863 51158
rect 434416 51128 434896 51158
rect 327677 50944 331098 50946
rect 327677 50888 327682 50944
rect 327738 50888 331098 50944
rect 327677 50886 331098 50888
rect 327677 50883 327743 50886
rect 233561 50808 237074 50810
rect 233561 50752 233566 50808
rect 233622 50752 237074 50808
rect 233561 50750 237074 50752
rect 233561 50747 233627 50750
rect 187285 50676 187351 50677
rect 187285 50674 187332 50676
rect 139721 50672 143050 50674
rect 139721 50616 139726 50672
rect 139782 50616 143050 50672
rect 139721 50614 143050 50616
rect 187240 50672 187332 50674
rect 187240 50616 187290 50672
rect 187240 50614 187332 50616
rect 93629 50611 93695 50612
rect 139721 50611 139787 50614
rect 187285 50612 187332 50614
rect 187396 50612 187402 50676
rect 280430 50612 280436 50676
rect 280500 50674 280506 50676
rect 281309 50674 281375 50677
rect 280500 50672 281375 50674
rect 280500 50616 281314 50672
rect 281370 50616 281375 50672
rect 280500 50614 281375 50616
rect 280500 50612 280506 50614
rect 187285 50611 187351 50612
rect 281309 50611 281375 50614
rect 139629 50402 139695 50405
rect 174037 50402 174103 50405
rect 139629 50400 143020 50402
rect 76382 50266 76442 50372
rect 139629 50344 139634 50400
rect 139690 50344 143020 50400
rect 139629 50342 143020 50344
rect 170804 50400 174103 50402
rect 170804 50344 174042 50400
rect 174098 50344 174103 50400
rect 170804 50342 174103 50344
rect 139629 50339 139695 50342
rect 174037 50339 174103 50342
rect 191374 50340 191380 50404
rect 191444 50402 191450 50404
rect 191977 50402 192043 50405
rect 191444 50400 192043 50402
rect 191444 50344 191982 50400
rect 192038 50344 192043 50400
rect 191444 50342 192043 50344
rect 191444 50340 191450 50342
rect 191977 50339 192043 50342
rect 233469 50402 233535 50405
rect 266589 50402 266655 50405
rect 233469 50400 237044 50402
rect 233469 50344 233474 50400
rect 233530 50344 237044 50400
rect 233469 50342 237044 50344
rect 264828 50400 266655 50402
rect 264828 50344 266594 50400
rect 266650 50344 266655 50400
rect 264828 50342 266655 50344
rect 233469 50339 233535 50342
rect 266589 50339 266655 50342
rect 328413 50402 328479 50405
rect 328413 50400 331068 50402
rect 328413 50344 328418 50400
rect 328474 50344 331068 50400
rect 328413 50342 331068 50344
rect 328413 50339 328479 50342
rect 78909 50266 78975 50269
rect 107521 50268 107587 50269
rect 76382 50264 78975 50266
rect 76382 50208 78914 50264
rect 78970 50208 78975 50264
rect 76382 50206 78975 50208
rect 78909 50203 78975 50206
rect 107470 50204 107476 50268
rect 107540 50266 107587 50268
rect 107540 50264 107632 50266
rect 107582 50208 107632 50264
rect 107540 50206 107632 50208
rect 107540 50204 107587 50206
rect 109310 50204 109316 50268
rect 109380 50266 109386 50268
rect 109453 50266 109519 50269
rect 109380 50264 109519 50266
rect 109380 50208 109458 50264
rect 109514 50208 109519 50264
rect 109380 50206 109519 50208
rect 109380 50204 109386 50206
rect 107521 50203 107587 50204
rect 109453 50203 109519 50206
rect 199061 50266 199127 50269
rect 199654 50266 199660 50268
rect 199061 50264 199660 50266
rect 199061 50208 199066 50264
rect 199122 50208 199660 50264
rect 199061 50206 199660 50208
rect 199061 50203 199127 50206
rect 199654 50204 199660 50206
rect 199724 50204 199730 50268
rect 274961 49996 275027 49997
rect 274910 49932 274916 49996
rect 274980 49994 275027 49996
rect 327217 49994 327283 49997
rect 330846 49994 330852 49996
rect 274980 49992 275072 49994
rect 275022 49936 275072 49992
rect 274980 49934 275072 49936
rect 327217 49992 330852 49994
rect 327217 49936 327222 49992
rect 327278 49936 330852 49992
rect 327217 49934 330852 49936
rect 274980 49932 275027 49934
rect 274961 49931 275027 49932
rect 327217 49931 327283 49934
rect 330846 49932 330852 49934
rect 330916 49932 330922 49996
rect 76382 49178 76442 49284
rect 87230 49252 87236 49316
rect 87300 49314 87306 49316
rect 87465 49314 87531 49317
rect 87300 49312 87531 49314
rect 87300 49256 87470 49312
rect 87526 49256 87531 49312
rect 87300 49254 87531 49256
rect 87300 49252 87306 49254
rect 87465 49251 87531 49254
rect 105129 49314 105195 49317
rect 105262 49314 105268 49316
rect 105129 49312 105268 49314
rect 105129 49256 105134 49312
rect 105190 49256 105268 49312
rect 105129 49254 105268 49256
rect 105129 49251 105195 49254
rect 105262 49252 105268 49254
rect 105332 49252 105338 49316
rect 173301 49314 173367 49317
rect 181857 49316 181923 49317
rect 181806 49314 181812 49316
rect 170804 49312 173367 49314
rect 170804 49256 173306 49312
rect 173362 49256 173367 49312
rect 170804 49254 173367 49256
rect 181766 49254 181812 49314
rect 181876 49312 181923 49316
rect 181918 49256 181923 49312
rect 173301 49251 173367 49254
rect 181806 49252 181812 49254
rect 181876 49252 181923 49256
rect 181857 49251 181923 49252
rect 203753 49314 203819 49317
rect 204254 49314 204260 49316
rect 203753 49312 204260 49314
rect 203753 49256 203758 49312
rect 203814 49256 204260 49312
rect 203753 49254 204260 49256
rect 203753 49251 203819 49254
rect 204254 49252 204260 49254
rect 204324 49252 204330 49316
rect 266589 49314 266655 49317
rect 264828 49312 266655 49314
rect 264828 49256 266594 49312
rect 266650 49256 266655 49312
rect 264828 49254 266655 49256
rect 266589 49251 266655 49254
rect 274910 49252 274916 49316
rect 274980 49314 274986 49316
rect 275053 49314 275119 49317
rect 274980 49312 275119 49314
rect 274980 49256 275058 49312
rect 275114 49256 275119 49312
rect 274980 49254 275119 49256
rect 274980 49252 274986 49254
rect 275053 49251 275119 49254
rect 78909 49178 78975 49181
rect 76382 49176 78975 49178
rect 76382 49120 78914 49176
rect 78970 49120 78975 49176
rect 76382 49118 78975 49120
rect 78909 49115 78975 49118
rect 140549 49042 140615 49045
rect 142990 49042 143050 49216
rect 140549 49040 143050 49042
rect 140549 48984 140554 49040
rect 140610 48984 143050 49040
rect 140549 48982 143050 48984
rect 233469 49042 233535 49045
rect 237014 49042 237074 49216
rect 233469 49040 237074 49042
rect 233469 48984 233474 49040
rect 233530 48984 237074 49040
rect 233469 48982 237074 48984
rect 328505 49042 328571 49045
rect 331038 49042 331098 49216
rect 328505 49040 331098 49042
rect 328505 48984 328510 49040
rect 328566 48984 331098 49040
rect 328505 48982 331098 48984
rect 140549 48979 140615 48982
rect 233469 48979 233535 48982
rect 328505 48979 328571 48982
rect 174037 48362 174103 48365
rect 266589 48362 266655 48365
rect 170804 48360 174103 48362
rect 67869 48090 67935 48093
rect 73246 48090 73252 48092
rect 67869 48088 73252 48090
rect 67869 48032 67874 48088
rect 67930 48032 73252 48088
rect 67869 48030 73252 48032
rect 67869 48027 67935 48030
rect 73246 48028 73252 48030
rect 73316 48028 73322 48092
rect 74309 48090 74375 48093
rect 75086 48090 75092 48092
rect 74309 48088 75092 48090
rect 74309 48032 74314 48088
rect 74370 48032 75092 48088
rect 74309 48030 75092 48032
rect 74309 48027 74375 48030
rect 75086 48028 75092 48030
rect 75156 48028 75162 48092
rect 76382 48090 76442 48332
rect 170804 48304 174042 48360
rect 174098 48304 174103 48360
rect 170804 48302 174103 48304
rect 264828 48360 266655 48362
rect 264828 48304 266594 48360
rect 266650 48304 266655 48360
rect 264828 48302 266655 48304
rect 174037 48299 174103 48302
rect 266589 48299 266655 48302
rect 87097 48090 87163 48093
rect 76382 48088 87163 48090
rect 76382 48032 87102 48088
rect 87158 48032 87163 48088
rect 76382 48030 87163 48032
rect 87097 48027 87163 48030
rect 87230 48028 87236 48092
rect 87300 48090 87306 48092
rect 88293 48090 88359 48093
rect 105129 48090 105195 48093
rect 87300 48088 105195 48090
rect 87300 48032 88298 48088
rect 88354 48032 105134 48088
rect 105190 48032 105195 48088
rect 87300 48030 105195 48032
rect 87300 48028 87306 48030
rect 88293 48027 88359 48030
rect 105129 48027 105195 48030
rect 139997 48090 140063 48093
rect 142990 48090 143050 48264
rect 139997 48088 143050 48090
rect 139997 48032 140002 48088
rect 140058 48032 143050 48088
rect 139997 48030 143050 48032
rect 147725 48090 147791 48093
rect 147950 48090 147956 48092
rect 147725 48088 147956 48090
rect 147725 48032 147730 48088
rect 147786 48032 147956 48088
rect 147725 48030 147956 48032
rect 139997 48027 140063 48030
rect 147725 48027 147791 48030
rect 147950 48028 147956 48030
rect 148020 48028 148026 48092
rect 153981 48090 154047 48093
rect 154758 48090 154764 48092
rect 153981 48088 154764 48090
rect 153981 48032 153986 48088
rect 154042 48032 154764 48088
rect 153981 48030 154764 48032
rect 153981 48027 154047 48030
rect 154758 48028 154764 48030
rect 154828 48028 154834 48092
rect 167597 48090 167663 48093
rect 168006 48090 168012 48092
rect 167597 48088 168012 48090
rect 167597 48032 167602 48088
rect 167658 48032 168012 48088
rect 167597 48030 168012 48032
rect 167597 48027 167663 48030
rect 168006 48028 168012 48030
rect 168076 48028 168082 48092
rect 160053 47956 160119 47957
rect 72510 47892 72516 47956
rect 72580 47954 72586 47956
rect 75270 47954 75276 47956
rect 72580 47894 75276 47954
rect 72580 47892 72586 47894
rect 75270 47892 75276 47894
rect 75340 47892 75346 47956
rect 144822 47892 144828 47956
rect 144892 47954 144898 47956
rect 147766 47954 147772 47956
rect 144892 47894 147772 47954
rect 144892 47892 144898 47894
rect 147766 47892 147772 47894
rect 147836 47892 147842 47956
rect 160053 47952 160100 47956
rect 160164 47954 160170 47956
rect 160053 47896 160058 47952
rect 160053 47892 160100 47896
rect 160164 47894 160210 47954
rect 160164 47892 160170 47894
rect 168742 47892 168748 47956
rect 168812 47954 168818 47956
rect 168885 47954 168951 47957
rect 182225 47956 182291 47957
rect 182174 47954 182180 47956
rect 168812 47952 168951 47954
rect 168812 47896 168890 47952
rect 168946 47896 168951 47952
rect 168812 47894 168951 47896
rect 182134 47894 182180 47954
rect 182244 47952 182291 47956
rect 182286 47896 182291 47952
rect 168812 47892 168818 47894
rect 160053 47891 160119 47892
rect 168885 47891 168951 47894
rect 182174 47892 182180 47894
rect 182244 47892 182291 47896
rect 182225 47891 182291 47892
rect 166401 47818 166467 47821
rect 169662 47818 169668 47820
rect 166401 47816 169668 47818
rect 166401 47760 166406 47816
rect 166462 47760 169668 47816
rect 166401 47758 169668 47760
rect 166401 47755 166467 47758
rect 169662 47756 169668 47758
rect 169732 47756 169738 47820
rect 233469 47818 233535 47821
rect 237014 47818 237074 48264
rect 237558 48028 237564 48092
rect 237628 48090 237634 48092
rect 241105 48090 241171 48093
rect 237628 48088 241171 48090
rect 237628 48032 241110 48088
rect 241166 48032 241171 48088
rect 237628 48030 241171 48032
rect 237628 48028 237634 48030
rect 241105 48027 241171 48030
rect 262398 48028 262404 48092
rect 262468 48090 262474 48092
rect 262909 48090 262975 48093
rect 262468 48088 262975 48090
rect 262468 48032 262914 48088
rect 262970 48032 262975 48088
rect 262468 48030 262975 48032
rect 262468 48028 262474 48030
rect 262909 48027 262975 48030
rect 263870 48028 263876 48092
rect 263940 48090 263946 48092
rect 264473 48090 264539 48093
rect 283701 48090 283767 48093
rect 263940 48088 283767 48090
rect 263940 48032 264478 48088
rect 264534 48032 283706 48088
rect 283762 48032 283767 48088
rect 263940 48030 283767 48032
rect 263940 48028 263946 48030
rect 264473 48027 264539 48030
rect 283701 48027 283767 48030
rect 244877 47954 244943 47957
rect 253985 47956 254051 47957
rect 248598 47954 248604 47956
rect 244877 47952 248604 47954
rect 244877 47896 244882 47952
rect 244938 47896 248604 47952
rect 244877 47894 248604 47896
rect 244877 47891 244943 47894
rect 248598 47892 248604 47894
rect 248668 47892 248674 47956
rect 253934 47954 253940 47956
rect 253894 47894 253940 47954
rect 254004 47952 254051 47956
rect 254046 47896 254051 47952
rect 253934 47892 253940 47894
rect 254004 47892 254051 47896
rect 274910 47892 274916 47956
rect 274980 47954 274986 47956
rect 275789 47954 275855 47957
rect 274980 47952 275855 47954
rect 274980 47896 275794 47952
rect 275850 47896 275855 47952
rect 274980 47894 275855 47896
rect 274980 47892 274986 47894
rect 253985 47891 254051 47892
rect 275789 47891 275855 47894
rect 328045 47954 328111 47957
rect 331038 47954 331098 48264
rect 328045 47952 331098 47954
rect 328045 47896 328050 47952
rect 328106 47896 331098 47952
rect 328045 47894 331098 47896
rect 328045 47891 328111 47894
rect 233469 47816 237074 47818
rect 233469 47760 233474 47816
rect 233530 47760 237074 47816
rect 233469 47758 237074 47760
rect 233469 47755 233535 47758
rect 113593 47548 113659 47549
rect 74166 47484 74172 47548
rect 74236 47546 74242 47548
rect 75454 47546 75460 47548
rect 74236 47486 75460 47546
rect 74236 47484 74242 47486
rect 75454 47484 75460 47486
rect 75524 47484 75530 47548
rect 113542 47546 113548 47548
rect 113502 47486 113548 47546
rect 113612 47544 113659 47548
rect 113654 47488 113659 47544
rect 113542 47484 113548 47486
rect 113612 47484 113659 47488
rect 113593 47483 113659 47484
rect 72561 47412 72627 47413
rect 72510 47410 72516 47412
rect 72470 47350 72516 47410
rect 72580 47408 72627 47412
rect 72622 47352 72627 47408
rect 72510 47348 72516 47350
rect 72580 47348 72627 47352
rect 74166 47348 74172 47412
rect 74236 47410 74242 47412
rect 74677 47410 74743 47413
rect 74236 47408 74743 47410
rect 74236 47352 74682 47408
rect 74738 47352 74743 47408
rect 74236 47350 74743 47352
rect 74236 47348 74242 47350
rect 72561 47347 72627 47348
rect 74677 47347 74743 47350
rect 106601 47410 106667 47413
rect 107470 47410 107476 47412
rect 106601 47408 107476 47410
rect 106601 47352 106606 47408
rect 106662 47352 107476 47408
rect 106601 47350 107476 47352
rect 106601 47347 106667 47350
rect 107470 47348 107476 47350
rect 107540 47348 107546 47412
rect 263870 47348 263876 47412
rect 263940 47410 263946 47412
rect 264422 47410 264428 47412
rect 263940 47350 264428 47410
rect 263940 47348 263946 47350
rect 264422 47348 264428 47350
rect 264492 47410 264498 47412
rect 285909 47410 285975 47413
rect 264492 47408 285975 47410
rect 264492 47352 285914 47408
rect 285970 47352 285975 47408
rect 264492 47350 285975 47352
rect 264492 47348 264498 47350
rect 285909 47347 285975 47350
rect 109310 47212 109316 47276
rect 109380 47274 109386 47276
rect 109453 47274 109519 47277
rect 110414 47274 110420 47276
rect 109380 47272 110420 47274
rect 109380 47216 109458 47272
rect 109514 47216 110420 47272
rect 109380 47214 110420 47216
rect 109380 47212 109386 47214
rect 109453 47211 109519 47214
rect 110414 47212 110420 47214
rect 110484 47212 110490 47276
rect 162854 47212 162860 47276
rect 162924 47274 162930 47276
rect 162997 47274 163063 47277
rect 162924 47272 163063 47274
rect 162924 47216 163002 47272
rect 163058 47216 163063 47272
rect 162924 47214 163063 47216
rect 162924 47212 162930 47214
rect 162997 47211 163063 47214
rect 248005 47274 248071 47277
rect 248598 47274 248604 47276
rect 248005 47272 248604 47274
rect 248005 47216 248010 47272
rect 248066 47216 248604 47272
rect 248005 47214 248604 47216
rect 248005 47211 248071 47214
rect 248598 47212 248604 47214
rect 248668 47212 248674 47276
rect 181070 46532 181076 46596
rect 181140 46594 181146 46596
rect 182133 46594 182199 46597
rect 260333 46596 260399 46597
rect 275881 46596 275947 46597
rect 260333 46594 260380 46596
rect 181140 46592 182199 46594
rect 181140 46536 182138 46592
rect 182194 46536 182199 46592
rect 181140 46534 182199 46536
rect 260288 46592 260380 46594
rect 260288 46536 260338 46592
rect 260288 46534 260380 46536
rect 181140 46532 181146 46534
rect 182133 46531 182199 46534
rect 260333 46532 260380 46534
rect 260444 46532 260450 46596
rect 275830 46532 275836 46596
rect 275900 46594 275947 46596
rect 275900 46592 275992 46594
rect 275942 46536 275992 46592
rect 275900 46534 275992 46536
rect 275900 46532 275947 46534
rect 260333 46531 260399 46532
rect 275881 46531 275947 46532
rect 9896 46458 10376 46488
rect 13037 46458 13103 46461
rect 9896 46456 13103 46458
rect 9896 46400 13042 46456
rect 13098 46400 13103 46456
rect 9896 46398 13103 46400
rect 9896 46368 10376 46398
rect 13037 46395 13103 46398
rect 158990 45988 158996 46052
rect 159060 46050 159066 46052
rect 168885 46050 168951 46053
rect 159060 46048 168951 46050
rect 159060 45992 168890 46048
rect 168946 45992 168951 46048
rect 159060 45990 168951 45992
rect 159060 45988 159066 45990
rect 168885 45987 168951 45990
rect 252646 45988 252652 46052
rect 252716 46050 252722 46052
rect 256929 46050 256995 46053
rect 252716 46048 256995 46050
rect 252716 45992 256934 46048
rect 256990 45992 256995 46048
rect 252716 45990 256995 45992
rect 252716 45988 252722 45990
rect 256929 45987 256995 45990
rect 263185 46050 263251 46053
rect 263502 46050 263508 46052
rect 263185 46048 263508 46050
rect 263185 45992 263190 46048
rect 263246 45992 263508 46048
rect 263185 45990 263508 45992
rect 263185 45987 263251 45990
rect 263502 45988 263508 45990
rect 263572 45988 263578 46052
rect 346629 46050 346695 46053
rect 356790 46050 356796 46052
rect 346629 46048 356796 46050
rect 346629 45992 346634 46048
rect 346690 45992 356796 46048
rect 346629 45990 356796 45992
rect 346629 45987 346695 45990
rect 356790 45988 356796 45990
rect 356860 45988 356866 46052
rect 64189 45914 64255 45917
rect 73246 45914 73252 45916
rect 64189 45912 73252 45914
rect 64189 45856 64194 45912
rect 64250 45856 73252 45912
rect 64189 45854 73252 45856
rect 64189 45851 64255 45854
rect 73246 45852 73252 45854
rect 73316 45852 73322 45916
rect 157518 45852 157524 45916
rect 157588 45914 157594 45916
rect 165941 45914 166007 45917
rect 157588 45912 166007 45914
rect 157588 45856 165946 45912
rect 166002 45856 166007 45912
rect 157588 45854 166007 45856
rect 157588 45852 157594 45854
rect 165941 45851 166007 45854
rect 147950 45716 147956 45780
rect 148020 45778 148026 45780
rect 162997 45778 163063 45781
rect 148020 45776 163063 45778
rect 148020 45720 163002 45776
rect 163058 45720 163063 45776
rect 148020 45718 163063 45720
rect 148020 45716 148026 45718
rect 162997 45715 163063 45718
rect 251133 45778 251199 45781
rect 263318 45778 263324 45780
rect 251133 45776 263324 45778
rect 251133 45720 251138 45776
rect 251194 45720 263324 45776
rect 251133 45718 263324 45720
rect 251133 45715 251199 45718
rect 263318 45716 263324 45718
rect 263388 45716 263394 45780
rect 331398 45308 331404 45372
rect 331468 45370 331474 45372
rect 338349 45370 338415 45373
rect 331468 45368 338415 45370
rect 331468 45312 338354 45368
rect 338410 45312 338415 45368
rect 331468 45310 338415 45312
rect 331468 45308 331474 45310
rect 338349 45307 338415 45310
rect 169713 44828 169779 44829
rect 169662 44764 169668 44828
rect 169732 44826 169779 44828
rect 169732 44824 169824 44826
rect 169774 44768 169824 44824
rect 169732 44766 169824 44768
rect 169732 44764 169779 44766
rect 169713 44763 169779 44764
rect 118142 44628 118148 44692
rect 118212 44690 118218 44692
rect 118653 44690 118719 44693
rect 118212 44688 118719 44690
rect 118212 44632 118658 44688
rect 118714 44632 118719 44688
rect 118212 44630 118719 44632
rect 118212 44628 118218 44630
rect 118653 44627 118719 44630
rect 211982 43404 211988 43468
rect 212052 43466 212058 43468
rect 212585 43466 212651 43469
rect 212052 43464 212651 43466
rect 212052 43408 212590 43464
rect 212646 43408 212651 43464
rect 212052 43406 212651 43408
rect 212052 43404 212058 43406
rect 212585 43403 212651 43406
rect 207525 39114 207591 39117
rect 301549 39116 301615 39117
rect 207750 39114 207756 39116
rect 207525 39112 207756 39114
rect 207525 39056 207530 39112
rect 207586 39056 207756 39112
rect 207525 39054 207756 39056
rect 207525 39051 207591 39054
rect 207750 39052 207756 39054
rect 207820 39052 207826 39116
rect 301549 39114 301596 39116
rect 301504 39112 301596 39114
rect 301504 39056 301554 39112
rect 301504 39054 301596 39056
rect 301549 39052 301596 39054
rect 301660 39052 301666 39116
rect 428693 39114 428759 39117
rect 434416 39114 434896 39144
rect 428693 39112 434896 39114
rect 428693 39056 428698 39112
rect 428754 39056 434896 39112
rect 428693 39054 434896 39056
rect 301549 39051 301615 39052
rect 428693 39051 428759 39054
rect 434416 39024 434896 39054
rect 306609 37754 306675 37757
rect 307110 37754 307116 37756
rect 306609 37752 307116 37754
rect 306609 37696 306614 37752
rect 306670 37696 307116 37752
rect 306609 37694 307116 37696
rect 306609 37691 306675 37694
rect 307110 37692 307116 37694
rect 307180 37692 307186 37756
rect 9896 35714 10376 35744
rect 12853 35714 12919 35717
rect 9896 35712 12919 35714
rect 9896 35656 12858 35712
rect 12914 35656 12919 35712
rect 9896 35654 12919 35656
rect 9896 35624 10376 35654
rect 12853 35651 12919 35654
rect 88109 33674 88175 33677
rect 181949 33674 182015 33677
rect 275789 33674 275855 33677
rect 88109 33672 90058 33674
rect 88109 33616 88114 33672
rect 88170 33616 90058 33672
rect 88109 33614 90058 33616
rect 88109 33611 88175 33614
rect 89998 33444 90058 33614
rect 181949 33672 184082 33674
rect 181949 33616 181954 33672
rect 182010 33616 184082 33672
rect 181949 33614 184082 33616
rect 181949 33611 182015 33614
rect 184022 33444 184082 33614
rect 275789 33672 278106 33674
rect 275789 33616 275794 33672
rect 275850 33616 278106 33672
rect 275789 33614 278106 33616
rect 275789 33611 275855 33614
rect 278046 33444 278106 33614
rect 88201 30818 88267 30821
rect 182041 30818 182107 30821
rect 275881 30818 275947 30821
rect 88201 30816 90058 30818
rect 88201 30760 88206 30816
rect 88262 30760 90058 30816
rect 88201 30758 90058 30760
rect 88201 30755 88267 30758
rect 89998 30724 90058 30758
rect 182041 30816 184082 30818
rect 182041 30760 182046 30816
rect 182102 30760 184082 30816
rect 182041 30758 184082 30760
rect 182041 30755 182107 30758
rect 184022 30724 184082 30758
rect 275881 30816 278106 30818
rect 275881 30760 275886 30816
rect 275942 30760 278106 30816
rect 275881 30758 278106 30760
rect 275881 30755 275947 30758
rect 278046 30724 278106 30758
rect 88293 28098 88359 28101
rect 89998 28098 90058 28136
rect 88293 28096 90058 28098
rect 88293 28040 88298 28096
rect 88354 28040 90058 28096
rect 88293 28038 90058 28040
rect 182133 28098 182199 28101
rect 184022 28098 184082 28136
rect 182133 28096 184082 28098
rect 182133 28040 182138 28096
rect 182194 28040 184082 28096
rect 182133 28038 184082 28040
rect 275973 28098 276039 28101
rect 278046 28098 278106 28136
rect 275973 28096 278106 28098
rect 275973 28040 275978 28096
rect 276034 28040 278106 28096
rect 275973 28038 278106 28040
rect 88293 28035 88359 28038
rect 182133 28035 182199 28038
rect 275973 28035 276039 28038
rect 429429 27010 429495 27013
rect 434416 27010 434896 27040
rect 429429 27008 434896 27010
rect 429429 26952 429434 27008
rect 429490 26952 434896 27008
rect 429429 26950 434896 26952
rect 429429 26947 429495 26950
rect 434416 26920 434896 26950
rect 88385 26058 88451 26061
rect 182225 26058 182291 26061
rect 276065 26058 276131 26061
rect 88385 26056 90058 26058
rect 88385 26000 88390 26056
rect 88446 26000 90058 26056
rect 88385 25998 90058 26000
rect 88385 25995 88451 25998
rect 89998 25420 90058 25998
rect 182225 26056 184082 26058
rect 182225 26000 182230 26056
rect 182286 26000 184082 26056
rect 182225 25998 184082 26000
rect 182225 25995 182291 25998
rect 184022 25420 184082 25998
rect 276065 26056 278106 26058
rect 276065 26000 276070 26056
rect 276126 26000 278106 26056
rect 276065 25998 278106 26000
rect 276065 25995 276131 25998
rect 278046 25420 278106 25998
rect 9896 24970 10376 25000
rect 12669 24970 12735 24973
rect 9896 24968 12735 24970
rect 9896 24912 12674 24968
rect 12730 24912 12735 24968
rect 9896 24910 12735 24912
rect 9896 24880 10376 24910
rect 12669 24907 12735 24910
rect 88017 23338 88083 23341
rect 181857 23338 181923 23341
rect 275605 23338 275671 23341
rect 88017 23336 90058 23338
rect 88017 23280 88022 23336
rect 88078 23280 90058 23336
rect 88017 23278 90058 23280
rect 88017 23275 88083 23278
rect 89998 22700 90058 23278
rect 181857 23336 184082 23338
rect 181857 23280 181862 23336
rect 181918 23280 184082 23336
rect 181857 23278 184082 23280
rect 181857 23275 181923 23278
rect 184022 22700 184082 23278
rect 275605 23336 278106 23338
rect 275605 23280 275610 23336
rect 275666 23280 278106 23336
rect 275605 23278 278106 23280
rect 275605 23275 275671 23278
rect 278046 22700 278106 23278
rect 88477 20754 88543 20757
rect 182317 20754 182383 20757
rect 276157 20754 276223 20757
rect 88477 20752 90058 20754
rect 88477 20696 88482 20752
rect 88538 20696 90058 20752
rect 88477 20694 90058 20696
rect 88477 20691 88543 20694
rect 89998 20116 90058 20694
rect 182317 20752 184082 20754
rect 182317 20696 182322 20752
rect 182378 20696 184082 20752
rect 182317 20694 184082 20696
rect 182317 20691 182383 20694
rect 184022 20116 184082 20694
rect 276157 20752 278106 20754
rect 276157 20696 276162 20752
rect 276218 20696 278106 20752
rect 276157 20694 278106 20696
rect 276157 20691 276223 20694
rect 278046 20116 278106 20694
rect 429429 14906 429495 14909
rect 434416 14906 434896 14936
rect 429429 14904 434896 14906
rect 429429 14848 429434 14904
rect 429490 14848 434896 14904
rect 429429 14846 434896 14848
rect 429429 14843 429495 14846
rect 434416 14816 434896 14846
rect 9896 14226 10376 14256
rect 12669 14226 12735 14229
rect 9896 14224 12735 14226
rect 9896 14168 12674 14224
rect 12730 14168 12735 14224
rect 9896 14166 12735 14168
rect 9896 14136 10376 14166
rect 12669 14163 12735 14166
<< via3 >>
rect 341708 393740 341772 393804
rect 191196 359332 191260 359396
rect 284484 356536 284548 356540
rect 284484 356480 284534 356536
rect 284534 356480 284548 356536
rect 284484 356476 284548 356480
rect 96804 355312 96868 355316
rect 96804 355256 96854 355312
rect 96854 355256 96868 355312
rect 96804 355252 96868 355256
rect 191196 351912 191260 351916
rect 191196 351856 191246 351912
rect 191246 351856 191260 351912
rect 191196 351852 191260 351856
rect 96804 351640 96868 351644
rect 96804 351584 96818 351640
rect 96818 351584 96868 351640
rect 96804 351580 96868 351584
rect 284484 351640 284548 351644
rect 284484 351584 284534 351640
rect 284534 351584 284548 351640
rect 284484 351580 284548 351584
rect 104900 333764 104964 333828
rect 212172 333492 212236 333556
rect 295524 333084 295588 333148
rect 137284 332132 137348 332196
rect 201684 332132 201748 332196
rect 230940 332192 231004 332196
rect 230940 332136 230954 332192
rect 230954 332136 231004 332192
rect 230940 332132 231004 332136
rect 204444 331588 204508 331652
rect 230940 331588 231004 331652
rect 299388 331452 299452 331516
rect 137284 330772 137348 330836
rect 231308 330772 231372 330836
rect 292764 330772 292828 330836
rect 158628 330152 158692 330156
rect 158628 330096 158642 330152
rect 158642 330096 158692 330152
rect 158628 330092 158692 330096
rect 159548 330152 159612 330156
rect 159548 330096 159598 330152
rect 159598 330096 159612 330152
rect 159548 330092 159612 330096
rect 251916 330152 251980 330156
rect 251916 330096 251966 330152
rect 251966 330096 251980 330152
rect 251916 330092 251980 330096
rect 252652 330152 252716 330156
rect 252652 330096 252666 330152
rect 252666 330096 252716 330152
rect 252652 330092 252716 330096
rect 137468 328732 137532 328796
rect 161756 328792 161820 328796
rect 161756 328736 161770 328792
rect 161770 328736 161820 328792
rect 161756 328732 161820 328736
rect 230940 328792 231004 328796
rect 230940 328736 230990 328792
rect 230990 328736 231004 328792
rect 230940 328732 231004 328736
rect 231860 328732 231924 328796
rect 253388 328732 253452 328796
rect 137468 328052 137532 328116
rect 160652 328112 160716 328116
rect 160652 328056 160702 328112
rect 160702 328056 160716 328112
rect 160652 328052 160716 328056
rect 208676 328112 208740 328116
rect 208676 328056 208726 328112
rect 208726 328056 208740 328112
rect 208676 328052 208740 328056
rect 339500 327372 339564 327436
rect 340972 327372 341036 327436
rect 336372 326828 336436 326892
rect 52644 326284 52708 326348
rect 54668 326284 54732 326348
rect 55036 326344 55100 326348
rect 55036 326288 55086 326344
rect 55086 326288 55100 326344
rect 55036 326284 55100 326288
rect 55956 326284 56020 326348
rect 353300 320164 353364 320228
rect 246212 316960 246276 316964
rect 246212 316904 246226 316960
rect 246226 316904 246276 316960
rect 246212 316900 246276 316904
rect 345572 316492 345636 316556
rect 55956 315812 56020 315876
rect 355692 315268 355756 315332
rect 345572 315132 345636 315196
rect 340972 314860 341036 314924
rect 351828 314860 351892 314924
rect 339500 314588 339564 314652
rect 352012 314588 352076 314652
rect 54852 310916 54916 310980
rect 55036 310916 55100 310980
rect 55036 308196 55100 308260
rect 73436 308196 73500 308260
rect 54668 306156 54732 306220
rect 429476 305748 429540 305812
rect 55036 300912 55100 300916
rect 55036 300856 55086 300912
rect 55086 300856 55100 300912
rect 55036 300852 55100 300856
rect 52644 300580 52708 300644
rect 74540 298676 74604 298740
rect 134708 298132 134772 298196
rect 322756 295412 322820 295476
rect 136916 295276 136980 295340
rect 230756 295276 230820 295340
rect 322756 293372 322820 293436
rect 137836 292692 137900 292756
rect 322756 292284 322820 292348
rect 229284 292148 229348 292212
rect 55036 292012 55100 292076
rect 165620 291876 165684 291940
rect 178684 291876 178748 291940
rect 259460 291876 259524 291940
rect 272708 291876 272772 291940
rect 74172 291664 74236 291668
rect 74172 291608 74222 291664
rect 74222 291608 74236 291664
rect 74172 291604 74236 291608
rect 229284 291332 229348 291396
rect 231860 291332 231924 291396
rect 258724 291332 258788 291396
rect 263692 291332 263756 291396
rect 228732 289564 228796 289628
rect 322756 289564 322820 289628
rect 55036 288986 55100 289050
rect 74356 289080 74420 289084
rect 74356 289024 74406 289080
rect 74406 289024 74420 289080
rect 137836 289292 137900 289356
rect 74356 289020 74420 289024
rect 236092 289080 236156 289084
rect 236092 289024 236106 289080
rect 236106 289024 236156 289080
rect 236092 289020 236156 289024
rect 74172 288884 74236 288948
rect 74356 288808 74420 288812
rect 74356 288752 74370 288808
rect 74370 288752 74420 288808
rect 74356 288748 74420 288752
rect 54484 287524 54548 287588
rect 55036 287524 55100 287588
rect 353668 285272 353732 285276
rect 353668 285216 353718 285272
rect 353718 285216 353732 285272
rect 353668 285212 353732 285216
rect 138572 284804 138636 284868
rect 84476 284592 84540 284596
rect 84476 284536 84526 284592
rect 84526 284536 84540 284592
rect 84476 284532 84540 284536
rect 13636 283580 13700 283644
rect 73620 282764 73684 282828
rect 84660 282764 84724 282828
rect 137284 282220 137348 282284
rect 84660 281872 84724 281876
rect 84660 281816 84674 281872
rect 84674 281816 84724 281872
rect 84660 281812 84724 281816
rect 84660 281132 84724 281196
rect 352748 279636 352812 279700
rect 74172 279364 74236 279428
rect 74356 279364 74420 279428
rect 54668 279228 54732 279292
rect 54668 278956 54732 279020
rect 138572 278200 138636 278204
rect 138572 278144 138622 278200
rect 138622 278144 138636 278200
rect 138572 278140 138636 278144
rect 415124 277188 415188 277252
rect 167828 274604 167892 274668
rect 247868 274664 247932 274668
rect 247868 274608 247918 274664
rect 247918 274608 247932 274664
rect 247868 274604 247932 274608
rect 149060 274468 149124 274532
rect 168564 274468 168628 274532
rect 262404 274468 262468 274532
rect 169116 274332 169180 274396
rect 247868 274332 247932 274396
rect 262956 274332 263020 274396
rect 136916 273788 136980 273852
rect 242348 273788 242412 273852
rect 241980 273652 242044 273716
rect 246212 273652 246276 273716
rect 54484 272292 54548 272356
rect 55036 272292 55100 272356
rect 261852 272156 261916 272220
rect 138572 269768 138636 269772
rect 138572 269712 138622 269768
rect 138622 269712 138636 269768
rect 138572 269708 138636 269712
rect 276756 269436 276820 269500
rect 219716 268348 219780 268412
rect 261852 268212 261916 268276
rect 262220 268212 262284 268276
rect 52644 266716 52708 266780
rect 54668 266716 54732 266780
rect 55036 266716 55100 266780
rect 55956 266716 56020 266780
rect 351828 266716 351892 266780
rect 352012 266580 352076 266644
rect 74356 266036 74420 266100
rect 75276 266036 75340 266100
rect 73436 265900 73500 265964
rect 74356 265900 74420 265964
rect 73988 263452 74052 263516
rect 74356 263452 74420 263516
rect 74540 263452 74604 263516
rect 75644 263452 75708 263516
rect 237196 263452 237260 263516
rect 242348 263452 242412 263516
rect 144092 263316 144156 263380
rect 149060 263316 149124 263380
rect 237564 263316 237628 263380
rect 241980 263316 242044 263380
rect 138572 262772 138636 262836
rect 138756 262500 138820 262564
rect 138756 259976 138820 259980
rect 138756 259920 138806 259976
rect 138806 259920 138820 259976
rect 138756 259916 138820 259920
rect 48596 255972 48660 256036
rect 358636 255836 358700 255900
rect 236644 254068 236708 254132
rect 237196 254068 237260 254132
rect 360476 252844 360540 252908
rect 49148 252300 49212 252364
rect 138940 250396 139004 250460
rect 325148 250260 325212 250324
rect 49148 249172 49212 249236
rect 358636 249172 358700 249236
rect 48412 246588 48476 246652
rect 138940 243596 139004 243660
rect 49148 243324 49212 243388
rect 138756 243324 138820 243388
rect 96068 241692 96132 241756
rect 104900 241692 104964 241756
rect 76564 241012 76628 241076
rect 93860 241012 93924 241076
rect 106556 240332 106620 240396
rect 118700 240332 118764 240396
rect 303804 240332 303868 240396
rect 125876 240196 125940 240260
rect 128636 240196 128700 240260
rect 49148 239788 49212 239852
rect 95148 239712 95212 239716
rect 95148 239656 95198 239712
rect 95198 239656 95212 239712
rect 95148 239652 95212 239656
rect 187884 239652 187948 239716
rect 211252 239652 211316 239716
rect 290556 239712 290620 239716
rect 290556 239656 290570 239712
rect 290570 239656 290620 239712
rect 290556 239652 290620 239656
rect 92572 239380 92636 239444
rect 284300 239380 284364 239444
rect 230940 239032 231004 239036
rect 230940 238976 230990 239032
rect 230990 238976 231004 239032
rect 230940 238972 231004 238976
rect 325332 238972 325396 239036
rect 102324 238564 102388 238628
rect 142804 238352 142868 238356
rect 142804 238296 142818 238352
rect 142818 238296 142868 238352
rect 142804 238292 142868 238296
rect 200028 238292 200092 238356
rect 231860 238292 231924 238356
rect 286876 238352 286940 238356
rect 286876 238296 286926 238352
rect 286926 238296 286940 238352
rect 286876 238292 286940 238296
rect 219716 237808 219780 237812
rect 219716 237752 219766 237808
rect 219766 237752 219780 237808
rect 219716 237748 219780 237752
rect 183836 236932 183900 236996
rect 73988 236388 74052 236452
rect 74172 236388 74236 236452
rect 74172 236252 74236 236316
rect 75828 236252 75892 236316
rect 149244 236252 149308 236316
rect 153476 236252 153540 236316
rect 162860 236252 162924 236316
rect 149612 236116 149676 236180
rect 238116 236116 238180 236180
rect 248788 236116 248852 236180
rect 148692 236040 148756 236044
rect 148692 235984 148706 236040
rect 148706 235984 148756 236040
rect 148692 235980 148756 235984
rect 147956 235844 148020 235908
rect 262036 235844 262100 235908
rect 110420 235708 110484 235772
rect 262404 235708 262468 235772
rect 74724 235632 74788 235636
rect 74724 235576 74738 235632
rect 74738 235576 74788 235632
rect 74724 235572 74788 235576
rect 75828 235572 75892 235636
rect 74540 235028 74604 235092
rect 136916 235088 136980 235092
rect 136916 235032 136966 235088
rect 136966 235032 136980 235088
rect 136916 235028 136980 235032
rect 74540 234892 74604 234956
rect 137836 234892 137900 234956
rect 145012 234892 145076 234956
rect 152004 234952 152068 234956
rect 152004 234896 152054 234952
rect 152054 234896 152068 234952
rect 152004 234892 152068 234896
rect 207204 234952 207268 234956
rect 207204 234896 207254 234952
rect 207254 234896 207268 234952
rect 207204 234892 207268 234896
rect 231860 234952 231924 234956
rect 231860 234896 231874 234952
rect 231874 234896 231924 234952
rect 231860 234892 231924 234896
rect 234804 234892 234868 234956
rect 237748 234892 237812 234956
rect 244372 234892 244436 234956
rect 301044 234892 301108 234956
rect 284300 234348 284364 234412
rect 141148 234212 141212 234276
rect 147772 234212 147836 234276
rect 147956 234212 148020 234276
rect 153108 234212 153172 234276
rect 246028 234272 246092 234276
rect 246028 234216 246042 234272
rect 246042 234216 246092 234272
rect 246028 234212 246092 234216
rect 73804 233940 73868 234004
rect 73436 233804 73500 233868
rect 75460 233804 75524 233868
rect 73436 233668 73500 233732
rect 73804 233668 73868 233732
rect 169116 233668 169180 233732
rect 153108 233532 153172 233596
rect 167828 233532 167892 233596
rect 249892 233532 249956 233596
rect 290004 233532 290068 233596
rect 297548 233532 297612 233596
rect 262956 233396 263020 233460
rect 259644 232852 259708 232916
rect 269212 232852 269276 232916
rect 282644 232852 282708 232916
rect 285220 232852 285284 232916
rect 52644 232444 52708 232508
rect 54668 232444 54732 232508
rect 351644 232444 351708 232508
rect 351828 232444 351892 232508
rect 55404 230948 55468 231012
rect 74172 231008 74236 231012
rect 74172 230952 74222 231008
rect 74222 230952 74236 231008
rect 74172 230948 74236 230952
rect 55588 229648 55652 229652
rect 55588 229592 55602 229648
rect 55602 229592 55652 229648
rect 55588 229588 55652 229592
rect 73988 229044 74052 229108
rect 74356 229044 74420 229108
rect 73988 228908 74052 228972
rect 74540 228908 74604 228972
rect 324596 228228 324660 228292
rect 325516 228228 325580 228292
rect 276756 226596 276820 226660
rect 92572 226460 92636 226524
rect 355692 225372 355756 225436
rect 324964 224284 325028 224348
rect 55404 221972 55468 222036
rect 358636 221972 358700 222036
rect 405924 221972 405988 222036
rect 74356 221428 74420 221492
rect 55588 221292 55652 221356
rect 56324 221292 56388 221356
rect 322940 217076 323004 217140
rect 242716 216940 242780 217004
rect 258724 216940 258788 217004
rect 272708 216940 272772 217004
rect 336924 216940 336988 217004
rect 352748 216940 352812 217004
rect 148692 216532 148756 216596
rect 164884 216532 164948 216596
rect 177580 216532 177644 216596
rect 228916 216532 228980 216596
rect 242716 216532 242780 216596
rect 258724 216532 258788 216596
rect 272708 216532 272772 216596
rect 322940 216532 323004 216596
rect 336740 216532 336804 216596
rect 352748 216532 352812 216596
rect 357532 215852 357596 215916
rect 405924 215852 405988 215916
rect 73436 214492 73500 214556
rect 73804 214492 73868 214556
rect 74172 213192 74236 213196
rect 74172 213136 74222 213192
rect 74222 213136 74236 213192
rect 74172 213132 74236 213136
rect 74356 211696 74420 211700
rect 74356 211640 74406 211696
rect 74406 211640 74420 211696
rect 74356 211636 74420 211640
rect 54668 210956 54732 211020
rect 147036 208236 147100 208300
rect 231860 207692 231924 207756
rect 52644 206740 52708 206804
rect 73988 206604 74052 206668
rect 74356 205440 74420 205444
rect 74356 205384 74406 205440
rect 74406 205384 74420 205440
rect 74356 205380 74420 205384
rect 73436 204972 73500 205036
rect 134708 204972 134772 205036
rect 73436 204836 73500 204900
rect 73988 204836 74052 204900
rect 73620 204428 73684 204492
rect 84660 204428 84724 204492
rect 73620 203204 73684 203268
rect 137836 200892 137900 200956
rect 322756 200892 322820 200956
rect 230756 200620 230820 200684
rect 74356 200544 74420 200548
rect 74356 200488 74370 200544
rect 74370 200488 74420 200544
rect 74356 200484 74420 200488
rect 73804 199320 73868 199324
rect 73804 199264 73818 199320
rect 73818 199264 73868 199320
rect 73804 199260 73868 199264
rect 74172 199260 74236 199324
rect 74540 199124 74604 199188
rect 322756 198716 322820 198780
rect 138020 198172 138084 198236
rect 230756 198232 230820 198236
rect 230756 198176 230770 198232
rect 230770 198176 230820 198232
rect 230756 198172 230820 198176
rect 73988 197900 74052 197964
rect 74540 197900 74604 197964
rect 74172 195180 74236 195244
rect 74540 195180 74604 195244
rect 138020 194636 138084 194700
rect 322756 194772 322820 194836
rect 236092 194500 236156 194564
rect 228732 194364 228796 194428
rect 352748 191372 352812 191436
rect 74356 191024 74420 191028
rect 74356 190968 74370 191024
rect 74370 190968 74420 191024
rect 74356 190964 74420 190968
rect 73804 189528 73868 189532
rect 73804 189472 73818 189528
rect 73818 189472 73868 189528
rect 73804 189468 73868 189472
rect 74540 187080 74604 187084
rect 74540 187024 74554 187080
rect 74554 187024 74604 187080
rect 74540 187020 74604 187024
rect 74540 186884 74604 186948
rect 351644 184028 351708 184092
rect 242532 183076 242596 183140
rect 271420 182124 271484 182188
rect 323124 182124 323188 182188
rect 174820 181988 174884 182052
rect 228732 181988 228796 182052
rect 323492 181988 323556 182052
rect 74356 181232 74420 181236
rect 74356 181176 74406 181232
rect 74406 181176 74420 181232
rect 74356 181172 74420 181176
rect 147036 181172 147100 181236
rect 267556 181232 267620 181236
rect 267556 181176 267570 181232
rect 267570 181176 267620 181232
rect 267556 181172 267620 181176
rect 168564 181036 168628 181100
rect 167828 180900 167892 180964
rect 169300 180764 169364 180828
rect 261668 180764 261732 180828
rect 167644 180628 167708 180692
rect 262404 180628 262468 180692
rect 141516 180492 141580 180556
rect 262956 180492 263020 180556
rect 242348 180220 242412 180284
rect 241796 180084 241860 180148
rect 73804 180008 73868 180012
rect 73804 179952 73818 180008
rect 73818 179952 73868 180008
rect 73804 179948 73868 179952
rect 74172 179948 74236 180012
rect 242532 179948 242596 180012
rect 309876 179268 309940 179332
rect 312636 179268 312700 179332
rect 311164 179132 311228 179196
rect 313740 179132 313804 179196
rect 74540 175732 74604 175796
rect 75092 175732 75156 175796
rect 219716 175460 219780 175524
rect 182916 174976 182980 174980
rect 182916 174920 182966 174976
rect 182966 174920 182980 174976
rect 182916 174916 182980 174920
rect 241796 173964 241860 174028
rect 242532 173964 242596 174028
rect 148692 173072 148756 173076
rect 148692 173016 148742 173072
rect 148742 173016 148756 173072
rect 148692 173012 148756 173016
rect 55588 172936 55652 172940
rect 55588 172880 55602 172936
rect 55602 172880 55652 172936
rect 55588 172876 55652 172880
rect 169300 172876 169364 172940
rect 55404 172740 55468 172804
rect 168748 172740 168812 172804
rect 351644 172876 351708 172940
rect 351828 172876 351892 172940
rect 52644 171652 52708 171716
rect 54668 171652 54732 171716
rect 74356 171712 74420 171716
rect 74356 171656 74406 171712
rect 74406 171656 74420 171712
rect 74356 171652 74420 171656
rect 75644 169748 75708 169812
rect 73988 169612 74052 169676
rect 75460 169612 75524 169676
rect 73436 169536 73500 169540
rect 73436 169480 73486 169536
rect 73486 169480 73500 169536
rect 73436 169476 73500 169480
rect 76012 169476 76076 169540
rect 237380 169476 237444 169540
rect 243452 169476 243516 169540
rect 73804 169204 73868 169268
rect 74724 169204 74788 169268
rect 144092 169204 144156 169268
rect 148692 169204 148756 169268
rect 238116 169204 238180 169268
rect 242348 169204 242412 169268
rect 242532 169204 242596 169268
rect 247132 169204 247196 169268
rect 49148 162268 49212 162332
rect 49148 158324 49212 158388
rect 49148 155332 49212 155396
rect 49148 152884 49212 152948
rect 49148 148940 49212 149004
rect 49148 146084 49212 146148
rect 98828 145192 98892 145196
rect 98828 145136 98878 145192
rect 98878 145136 98892 145192
rect 98828 145132 98892 145136
rect 197636 144588 197700 144652
rect 292580 144588 292644 144652
rect 95148 144512 95212 144516
rect 95148 144456 95198 144512
rect 95198 144456 95212 144512
rect 95148 144452 95212 144456
rect 187884 144452 187948 144516
rect 282460 143772 282524 143836
rect 283748 143772 283812 143836
rect 302332 143772 302396 143836
rect 203156 143228 203220 143292
rect 231676 143228 231740 143292
rect 109684 143152 109748 143156
rect 109684 143096 109734 143152
rect 109734 143096 109748 143152
rect 109684 143092 109748 143096
rect 231124 143092 231188 143156
rect 297732 143152 297796 143156
rect 297732 143096 297782 143152
rect 297782 143096 297796 143152
rect 297732 143092 297796 143096
rect 106004 142548 106068 142612
rect 73988 142412 74052 142476
rect 74908 142412 74972 142476
rect 147036 142412 147100 142476
rect 150348 142412 150412 142476
rect 74172 142276 74236 142340
rect 77116 142276 77180 142340
rect 144092 142140 144156 142204
rect 167828 142200 167892 142204
rect 167828 142144 167842 142200
rect 167842 142144 167892 142200
rect 167828 142140 167892 142144
rect 76380 142004 76444 142068
rect 77668 142004 77732 142068
rect 147772 142004 147836 142068
rect 148324 142004 148388 142068
rect 219716 142064 219780 142068
rect 242900 142412 242964 142476
rect 247316 142412 247380 142476
rect 249892 142412 249956 142476
rect 250444 142412 250508 142476
rect 255228 142412 255292 142476
rect 290004 142412 290068 142476
rect 242532 142200 242596 142204
rect 242532 142144 242546 142200
rect 242546 142144 242596 142200
rect 242532 142140 242596 142144
rect 219716 142008 219730 142064
rect 219730 142008 219780 142064
rect 219716 142004 219780 142008
rect 246396 142004 246460 142068
rect 106004 141868 106068 141932
rect 74356 141792 74420 141796
rect 74356 141736 74370 141792
rect 74370 141736 74420 141792
rect 74356 141732 74420 141736
rect 75644 141596 75708 141660
rect 76012 141460 76076 141524
rect 73804 141324 73868 141388
rect 74724 141324 74788 141388
rect 74540 141188 74604 141252
rect 76380 141188 76444 141252
rect 137468 141052 137532 141116
rect 146484 141052 146548 141116
rect 149060 141112 149124 141116
rect 149060 141056 149110 141112
rect 149110 141056 149124 141112
rect 149060 141052 149124 141056
rect 152004 141112 152068 141116
rect 152004 141056 152054 141112
rect 152054 141056 152068 141112
rect 152004 141052 152068 141056
rect 207572 141052 207636 141116
rect 301964 141112 302028 141116
rect 301964 141056 302014 141112
rect 302014 141056 302028 141112
rect 301964 141052 302028 141056
rect 197268 140508 197332 140572
rect 137652 140432 137716 140436
rect 137652 140376 137666 140432
rect 137666 140376 137716 140432
rect 137652 140372 137716 140376
rect 231676 139964 231740 140028
rect 141516 139828 141580 139892
rect 148508 139828 148572 139892
rect 251364 139828 251428 139892
rect 238116 139692 238180 139756
rect 52644 139556 52708 139620
rect 54668 139556 54732 139620
rect 73804 139556 73868 139620
rect 74540 139556 74604 139620
rect 245292 139616 245356 139620
rect 245292 139560 245342 139616
rect 245342 139560 245356 139616
rect 245292 139556 245356 139560
rect 262956 139556 263020 139620
rect 351644 139556 351708 139620
rect 351828 139556 351892 139620
rect 73988 138876 74052 138940
rect 74724 138876 74788 138940
rect 249156 137304 249220 137308
rect 249156 137248 249170 137304
rect 249170 137248 249220 137304
rect 249156 137244 249220 137248
rect 137100 134388 137164 134452
rect 249708 133088 249772 133092
rect 249708 133032 249722 133088
rect 249722 133032 249772 133088
rect 249708 133028 249772 133032
rect 55404 132348 55468 132412
rect 197636 132484 197700 132548
rect 198556 132484 198620 132548
rect 54116 131532 54180 131596
rect 246212 130172 246276 130236
rect 55404 127180 55468 127244
rect 248604 126772 248668 126836
rect 249708 126772 249772 126836
rect 322756 124052 322820 124116
rect 54116 122692 54180 122756
rect 242716 122556 242780 122620
rect 258724 122556 258788 122620
rect 272708 122556 272772 122620
rect 148692 122284 148756 122348
rect 148876 122148 148940 122212
rect 177580 117796 177644 117860
rect 178684 117796 178748 117860
rect 54668 117116 54732 117180
rect 136916 116572 136980 116636
rect 138204 116572 138268 116636
rect 145012 116572 145076 116636
rect 228732 116436 228796 116500
rect 177580 114940 177644 115004
rect 147772 113580 147836 113644
rect 52644 113036 52708 113100
rect 230756 112900 230820 112964
rect 73436 112764 73500 112828
rect 147772 112492 147836 112556
rect 78036 110860 78100 110924
rect 134708 109772 134772 109836
rect 240140 109832 240204 109836
rect 240140 109776 240154 109832
rect 240154 109776 240204 109832
rect 240140 109772 240204 109776
rect 322756 109772 322820 109836
rect 84660 109636 84724 109700
rect 74540 109500 74604 109564
rect 148692 108820 148756 108884
rect 148876 108820 148940 108884
rect 230940 107384 231004 107388
rect 230940 107328 230954 107384
rect 230954 107328 231004 107384
rect 136916 107052 136980 107116
rect 230940 107324 231004 107328
rect 228732 106780 228796 106844
rect 177764 105420 177828 105484
rect 242164 105420 242228 105484
rect 242532 105420 242596 105484
rect 352748 105208 352812 105212
rect 352748 105152 352798 105208
rect 352798 105152 352812 105208
rect 352748 105148 352812 105152
rect 74172 102020 74236 102084
rect 136916 100932 136980 100996
rect 228732 100796 228796 100860
rect 164884 100660 164948 100724
rect 178132 100660 178196 100724
rect 258908 100660 258972 100724
rect 272708 100660 272772 100724
rect 323124 100932 323188 100996
rect 322756 100388 322820 100452
rect 176108 100252 176172 100316
rect 177028 100252 177092 100316
rect 263140 100252 263204 100316
rect 264428 100252 264492 100316
rect 73620 98212 73684 98276
rect 352748 97592 352812 97596
rect 352748 97536 352798 97592
rect 352798 97536 352812 97592
rect 352748 97532 352812 97536
rect 148692 95492 148756 95556
rect 148876 95492 148940 95556
rect 242532 95356 242596 95420
rect 148508 95220 148572 95284
rect 164884 95220 164948 95284
rect 178684 95220 178748 95284
rect 258724 95220 258788 95284
rect 272708 95220 272772 95284
rect 229100 94812 229164 94876
rect 322756 94404 322820 94468
rect 152188 90052 152252 90116
rect 155316 90052 155380 90116
rect 246212 90052 246276 90116
rect 249156 90052 249220 90116
rect 351644 90052 351708 90116
rect 155316 89160 155380 89164
rect 155316 89104 155366 89160
rect 155366 89104 155380 89160
rect 155316 89100 155380 89104
rect 245844 89100 245908 89164
rect 249156 88828 249220 88892
rect 249156 88480 249220 88484
rect 249156 88424 249170 88480
rect 249170 88424 249220 88480
rect 249156 88420 249220 88424
rect 72516 88344 72580 88348
rect 72516 88288 72566 88344
rect 72566 88288 72580 88344
rect 72516 88284 72580 88288
rect 252100 88072 252164 88076
rect 252100 88016 252150 88072
rect 252150 88016 252164 88072
rect 252100 88012 252164 88016
rect 261668 87468 261732 87532
rect 163780 87332 163844 87396
rect 167644 87332 167708 87396
rect 356796 87332 356860 87396
rect 148508 87060 148572 87124
rect 168748 87060 168812 87124
rect 169300 86924 169364 86988
rect 262772 86924 262836 86988
rect 168012 86788 168076 86852
rect 263508 86788 263572 86852
rect 169116 86652 169180 86716
rect 263140 86652 263204 86716
rect 73988 86380 74052 86444
rect 73252 86244 73316 86308
rect 72700 86108 72764 86172
rect 74356 86108 74420 86172
rect 252652 86108 252716 86172
rect 242532 85972 242596 86036
rect 72700 85836 72764 85900
rect 182548 83720 182612 83724
rect 182548 83664 182562 83720
rect 182562 83664 182612 83720
rect 182548 83660 182612 83664
rect 52644 79036 52708 79100
rect 54668 79036 54732 79100
rect 55404 79036 55468 79100
rect 54116 78900 54180 78964
rect 351644 77812 351708 77876
rect 351828 77812 351892 77876
rect 73068 76452 73132 76516
rect 242716 76452 242780 76516
rect 73068 76316 73132 76380
rect 73068 76044 73132 76108
rect 73252 75364 73316 75428
rect 73804 75364 73868 75428
rect 155316 75560 155380 75564
rect 155316 75504 155366 75560
rect 155366 75504 155380 75560
rect 155316 75500 155380 75504
rect 249156 75560 249220 75564
rect 249156 75504 249206 75560
rect 249206 75504 249220 75560
rect 249156 75500 249220 75504
rect 252652 75364 252716 75428
rect 261852 75364 261916 75428
rect 307116 53332 307180 53396
rect 118148 53120 118212 53124
rect 118148 53064 118198 53120
rect 118198 53064 118212 53120
rect 118148 53060 118212 53064
rect 211988 53120 212052 53124
rect 211988 53064 212038 53120
rect 212038 53064 212052 53120
rect 211988 53060 212052 53064
rect 78956 52788 79020 52852
rect 173900 52380 173964 52444
rect 266636 52380 266700 52444
rect 134156 51700 134220 51764
rect 227996 51700 228060 51764
rect 321836 51700 321900 51764
rect 102508 51292 102572 51356
rect 142804 51080 142868 51084
rect 142804 51024 142854 51080
rect 142854 51024 142868 51080
rect 142804 51020 142868 51024
rect 93676 50672 93740 50676
rect 93676 50616 93690 50672
rect 93690 50616 93740 50672
rect 93676 50612 93740 50616
rect 187332 50672 187396 50676
rect 187332 50616 187346 50672
rect 187346 50616 187396 50672
rect 187332 50612 187396 50616
rect 280436 50612 280500 50676
rect 191380 50340 191444 50404
rect 107476 50264 107540 50268
rect 107476 50208 107526 50264
rect 107526 50208 107540 50264
rect 107476 50204 107540 50208
rect 109316 50204 109380 50268
rect 199660 50204 199724 50268
rect 274916 49992 274980 49996
rect 274916 49936 274966 49992
rect 274966 49936 274980 49992
rect 274916 49932 274980 49936
rect 330852 49932 330916 49996
rect 87236 49252 87300 49316
rect 105268 49252 105332 49316
rect 181812 49312 181876 49316
rect 181812 49256 181862 49312
rect 181862 49256 181876 49312
rect 181812 49252 181876 49256
rect 204260 49252 204324 49316
rect 274916 49252 274980 49316
rect 73252 48028 73316 48092
rect 75092 48028 75156 48092
rect 87236 48028 87300 48092
rect 147956 48028 148020 48092
rect 154764 48028 154828 48092
rect 168012 48028 168076 48092
rect 72516 47892 72580 47956
rect 75276 47892 75340 47956
rect 144828 47892 144892 47956
rect 147772 47892 147836 47956
rect 160100 47952 160164 47956
rect 160100 47896 160114 47952
rect 160114 47896 160164 47952
rect 160100 47892 160164 47896
rect 168748 47892 168812 47956
rect 182180 47952 182244 47956
rect 182180 47896 182230 47952
rect 182230 47896 182244 47952
rect 182180 47892 182244 47896
rect 169668 47756 169732 47820
rect 237564 48028 237628 48092
rect 262404 48028 262468 48092
rect 263876 48028 263940 48092
rect 248604 47892 248668 47956
rect 253940 47952 254004 47956
rect 253940 47896 253990 47952
rect 253990 47896 254004 47952
rect 253940 47892 254004 47896
rect 274916 47892 274980 47956
rect 74172 47484 74236 47548
rect 75460 47484 75524 47548
rect 113548 47544 113612 47548
rect 113548 47488 113598 47544
rect 113598 47488 113612 47544
rect 113548 47484 113612 47488
rect 72516 47408 72580 47412
rect 72516 47352 72566 47408
rect 72566 47352 72580 47408
rect 72516 47348 72580 47352
rect 74172 47348 74236 47412
rect 107476 47348 107540 47412
rect 263876 47348 263940 47412
rect 264428 47348 264492 47412
rect 109316 47212 109380 47276
rect 110420 47212 110484 47276
rect 162860 47212 162924 47276
rect 248604 47212 248668 47276
rect 181076 46532 181140 46596
rect 260380 46592 260444 46596
rect 260380 46536 260394 46592
rect 260394 46536 260444 46592
rect 260380 46532 260444 46536
rect 275836 46592 275900 46596
rect 275836 46536 275886 46592
rect 275886 46536 275900 46592
rect 275836 46532 275900 46536
rect 158996 45988 159060 46052
rect 252652 45988 252716 46052
rect 263508 45988 263572 46052
rect 356796 45988 356860 46052
rect 73252 45852 73316 45916
rect 157524 45852 157588 45916
rect 147956 45716 148020 45780
rect 263324 45716 263388 45780
rect 331404 45308 331468 45372
rect 169668 44824 169732 44828
rect 169668 44768 169718 44824
rect 169718 44768 169732 44824
rect 169668 44764 169732 44768
rect 118148 44628 118212 44692
rect 211988 43404 212052 43468
rect 207756 39052 207820 39116
rect 301596 39112 301660 39116
rect 301596 39056 301610 39112
rect 301610 39056 301660 39112
rect 301596 39052 301660 39056
rect 307116 37692 307180 37756
<< metal4 >>
rect 0 405398 4000 405520
rect 0 405162 122 405398
rect 358 405162 442 405398
rect 678 405162 762 405398
rect 998 405162 1082 405398
rect 1318 405162 1402 405398
rect 1638 405162 1722 405398
rect 1958 405162 2042 405398
rect 2278 405162 2362 405398
rect 2598 405162 2682 405398
rect 2918 405162 3002 405398
rect 3238 405162 3322 405398
rect 3558 405162 3642 405398
rect 3878 405162 4000 405398
rect 0 405078 4000 405162
rect 0 404842 122 405078
rect 358 404842 442 405078
rect 678 404842 762 405078
rect 998 404842 1082 405078
rect 1318 404842 1402 405078
rect 1638 404842 1722 405078
rect 1958 404842 2042 405078
rect 2278 404842 2362 405078
rect 2598 404842 2682 405078
rect 2918 404842 3002 405078
rect 3238 404842 3322 405078
rect 3558 404842 3642 405078
rect 3878 404842 4000 405078
rect 0 404758 4000 404842
rect 0 404522 122 404758
rect 358 404522 442 404758
rect 678 404522 762 404758
rect 998 404522 1082 404758
rect 1318 404522 1402 404758
rect 1638 404522 1722 404758
rect 1958 404522 2042 404758
rect 2278 404522 2362 404758
rect 2598 404522 2682 404758
rect 2918 404522 3002 404758
rect 3238 404522 3322 404758
rect 3558 404522 3642 404758
rect 3878 404522 4000 404758
rect 0 404438 4000 404522
rect 0 404202 122 404438
rect 358 404202 442 404438
rect 678 404202 762 404438
rect 998 404202 1082 404438
rect 1318 404202 1402 404438
rect 1638 404202 1722 404438
rect 1958 404202 2042 404438
rect 2278 404202 2362 404438
rect 2598 404202 2682 404438
rect 2918 404202 3002 404438
rect 3238 404202 3322 404438
rect 3558 404202 3642 404438
rect 3878 404202 4000 404438
rect 0 404118 4000 404202
rect 0 403882 122 404118
rect 358 403882 442 404118
rect 678 403882 762 404118
rect 998 403882 1082 404118
rect 1318 403882 1402 404118
rect 1638 403882 1722 404118
rect 1958 403882 2042 404118
rect 2278 403882 2362 404118
rect 2598 403882 2682 404118
rect 2918 403882 3002 404118
rect 3238 403882 3322 404118
rect 3558 403882 3642 404118
rect 3878 403882 4000 404118
rect 0 403798 4000 403882
rect 0 403562 122 403798
rect 358 403562 442 403798
rect 678 403562 762 403798
rect 998 403562 1082 403798
rect 1318 403562 1402 403798
rect 1638 403562 1722 403798
rect 1958 403562 2042 403798
rect 2278 403562 2362 403798
rect 2598 403562 2682 403798
rect 2918 403562 3002 403798
rect 3238 403562 3322 403798
rect 3558 403562 3642 403798
rect 3878 403562 4000 403798
rect 0 403478 4000 403562
rect 0 403242 122 403478
rect 358 403242 442 403478
rect 678 403242 762 403478
rect 998 403242 1082 403478
rect 1318 403242 1402 403478
rect 1638 403242 1722 403478
rect 1958 403242 2042 403478
rect 2278 403242 2362 403478
rect 2598 403242 2682 403478
rect 2918 403242 3002 403478
rect 3238 403242 3322 403478
rect 3558 403242 3642 403478
rect 3878 403242 4000 403478
rect 0 403158 4000 403242
rect 0 402922 122 403158
rect 358 402922 442 403158
rect 678 402922 762 403158
rect 998 402922 1082 403158
rect 1318 402922 1402 403158
rect 1638 402922 1722 403158
rect 1958 402922 2042 403158
rect 2278 402922 2362 403158
rect 2598 402922 2682 403158
rect 2918 402922 3002 403158
rect 3238 402922 3322 403158
rect 3558 402922 3642 403158
rect 3878 402922 4000 403158
rect 0 402838 4000 402922
rect 0 402602 122 402838
rect 358 402602 442 402838
rect 678 402602 762 402838
rect 998 402602 1082 402838
rect 1318 402602 1402 402838
rect 1638 402602 1722 402838
rect 1958 402602 2042 402838
rect 2278 402602 2362 402838
rect 2598 402602 2682 402838
rect 2918 402602 3002 402838
rect 3238 402602 3322 402838
rect 3558 402602 3642 402838
rect 3878 402602 4000 402838
rect 0 402518 4000 402602
rect 0 402282 122 402518
rect 358 402282 442 402518
rect 678 402282 762 402518
rect 998 402282 1082 402518
rect 1318 402282 1402 402518
rect 1638 402282 1722 402518
rect 1958 402282 2042 402518
rect 2278 402282 2362 402518
rect 2598 402282 2682 402518
rect 2918 402282 3002 402518
rect 3238 402282 3322 402518
rect 3558 402282 3642 402518
rect 3878 402282 4000 402518
rect 0 402198 4000 402282
rect 0 401962 122 402198
rect 358 401962 442 402198
rect 678 401962 762 402198
rect 998 401962 1082 402198
rect 1318 401962 1402 402198
rect 1638 401962 1722 402198
rect 1958 401962 2042 402198
rect 2278 401962 2362 402198
rect 2598 401962 2682 402198
rect 2918 401962 3002 402198
rect 3238 401962 3322 402198
rect 3558 401962 3642 402198
rect 3878 401962 4000 402198
rect 0 401878 4000 401962
rect 0 401642 122 401878
rect 358 401642 442 401878
rect 678 401642 762 401878
rect 998 401642 1082 401878
rect 1318 401642 1402 401878
rect 1638 401642 1722 401878
rect 1958 401642 2042 401878
rect 2278 401642 2362 401878
rect 2598 401642 2682 401878
rect 2918 401642 3002 401878
rect 3238 401642 3322 401878
rect 3558 401642 3642 401878
rect 3878 401642 4000 401878
rect 0 366762 4000 401642
rect 440740 405398 444740 405520
rect 440740 405162 440862 405398
rect 441098 405162 441182 405398
rect 441418 405162 441502 405398
rect 441738 405162 441822 405398
rect 442058 405162 442142 405398
rect 442378 405162 442462 405398
rect 442698 405162 442782 405398
rect 443018 405162 443102 405398
rect 443338 405162 443422 405398
rect 443658 405162 443742 405398
rect 443978 405162 444062 405398
rect 444298 405162 444382 405398
rect 444618 405162 444740 405398
rect 440740 405078 444740 405162
rect 440740 404842 440862 405078
rect 441098 404842 441182 405078
rect 441418 404842 441502 405078
rect 441738 404842 441822 405078
rect 442058 404842 442142 405078
rect 442378 404842 442462 405078
rect 442698 404842 442782 405078
rect 443018 404842 443102 405078
rect 443338 404842 443422 405078
rect 443658 404842 443742 405078
rect 443978 404842 444062 405078
rect 444298 404842 444382 405078
rect 444618 404842 444740 405078
rect 440740 404758 444740 404842
rect 440740 404522 440862 404758
rect 441098 404522 441182 404758
rect 441418 404522 441502 404758
rect 441738 404522 441822 404758
rect 442058 404522 442142 404758
rect 442378 404522 442462 404758
rect 442698 404522 442782 404758
rect 443018 404522 443102 404758
rect 443338 404522 443422 404758
rect 443658 404522 443742 404758
rect 443978 404522 444062 404758
rect 444298 404522 444382 404758
rect 444618 404522 444740 404758
rect 440740 404438 444740 404522
rect 440740 404202 440862 404438
rect 441098 404202 441182 404438
rect 441418 404202 441502 404438
rect 441738 404202 441822 404438
rect 442058 404202 442142 404438
rect 442378 404202 442462 404438
rect 442698 404202 442782 404438
rect 443018 404202 443102 404438
rect 443338 404202 443422 404438
rect 443658 404202 443742 404438
rect 443978 404202 444062 404438
rect 444298 404202 444382 404438
rect 444618 404202 444740 404438
rect 440740 404118 444740 404202
rect 440740 403882 440862 404118
rect 441098 403882 441182 404118
rect 441418 403882 441502 404118
rect 441738 403882 441822 404118
rect 442058 403882 442142 404118
rect 442378 403882 442462 404118
rect 442698 403882 442782 404118
rect 443018 403882 443102 404118
rect 443338 403882 443422 404118
rect 443658 403882 443742 404118
rect 443978 403882 444062 404118
rect 444298 403882 444382 404118
rect 444618 403882 444740 404118
rect 440740 403798 444740 403882
rect 440740 403562 440862 403798
rect 441098 403562 441182 403798
rect 441418 403562 441502 403798
rect 441738 403562 441822 403798
rect 442058 403562 442142 403798
rect 442378 403562 442462 403798
rect 442698 403562 442782 403798
rect 443018 403562 443102 403798
rect 443338 403562 443422 403798
rect 443658 403562 443742 403798
rect 443978 403562 444062 403798
rect 444298 403562 444382 403798
rect 444618 403562 444740 403798
rect 440740 403478 444740 403562
rect 440740 403242 440862 403478
rect 441098 403242 441182 403478
rect 441418 403242 441502 403478
rect 441738 403242 441822 403478
rect 442058 403242 442142 403478
rect 442378 403242 442462 403478
rect 442698 403242 442782 403478
rect 443018 403242 443102 403478
rect 443338 403242 443422 403478
rect 443658 403242 443742 403478
rect 443978 403242 444062 403478
rect 444298 403242 444382 403478
rect 444618 403242 444740 403478
rect 440740 403158 444740 403242
rect 440740 402922 440862 403158
rect 441098 402922 441182 403158
rect 441418 402922 441502 403158
rect 441738 402922 441822 403158
rect 442058 402922 442142 403158
rect 442378 402922 442462 403158
rect 442698 402922 442782 403158
rect 443018 402922 443102 403158
rect 443338 402922 443422 403158
rect 443658 402922 443742 403158
rect 443978 402922 444062 403158
rect 444298 402922 444382 403158
rect 444618 402922 444740 403158
rect 440740 402838 444740 402922
rect 440740 402602 440862 402838
rect 441098 402602 441182 402838
rect 441418 402602 441502 402838
rect 441738 402602 441822 402838
rect 442058 402602 442142 402838
rect 442378 402602 442462 402838
rect 442698 402602 442782 402838
rect 443018 402602 443102 402838
rect 443338 402602 443422 402838
rect 443658 402602 443742 402838
rect 443978 402602 444062 402838
rect 444298 402602 444382 402838
rect 444618 402602 444740 402838
rect 440740 402518 444740 402602
rect 440740 402282 440862 402518
rect 441098 402282 441182 402518
rect 441418 402282 441502 402518
rect 441738 402282 441822 402518
rect 442058 402282 442142 402518
rect 442378 402282 442462 402518
rect 442698 402282 442782 402518
rect 443018 402282 443102 402518
rect 443338 402282 443422 402518
rect 443658 402282 443742 402518
rect 443978 402282 444062 402518
rect 444298 402282 444382 402518
rect 444618 402282 444740 402518
rect 440740 402198 444740 402282
rect 440740 401962 440862 402198
rect 441098 401962 441182 402198
rect 441418 401962 441502 402198
rect 441738 401962 441822 402198
rect 442058 401962 442142 402198
rect 442378 401962 442462 402198
rect 442698 401962 442782 402198
rect 443018 401962 443102 402198
rect 443338 401962 443422 402198
rect 443658 401962 443742 402198
rect 443978 401962 444062 402198
rect 444298 401962 444382 402198
rect 444618 401962 444740 402198
rect 440740 401878 444740 401962
rect 440740 401642 440862 401878
rect 441098 401642 441182 401878
rect 441418 401642 441502 401878
rect 441738 401642 441822 401878
rect 442058 401642 442142 401878
rect 442378 401642 442462 401878
rect 442698 401642 442782 401878
rect 443018 401642 443102 401878
rect 443338 401642 443422 401878
rect 443658 401642 443742 401878
rect 443978 401642 444062 401878
rect 444298 401642 444382 401878
rect 444618 401642 444740 401878
rect 0 366526 122 366762
rect 358 366526 442 366762
rect 678 366526 762 366762
rect 998 366526 1082 366762
rect 1318 366526 1402 366762
rect 1638 366526 1722 366762
rect 1958 366526 2042 366762
rect 2278 366526 2362 366762
rect 2598 366526 2682 366762
rect 2918 366526 3002 366762
rect 3238 366526 3322 366762
rect 3558 366526 3642 366762
rect 3878 366526 4000 366762
rect 0 336126 4000 366526
rect 0 335890 122 336126
rect 358 335890 442 336126
rect 678 335890 762 336126
rect 998 335890 1082 336126
rect 1318 335890 1402 336126
rect 1638 335890 1722 336126
rect 1958 335890 2042 336126
rect 2278 335890 2362 336126
rect 2598 335890 2682 336126
rect 2918 335890 3002 336126
rect 3238 335890 3322 336126
rect 3558 335890 3642 336126
rect 3878 335890 4000 336126
rect 0 305490 4000 335890
rect 0 305254 122 305490
rect 358 305254 442 305490
rect 678 305254 762 305490
rect 998 305254 1082 305490
rect 1318 305254 1402 305490
rect 1638 305254 1722 305490
rect 1958 305254 2042 305490
rect 2278 305254 2362 305490
rect 2598 305254 2682 305490
rect 2918 305254 3002 305490
rect 3238 305254 3322 305490
rect 3558 305254 3642 305490
rect 3878 305254 4000 305490
rect 0 274854 4000 305254
rect 0 274618 122 274854
rect 358 274618 442 274854
rect 678 274618 762 274854
rect 998 274618 1082 274854
rect 1318 274618 1402 274854
rect 1638 274618 1722 274854
rect 1958 274618 2042 274854
rect 2278 274618 2362 274854
rect 2598 274618 2682 274854
rect 2918 274618 3002 274854
rect 3238 274618 3322 274854
rect 3558 274618 3642 274854
rect 3878 274618 4000 274854
rect 0 244218 4000 274618
rect 0 243982 122 244218
rect 358 243982 442 244218
rect 678 243982 762 244218
rect 998 243982 1082 244218
rect 1318 243982 1402 244218
rect 1638 243982 1722 244218
rect 1958 243982 2042 244218
rect 2278 243982 2362 244218
rect 2598 243982 2682 244218
rect 2918 243982 3002 244218
rect 3238 243982 3322 244218
rect 3558 243982 3642 244218
rect 3878 243982 4000 244218
rect 0 213582 4000 243982
rect 0 213346 122 213582
rect 358 213346 442 213582
rect 678 213346 762 213582
rect 998 213346 1082 213582
rect 1318 213346 1402 213582
rect 1638 213346 1722 213582
rect 1958 213346 2042 213582
rect 2278 213346 2362 213582
rect 2598 213346 2682 213582
rect 2918 213346 3002 213582
rect 3238 213346 3322 213582
rect 3558 213346 3642 213582
rect 3878 213346 4000 213582
rect 0 182946 4000 213346
rect 0 182710 122 182946
rect 358 182710 442 182946
rect 678 182710 762 182946
rect 998 182710 1082 182946
rect 1318 182710 1402 182946
rect 1638 182710 1722 182946
rect 1958 182710 2042 182946
rect 2278 182710 2362 182946
rect 2598 182710 2682 182946
rect 2918 182710 3002 182946
rect 3238 182710 3322 182946
rect 3558 182710 3642 182946
rect 3878 182710 4000 182946
rect 0 152310 4000 182710
rect 0 152074 122 152310
rect 358 152074 442 152310
rect 678 152074 762 152310
rect 998 152074 1082 152310
rect 1318 152074 1402 152310
rect 1638 152074 1722 152310
rect 1958 152074 2042 152310
rect 2278 152074 2362 152310
rect 2598 152074 2682 152310
rect 2918 152074 3002 152310
rect 3238 152074 3322 152310
rect 3558 152074 3642 152310
rect 3878 152074 4000 152310
rect 0 121674 4000 152074
rect 0 121438 122 121674
rect 358 121438 442 121674
rect 678 121438 762 121674
rect 998 121438 1082 121674
rect 1318 121438 1402 121674
rect 1638 121438 1722 121674
rect 1958 121438 2042 121674
rect 2278 121438 2362 121674
rect 2598 121438 2682 121674
rect 2918 121438 3002 121674
rect 3238 121438 3322 121674
rect 3558 121438 3642 121674
rect 3878 121438 4000 121674
rect 0 91038 4000 121438
rect 0 90802 122 91038
rect 358 90802 442 91038
rect 678 90802 762 91038
rect 998 90802 1082 91038
rect 1318 90802 1402 91038
rect 1638 90802 1722 91038
rect 1958 90802 2042 91038
rect 2278 90802 2362 91038
rect 2598 90802 2682 91038
rect 2918 90802 3002 91038
rect 3238 90802 3322 91038
rect 3558 90802 3642 91038
rect 3878 90802 4000 91038
rect 0 60402 4000 90802
rect 0 60166 122 60402
rect 358 60166 442 60402
rect 678 60166 762 60402
rect 998 60166 1082 60402
rect 1318 60166 1402 60402
rect 1638 60166 1722 60402
rect 1958 60166 2042 60402
rect 2278 60166 2362 60402
rect 2598 60166 2682 60402
rect 2918 60166 3002 60402
rect 3238 60166 3322 60402
rect 3558 60166 3642 60402
rect 3878 60166 4000 60402
rect 0 29766 4000 60166
rect 0 29530 122 29766
rect 358 29530 442 29766
rect 678 29530 762 29766
rect 998 29530 1082 29766
rect 1318 29530 1402 29766
rect 1638 29530 1722 29766
rect 1958 29530 2042 29766
rect 2278 29530 2362 29766
rect 2598 29530 2682 29766
rect 2918 29530 3002 29766
rect 3238 29530 3322 29766
rect 3558 29530 3642 29766
rect 3878 29530 4000 29766
rect 0 3878 4000 29530
rect 5000 400398 9000 400520
rect 5000 400162 5122 400398
rect 5358 400162 5442 400398
rect 5678 400162 5762 400398
rect 5998 400162 6082 400398
rect 6318 400162 6402 400398
rect 6638 400162 6722 400398
rect 6958 400162 7042 400398
rect 7278 400162 7362 400398
rect 7598 400162 7682 400398
rect 7918 400162 8002 400398
rect 8238 400162 8322 400398
rect 8558 400162 8642 400398
rect 8878 400162 9000 400398
rect 5000 400078 9000 400162
rect 5000 399842 5122 400078
rect 5358 399842 5442 400078
rect 5678 399842 5762 400078
rect 5998 399842 6082 400078
rect 6318 399842 6402 400078
rect 6638 399842 6722 400078
rect 6958 399842 7042 400078
rect 7278 399842 7362 400078
rect 7598 399842 7682 400078
rect 7918 399842 8002 400078
rect 8238 399842 8322 400078
rect 8558 399842 8642 400078
rect 8878 399842 9000 400078
rect 5000 399758 9000 399842
rect 5000 399522 5122 399758
rect 5358 399522 5442 399758
rect 5678 399522 5762 399758
rect 5998 399522 6082 399758
rect 6318 399522 6402 399758
rect 6638 399522 6722 399758
rect 6958 399522 7042 399758
rect 7278 399522 7362 399758
rect 7598 399522 7682 399758
rect 7918 399522 8002 399758
rect 8238 399522 8322 399758
rect 8558 399522 8642 399758
rect 8878 399522 9000 399758
rect 5000 399438 9000 399522
rect 5000 399202 5122 399438
rect 5358 399202 5442 399438
rect 5678 399202 5762 399438
rect 5998 399202 6082 399438
rect 6318 399202 6402 399438
rect 6638 399202 6722 399438
rect 6958 399202 7042 399438
rect 7278 399202 7362 399438
rect 7598 399202 7682 399438
rect 7918 399202 8002 399438
rect 8238 399202 8322 399438
rect 8558 399202 8642 399438
rect 8878 399202 9000 399438
rect 5000 399118 9000 399202
rect 5000 398882 5122 399118
rect 5358 398882 5442 399118
rect 5678 398882 5762 399118
rect 5998 398882 6082 399118
rect 6318 398882 6402 399118
rect 6638 398882 6722 399118
rect 6958 398882 7042 399118
rect 7278 398882 7362 399118
rect 7598 398882 7682 399118
rect 7918 398882 8002 399118
rect 8238 398882 8322 399118
rect 8558 398882 8642 399118
rect 8878 398882 9000 399118
rect 5000 398798 9000 398882
rect 5000 398562 5122 398798
rect 5358 398562 5442 398798
rect 5678 398562 5762 398798
rect 5998 398562 6082 398798
rect 6318 398562 6402 398798
rect 6638 398562 6722 398798
rect 6958 398562 7042 398798
rect 7278 398562 7362 398798
rect 7598 398562 7682 398798
rect 7918 398562 8002 398798
rect 8238 398562 8322 398798
rect 8558 398562 8642 398798
rect 8878 398562 9000 398798
rect 5000 398478 9000 398562
rect 5000 398242 5122 398478
rect 5358 398242 5442 398478
rect 5678 398242 5762 398478
rect 5998 398242 6082 398478
rect 6318 398242 6402 398478
rect 6638 398242 6722 398478
rect 6958 398242 7042 398478
rect 7278 398242 7362 398478
rect 7598 398242 7682 398478
rect 7918 398242 8002 398478
rect 8238 398242 8322 398478
rect 8558 398242 8642 398478
rect 8878 398242 9000 398478
rect 5000 398158 9000 398242
rect 5000 397922 5122 398158
rect 5358 397922 5442 398158
rect 5678 397922 5762 398158
rect 5998 397922 6082 398158
rect 6318 397922 6402 398158
rect 6638 397922 6722 398158
rect 6958 397922 7042 398158
rect 7278 397922 7362 398158
rect 7598 397922 7682 398158
rect 7918 397922 8002 398158
rect 8238 397922 8322 398158
rect 8558 397922 8642 398158
rect 8878 397922 9000 398158
rect 5000 397838 9000 397922
rect 5000 397602 5122 397838
rect 5358 397602 5442 397838
rect 5678 397602 5762 397838
rect 5998 397602 6082 397838
rect 6318 397602 6402 397838
rect 6638 397602 6722 397838
rect 6958 397602 7042 397838
rect 7278 397602 7362 397838
rect 7598 397602 7682 397838
rect 7918 397602 8002 397838
rect 8238 397602 8322 397838
rect 8558 397602 8642 397838
rect 8878 397602 9000 397838
rect 5000 397518 9000 397602
rect 5000 397282 5122 397518
rect 5358 397282 5442 397518
rect 5678 397282 5762 397518
rect 5998 397282 6082 397518
rect 6318 397282 6402 397518
rect 6638 397282 6722 397518
rect 6958 397282 7042 397518
rect 7278 397282 7362 397518
rect 7598 397282 7682 397518
rect 7918 397282 8002 397518
rect 8238 397282 8322 397518
rect 8558 397282 8642 397518
rect 8878 397282 9000 397518
rect 5000 397198 9000 397282
rect 5000 396962 5122 397198
rect 5358 396962 5442 397198
rect 5678 396962 5762 397198
rect 5998 396962 6082 397198
rect 6318 396962 6402 397198
rect 6638 396962 6722 397198
rect 6958 396962 7042 397198
rect 7278 396962 7362 397198
rect 7598 396962 7682 397198
rect 7918 396962 8002 397198
rect 8238 396962 8322 397198
rect 8558 396962 8642 397198
rect 8878 396962 9000 397198
rect 5000 396878 9000 396962
rect 5000 396642 5122 396878
rect 5358 396642 5442 396878
rect 5678 396642 5762 396878
rect 5998 396642 6082 396878
rect 6318 396642 6402 396878
rect 6638 396642 6722 396878
rect 6958 396642 7042 396878
rect 7278 396642 7362 396878
rect 7598 396642 7682 396878
rect 7918 396642 8002 396878
rect 8238 396642 8322 396878
rect 8558 396642 8642 396878
rect 8878 396642 9000 396878
rect 5000 382080 9000 396642
rect 435740 400398 439740 400520
rect 435740 400162 435862 400398
rect 436098 400162 436182 400398
rect 436418 400162 436502 400398
rect 436738 400162 436822 400398
rect 437058 400162 437142 400398
rect 437378 400162 437462 400398
rect 437698 400162 437782 400398
rect 438018 400162 438102 400398
rect 438338 400162 438422 400398
rect 438658 400162 438742 400398
rect 438978 400162 439062 400398
rect 439298 400162 439382 400398
rect 439618 400162 439740 400398
rect 435740 400078 439740 400162
rect 435740 399842 435862 400078
rect 436098 399842 436182 400078
rect 436418 399842 436502 400078
rect 436738 399842 436822 400078
rect 437058 399842 437142 400078
rect 437378 399842 437462 400078
rect 437698 399842 437782 400078
rect 438018 399842 438102 400078
rect 438338 399842 438422 400078
rect 438658 399842 438742 400078
rect 438978 399842 439062 400078
rect 439298 399842 439382 400078
rect 439618 399842 439740 400078
rect 435740 399758 439740 399842
rect 435740 399522 435862 399758
rect 436098 399522 436182 399758
rect 436418 399522 436502 399758
rect 436738 399522 436822 399758
rect 437058 399522 437142 399758
rect 437378 399522 437462 399758
rect 437698 399522 437782 399758
rect 438018 399522 438102 399758
rect 438338 399522 438422 399758
rect 438658 399522 438742 399758
rect 438978 399522 439062 399758
rect 439298 399522 439382 399758
rect 439618 399522 439740 399758
rect 435740 399438 439740 399522
rect 435740 399202 435862 399438
rect 436098 399202 436182 399438
rect 436418 399202 436502 399438
rect 436738 399202 436822 399438
rect 437058 399202 437142 399438
rect 437378 399202 437462 399438
rect 437698 399202 437782 399438
rect 438018 399202 438102 399438
rect 438338 399202 438422 399438
rect 438658 399202 438742 399438
rect 438978 399202 439062 399438
rect 439298 399202 439382 399438
rect 439618 399202 439740 399438
rect 435740 399118 439740 399202
rect 435740 398882 435862 399118
rect 436098 398882 436182 399118
rect 436418 398882 436502 399118
rect 436738 398882 436822 399118
rect 437058 398882 437142 399118
rect 437378 398882 437462 399118
rect 437698 398882 437782 399118
rect 438018 398882 438102 399118
rect 438338 398882 438422 399118
rect 438658 398882 438742 399118
rect 438978 398882 439062 399118
rect 439298 398882 439382 399118
rect 439618 398882 439740 399118
rect 435740 398798 439740 398882
rect 435740 398562 435862 398798
rect 436098 398562 436182 398798
rect 436418 398562 436502 398798
rect 436738 398562 436822 398798
rect 437058 398562 437142 398798
rect 437378 398562 437462 398798
rect 437698 398562 437782 398798
rect 438018 398562 438102 398798
rect 438338 398562 438422 398798
rect 438658 398562 438742 398798
rect 438978 398562 439062 398798
rect 439298 398562 439382 398798
rect 439618 398562 439740 398798
rect 435740 398478 439740 398562
rect 435740 398242 435862 398478
rect 436098 398242 436182 398478
rect 436418 398242 436502 398478
rect 436738 398242 436822 398478
rect 437058 398242 437142 398478
rect 437378 398242 437462 398478
rect 437698 398242 437782 398478
rect 438018 398242 438102 398478
rect 438338 398242 438422 398478
rect 438658 398242 438742 398478
rect 438978 398242 439062 398478
rect 439298 398242 439382 398478
rect 439618 398242 439740 398478
rect 435740 398158 439740 398242
rect 435740 397922 435862 398158
rect 436098 397922 436182 398158
rect 436418 397922 436502 398158
rect 436738 397922 436822 398158
rect 437058 397922 437142 398158
rect 437378 397922 437462 398158
rect 437698 397922 437782 398158
rect 438018 397922 438102 398158
rect 438338 397922 438422 398158
rect 438658 397922 438742 398158
rect 438978 397922 439062 398158
rect 439298 397922 439382 398158
rect 439618 397922 439740 398158
rect 435740 397838 439740 397922
rect 435740 397602 435862 397838
rect 436098 397602 436182 397838
rect 436418 397602 436502 397838
rect 436738 397602 436822 397838
rect 437058 397602 437142 397838
rect 437378 397602 437462 397838
rect 437698 397602 437782 397838
rect 438018 397602 438102 397838
rect 438338 397602 438422 397838
rect 438658 397602 438742 397838
rect 438978 397602 439062 397838
rect 439298 397602 439382 397838
rect 439618 397602 439740 397838
rect 435740 397518 439740 397602
rect 435740 397282 435862 397518
rect 436098 397282 436182 397518
rect 436418 397282 436502 397518
rect 436738 397282 436822 397518
rect 437058 397282 437142 397518
rect 437378 397282 437462 397518
rect 437698 397282 437782 397518
rect 438018 397282 438102 397518
rect 438338 397282 438422 397518
rect 438658 397282 438742 397518
rect 438978 397282 439062 397518
rect 439298 397282 439382 397518
rect 439618 397282 439740 397518
rect 435740 397198 439740 397282
rect 435740 396962 435862 397198
rect 436098 396962 436182 397198
rect 436418 396962 436502 397198
rect 436738 396962 436822 397198
rect 437058 396962 437142 397198
rect 437378 396962 437462 397198
rect 437698 396962 437782 397198
rect 438018 396962 438102 397198
rect 438338 396962 438422 397198
rect 438658 396962 438742 397198
rect 438978 396962 439062 397198
rect 439298 396962 439382 397198
rect 439618 396962 439740 397198
rect 435740 396878 439740 396962
rect 435740 396642 435862 396878
rect 436098 396642 436182 396878
rect 436418 396642 436502 396878
rect 436738 396642 436822 396878
rect 437058 396642 437142 396878
rect 437378 396642 437462 396878
rect 437698 396642 437782 396878
rect 438018 396642 438102 396878
rect 438338 396642 438422 396878
rect 438658 396642 438742 396878
rect 438978 396642 439062 396878
rect 439298 396642 439382 396878
rect 439618 396642 439740 396878
rect 341707 393804 341773 393805
rect 341707 393740 341708 393804
rect 341772 393740 341773 393804
rect 341707 393739 341773 393740
rect 5000 381844 5122 382080
rect 5358 381844 5442 382080
rect 5678 381844 5762 382080
rect 5998 381844 6082 382080
rect 6318 381844 6402 382080
rect 6638 381844 6722 382080
rect 6958 381844 7042 382080
rect 7278 381844 7362 382080
rect 7598 381844 7682 382080
rect 7918 381844 8002 382080
rect 8238 381844 8322 382080
rect 8558 381844 8642 382080
rect 8878 381844 9000 382080
rect 5000 351444 9000 381844
rect 191195 359396 191261 359397
rect 191195 359332 191196 359396
rect 191260 359332 191261 359396
rect 191195 359331 191261 359332
rect 96803 355316 96869 355317
rect 96803 355252 96804 355316
rect 96868 355252 96869 355316
rect 96803 355251 96869 355252
rect 96806 351645 96866 355251
rect 191198 351917 191258 359331
rect 284483 356540 284549 356541
rect 284483 356476 284484 356540
rect 284548 356476 284549 356540
rect 284483 356475 284549 356476
rect 191195 351916 191261 351917
rect 191195 351852 191196 351916
rect 191260 351852 191261 351916
rect 191195 351851 191261 351852
rect 284486 351645 284546 356475
rect 341710 356082 341770 393739
rect 435740 382080 439740 396642
rect 435740 381844 435862 382080
rect 436098 381844 436182 382080
rect 436418 381844 436502 382080
rect 436738 381844 436822 382080
rect 437058 381844 437142 382080
rect 437378 381844 437462 382080
rect 437698 381844 437782 382080
rect 438018 381844 438102 382080
rect 438338 381844 438422 382080
rect 438658 381844 438742 382080
rect 438978 381844 439062 382080
rect 439298 381844 439382 382080
rect 439618 381844 439740 382080
rect 96803 351644 96869 351645
rect 96803 351580 96804 351644
rect 96868 351580 96869 351644
rect 96803 351579 96869 351580
rect 284483 351644 284549 351645
rect 284483 351580 284484 351644
rect 284548 351580 284549 351644
rect 284483 351579 284549 351580
rect 5000 351208 5122 351444
rect 5358 351208 5442 351444
rect 5678 351208 5762 351444
rect 5998 351208 6082 351444
rect 6318 351208 6402 351444
rect 6638 351208 6722 351444
rect 6958 351208 7042 351444
rect 7278 351208 7362 351444
rect 7598 351208 7682 351444
rect 7918 351208 8002 351444
rect 8238 351208 8322 351444
rect 8558 351208 8642 351444
rect 8878 351208 9000 351444
rect 5000 320808 9000 351208
rect 332142 349962 332202 355846
rect 435740 351444 439740 381844
rect 435740 351208 435862 351444
rect 436098 351208 436182 351444
rect 436418 351208 436502 351444
rect 436738 351208 436822 351444
rect 437058 351208 437142 351444
rect 437378 351208 437462 351444
rect 437698 351208 437782 351444
rect 438018 351208 438102 351444
rect 438338 351208 438422 351444
rect 438658 351208 438742 351444
rect 438978 351208 439062 351444
rect 439298 351208 439382 351444
rect 439618 351208 439740 351444
rect 341158 335002 341218 336806
rect 104899 333828 104965 333829
rect 104899 333764 104900 333828
rect 104964 333764 104965 333828
rect 104899 333763 104965 333764
rect 52643 326348 52709 326349
rect 52643 326284 52644 326348
rect 52708 326284 52709 326348
rect 52643 326283 52709 326284
rect 54667 326348 54733 326349
rect 54667 326284 54668 326348
rect 54732 326284 54733 326348
rect 54667 326283 54733 326284
rect 55035 326348 55101 326349
rect 55035 326284 55036 326348
rect 55100 326284 55101 326348
rect 55035 326283 55101 326284
rect 55955 326348 56021 326349
rect 55955 326284 55956 326348
rect 56020 326284 56021 326348
rect 55955 326283 56021 326284
rect 5000 320572 5122 320808
rect 5358 320572 5442 320808
rect 5678 320572 5762 320808
rect 5998 320572 6082 320808
rect 6318 320572 6402 320808
rect 6638 320572 6722 320808
rect 6958 320572 7042 320808
rect 7278 320572 7362 320808
rect 7598 320572 7682 320808
rect 7918 320572 8002 320808
rect 8238 320572 8322 320808
rect 8558 320572 8642 320808
rect 8878 320572 9000 320808
rect 5000 290172 9000 320572
rect 52646 300645 52706 326283
rect 54670 306221 54730 326283
rect 55038 311114 55098 326283
rect 55958 315877 56018 326283
rect 104902 319954 104962 333763
rect 212171 333556 212237 333557
rect 212171 333492 212172 333556
rect 212236 333492 212237 333556
rect 212171 333491 212237 333492
rect 204443 331652 204509 331653
rect 204443 331588 204444 331652
rect 204508 331588 204509 331652
rect 204443 331587 204509 331588
rect 158630 330157 158690 331366
rect 204446 330922 204506 331587
rect 159550 330157 159610 330686
rect 158627 330156 158693 330157
rect 158627 330092 158628 330156
rect 158692 330092 158693 330156
rect 158627 330091 158693 330092
rect 159547 330156 159613 330157
rect 159547 330092 159548 330156
rect 159612 330092 159613 330156
rect 159547 330091 159613 330092
rect 212174 329562 212234 333491
rect 295523 333148 295589 333149
rect 295523 333084 295524 333148
rect 295588 333084 295589 333148
rect 295523 333083 295589 333084
rect 295526 332282 295586 333083
rect 230939 331652 231005 331653
rect 230939 331588 230940 331652
rect 231004 331588 231005 331652
rect 230939 331587 231005 331588
rect 230942 328797 231002 331587
rect 299387 331516 299453 331517
rect 299387 331452 299388 331516
rect 299452 331452 299453 331516
rect 299387 331451 299453 331452
rect 251918 330157 251978 330686
rect 252654 330157 252714 331366
rect 251915 330156 251981 330157
rect 251915 330092 251916 330156
rect 251980 330092 251981 330156
rect 251915 330091 251981 330092
rect 252651 330156 252717 330157
rect 252651 330092 252652 330156
rect 252716 330092 252717 330156
rect 252651 330091 252717 330092
rect 299390 329562 299450 331451
rect 230939 328796 231005 328797
rect 230939 328732 230940 328796
rect 231004 328732 231005 328796
rect 230939 328731 231005 328732
rect 336374 326893 336434 331366
rect 339499 327436 339565 327437
rect 339499 327372 339500 327436
rect 339564 327372 339565 327436
rect 339499 327371 339565 327372
rect 340971 327436 341037 327437
rect 340971 327372 340972 327436
rect 341036 327372 341037 327436
rect 340971 327371 341037 327372
rect 336371 326892 336437 326893
rect 336371 326828 336372 326892
rect 336436 326828 336437 326892
rect 336371 326827 336437 326828
rect 104902 319894 105182 319954
rect 246211 316964 246277 316965
rect 246211 316900 246212 316964
rect 246276 316900 246277 316964
rect 246211 316899 246277 316900
rect 55955 315876 56021 315877
rect 55955 315812 55956 315876
rect 56020 315812 56021 315876
rect 55955 315811 56021 315812
rect 54854 311054 55098 311114
rect 54854 310981 54914 311054
rect 54851 310980 54917 310981
rect 54851 310916 54852 310980
rect 54916 310916 54917 310980
rect 54851 310915 54917 310916
rect 55035 310980 55101 310981
rect 55035 310916 55036 310980
rect 55100 310916 55101 310980
rect 55035 310915 55101 310916
rect 55038 308261 55098 310915
rect 55035 308260 55101 308261
rect 55035 308196 55036 308260
rect 55100 308196 55101 308260
rect 55035 308195 55101 308196
rect 54667 306220 54733 306221
rect 54667 306156 54668 306220
rect 54732 306156 54733 306220
rect 54667 306155 54733 306156
rect 52643 300644 52709 300645
rect 52643 300580 52644 300644
rect 52708 300580 52709 300644
rect 52643 300579 52709 300580
rect 5000 289936 5122 290172
rect 5358 289936 5442 290172
rect 5678 289936 5762 290172
rect 5998 289936 6082 290172
rect 6318 289936 6402 290172
rect 6638 289936 6722 290172
rect 6958 289936 7042 290172
rect 7278 289936 7362 290172
rect 7598 289936 7682 290172
rect 7918 289936 8002 290172
rect 8238 289936 8322 290172
rect 8558 289936 8642 290172
rect 8878 289936 9000 290172
rect 5000 259536 9000 289936
rect 38662 284002 38722 286486
rect 13638 283645 13698 283766
rect 13635 283644 13701 283645
rect 13635 283580 13636 283644
rect 13700 283580 13701 283644
rect 13635 283579 13701 283580
rect 52646 266781 52706 300579
rect 54483 287588 54549 287589
rect 54483 287524 54484 287588
rect 54548 287524 54549 287588
rect 54483 287523 54549 287524
rect 54486 272357 54546 287523
rect 54670 279293 54730 306155
rect 55035 300916 55101 300917
rect 55035 300852 55036 300916
rect 55100 300914 55101 300916
rect 55100 300854 55282 300914
rect 55100 300852 55101 300854
rect 55035 300851 55101 300852
rect 55035 292076 55101 292077
rect 55035 292012 55036 292076
rect 55100 292074 55101 292076
rect 55222 292074 55282 300854
rect 55100 292014 55282 292074
rect 55100 292012 55101 292014
rect 55035 292011 55101 292012
rect 55035 289050 55101 289051
rect 55035 288986 55036 289050
rect 55100 288986 55101 289050
rect 55035 288985 55101 288986
rect 55038 287589 55098 288985
rect 55035 287588 55101 287589
rect 55035 287524 55036 287588
rect 55100 287524 55101 287588
rect 55035 287523 55101 287524
rect 54667 279292 54733 279293
rect 54667 279228 54668 279292
rect 54732 279228 54733 279292
rect 54667 279227 54733 279228
rect 54667 279020 54733 279021
rect 54667 278956 54668 279020
rect 54732 278956 54733 279020
rect 54667 278955 54733 278956
rect 54483 272356 54549 272357
rect 54483 272292 54484 272356
rect 54548 272292 54549 272356
rect 54483 272291 54549 272292
rect 54670 266781 54730 278955
rect 55035 272356 55101 272357
rect 55035 272292 55036 272356
rect 55100 272292 55101 272356
rect 55035 272291 55101 272292
rect 55038 266781 55098 272291
rect 55958 266781 56018 315811
rect 73435 308260 73501 308261
rect 73435 308196 73436 308260
rect 73500 308196 73501 308260
rect 73435 308195 73501 308196
rect 52643 266780 52709 266781
rect 52643 266716 52644 266780
rect 52708 266716 52709 266780
rect 52643 266715 52709 266716
rect 54667 266780 54733 266781
rect 54667 266716 54668 266780
rect 54732 266716 54733 266780
rect 54667 266715 54733 266716
rect 55035 266780 55101 266781
rect 55035 266716 55036 266780
rect 55100 266716 55101 266780
rect 55035 266715 55101 266716
rect 55955 266780 56021 266781
rect 55955 266716 55956 266780
rect 56020 266716 56021 266780
rect 55955 266715 56021 266716
rect 73438 265965 73498 308195
rect 104534 307034 104594 307566
rect 104534 306974 104778 307034
rect 104718 305532 104778 306974
rect 104464 305490 104784 305532
rect 104464 305254 104506 305490
rect 104742 305254 104784 305490
rect 104464 305212 104784 305254
rect 198464 305490 198784 305532
rect 198464 305254 198506 305490
rect 198742 305254 198784 305490
rect 198464 305212 198784 305254
rect 104718 303634 104778 305212
rect 104534 303574 104778 303634
rect 104534 303042 104594 303574
rect 246214 298962 246274 316899
rect 339502 314653 339562 327371
rect 340974 314925 341034 327371
rect 435740 320808 439740 351208
rect 435740 320572 435862 320808
rect 436098 320572 436182 320808
rect 436418 320572 436502 320808
rect 436738 320572 436822 320808
rect 437058 320572 437142 320808
rect 437378 320572 437462 320808
rect 437698 320572 437782 320808
rect 438018 320572 438102 320808
rect 438338 320572 438422 320808
rect 438658 320572 438742 320808
rect 438978 320572 439062 320808
rect 439298 320572 439382 320808
rect 439618 320572 439740 320808
rect 353299 320228 353365 320229
rect 353299 320164 353300 320228
rect 353364 320164 353365 320228
rect 353299 320163 353365 320164
rect 345571 316556 345637 316557
rect 345571 316492 345572 316556
rect 345636 316492 345637 316556
rect 345571 316491 345637 316492
rect 345574 315197 345634 316491
rect 345571 315196 345637 315197
rect 345571 315132 345572 315196
rect 345636 315132 345637 315196
rect 345571 315131 345637 315132
rect 340971 314924 341037 314925
rect 340971 314860 340972 314924
rect 341036 314860 341037 314924
rect 340971 314859 341037 314860
rect 351827 314924 351893 314925
rect 351827 314860 351828 314924
rect 351892 314860 351893 314924
rect 351827 314859 351893 314860
rect 339499 314652 339565 314653
rect 339499 314588 339500 314652
rect 339564 314588 339565 314652
rect 339499 314587 339565 314588
rect 292464 305490 292784 305532
rect 292464 305254 292506 305490
rect 292742 305254 292784 305490
rect 292464 305212 292784 305254
rect 74539 298740 74605 298741
rect 74539 298676 74540 298740
rect 74604 298676 74605 298740
rect 74539 298675 74605 298676
rect 74171 291668 74237 291669
rect 74171 291604 74172 291668
rect 74236 291604 74237 291668
rect 74171 291603 74237 291604
rect 74174 288949 74234 291603
rect 74355 289084 74421 289085
rect 74355 289020 74356 289084
rect 74420 289020 74421 289084
rect 74355 289019 74421 289020
rect 74171 288948 74237 288949
rect 74171 288884 74172 288948
rect 74236 288884 74237 288948
rect 74171 288883 74237 288884
rect 74358 288813 74418 289019
rect 74355 288812 74421 288813
rect 74355 288748 74356 288812
rect 74420 288748 74421 288812
rect 74355 288747 74421 288748
rect 73619 282828 73685 282829
rect 73619 282764 73620 282828
rect 73684 282764 73685 282828
rect 73619 282763 73685 282764
rect 73435 265964 73501 265965
rect 73435 265900 73436 265964
rect 73500 265900 73501 265964
rect 73435 265899 73501 265900
rect 5000 259300 5122 259536
rect 5358 259300 5442 259536
rect 5678 259300 5762 259536
rect 5998 259300 6082 259536
rect 6318 259300 6402 259536
rect 6638 259300 6722 259536
rect 6958 259300 7042 259536
rect 7278 259300 7362 259536
rect 7598 259300 7682 259536
rect 7918 259300 8002 259536
rect 8238 259300 8322 259536
rect 8558 259300 8642 259536
rect 8878 259300 9000 259536
rect 5000 228900 9000 259300
rect 49147 252364 49213 252365
rect 49147 252300 49148 252364
rect 49212 252300 49213 252364
rect 49147 252299 49213 252300
rect 49150 252042 49210 252299
rect 48411 246652 48477 246653
rect 48411 246588 48412 246652
rect 48476 246588 48477 246652
rect 48411 246587 48477 246588
rect 48414 242522 48474 246587
rect 49147 243388 49213 243389
rect 49147 243324 49148 243388
rect 49212 243324 49213 243388
rect 49147 243323 49213 243324
rect 49150 243202 49210 243323
rect 49147 239852 49213 239853
rect 49147 239802 49148 239852
rect 49212 239802 49213 239852
rect 73622 237674 73682 282763
rect 74171 279428 74237 279429
rect 74171 279364 74172 279428
rect 74236 279364 74237 279428
rect 74171 279363 74237 279364
rect 74355 279428 74421 279429
rect 74355 279364 74356 279428
rect 74420 279364 74421 279428
rect 74355 279363 74421 279364
rect 73987 263516 74053 263517
rect 73987 263452 73988 263516
rect 74052 263452 74053 263516
rect 73987 263451 74053 263452
rect 73990 251362 74050 263451
rect 74174 252634 74234 279363
rect 74358 266101 74418 279363
rect 74355 266100 74421 266101
rect 74355 266036 74356 266100
rect 74420 266036 74421 266100
rect 74355 266035 74421 266036
rect 74355 265964 74421 265965
rect 74355 265900 74356 265964
rect 74420 265900 74421 265964
rect 74355 265899 74421 265900
rect 74358 263517 74418 265899
rect 74542 263517 74602 298675
rect 136918 295341 136978 297366
rect 230758 295341 230818 297366
rect 136915 295340 136981 295341
rect 136915 295276 136916 295340
rect 136980 295276 136981 295340
rect 136915 295275 136981 295276
rect 230755 295340 230821 295341
rect 230755 295276 230756 295340
rect 230820 295276 230821 295340
rect 230755 295275 230821 295276
rect 89104 290172 89424 290214
rect 89104 289936 89146 290172
rect 89382 289936 89424 290172
rect 89104 289894 89424 289936
rect 104718 289442 104778 291246
rect 136918 290034 136978 295275
rect 165619 291940 165685 291941
rect 165619 291876 165620 291940
rect 165684 291876 165685 291940
rect 165619 291875 165685 291876
rect 178683 291940 178749 291941
rect 178683 291876 178684 291940
rect 178748 291876 178749 291940
rect 178683 291875 178749 291876
rect 136918 289974 137162 290034
rect 84659 282828 84725 282829
rect 84659 282764 84660 282828
rect 84724 282764 84725 282828
rect 84659 282763 84725 282764
rect 84662 282642 84722 282763
rect 134710 282642 134770 285126
rect 137102 284866 137162 289974
rect 165622 289442 165682 291875
rect 178686 291482 178746 291875
rect 183104 290172 183424 290214
rect 183104 289936 183146 290172
rect 183382 289936 183424 290172
rect 183104 289894 183424 289936
rect 228734 289629 228794 293286
rect 229286 292213 229346 293966
rect 229283 292212 229349 292213
rect 229283 292148 229284 292212
rect 229348 292148 229349 292212
rect 229283 292147 229349 292148
rect 229286 291397 229346 292147
rect 229283 291396 229349 291397
rect 229283 291332 229284 291396
rect 229348 291332 229349 291396
rect 229283 291331 229349 291332
rect 228731 289628 228797 289629
rect 228731 289564 228732 289628
rect 228796 289564 228797 289628
rect 228731 289563 228797 289564
rect 236094 289085 236154 289206
rect 236091 289084 236157 289085
rect 236091 289020 236092 289084
rect 236156 289020 236157 289084
rect 236091 289019 236157 289020
rect 138571 284868 138637 284869
rect 137102 284806 137346 284866
rect 137286 284682 137346 284806
rect 138571 284804 138572 284868
rect 138636 284804 138637 284868
rect 138571 284803 138637 284804
rect 137286 282285 137346 284446
rect 138574 282642 138634 284803
rect 137283 282284 137349 282285
rect 137283 282220 137284 282284
rect 137348 282220 137349 282284
rect 137283 282219 137349 282220
rect 138574 278205 138634 282406
rect 138571 278204 138637 278205
rect 138571 278140 138572 278204
rect 138636 278140 138637 278204
rect 138571 278139 138637 278140
rect 104464 274854 104784 274896
rect 104464 274618 104506 274854
rect 104742 274618 104784 274854
rect 198464 274854 198784 274896
rect 104464 274576 104784 274618
rect 167827 274668 167893 274669
rect 167827 274604 167828 274668
rect 167892 274604 167893 274668
rect 167827 274603 167893 274604
rect 198464 274618 198506 274854
rect 198742 274618 198784 274854
rect 149059 274532 149125 274533
rect 149059 274468 149060 274532
rect 149124 274468 149125 274532
rect 149059 274467 149125 274468
rect 136915 273852 136981 273853
rect 136915 273788 136916 273852
rect 136980 273788 136981 273852
rect 136915 273787 136981 273788
rect 75275 266100 75341 266101
rect 75275 266036 75276 266100
rect 75340 266036 75341 266100
rect 75275 266035 75341 266036
rect 74355 263516 74421 263517
rect 74355 263452 74356 263516
rect 74420 263452 74421 263516
rect 74355 263451 74421 263452
rect 74539 263516 74605 263517
rect 74539 263452 74540 263516
rect 74604 263452 74605 263516
rect 74539 263451 74605 263452
rect 75278 258754 75338 266035
rect 75643 263516 75709 263517
rect 75643 263452 75644 263516
rect 75708 263452 75709 263516
rect 75643 263451 75709 263452
rect 74910 258694 75338 258754
rect 74174 252574 74418 252634
rect 74358 247962 74418 252574
rect 74910 251954 74970 258694
rect 75646 256034 75706 263451
rect 75646 255974 76110 256034
rect 74910 251894 75190 251954
rect 75278 251274 75338 251806
rect 76198 251362 76258 255886
rect 75278 251214 75890 251274
rect 73990 237674 74050 245006
rect 74358 244474 74418 247726
rect 74910 245154 74970 251126
rect 75278 249234 75338 250446
rect 74174 244414 74418 244474
rect 74726 245094 74970 245154
rect 75094 249174 75338 249234
rect 74174 239122 74234 244414
rect 74726 243114 74786 245094
rect 74358 243054 74786 243114
rect 74358 239714 74418 243054
rect 75094 242434 75154 249174
rect 75830 248554 75890 251214
rect 75646 248494 75890 248554
rect 75646 245242 75706 248494
rect 74726 242374 75154 242434
rect 74358 239654 74602 239714
rect 73402 237614 73682 237674
rect 73435 233868 73501 233869
rect 73435 233804 73436 233868
rect 73500 233804 73501 233868
rect 73435 233803 73501 233804
rect 73438 233733 73498 233803
rect 73435 233732 73501 233733
rect 73435 233668 73436 233732
rect 73500 233668 73501 233732
rect 73435 233667 73501 233668
rect 52643 232508 52709 232509
rect 52643 232444 52644 232508
rect 52708 232444 52709 232508
rect 52643 232443 52709 232444
rect 54667 232508 54733 232509
rect 54667 232444 54668 232508
rect 54732 232444 54733 232508
rect 54667 232443 54733 232444
rect 5000 228664 5122 228900
rect 5358 228664 5442 228900
rect 5678 228664 5762 228900
rect 5998 228664 6082 228900
rect 6318 228664 6402 228900
rect 6638 228664 6722 228900
rect 6958 228664 7042 228900
rect 7278 228664 7362 228900
rect 7598 228664 7682 228900
rect 7918 228664 8002 228900
rect 8238 228664 8322 228900
rect 8558 228664 8642 228900
rect 8878 228664 9000 228900
rect 5000 198264 9000 228664
rect 52646 206805 52706 232443
rect 54670 211021 54730 232443
rect 55403 231012 55469 231013
rect 55403 230948 55404 231012
rect 55468 230948 55469 231012
rect 55403 230947 55469 230948
rect 55406 222037 55466 230947
rect 55587 229652 55653 229653
rect 55587 229588 55588 229652
rect 55652 229588 55653 229652
rect 55587 229587 55653 229588
rect 55403 222036 55469 222037
rect 55403 221972 55404 222036
rect 55468 221972 55469 222036
rect 55403 221971 55469 221972
rect 55406 217954 55466 221971
rect 55590 221357 55650 229587
rect 55587 221356 55653 221357
rect 55587 221292 55588 221356
rect 55652 221292 55653 221356
rect 55587 221291 55653 221292
rect 56323 221356 56389 221357
rect 56323 221292 56324 221356
rect 56388 221292 56389 221356
rect 56323 221291 56389 221292
rect 55406 217894 55834 217954
rect 55774 215234 55834 217894
rect 55406 215174 55834 215234
rect 54667 211020 54733 211021
rect 54667 210956 54668 211020
rect 54732 210956 54733 211020
rect 54667 210955 54733 210956
rect 52643 206804 52709 206805
rect 52643 206740 52644 206804
rect 52708 206740 52709 206804
rect 52643 206739 52709 206740
rect 5000 198028 5122 198264
rect 5358 198028 5442 198264
rect 5678 198028 5762 198264
rect 5998 198028 6082 198264
rect 6318 198028 6402 198264
rect 6638 198028 6722 198264
rect 6958 198028 7042 198264
rect 7278 198028 7362 198264
rect 7598 198028 7682 198264
rect 7918 198028 8002 198264
rect 8238 198028 8322 198264
rect 8558 198028 8642 198264
rect 8878 198028 9000 198264
rect 5000 167628 9000 198028
rect 52646 171717 52706 206739
rect 54670 171717 54730 210955
rect 55406 172805 55466 215174
rect 56326 213874 56386 221291
rect 73435 214556 73501 214557
rect 73435 214492 73436 214556
rect 73500 214492 73501 214556
rect 73435 214491 73501 214492
rect 55590 213814 56386 213874
rect 55590 172941 55650 213814
rect 73438 205037 73498 214491
rect 73435 205036 73501 205037
rect 73435 204972 73436 205036
rect 73500 204972 73501 205036
rect 73435 204971 73501 204972
rect 73435 204900 73501 204901
rect 73435 204836 73436 204900
rect 73500 204836 73501 204900
rect 73435 204835 73501 204836
rect 55587 172940 55653 172941
rect 55587 172876 55588 172940
rect 55652 172876 55653 172940
rect 55587 172875 55653 172876
rect 55403 172804 55469 172805
rect 55403 172740 55404 172804
rect 55468 172740 55469 172804
rect 55403 172739 55469 172740
rect 52643 171716 52709 171717
rect 52643 171652 52644 171716
rect 52708 171652 52709 171716
rect 52643 171651 52709 171652
rect 54667 171716 54733 171717
rect 54667 171652 54668 171716
rect 54732 171652 54733 171716
rect 54667 171651 54733 171652
rect 73438 169541 73498 204835
rect 73622 204493 73682 237614
rect 73806 237614 74050 237674
rect 74128 238886 74132 239034
rect 73806 234005 73866 237614
rect 74128 236994 74188 238886
rect 74128 236934 74234 236994
rect 74174 236453 74234 236934
rect 73987 236452 74053 236453
rect 73987 236388 73988 236452
rect 74052 236388 74053 236452
rect 73987 236387 74053 236388
rect 74171 236452 74237 236453
rect 74171 236388 74172 236452
rect 74236 236388 74237 236452
rect 74171 236387 74237 236388
rect 73803 234004 73869 234005
rect 73803 233940 73804 234004
rect 73868 233940 73869 234004
rect 73803 233939 73869 233940
rect 73803 233732 73869 233733
rect 73803 233668 73804 233732
rect 73868 233668 73869 233732
rect 73803 233667 73869 233668
rect 73806 214557 73866 233667
rect 73990 229109 74050 236387
rect 74171 236316 74237 236317
rect 74171 236252 74172 236316
rect 74236 236252 74237 236316
rect 74171 236251 74237 236252
rect 74174 231013 74234 236251
rect 74542 235093 74602 239654
rect 74726 235637 74786 242374
rect 74723 235636 74789 235637
rect 74723 235572 74724 235636
rect 74788 235572 74789 235636
rect 74723 235571 74789 235572
rect 74539 235092 74605 235093
rect 74539 235028 74540 235092
rect 74604 235028 74605 235092
rect 74539 235027 74605 235028
rect 74539 234956 74605 234957
rect 74539 234892 74540 234956
rect 74604 234892 74605 234956
rect 74539 234891 74605 234892
rect 74171 231012 74237 231013
rect 74171 230948 74172 231012
rect 74236 230948 74237 231012
rect 74171 230947 74237 230948
rect 73987 229108 74053 229109
rect 73987 229044 73988 229108
rect 74052 229044 74053 229108
rect 73987 229043 74053 229044
rect 74355 229108 74421 229109
rect 74355 229044 74356 229108
rect 74420 229044 74421 229108
rect 74355 229043 74421 229044
rect 73987 228972 74053 228973
rect 73987 228908 73988 228972
rect 74052 228908 74053 228972
rect 73987 228907 74053 228908
rect 73803 214556 73869 214557
rect 73803 214492 73804 214556
rect 73868 214492 73869 214556
rect 73803 214491 73869 214492
rect 73990 206669 74050 228907
rect 74358 228834 74418 229043
rect 74542 228973 74602 234891
rect 75462 233869 75522 240246
rect 75830 239802 75890 242966
rect 136918 241842 136978 273787
rect 138571 269772 138637 269773
rect 138571 269708 138572 269772
rect 138636 269708 138637 269772
rect 138571 269707 138637 269708
rect 138574 262837 138634 269707
rect 149062 263381 149122 274467
rect 144091 263380 144157 263381
rect 144091 263316 144092 263380
rect 144156 263316 144157 263380
rect 144091 263315 144157 263316
rect 149059 263380 149125 263381
rect 149059 263316 149060 263380
rect 149124 263316 149125 263380
rect 149059 263315 149125 263316
rect 138571 262836 138637 262837
rect 138571 262772 138572 262836
rect 138636 262772 138637 262836
rect 138571 262771 138637 262772
rect 138755 262564 138821 262565
rect 138755 262500 138756 262564
rect 138820 262500 138821 262564
rect 138755 262499 138821 262500
rect 138758 259981 138818 262499
rect 138755 259980 138821 259981
rect 138755 259916 138756 259980
rect 138820 259916 138821 259980
rect 138755 259915 138821 259916
rect 144094 257482 144154 263315
rect 138939 250460 139005 250461
rect 138939 250396 138940 250460
rect 139004 250396 139005 250460
rect 138939 250395 139005 250396
rect 138942 243661 139002 250395
rect 138939 243660 139005 243661
rect 138939 243596 138940 243660
rect 139004 243596 139005 243660
rect 138939 243595 139005 243596
rect 138755 243388 138821 243389
rect 138755 243324 138756 243388
rect 138820 243324 138821 243388
rect 138755 243323 138821 243324
rect 96067 241756 96133 241757
rect 96067 241692 96068 241756
rect 96132 241692 96133 241756
rect 96067 241691 96133 241692
rect 104899 241756 104965 241757
rect 104899 241692 104900 241756
rect 104964 241692 104965 241756
rect 104899 241691 104965 241692
rect 96070 241162 96130 241691
rect 76563 241076 76629 241077
rect 76563 241074 76564 241076
rect 76198 241014 76564 241074
rect 76198 240482 76258 241014
rect 76563 241012 76564 241014
rect 76628 241012 76629 241076
rect 76563 241011 76629 241012
rect 104902 240482 104962 241691
rect 125875 240196 125876 240246
rect 125940 240196 125941 240246
rect 125875 240195 125941 240196
rect 128635 240196 128636 240246
rect 128700 240196 128701 240246
rect 128635 240195 128701 240196
rect 75830 236317 75890 239566
rect 92571 239444 92637 239445
rect 92571 239380 92572 239444
rect 92636 239380 92637 239444
rect 92571 239379 92637 239380
rect 75827 236316 75893 236317
rect 75827 236252 75828 236316
rect 75892 236252 75893 236316
rect 75827 236251 75893 236252
rect 75459 233868 75525 233869
rect 75459 233804 75460 233868
rect 75524 233804 75525 233868
rect 75459 233803 75525 233804
rect 74539 228972 74605 228973
rect 74539 228908 74540 228972
rect 74604 228908 74605 228972
rect 74539 228907 74605 228908
rect 74358 228774 74602 228834
rect 74355 221492 74421 221493
rect 74355 221428 74356 221492
rect 74420 221428 74421 221492
rect 74355 221427 74421 221428
rect 74171 213196 74237 213197
rect 74171 213132 74172 213196
rect 74236 213132 74237 213196
rect 74171 213131 74237 213132
rect 73987 206668 74053 206669
rect 73987 206604 73988 206668
rect 74052 206604 74053 206668
rect 73987 206603 74053 206604
rect 74174 205170 74234 213131
rect 74358 211701 74418 221427
rect 74355 211700 74421 211701
rect 74355 211636 74356 211700
rect 74420 211636 74421 211700
rect 74355 211635 74421 211636
rect 74355 205444 74421 205445
rect 74355 205380 74356 205444
rect 74420 205380 74421 205444
rect 74355 205379 74421 205380
rect 73990 205110 74234 205170
rect 73990 204901 74050 205110
rect 73987 204900 74053 204901
rect 73987 204836 73988 204900
rect 74052 204836 74053 204900
rect 73987 204835 74053 204836
rect 73619 204492 73685 204493
rect 73619 204428 73620 204492
rect 73684 204428 73685 204492
rect 73619 204427 73685 204428
rect 73619 203268 73685 203269
rect 73619 203204 73620 203268
rect 73684 203204 73685 203268
rect 73619 203203 73685 203204
rect 73435 169540 73501 169541
rect 73435 169476 73436 169540
rect 73500 169476 73501 169540
rect 73435 169475 73501 169476
rect 73622 168402 73682 203203
rect 74358 200549 74418 205379
rect 74355 200548 74421 200549
rect 74355 200484 74356 200548
rect 74420 200484 74421 200548
rect 74355 200483 74421 200484
rect 73803 199324 73869 199325
rect 73803 199260 73804 199324
rect 73868 199260 73869 199324
rect 73803 199259 73869 199260
rect 74171 199324 74237 199325
rect 74171 199260 74172 199324
rect 74236 199260 74237 199324
rect 74171 199259 74237 199260
rect 73806 189533 73866 199259
rect 73987 197964 74053 197965
rect 73987 197900 73988 197964
rect 74052 197900 74053 197964
rect 73987 197899 74053 197900
rect 73803 189532 73869 189533
rect 73803 189468 73804 189532
rect 73868 189468 73869 189532
rect 73803 189467 73869 189468
rect 73803 180012 73869 180013
rect 73803 179948 73804 180012
rect 73868 179948 73869 180012
rect 73803 179947 73869 179948
rect 73806 169269 73866 179947
rect 73990 169677 74050 197899
rect 74174 195245 74234 199259
rect 74542 199189 74602 228774
rect 92574 226525 92634 239379
rect 102323 238628 102389 238629
rect 102323 238564 102324 238628
rect 102388 238564 102389 238628
rect 102323 238563 102389 238564
rect 102326 238442 102386 238563
rect 110419 235772 110485 235773
rect 110419 235722 110420 235772
rect 110484 235722 110485 235772
rect 136918 235093 136978 241606
rect 138758 239802 138818 243323
rect 143726 239802 143786 241606
rect 144094 237082 144154 248406
rect 167830 240482 167890 274603
rect 198464 274576 198784 274618
rect 168563 274532 168629 274533
rect 168563 274468 168564 274532
rect 168628 274468 168629 274532
rect 168563 274467 168629 274468
rect 147958 235909 148018 237526
rect 148694 236045 148754 236846
rect 149246 236317 149306 237526
rect 149243 236316 149309 236317
rect 149243 236252 149244 236316
rect 149308 236252 149309 236316
rect 149243 236251 149309 236252
rect 149611 236116 149612 236166
rect 149676 236116 149677 236166
rect 149611 236115 149677 236116
rect 148691 236044 148757 236045
rect 148691 235980 148692 236044
rect 148756 235980 148757 236044
rect 148691 235979 148757 235980
rect 147955 235908 148021 235909
rect 147955 235844 147956 235908
rect 148020 235844 148021 235908
rect 147955 235843 148021 235844
rect 136915 235092 136981 235093
rect 136915 235028 136916 235092
rect 136980 235028 136981 235092
rect 136915 235027 136981 235028
rect 141150 234277 141210 234806
rect 141147 234276 141213 234277
rect 141147 234212 141148 234276
rect 141212 234212 141213 234276
rect 141147 234211 141213 234212
rect 147771 234276 147837 234277
rect 147771 234212 147772 234276
rect 147836 234274 147837 234276
rect 147955 234276 148021 234277
rect 147955 234274 147956 234276
rect 147836 234214 147956 234274
rect 147836 234212 147837 234214
rect 147771 234211 147837 234212
rect 147955 234212 147956 234214
rect 148020 234212 148021 234276
rect 147955 234211 148021 234212
rect 153107 234276 153173 234277
rect 153107 234212 153108 234276
rect 153172 234212 153173 234276
rect 153107 234211 153173 234212
rect 153110 233597 153170 234211
rect 167830 233597 167890 240246
rect 168566 235042 168626 274467
rect 169115 274396 169181 274397
rect 169115 274332 169116 274396
rect 169180 274332 169181 274396
rect 169115 274331 169181 274332
rect 169118 238442 169178 274331
rect 219715 268412 219781 268413
rect 219715 268348 219716 268412
rect 219780 268348 219781 268412
rect 219715 268347 219781 268348
rect 169118 233733 169178 238206
rect 219718 237813 219778 268347
rect 219715 237812 219781 237813
rect 219715 237748 219716 237812
rect 219780 237748 219781 237812
rect 219715 237747 219781 237748
rect 169115 233732 169181 233733
rect 169115 233668 169116 233732
rect 169180 233668 169181 233732
rect 169115 233667 169181 233668
rect 153107 233596 153173 233597
rect 153107 233532 153108 233596
rect 153172 233532 153173 233596
rect 153107 233531 153173 233532
rect 167827 233596 167893 233597
rect 167827 233532 167828 233596
rect 167892 233532 167893 233596
rect 167827 233531 167893 233532
rect 92571 226524 92637 226525
rect 92571 226460 92572 226524
rect 92636 226460 92637 226524
rect 92571 226459 92637 226460
rect 164883 216596 164949 216597
rect 164883 216532 164884 216596
rect 164948 216532 164949 216596
rect 164883 216531 164949 216532
rect 228918 216597 228978 217126
rect 164886 215322 164946 216531
rect 228915 216596 228981 216597
rect 228915 216532 228916 216596
rect 228980 216532 228981 216596
rect 228915 216531 228981 216532
rect 104464 213582 104784 213624
rect 104464 213346 104506 213582
rect 104742 213346 104784 213582
rect 104464 213304 104784 213346
rect 198464 213582 198784 213624
rect 198464 213346 198506 213582
rect 198742 213346 198784 213582
rect 198464 213304 198784 213346
rect 147035 208300 147101 208301
rect 147035 208236 147036 208300
rect 147100 208236 147101 208300
rect 147035 208235 147101 208236
rect 84659 204492 84725 204493
rect 84659 204442 84660 204492
rect 84724 204442 84725 204492
rect 74539 199188 74605 199189
rect 74539 199124 74540 199188
rect 74604 199124 74605 199188
rect 74539 199123 74605 199124
rect 74542 197965 74602 199123
rect 89104 198264 89424 198306
rect 89104 198028 89146 198264
rect 89382 198028 89424 198264
rect 138022 198237 138082 198766
rect 138019 198236 138085 198237
rect 138019 198172 138020 198236
rect 138084 198172 138085 198236
rect 138019 198171 138085 198172
rect 89104 197986 89424 198028
rect 74539 197964 74605 197965
rect 74539 197900 74540 197964
rect 74604 197900 74605 197964
rect 74539 197899 74605 197900
rect 74171 195244 74237 195245
rect 74171 195180 74172 195244
rect 74236 195180 74237 195244
rect 74171 195179 74237 195180
rect 74539 195244 74605 195245
rect 74539 195180 74540 195244
rect 74604 195180 74605 195244
rect 74539 195179 74605 195180
rect 74355 191028 74421 191029
rect 74355 190964 74356 191028
rect 74420 190964 74421 191028
rect 74355 190963 74421 190964
rect 74358 181237 74418 190963
rect 74542 187085 74602 195179
rect 138019 194700 138085 194701
rect 138019 194636 138020 194700
rect 138084 194636 138085 194700
rect 138019 194635 138085 194636
rect 138022 194242 138082 194635
rect 74539 187084 74605 187085
rect 74539 187020 74540 187084
rect 74604 187020 74605 187084
rect 74539 187019 74605 187020
rect 74539 186948 74605 186949
rect 74539 186884 74540 186948
rect 74604 186884 74605 186948
rect 74539 186883 74605 186884
rect 74355 181236 74421 181237
rect 74355 181172 74356 181236
rect 74420 181172 74421 181236
rect 74355 181171 74421 181172
rect 74171 180012 74237 180013
rect 74171 179948 74172 180012
rect 74236 179948 74237 180012
rect 74171 179947 74237 179948
rect 73987 169676 74053 169677
rect 73987 169612 73988 169676
rect 74052 169612 74053 169676
rect 73987 169611 74053 169612
rect 74174 169402 74234 179947
rect 74542 175797 74602 186883
rect 104464 182946 104784 182988
rect 104464 182710 104506 182946
rect 104742 182710 104784 182946
rect 104464 182668 104784 182710
rect 147038 181237 147098 208235
rect 230758 200685 230818 200806
rect 230755 200684 230821 200685
rect 230755 200620 230756 200684
rect 230820 200620 230821 200684
rect 230755 200619 230821 200620
rect 183104 198264 183424 198306
rect 183104 198028 183146 198264
rect 183382 198028 183424 198264
rect 230758 198237 230818 198766
rect 230755 198236 230821 198237
rect 230755 198172 230756 198236
rect 230820 198172 230821 198236
rect 230755 198171 230821 198172
rect 183104 197986 183424 198028
rect 236094 194922 236154 289019
rect 246214 282642 246274 298046
rect 322758 295477 322818 297366
rect 322755 295476 322821 295477
rect 322755 295412 322756 295476
rect 322820 295412 322821 295476
rect 322755 295411 322821 295412
rect 322758 292349 322818 293286
rect 322755 292348 322821 292349
rect 322755 292284 322756 292348
rect 322820 292284 322821 292348
rect 322755 292283 322821 292284
rect 259459 291940 259525 291941
rect 259459 291876 259460 291940
rect 259524 291876 259525 291940
rect 259459 291875 259525 291876
rect 272707 291940 272773 291941
rect 272707 291876 272708 291940
rect 272772 291876 272773 291940
rect 272707 291875 272773 291876
rect 258723 291396 258789 291397
rect 258723 291394 258724 291396
rect 257954 291334 258724 291394
rect 258723 291332 258724 291334
rect 258788 291332 258789 291396
rect 258723 291331 258789 291332
rect 259462 289442 259522 291875
rect 272710 291482 272770 291875
rect 277104 290172 277424 290214
rect 277104 289936 277146 290172
rect 277382 289936 277424 290172
rect 277104 289894 277424 289936
rect 322758 289629 322818 291246
rect 322755 289628 322821 289629
rect 322755 289564 322756 289628
rect 322820 289564 322821 289628
rect 322755 289563 322821 289564
rect 351830 285362 351890 314859
rect 352011 314652 352077 314653
rect 352011 314588 352012 314652
rect 352076 314588 352077 314652
rect 353302 314602 353362 320163
rect 355691 315332 355757 315333
rect 355691 315268 355692 315332
rect 355756 315268 355757 315332
rect 355691 315267 355757 315268
rect 352011 314587 352077 314588
rect 352014 311794 352074 314587
rect 352014 311734 352258 311794
rect 352198 310434 352258 311734
rect 352014 310374 352258 310434
rect 352014 292754 352074 310374
rect 352014 292694 352626 292754
rect 352566 286634 352626 292694
rect 352382 286574 352626 286634
rect 351830 284594 351890 285126
rect 351830 284534 352074 284594
rect 352014 281194 352074 284534
rect 351830 281134 352074 281194
rect 242347 273852 242413 273853
rect 242347 273788 242348 273852
rect 242412 273788 242413 273852
rect 242347 273787 242413 273788
rect 241979 273716 242045 273717
rect 241979 273652 241980 273716
rect 242044 273652 242045 273716
rect 241979 273651 242045 273652
rect 237195 263516 237261 263517
rect 237195 263452 237196 263516
rect 237260 263452 237261 263516
rect 237195 263451 237261 263452
rect 237198 254133 237258 263451
rect 241982 263381 242042 273651
rect 242350 263517 242410 273787
rect 246214 273717 246274 279006
rect 292464 274854 292784 274896
rect 247867 274668 247933 274669
rect 247867 274604 247868 274668
rect 247932 274604 247933 274668
rect 247867 274603 247933 274604
rect 292464 274618 292506 274854
rect 292742 274618 292784 274854
rect 247870 274397 247930 274603
rect 292464 274576 292784 274618
rect 262403 274532 262469 274533
rect 262403 274468 262404 274532
rect 262468 274468 262469 274532
rect 262403 274467 262469 274468
rect 247867 274396 247933 274397
rect 247867 274332 247868 274396
rect 247932 274332 247933 274396
rect 247867 274331 247933 274332
rect 246211 273716 246277 273717
rect 246211 273652 246212 273716
rect 246276 273652 246277 273716
rect 246211 273651 246277 273652
rect 242347 263516 242413 263517
rect 242347 263452 242348 263516
rect 242412 263452 242413 263516
rect 242347 263451 242413 263452
rect 237563 263380 237629 263381
rect 237563 263316 237564 263380
rect 237628 263316 237629 263380
rect 237563 263315 237629 263316
rect 241979 263380 242045 263381
rect 241979 263316 241980 263380
rect 242044 263316 242045 263380
rect 241979 263315 242045 263316
rect 236643 254132 236709 254133
rect 236643 254068 236644 254132
rect 236708 254068 236709 254132
rect 236643 254067 236709 254068
rect 237195 254132 237261 254133
rect 237195 254068 237196 254132
rect 237260 254068 237261 254132
rect 237195 254067 237261 254068
rect 236646 249322 236706 254067
rect 237566 253994 237626 263315
rect 247870 262242 247930 274331
rect 261851 272220 261917 272221
rect 261851 272156 261852 272220
rect 261916 272156 261917 272220
rect 261851 272155 261917 272156
rect 261854 268277 261914 272155
rect 261851 268276 261917 268277
rect 261851 268212 261852 268276
rect 261916 268212 261917 268276
rect 261851 268211 261917 268212
rect 262219 268276 262285 268277
rect 262219 268212 262220 268276
rect 262284 268212 262285 268276
rect 262219 268211 262285 268212
rect 238118 257482 238178 259966
rect 262222 258754 262282 268211
rect 261670 258694 262282 258754
rect 237382 253934 237626 253994
rect 237382 245154 237442 253934
rect 237382 245094 237810 245154
rect 237014 242522 237074 245006
rect 237750 234957 237810 245094
rect 238118 238442 238178 249086
rect 261670 240482 261730 258694
rect 262038 238442 262098 241606
rect 238118 236181 238178 238206
rect 248790 236181 248850 237526
rect 238115 236180 238181 236181
rect 238115 236116 238116 236180
rect 238180 236116 238181 236180
rect 238115 236115 238181 236116
rect 248787 236180 248853 236181
rect 248787 236116 248788 236180
rect 248852 236116 248853 236180
rect 248787 236115 248853 236116
rect 262038 235909 262098 238206
rect 262035 235908 262101 235909
rect 262035 235844 262036 235908
rect 262100 235844 262101 235908
rect 262035 235843 262101 235844
rect 262406 235773 262466 274467
rect 262955 274396 263021 274397
rect 262955 274332 262956 274396
rect 263020 274332 263021 274396
rect 262955 274331 263021 274332
rect 262958 239802 263018 274331
rect 276755 269500 276821 269501
rect 276755 269436 276756 269500
rect 276820 269436 276821 269500
rect 276755 269435 276821 269436
rect 262403 235772 262469 235773
rect 262403 235708 262404 235772
rect 262468 235708 262469 235772
rect 262403 235707 262469 235708
rect 237747 234956 237813 234957
rect 237747 234892 237748 234956
rect 237812 234892 237813 234956
rect 237747 234891 237813 234892
rect 244371 234956 244437 234957
rect 244371 234892 244372 234956
rect 244436 234892 244437 234956
rect 244371 234891 244437 234892
rect 244374 234362 244434 234891
rect 249894 233597 249954 234806
rect 249891 233596 249957 233597
rect 249891 233532 249892 233596
rect 249956 233532 249957 233596
rect 249891 233531 249957 233532
rect 262958 233461 263018 239566
rect 262955 233460 263021 233461
rect 262955 233396 262956 233460
rect 263020 233396 263021 233460
rect 262955 233395 263021 233396
rect 269214 232917 269274 233446
rect 269211 232916 269277 232917
rect 269211 232852 269212 232916
rect 269276 232852 269277 232916
rect 269211 232851 269277 232852
rect 276758 226661 276818 269435
rect 351830 266781 351890 281134
rect 352382 280514 352442 286574
rect 352198 280454 352442 280514
rect 352198 279698 352258 280454
rect 352747 279700 352813 279701
rect 352747 279698 352748 279700
rect 352198 279638 352748 279698
rect 352198 272354 352258 279638
rect 352747 279636 352748 279638
rect 352812 279636 352813 279700
rect 352747 279635 352813 279636
rect 352014 272294 352258 272354
rect 351827 266780 351893 266781
rect 351827 266716 351828 266780
rect 351892 266716 351893 266780
rect 351827 266715 351893 266716
rect 352014 266645 352074 272294
rect 352011 266644 352077 266645
rect 352011 266580 352012 266644
rect 352076 266580 352077 266644
rect 352011 266579 352077 266580
rect 355694 256122 355754 315267
rect 412182 308482 412242 314366
rect 412182 282642 412242 306206
rect 429478 305813 429538 306206
rect 429475 305812 429541 305813
rect 429475 305748 429476 305812
rect 429540 305748 429541 305812
rect 429475 305747 429541 305748
rect 435740 290172 439740 320572
rect 435740 289936 435862 290172
rect 436098 289936 436182 290172
rect 436418 289936 436502 290172
rect 436738 289936 436822 290172
rect 437058 289936 437142 290172
rect 437378 289936 437462 290172
rect 437698 289936 437782 290172
rect 438018 289936 438102 290172
rect 438338 289936 438422 290172
rect 438658 289936 438742 290172
rect 438978 289936 439062 290172
rect 439298 289936 439382 290172
rect 439618 289936 439740 290172
rect 415126 277253 415186 278326
rect 415123 277252 415189 277253
rect 415123 277188 415124 277252
rect 415188 277188 415189 277252
rect 415123 277187 415189 277188
rect 435740 259536 439740 289936
rect 435740 259300 435862 259536
rect 436098 259300 436182 259536
rect 436418 259300 436502 259536
rect 436738 259300 436822 259536
rect 437058 259300 437142 259536
rect 437378 259300 437462 259536
rect 437698 259300 437782 259536
rect 438018 259300 438102 259536
rect 438338 259300 438422 259536
rect 438658 259300 438742 259536
rect 438978 259300 439062 259536
rect 439298 259300 439382 259536
rect 439618 259300 439740 259536
rect 325147 250324 325213 250325
rect 325147 250260 325148 250324
rect 325212 250260 325213 250324
rect 325147 250259 325213 250260
rect 325150 249322 325210 250259
rect 325150 239714 325210 249086
rect 325150 239654 325614 239714
rect 284299 239444 284365 239445
rect 284299 239380 284300 239444
rect 284364 239380 284365 239444
rect 284299 239379 284365 239380
rect 284302 235042 284362 239379
rect 284302 234413 284362 234806
rect 284299 234412 284365 234413
rect 284299 234348 284300 234412
rect 284364 234348 284365 234412
rect 284299 234347 284365 234348
rect 297550 233597 297610 234806
rect 297547 233596 297613 233597
rect 297547 233532 297548 233596
rect 297612 233532 297613 233596
rect 297547 233531 297613 233532
rect 285222 232917 285282 233446
rect 285219 232916 285285 232917
rect 285219 232852 285220 232916
rect 285284 232852 285285 232916
rect 285219 232851 285285 232852
rect 325702 228834 325762 239566
rect 351643 232508 351709 232509
rect 351643 232444 351644 232508
rect 351708 232444 351709 232508
rect 351643 232443 351709 232444
rect 351827 232508 351893 232509
rect 351827 232444 351828 232508
rect 351892 232444 351893 232508
rect 351827 232443 351893 232444
rect 325518 228774 325762 228834
rect 325518 228293 325578 228774
rect 324595 228292 324661 228293
rect 324595 228228 324596 228292
rect 324660 228228 324661 228292
rect 324595 228227 324661 228228
rect 325515 228292 325581 228293
rect 325515 228228 325516 228292
rect 325580 228228 325581 228292
rect 325515 228227 325581 228228
rect 324598 228154 324658 228227
rect 324598 228094 325026 228154
rect 276755 226660 276821 226661
rect 276755 226596 276756 226660
rect 276820 226596 276821 226660
rect 276755 226595 276821 226596
rect 324966 224349 325026 228094
rect 324963 224348 325029 224349
rect 324963 224284 324964 224348
rect 325028 224284 325029 224348
rect 324963 224283 325029 224284
rect 242718 217005 242778 217126
rect 258726 217005 258786 217126
rect 272710 217005 272770 217126
rect 322939 217076 322940 217126
rect 323004 217076 323005 217126
rect 322939 217075 323005 217076
rect 336926 217005 336986 217126
rect 242715 217004 242781 217005
rect 242715 216940 242716 217004
rect 242780 216940 242781 217004
rect 242715 216939 242781 216940
rect 258723 217004 258789 217005
rect 258723 216940 258724 217004
rect 258788 216940 258789 217004
rect 258723 216939 258789 216940
rect 272707 217004 272773 217005
rect 272707 216940 272708 217004
rect 272772 216940 272773 217004
rect 272707 216939 272773 216940
rect 336923 217004 336989 217005
rect 336923 216940 336924 217004
rect 336988 216940 336989 217004
rect 336923 216939 336989 216940
rect 322939 216596 323005 216597
rect 322939 216532 322940 216596
rect 323004 216532 323005 216596
rect 322939 216531 323005 216532
rect 322942 216002 323002 216531
rect 292464 213582 292784 213624
rect 292464 213346 292506 213582
rect 292742 213346 292784 213582
rect 292464 213304 292784 213346
rect 236094 194565 236154 194686
rect 236091 194564 236157 194565
rect 236091 194500 236092 194564
rect 236156 194500 236157 194564
rect 236091 194499 236157 194500
rect 228731 194428 228797 194429
rect 228731 194364 228732 194428
rect 228796 194364 228797 194428
rect 228731 194363 228797 194364
rect 228734 194242 228794 194363
rect 242534 183141 242594 207606
rect 322755 198716 322756 198766
rect 322820 198716 322821 198766
rect 322755 198715 322821 198716
rect 277104 198264 277424 198306
rect 277104 198028 277146 198264
rect 277382 198028 277424 198264
rect 277104 197986 277424 198028
rect 351646 184093 351706 232443
rect 351830 191434 351890 232443
rect 355694 225437 355754 255886
rect 358635 255836 358636 255886
rect 358700 255836 358701 255886
rect 358635 255835 358701 255836
rect 360475 252908 360541 252909
rect 360475 252844 360476 252908
rect 360540 252844 360541 252908
rect 360475 252843 360541 252844
rect 360478 239122 360538 252843
rect 376840 228900 377160 228942
rect 376840 228664 376882 228900
rect 377118 228664 377160 228900
rect 376840 228622 377160 228664
rect 435740 228900 439740 259300
rect 435740 228664 435862 228900
rect 436098 228664 436182 228900
rect 436418 228664 436502 228900
rect 436738 228664 436822 228900
rect 437058 228664 437142 228900
rect 437378 228664 437462 228900
rect 437698 228664 437782 228900
rect 438018 228664 438102 228900
rect 438338 228664 438422 228900
rect 438658 228664 438742 228900
rect 438978 228664 439062 228900
rect 439298 228664 439382 228900
rect 439618 228664 439740 228900
rect 355691 225436 355757 225437
rect 355691 225372 355692 225436
rect 355756 225372 355757 225436
rect 355691 225371 355757 225372
rect 352750 217005 352810 217126
rect 352747 217004 352813 217005
rect 352747 216940 352748 217004
rect 352812 216940 352813 217004
rect 352747 216939 352813 216940
rect 435740 198264 439740 228664
rect 435740 198028 435862 198264
rect 436098 198028 436182 198264
rect 436418 198028 436502 198264
rect 436738 198028 436822 198264
rect 437058 198028 437142 198264
rect 437378 198028 437462 198264
rect 437698 198028 437782 198264
rect 438018 198028 438102 198264
rect 438338 198028 438422 198264
rect 438658 198028 438742 198264
rect 438978 198028 439062 198264
rect 439298 198028 439382 198264
rect 439618 198028 439740 198264
rect 352747 191436 352813 191437
rect 352747 191434 352748 191436
rect 351830 191374 352748 191434
rect 351643 184092 351709 184093
rect 351643 184028 351644 184092
rect 351708 184028 351709 184092
rect 351643 184027 351709 184028
rect 242531 183140 242597 183141
rect 242531 183076 242532 183140
rect 242596 183076 242597 183140
rect 242531 183075 242597 183076
rect 198464 182946 198784 182988
rect 198464 182710 198506 182946
rect 198742 182710 198784 182946
rect 198464 182668 198784 182710
rect 292464 182946 292784 182988
rect 292464 182710 292506 182946
rect 292742 182710 292784 182946
rect 292464 182668 292784 182710
rect 271419 182188 271485 182189
rect 271419 182124 271420 182188
rect 271484 182124 271485 182188
rect 271419 182123 271485 182124
rect 323123 182188 323189 182189
rect 323123 182124 323124 182188
rect 323188 182124 323189 182188
rect 323123 182123 323189 182124
rect 174819 182052 174885 182053
rect 174819 181988 174820 182052
rect 174884 181988 174885 182052
rect 174819 181987 174885 181988
rect 228731 182052 228797 182053
rect 228731 181988 228732 182052
rect 228796 181988 228797 182052
rect 271422 182002 271482 182123
rect 228731 181987 228797 181988
rect 174822 181322 174882 181987
rect 147035 181236 147101 181237
rect 147035 181172 147036 181236
rect 147100 181172 147101 181236
rect 147035 181171 147101 181172
rect 168563 181100 168629 181101
rect 168563 181036 168564 181100
rect 168628 181036 168629 181100
rect 168563 181035 168629 181036
rect 167827 180964 167893 180965
rect 167827 180900 167828 180964
rect 167892 180900 167893 180964
rect 167827 180899 167893 180900
rect 167643 180692 167709 180693
rect 167643 180628 167644 180692
rect 167708 180628 167709 180692
rect 167643 180627 167709 180628
rect 141515 180556 141581 180557
rect 141515 180492 141516 180556
rect 141580 180492 141581 180556
rect 141515 180491 141581 180492
rect 74539 175796 74605 175797
rect 74539 175732 74540 175796
rect 74604 175732 74605 175796
rect 74539 175731 74605 175732
rect 75091 175796 75157 175797
rect 75091 175732 75092 175796
rect 75156 175732 75157 175796
rect 75091 175731 75157 175732
rect 74355 171716 74421 171717
rect 74355 171652 74356 171716
rect 74420 171652 74421 171716
rect 74355 171651 74421 171652
rect 73990 169342 74234 169402
rect 73803 169268 73869 169269
rect 73803 169204 73804 169268
rect 73868 169204 73869 169268
rect 73803 169203 73869 169204
rect 5000 167392 5122 167628
rect 5358 167392 5442 167628
rect 5678 167392 5762 167628
rect 5998 167392 6082 167628
rect 6318 167392 6402 167628
rect 6638 167392 6722 167628
rect 6958 167392 7042 167628
rect 7278 167392 7362 167628
rect 7598 167392 7682 167628
rect 7918 167392 8002 167628
rect 8238 167392 8322 167628
rect 8558 167392 8642 167628
rect 8878 167392 9000 167628
rect 5000 136992 9000 167392
rect 49147 162332 49213 162333
rect 49147 162282 49148 162332
rect 49212 162282 49213 162332
rect 49147 158388 49213 158389
rect 49147 158324 49148 158388
rect 49212 158324 49213 158388
rect 49147 158323 49213 158324
rect 49150 158202 49210 158323
rect 73990 158114 74050 169342
rect 74358 163554 74418 171651
rect 74723 169268 74789 169269
rect 74723 169204 74724 169268
rect 74788 169204 74789 169268
rect 74723 169203 74789 169204
rect 74174 163494 74418 163554
rect 74174 161514 74234 163494
rect 74726 162282 74786 169203
rect 74174 161454 74970 161514
rect 74542 158794 74602 160686
rect 74542 158734 74786 158794
rect 73990 158054 74602 158114
rect 73806 155394 73866 157286
rect 73622 155334 73866 155394
rect 49150 152949 49210 153206
rect 49147 152948 49213 152949
rect 49147 152884 49148 152948
rect 49212 152884 49213 152948
rect 49147 152883 49213 152884
rect 49147 149004 49213 149005
rect 49147 148940 49148 149004
rect 49212 148940 49213 149004
rect 49147 148939 49213 148940
rect 49150 148682 49210 148939
rect 49147 146148 49213 146149
rect 49147 146084 49148 146148
rect 49212 146084 49213 146148
rect 49147 146083 49213 146084
rect 49150 145962 49210 146083
rect 73622 143834 73682 155334
rect 74542 154034 74602 158054
rect 73990 153974 74602 154034
rect 73990 153442 74050 153974
rect 73990 151994 74050 153206
rect 73990 151934 74418 151994
rect 74358 151402 74418 151934
rect 74726 150634 74786 158734
rect 74910 153354 74970 161454
rect 75094 154034 75154 175731
rect 75643 169812 75709 169813
rect 75643 169748 75644 169812
rect 75708 169748 75709 169812
rect 75643 169747 75709 169748
rect 75459 169676 75525 169677
rect 75459 169612 75460 169676
rect 75524 169612 75525 169676
rect 75459 169611 75525 169612
rect 75462 165594 75522 169611
rect 75646 166274 75706 169747
rect 76011 169540 76077 169541
rect 76011 169476 76012 169540
rect 76076 169476 76077 169540
rect 76011 169475 76077 169476
rect 76014 166954 76074 169475
rect 76014 166894 76442 166954
rect 75646 166214 76074 166274
rect 75462 165534 75706 165594
rect 75646 155482 75706 165534
rect 75094 153974 75522 154034
rect 74910 153294 75154 153354
rect 74358 150574 74786 150634
rect 74358 149954 74418 150574
rect 73990 149894 74418 149954
rect 73622 143774 73866 143834
rect 73806 141389 73866 143774
rect 73990 142477 74050 149894
rect 74358 148594 74418 149126
rect 74174 148534 74418 148594
rect 73987 142476 74053 142477
rect 73987 142412 73988 142476
rect 74052 142412 74053 142476
rect 73987 142411 74053 142412
rect 73803 141388 73869 141389
rect 73803 141324 73804 141388
rect 73868 141324 73869 141388
rect 73803 141323 73869 141324
rect 73806 139621 73866 141323
rect 52643 139620 52709 139621
rect 52643 139556 52644 139620
rect 52708 139556 52709 139620
rect 52643 139555 52709 139556
rect 54667 139620 54733 139621
rect 54667 139556 54668 139620
rect 54732 139556 54733 139620
rect 54667 139555 54733 139556
rect 73803 139620 73869 139621
rect 73803 139556 73804 139620
rect 73868 139556 73869 139620
rect 73803 139555 73869 139556
rect 5000 136756 5122 136992
rect 5358 136756 5442 136992
rect 5678 136756 5762 136992
rect 5998 136756 6082 136992
rect 6318 136756 6402 136992
rect 6638 136756 6722 136992
rect 6958 136756 7042 136992
rect 7278 136756 7362 136992
rect 7598 136756 7682 136992
rect 7918 136756 8002 136992
rect 8238 136756 8322 136992
rect 8558 136756 8642 136992
rect 8878 136756 9000 136992
rect 5000 106356 9000 136756
rect 52646 113101 52706 139555
rect 54115 131596 54181 131597
rect 54115 131532 54116 131596
rect 54180 131532 54181 131596
rect 54115 131531 54181 131532
rect 54118 122757 54178 131531
rect 54115 122756 54181 122757
rect 54115 122692 54116 122756
rect 54180 122692 54181 122756
rect 54115 122691 54181 122692
rect 52643 113100 52709 113101
rect 52643 113036 52644 113100
rect 52708 113036 52709 113100
rect 52643 113035 52709 113036
rect 5000 106120 5122 106356
rect 5358 106120 5442 106356
rect 5678 106120 5762 106356
rect 5998 106120 6082 106356
rect 6318 106120 6402 106356
rect 6638 106120 6722 106356
rect 6958 106120 7042 106356
rect 7278 106120 7362 106356
rect 7598 106120 7682 106356
rect 7918 106120 8002 106356
rect 8238 106120 8322 106356
rect 8558 106120 8642 106356
rect 8878 106120 9000 106356
rect 5000 75720 9000 106120
rect 52646 79101 52706 113035
rect 52643 79100 52709 79101
rect 52643 79036 52644 79100
rect 52708 79036 52709 79100
rect 52643 79035 52709 79036
rect 54118 78965 54178 122691
rect 54670 117181 54730 139555
rect 73990 139074 74050 142411
rect 74174 142341 74234 148534
rect 74726 147914 74786 149806
rect 75094 148682 75154 153294
rect 74726 147854 75154 147914
rect 75094 146554 75154 147854
rect 75462 146554 75522 153974
rect 74726 146494 75154 146554
rect 75278 146494 75522 146554
rect 74726 145874 74786 146494
rect 75278 145962 75338 146494
rect 74358 145814 74786 145874
rect 74171 142340 74237 142341
rect 74171 142276 74172 142340
rect 74236 142276 74237 142340
rect 74171 142275 74237 142276
rect 73438 139014 74050 139074
rect 55403 132412 55469 132413
rect 55403 132348 55404 132412
rect 55468 132348 55469 132412
rect 55403 132347 55469 132348
rect 55406 127245 55466 132347
rect 55403 127244 55469 127245
rect 55403 127180 55404 127244
rect 55468 127180 55469 127244
rect 55403 127179 55469 127180
rect 54667 117180 54733 117181
rect 54667 117116 54668 117180
rect 54732 117116 54733 117180
rect 54667 117115 54733 117116
rect 54670 79101 54730 117115
rect 55406 79101 55466 127179
rect 73438 112829 73498 139014
rect 73987 138940 74053 138941
rect 73987 138876 73988 138940
rect 74052 138876 74053 138940
rect 73987 138875 74053 138876
rect 73990 117994 74050 138875
rect 73806 117934 74050 117994
rect 73435 112828 73501 112829
rect 73435 112764 73436 112828
rect 73500 112764 73501 112828
rect 73435 112763 73501 112764
rect 73806 107794 73866 117934
rect 73622 107734 73866 107794
rect 73622 98277 73682 107734
rect 74174 102085 74234 142275
rect 74358 141797 74418 145814
rect 75278 143922 75338 145726
rect 74910 142477 74970 143006
rect 74907 142476 74973 142477
rect 74907 142412 74908 142476
rect 74972 142412 74973 142476
rect 74907 142411 74973 142412
rect 74355 141796 74421 141797
rect 74355 141732 74356 141796
rect 74420 141732 74421 141796
rect 74355 141731 74421 141732
rect 75646 141661 75706 155246
rect 75643 141660 75709 141661
rect 74726 141389 74786 141646
rect 75643 141596 75644 141660
rect 75708 141596 75709 141660
rect 75643 141595 75709 141596
rect 76014 141525 76074 166214
rect 76382 150042 76442 166894
rect 76750 158202 76810 168166
rect 77118 142341 77178 145046
rect 77670 144602 77730 148446
rect 77115 142340 77181 142341
rect 77115 142276 77116 142340
rect 77180 142276 77181 142340
rect 77115 142275 77181 142276
rect 77670 142069 77730 144366
rect 76379 142068 76445 142069
rect 76379 142004 76380 142068
rect 76444 142004 76445 142068
rect 76379 142003 76445 142004
rect 77667 142068 77733 142069
rect 77667 142004 77668 142068
rect 77732 142004 77733 142068
rect 77667 142003 77733 142004
rect 76011 141524 76077 141525
rect 76011 141460 76012 141524
rect 76076 141460 76077 141524
rect 76011 141459 76077 141460
rect 74723 141388 74789 141389
rect 74723 141324 74724 141388
rect 74788 141324 74789 141388
rect 74723 141323 74789 141324
rect 76382 141253 76442 142003
rect 74539 141252 74605 141253
rect 74539 141188 74540 141252
rect 74604 141188 74605 141252
rect 74539 141187 74605 141188
rect 76379 141252 76445 141253
rect 76379 141188 76380 141252
rect 76444 141188 76445 141252
rect 76379 141187 76445 141188
rect 74542 139754 74602 141187
rect 74542 139694 74786 139754
rect 74539 139620 74605 139621
rect 74539 139556 74540 139620
rect 74604 139556 74605 139620
rect 74539 139555 74605 139556
rect 74542 109565 74602 139555
rect 74726 138941 74786 139694
rect 74723 138940 74789 138941
rect 74723 138876 74724 138940
rect 74788 138876 74789 138940
rect 74723 138875 74789 138876
rect 78038 110925 78098 143686
rect 106003 142612 106069 142613
rect 106003 142548 106004 142612
rect 106068 142548 106069 142612
rect 106003 142547 106069 142548
rect 106006 141933 106066 142547
rect 106003 141932 106069 141933
rect 106003 141882 106004 141932
rect 106068 141882 106069 141932
rect 137102 134453 137162 143006
rect 141518 139893 141578 180491
rect 148691 173076 148757 173077
rect 148691 173012 148692 173076
rect 148756 173012 148757 173076
rect 148691 173011 148757 173012
rect 148694 169269 148754 173011
rect 144091 169268 144157 169269
rect 144091 169204 144092 169268
rect 144156 169204 144157 169268
rect 144091 169203 144157 169204
rect 148691 169268 148757 169269
rect 148691 169204 148692 169268
rect 148756 169204 148757 169268
rect 148691 169203 148757 169204
rect 144094 162282 144154 169203
rect 144094 151402 144154 160006
rect 144094 142205 144154 145046
rect 148326 143774 148938 143834
rect 147038 142477 147098 143006
rect 147035 142476 147101 142477
rect 147035 142412 147036 142476
rect 147100 142412 147101 142476
rect 147035 142411 147101 142412
rect 144091 142204 144157 142205
rect 144091 142140 144092 142204
rect 144156 142140 144157 142204
rect 144091 142139 144157 142140
rect 148326 142069 148386 143774
rect 148878 143242 148938 143774
rect 150350 142477 150410 143006
rect 150347 142476 150413 142477
rect 150347 142412 150348 142476
rect 150412 142412 150413 142476
rect 150347 142411 150413 142412
rect 147771 142068 147837 142069
rect 147771 142004 147772 142068
rect 147836 142004 147837 142068
rect 147771 142003 147837 142004
rect 148323 142068 148389 142069
rect 148323 142004 148324 142068
rect 148388 142004 148389 142068
rect 148323 142003 148389 142004
rect 141515 139892 141581 139893
rect 141515 139828 141516 139892
rect 141580 139828 141581 139892
rect 141515 139827 141581 139828
rect 137099 134452 137165 134453
rect 137099 134388 137100 134452
rect 137164 134388 137165 134452
rect 137099 134387 137165 134388
rect 104464 121674 104784 121716
rect 104464 121438 104506 121674
rect 104742 121438 104784 121674
rect 104464 121396 104784 121438
rect 145014 116637 145074 117166
rect 145011 116636 145077 116637
rect 145011 116572 145012 116636
rect 145076 116572 145077 116636
rect 145011 116571 145077 116572
rect 147774 113645 147834 142003
rect 149059 141116 149125 141117
rect 149059 141052 149060 141116
rect 149124 141052 149125 141116
rect 149059 141051 149125 141052
rect 149062 140522 149122 141051
rect 167646 140522 167706 180627
rect 167830 142205 167890 180899
rect 167827 142204 167893 142205
rect 167827 142140 167828 142204
rect 167892 142140 167893 142204
rect 167827 142139 167893 142140
rect 168566 141202 168626 181035
rect 169299 180828 169365 180829
rect 169299 180764 169300 180828
rect 169364 180764 169365 180828
rect 169299 180763 169365 180764
rect 169302 172941 169362 180763
rect 228734 180642 228794 181987
rect 323126 181322 323186 182123
rect 323491 182052 323557 182053
rect 323491 182002 323492 182052
rect 323556 182002 323557 182052
rect 261667 180828 261733 180829
rect 261667 180764 261668 180828
rect 261732 180764 261733 180828
rect 261667 180763 261733 180764
rect 242347 180284 242413 180285
rect 242347 180220 242348 180284
rect 242412 180220 242413 180284
rect 242347 180219 242413 180220
rect 241795 180148 241861 180149
rect 241795 180084 241796 180148
rect 241860 180084 241861 180148
rect 241795 180083 241861 180084
rect 219715 175524 219781 175525
rect 219715 175460 219716 175524
rect 219780 175460 219781 175524
rect 219715 175459 219781 175460
rect 182915 174980 182981 174981
rect 182915 174916 182916 174980
rect 182980 174916 182981 174980
rect 182915 174915 182981 174916
rect 169299 172940 169365 172941
rect 169299 172876 169300 172940
rect 169364 172876 169365 172940
rect 169299 172875 169365 172876
rect 168747 172804 168813 172805
rect 168747 172740 168748 172804
rect 168812 172740 168813 172804
rect 168747 172739 168813 172740
rect 168750 164234 168810 172739
rect 168750 164174 169362 164234
rect 169302 143922 169362 164174
rect 148507 139892 148573 139893
rect 148507 139828 148508 139892
rect 148572 139828 148573 139892
rect 148507 139827 148573 139828
rect 148510 118082 148570 139827
rect 182918 131682 182978 174915
rect 197635 144652 197701 144653
rect 197635 144588 197636 144652
rect 197700 144588 197701 144652
rect 197635 144587 197701 144588
rect 197267 140572 197333 140573
rect 197267 140522 197268 140572
rect 197332 140522 197333 140572
rect 197638 132549 197698 144587
rect 203158 143293 203218 143686
rect 203155 143292 203221 143293
rect 203155 143228 203156 143292
rect 203220 143228 203221 143292
rect 203155 143227 203221 143228
rect 219718 142069 219778 175459
rect 241798 174029 241858 180083
rect 241795 174028 241861 174029
rect 241795 173964 241796 174028
rect 241860 173964 241861 174028
rect 241795 173963 241861 173964
rect 237379 169540 237445 169541
rect 237379 169476 237380 169540
rect 237444 169476 237445 169540
rect 237379 169475 237445 169476
rect 237382 166362 237442 169475
rect 242350 169269 242410 180219
rect 242531 180012 242597 180013
rect 242531 179948 242532 180012
rect 242596 179948 242597 180012
rect 242531 179947 242597 179948
rect 242534 175794 242594 179947
rect 242534 175734 242778 175794
rect 242531 174028 242597 174029
rect 242531 173964 242532 174028
rect 242596 173964 242597 174028
rect 242531 173963 242597 173964
rect 242534 169269 242594 173963
rect 238115 169268 238181 169269
rect 238115 169204 238116 169268
rect 238180 169204 238181 169268
rect 238115 169203 238181 169204
rect 242347 169268 242413 169269
rect 242347 169204 242348 169268
rect 242412 169204 242413 169268
rect 242347 169203 242413 169204
rect 242531 169268 242597 169269
rect 242531 169204 242532 169268
rect 242596 169204 242597 169268
rect 242531 169203 242597 169204
rect 237382 150722 237442 157286
rect 237750 148002 237810 168166
rect 238118 147322 238178 169203
rect 242718 168402 242778 175734
rect 243451 169540 243517 169541
rect 243451 169476 243452 169540
rect 243516 169476 243517 169540
rect 243451 169475 243517 169476
rect 243454 168402 243514 169475
rect 247131 169268 247197 169269
rect 247131 169204 247132 169268
rect 247196 169204 247197 169268
rect 247131 169203 247197 169204
rect 247134 168402 247194 169203
rect 231675 143292 231741 143293
rect 231675 143228 231676 143292
rect 231740 143228 231741 143292
rect 231675 143227 231741 143228
rect 219715 142068 219781 142069
rect 219715 142004 219716 142068
rect 219780 142004 219781 142068
rect 219715 142003 219781 142004
rect 231678 140522 231738 143227
rect 231678 140029 231738 140286
rect 231675 140028 231741 140029
rect 231675 139964 231676 140028
rect 231740 139964 231741 140028
rect 231675 139963 231741 139964
rect 238118 139757 238178 146406
rect 261670 144602 261730 180763
rect 262403 180692 262469 180693
rect 262403 180628 262404 180692
rect 262468 180628 262469 180692
rect 262403 180627 262469 180628
rect 242902 142477 242962 143006
rect 242899 142476 242965 142477
rect 242899 142412 242900 142476
rect 242964 142412 242965 142476
rect 242899 142411 242965 142412
rect 242534 142205 242594 142326
rect 242531 142204 242597 142205
rect 242531 142140 242532 142204
rect 242596 142140 242597 142204
rect 242531 142139 242597 142140
rect 246398 142069 246458 143006
rect 247318 142477 247378 143006
rect 247315 142476 247381 142477
rect 247315 142412 247316 142476
rect 247380 142412 247381 142476
rect 247315 142411 247381 142412
rect 255227 142476 255293 142477
rect 255227 142412 255228 142476
rect 255292 142412 255293 142476
rect 255227 142411 255293 142412
rect 246395 142068 246461 142069
rect 246395 142004 246396 142068
rect 246460 142004 246461 142068
rect 246395 142003 246461 142004
rect 255230 141882 255290 142411
rect 262406 140522 262466 180627
rect 262955 180556 263021 180557
rect 262955 180492 262956 180556
rect 263020 180492 263021 180556
rect 262955 180491 263021 180492
rect 262958 143242 263018 180491
rect 309875 179332 309941 179333
rect 309875 179282 309876 179332
rect 309940 179282 309941 179332
rect 312635 179332 312701 179333
rect 312635 179282 312636 179332
rect 312700 179282 312701 179332
rect 351646 172941 351706 184027
rect 351830 172941 351890 191374
rect 352747 191372 352748 191374
rect 352812 191372 352813 191436
rect 352747 191371 352813 191372
rect 351643 172940 351709 172941
rect 351643 172876 351644 172940
rect 351708 172876 351709 172940
rect 351643 172875 351709 172876
rect 351827 172940 351893 172941
rect 351827 172876 351828 172940
rect 351892 172876 351893 172940
rect 351827 172875 351893 172876
rect 435740 167628 439740 198028
rect 435740 167392 435862 167628
rect 436098 167392 436182 167628
rect 436418 167392 436502 167628
rect 436738 167392 436822 167628
rect 437058 167392 437142 167628
rect 437378 167392 437462 167628
rect 437698 167392 437782 167628
rect 438018 167392 438102 167628
rect 438338 167392 438422 167628
rect 438658 167392 438742 167628
rect 438978 167392 439062 167628
rect 439298 167392 439382 167628
rect 439618 167392 439740 167628
rect 292579 144652 292645 144653
rect 292579 144588 292580 144652
rect 292644 144588 292645 144652
rect 292579 144587 292645 144588
rect 238115 139756 238181 139757
rect 238115 139692 238116 139756
rect 238180 139692 238181 139756
rect 238115 139691 238181 139692
rect 245294 139621 245354 140286
rect 251366 139893 251426 140286
rect 251363 139892 251429 139893
rect 251363 139828 251364 139892
rect 251428 139828 251429 139892
rect 251363 139827 251429 139828
rect 262958 139621 263018 143006
rect 245291 139620 245357 139621
rect 245291 139556 245292 139620
rect 245356 139556 245357 139620
rect 245291 139555 245357 139556
rect 262955 139620 263021 139621
rect 262955 139556 262956 139620
rect 263020 139556 263021 139620
rect 262955 139555 263021 139556
rect 249155 137308 249221 137309
rect 249155 137244 249156 137308
rect 249220 137244 249221 137308
rect 249155 137243 249221 137244
rect 197635 132548 197701 132549
rect 197635 132484 197636 132548
rect 197700 132484 197701 132548
rect 197635 132483 197701 132484
rect 198555 132548 198621 132549
rect 198555 132484 198556 132548
rect 198620 132484 198621 132548
rect 198555 132483 198621 132484
rect 148691 122348 148757 122349
rect 148691 122284 148692 122348
rect 148756 122284 148757 122348
rect 148691 122283 148757 122284
rect 148694 122074 148754 122283
rect 148875 122212 148941 122213
rect 148875 122148 148876 122212
rect 148940 122148 148941 122212
rect 148875 122147 148941 122148
rect 148878 122074 148938 122147
rect 148694 122014 148938 122074
rect 178686 117861 178746 123966
rect 198558 121716 198618 132483
rect 246211 130236 246277 130237
rect 246211 130172 246212 130236
rect 246276 130172 246277 130236
rect 246211 130171 246277 130172
rect 242715 122556 242716 122606
rect 242780 122556 242781 122606
rect 242715 122555 242781 122556
rect 198464 121674 198784 121716
rect 198464 121438 198506 121674
rect 198742 121438 198784 121674
rect 198464 121396 198784 121438
rect 198558 120122 198618 121396
rect 177579 117860 177645 117861
rect 177579 117796 177580 117860
rect 177644 117796 177645 117860
rect 177579 117795 177645 117796
rect 178683 117860 178749 117861
rect 178683 117796 178684 117860
rect 178748 117796 178749 117860
rect 178683 117795 178749 117796
rect 147771 113644 147837 113645
rect 147771 113580 147772 113644
rect 147836 113580 147837 113644
rect 147771 113579 147837 113580
rect 78035 110924 78101 110925
rect 78035 110860 78036 110924
rect 78100 110860 78101 110924
rect 78035 110859 78101 110860
rect 84659 109636 84660 109686
rect 84724 109636 84725 109686
rect 84659 109635 84725 109636
rect 74539 109564 74605 109565
rect 74539 109500 74540 109564
rect 74604 109500 74605 109564
rect 74539 109499 74605 109500
rect 148694 109094 148938 109154
rect 148694 108885 148754 109094
rect 148878 108885 148938 109094
rect 148691 108884 148757 108885
rect 148691 108820 148692 108884
rect 148756 108820 148757 108884
rect 148691 108819 148757 108820
rect 148875 108884 148941 108885
rect 148875 108820 148876 108884
rect 148940 108820 148941 108884
rect 148875 108819 148941 108820
rect 89104 106356 89424 106398
rect 89104 106120 89146 106356
rect 89382 106120 89424 106356
rect 89104 106078 89424 106120
rect 74171 102084 74237 102085
rect 74171 102020 74172 102084
rect 74236 102020 74237 102084
rect 74171 102019 74237 102020
rect 73619 98276 73685 98277
rect 73619 98212 73620 98276
rect 73684 98212 73685 98276
rect 73619 98211 73685 98212
rect 148691 95556 148757 95557
rect 148691 95492 148692 95556
rect 148756 95554 148757 95556
rect 148875 95556 148941 95557
rect 148875 95554 148876 95556
rect 148756 95494 148876 95554
rect 148756 95492 148757 95494
rect 148691 95491 148757 95492
rect 148875 95492 148876 95494
rect 148940 95492 148941 95556
rect 148875 95491 148941 95492
rect 148507 95284 148573 95285
rect 148507 95220 148508 95284
rect 148572 95220 148573 95284
rect 148507 95219 148573 95220
rect 148510 94962 148570 95219
rect 104464 91038 104784 91080
rect 104464 90802 104506 91038
rect 104742 90802 104784 91038
rect 104464 90760 104784 90802
rect 152190 90117 152250 112406
rect 163782 96322 163842 115806
rect 177582 115005 177642 117795
rect 245478 116722 245538 123286
rect 228731 116500 228797 116501
rect 228731 116436 228732 116500
rect 228796 116436 228797 116500
rect 228731 116435 228797 116436
rect 228734 116042 228794 116435
rect 177579 115004 177645 115005
rect 177579 114940 177580 115004
rect 177644 114940 177645 115004
rect 177579 114939 177645 114940
rect 245478 113914 245538 116486
rect 245110 113854 245538 113914
rect 245110 113234 245170 113854
rect 245846 113322 245906 123966
rect 244742 113174 245170 113234
rect 230755 112964 230821 112965
rect 230755 112900 230756 112964
rect 230820 112900 230821 112964
rect 230755 112899 230821 112900
rect 230758 112642 230818 112899
rect 230939 107388 231005 107389
rect 230939 107324 230940 107388
rect 231004 107324 231005 107388
rect 230939 107323 231005 107324
rect 230942 107202 231002 107323
rect 164886 100725 164946 106966
rect 228731 106844 228797 106845
rect 228731 106780 228732 106844
rect 228796 106780 228797 106844
rect 228731 106779 228797 106780
rect 183104 106356 183424 106398
rect 183104 106120 183146 106356
rect 183382 106120 183424 106356
rect 183104 106078 183424 106120
rect 177763 105484 177829 105485
rect 177763 105420 177764 105484
rect 177828 105420 177829 105484
rect 177763 105419 177829 105420
rect 164883 100724 164949 100725
rect 164883 100660 164884 100724
rect 164948 100660 164949 100724
rect 164883 100659 164949 100660
rect 177766 100314 177826 105419
rect 228734 102442 228794 106779
rect 242166 105485 242226 109686
rect 242163 105484 242229 105485
rect 242163 105420 242164 105484
rect 242228 105420 242229 105484
rect 242163 105419 242229 105420
rect 242531 105484 242597 105485
rect 242531 105420 242532 105484
rect 242596 105420 242597 105484
rect 242531 105419 242597 105420
rect 178134 100725 178194 100846
rect 228731 100796 228732 100846
rect 228796 100796 228797 100846
rect 228731 100795 228797 100796
rect 178131 100724 178197 100725
rect 178131 100660 178132 100724
rect 178196 100660 178197 100724
rect 178131 100659 178197 100660
rect 177766 100254 178194 100314
rect 178134 96322 178194 100254
rect 242534 95554 242594 105419
rect 244190 96322 244250 112406
rect 244742 99042 244802 113174
rect 246214 99634 246274 130171
rect 249158 127602 249218 137243
rect 249707 133092 249773 133093
rect 249707 133028 249708 133092
rect 249772 133028 249773 133092
rect 249707 133027 249773 133028
rect 249710 126837 249770 133027
rect 292582 131682 292642 144587
rect 351643 139620 351709 139621
rect 351643 139556 351644 139620
rect 351708 139556 351709 139620
rect 351643 139555 351709 139556
rect 351827 139620 351893 139621
rect 351827 139556 351828 139620
rect 351892 139556 351893 139620
rect 351827 139555 351893 139556
rect 249707 126836 249773 126837
rect 249707 126772 249708 126836
rect 249772 126772 249773 126836
rect 249707 126771 249773 126772
rect 258723 122556 258724 122606
rect 258788 122556 258789 122606
rect 258723 122555 258789 122556
rect 272707 122556 272708 122606
rect 272772 122556 272773 122606
rect 272707 122555 272773 122556
rect 292464 121674 292784 121716
rect 292464 121438 292506 121674
rect 292742 121438 292784 121674
rect 292464 121396 292784 121438
rect 258910 100725 258970 106966
rect 277104 106356 277424 106398
rect 277104 106120 277146 106356
rect 277382 106120 277424 106356
rect 277104 106078 277424 106120
rect 272710 100725 272770 100846
rect 258907 100724 258973 100725
rect 258907 100660 258908 100724
rect 258972 100660 258973 100724
rect 258907 100659 258973 100660
rect 272707 100724 272773 100725
rect 272707 100660 272708 100724
rect 272772 100660 272773 100724
rect 272707 100659 272773 100660
rect 322755 100452 322821 100453
rect 322755 100402 322756 100452
rect 322820 100402 322821 100452
rect 264427 100316 264493 100317
rect 264427 100252 264428 100316
rect 264492 100252 264493 100316
rect 264427 100251 264493 100252
rect 245662 99574 246274 99634
rect 245662 96914 245722 99574
rect 264430 99042 264490 100251
rect 245110 96854 245722 96914
rect 242534 95494 242962 95554
rect 242531 95420 242597 95421
rect 152187 90116 152253 90117
rect 152187 90052 152188 90116
rect 152252 90052 152253 90116
rect 152187 90051 152253 90052
rect 155315 90116 155381 90117
rect 155315 90052 155316 90116
rect 155380 90052 155381 90116
rect 155315 90051 155381 90052
rect 155318 89165 155378 90051
rect 155315 89164 155381 89165
rect 155315 89100 155316 89164
rect 155380 89100 155381 89164
rect 155315 89099 155381 89100
rect 72515 88348 72581 88349
rect 72515 88284 72516 88348
rect 72580 88284 72581 88348
rect 72515 88283 72581 88284
rect 54667 79100 54733 79101
rect 54667 79036 54668 79100
rect 54732 79036 54733 79100
rect 54667 79035 54733 79036
rect 55403 79100 55469 79101
rect 55403 79036 55404 79100
rect 55468 79036 55469 79100
rect 55403 79035 55469 79036
rect 54115 78964 54181 78965
rect 54115 78900 54116 78964
rect 54180 78900 54181 78964
rect 54115 78899 54181 78900
rect 5000 75484 5122 75720
rect 5358 75484 5442 75720
rect 5678 75484 5762 75720
rect 5998 75484 6082 75720
rect 6318 75484 6402 75720
rect 6638 75484 6722 75720
rect 6958 75484 7042 75720
rect 7278 75484 7362 75720
rect 7598 75484 7682 75720
rect 7918 75484 8002 75720
rect 8238 75484 8322 75720
rect 8558 75484 8642 75720
rect 8878 75484 9000 75720
rect 5000 45084 9000 75484
rect 72518 73882 72578 88283
rect 148507 87124 148573 87125
rect 148507 87060 148508 87124
rect 148572 87060 148573 87124
rect 148507 87059 148573 87060
rect 73987 86444 74053 86445
rect 73987 86380 73988 86444
rect 74052 86380 74053 86444
rect 73987 86379 74053 86380
rect 73251 86308 73317 86309
rect 73251 86244 73252 86308
rect 73316 86244 73317 86308
rect 73251 86243 73317 86244
rect 72699 86172 72765 86173
rect 72699 86108 72700 86172
rect 72764 86108 72765 86172
rect 72699 86107 72765 86108
rect 72702 85901 72762 86107
rect 72699 85900 72765 85901
rect 72699 85836 72700 85900
rect 72764 85836 72765 85900
rect 72699 85835 72765 85836
rect 73067 76516 73133 76517
rect 73067 76452 73068 76516
rect 73132 76452 73133 76516
rect 73067 76451 73133 76452
rect 73070 76381 73130 76451
rect 73067 76380 73133 76381
rect 73067 76316 73068 76380
rect 73132 76316 73133 76380
rect 73067 76315 73133 76316
rect 73067 76108 73133 76109
rect 73067 76044 73068 76108
rect 73132 76044 73133 76108
rect 73067 76043 73133 76044
rect 73070 73794 73130 76043
rect 73254 75429 73314 86243
rect 73251 75428 73317 75429
rect 73251 75364 73252 75428
rect 73316 75364 73317 75428
rect 73251 75363 73317 75364
rect 73803 75428 73869 75429
rect 73803 75364 73804 75428
rect 73868 75364 73869 75428
rect 73803 75363 73869 75364
rect 73070 73734 73498 73794
rect 73438 61642 73498 73734
rect 73806 60194 73866 75363
rect 73438 60134 73866 60194
rect 73438 49402 73498 60134
rect 73990 59602 74050 86379
rect 74355 86172 74421 86173
rect 74355 86108 74356 86172
rect 74420 86108 74421 86172
rect 74355 86107 74421 86108
rect 74358 57474 74418 86107
rect 148510 73882 148570 87059
rect 155318 75565 155378 89099
rect 163782 87397 163842 95406
rect 164883 95284 164949 95285
rect 164883 95220 164884 95284
rect 164948 95220 164949 95284
rect 164883 95219 164949 95220
rect 164886 93602 164946 95219
rect 178134 94194 178194 95406
rect 242531 95356 242532 95420
rect 242596 95356 242597 95420
rect 242531 95355 242597 95356
rect 178683 95284 178749 95285
rect 178683 95220 178684 95284
rect 178748 95220 178749 95284
rect 178683 95219 178749 95220
rect 178686 94962 178746 95219
rect 242534 94962 242594 95355
rect 178134 94134 178746 94194
rect 163779 87396 163845 87397
rect 163779 87332 163780 87396
rect 163844 87332 163845 87396
rect 163779 87331 163845 87332
rect 167643 87396 167709 87397
rect 167643 87332 167644 87396
rect 167708 87332 167709 87396
rect 167643 87331 167709 87332
rect 155315 75564 155381 75565
rect 155315 75500 155316 75564
rect 155380 75500 155381 75564
rect 155315 75499 155381 75500
rect 74726 62914 74786 68886
rect 74726 62854 75706 62914
rect 73990 57414 74418 57474
rect 74542 61494 75006 61554
rect 73990 56114 74050 57414
rect 73990 56054 74418 56114
rect 74358 51354 74418 56054
rect 74542 52034 74602 61494
rect 75646 60194 75706 62854
rect 74726 60134 75706 60194
rect 74726 53394 74786 60134
rect 74726 53334 75338 53394
rect 74542 51974 75154 52034
rect 74358 51294 74602 51354
rect 72886 49254 73350 49314
rect 72515 47956 72581 47957
rect 72515 47892 72516 47956
rect 72580 47892 72581 47956
rect 72886 47954 72946 49254
rect 74542 48722 74602 51294
rect 73254 48093 73314 48486
rect 75094 48093 75154 51974
rect 73251 48092 73317 48093
rect 73251 48028 73252 48092
rect 73316 48028 73317 48092
rect 73251 48027 73317 48028
rect 75091 48092 75157 48093
rect 75091 48028 75092 48092
rect 75156 48028 75157 48092
rect 75091 48027 75157 48028
rect 75278 47957 75338 53334
rect 75275 47956 75341 47957
rect 72886 47894 73314 47954
rect 72515 47891 72581 47892
rect 72518 47413 72578 47891
rect 72515 47412 72581 47413
rect 72515 47348 72516 47412
rect 72580 47348 72581 47412
rect 72515 47347 72581 47348
rect 73254 45917 73314 47894
rect 75275 47892 75276 47956
rect 75340 47892 75341 47956
rect 75275 47891 75341 47892
rect 75462 47549 75522 59366
rect 144830 54842 144890 63446
rect 78958 52853 79018 53246
rect 78955 52852 79021 52853
rect 78955 52788 78956 52852
rect 79020 52788 79021 52852
rect 78955 52787 79021 52788
rect 107475 50268 107541 50269
rect 107475 50204 107476 50268
rect 107540 50204 107541 50268
rect 107475 50203 107541 50204
rect 109315 50268 109381 50269
rect 109315 50204 109316 50268
rect 109380 50204 109381 50268
rect 109315 50203 109381 50204
rect 87238 48093 87298 48486
rect 87235 48092 87301 48093
rect 87235 48028 87236 48092
rect 87300 48028 87301 48092
rect 87235 48027 87301 48028
rect 74171 47548 74237 47549
rect 74171 47484 74172 47548
rect 74236 47484 74237 47548
rect 74171 47483 74237 47484
rect 75459 47548 75525 47549
rect 75459 47484 75460 47548
rect 75524 47484 75525 47548
rect 75459 47483 75525 47484
rect 74174 47413 74234 47483
rect 107478 47413 107538 50203
rect 74171 47412 74237 47413
rect 74171 47348 74172 47412
rect 74236 47348 74237 47412
rect 74171 47347 74237 47348
rect 107475 47412 107541 47413
rect 107475 47348 107476 47412
rect 107540 47348 107541 47412
rect 107475 47347 107541 47348
rect 107478 46682 107538 47347
rect 109318 47277 109378 50203
rect 113550 47549 113610 53246
rect 118147 53124 118213 53125
rect 118147 53060 118148 53124
rect 118212 53060 118213 53124
rect 118147 53059 118213 53060
rect 113547 47548 113613 47549
rect 113547 47484 113548 47548
rect 113612 47484 113613 47548
rect 113547 47483 113613 47484
rect 109315 47276 109381 47277
rect 109315 47212 109316 47276
rect 109380 47212 109381 47276
rect 109315 47211 109381 47212
rect 73251 45916 73317 45917
rect 73251 45852 73252 45916
rect 73316 45852 73317 45916
rect 73251 45851 73317 45852
rect 5000 44848 5122 45084
rect 5358 44848 5442 45084
rect 5678 44848 5762 45084
rect 5998 44848 6082 45084
rect 6318 44848 6402 45084
rect 6638 44848 6722 45084
rect 6958 44848 7042 45084
rect 7278 44848 7362 45084
rect 7598 44848 7682 45084
rect 7918 44848 8002 45084
rect 8238 44848 8322 45084
rect 8558 44848 8642 45084
rect 8878 44848 9000 45084
rect 5000 14448 9000 44848
rect 118150 44693 118210 53059
rect 134158 51765 134218 53246
rect 134155 51764 134221 51765
rect 134155 51700 134156 51764
rect 134220 51700 134221 51764
rect 134155 51699 134221 51700
rect 142806 51085 142866 51206
rect 142803 51084 142869 51085
rect 142803 51020 142804 51084
rect 142868 51020 142869 51084
rect 142803 51019 142869 51020
rect 144830 49402 144890 53926
rect 144830 47957 144890 49166
rect 147958 48093 148018 49166
rect 167646 48722 167706 87331
rect 168747 87124 168813 87125
rect 168747 87060 168748 87124
rect 168812 87060 168813 87124
rect 168747 87059 168813 87060
rect 168011 86852 168077 86853
rect 168011 86788 168012 86852
rect 168076 86788 168077 86852
rect 168011 86787 168077 86788
rect 168014 49402 168074 86787
rect 154766 48093 154826 48486
rect 168014 48093 168074 49166
rect 147955 48092 148021 48093
rect 147955 48028 147956 48092
rect 148020 48028 148021 48092
rect 147955 48027 148021 48028
rect 154763 48092 154829 48093
rect 154763 48028 154764 48092
rect 154828 48028 154829 48092
rect 168011 48092 168077 48093
rect 154763 48027 154829 48028
rect 144827 47956 144893 47957
rect 144827 47892 144828 47956
rect 144892 47892 144893 47956
rect 144827 47891 144893 47892
rect 147771 47956 147837 47957
rect 147771 47892 147772 47956
rect 147836 47954 147837 47956
rect 168011 48028 168012 48092
rect 168076 48028 168077 48092
rect 168011 48027 168077 48028
rect 168750 47957 168810 87059
rect 169299 86988 169365 86989
rect 169299 86924 169300 86988
rect 169364 86924 169365 86988
rect 169299 86923 169365 86924
rect 169115 86716 169181 86717
rect 169115 86652 169116 86716
rect 169180 86652 169181 86716
rect 169115 86651 169181 86652
rect 169118 48042 169178 86651
rect 169302 48634 169362 86923
rect 178686 86802 178746 94134
rect 242902 93514 242962 95494
rect 242534 93454 242962 93514
rect 198464 91038 198784 91080
rect 198464 90802 198506 91038
rect 198742 90802 198784 91038
rect 198464 90760 198784 90802
rect 242534 86037 242594 93454
rect 245110 88162 245170 96854
rect 245846 89165 245906 96086
rect 246214 90117 246274 98806
rect 258726 95285 258786 95406
rect 272710 95285 272770 95406
rect 258723 95284 258789 95285
rect 258723 95220 258724 95284
rect 258788 95220 258789 95284
rect 258723 95219 258789 95220
rect 272707 95284 272773 95285
rect 272707 95220 272708 95284
rect 272772 95220 272773 95284
rect 272707 95219 272773 95220
rect 322755 94468 322821 94469
rect 322755 94404 322756 94468
rect 322820 94404 322821 94468
rect 322755 94403 322821 94404
rect 322758 94282 322818 94403
rect 292464 91038 292784 91080
rect 292464 90802 292506 91038
rect 292742 90802 292784 91038
rect 292464 90760 292784 90802
rect 351646 90117 351706 139555
rect 351830 117314 351890 139555
rect 435740 136992 439740 167392
rect 435740 136756 435862 136992
rect 436098 136756 436182 136992
rect 436418 136756 436502 136992
rect 436738 136756 436822 136992
rect 437058 136756 437142 136992
rect 437378 136756 437462 136992
rect 437698 136756 437782 136992
rect 438018 136756 438102 136992
rect 438338 136756 438422 136992
rect 438658 136756 438742 136992
rect 438978 136756 439062 136992
rect 439298 136756 439382 136992
rect 439618 136756 439740 136992
rect 351830 117254 352810 117314
rect 352750 105213 352810 117254
rect 435740 106356 439740 136756
rect 435740 106120 435862 106356
rect 436098 106120 436182 106356
rect 436418 106120 436502 106356
rect 436738 106120 436822 106356
rect 437058 106120 437142 106356
rect 437378 106120 437462 106356
rect 437698 106120 437782 106356
rect 438018 106120 438102 106356
rect 438338 106120 438422 106356
rect 438658 106120 438742 106356
rect 438978 106120 439062 106356
rect 439298 106120 439382 106356
rect 439618 106120 439740 106356
rect 352747 105212 352813 105213
rect 352747 105148 352748 105212
rect 352812 105148 352813 105212
rect 352747 105147 352813 105148
rect 352747 97596 352813 97597
rect 352747 97594 352748 97596
rect 352566 97534 352748 97594
rect 352566 96234 352626 97534
rect 352747 97532 352748 97534
rect 352812 97532 352813 97596
rect 352747 97531 352813 97532
rect 352014 96174 352626 96234
rect 246211 90116 246277 90117
rect 246211 90052 246212 90116
rect 246276 90052 246277 90116
rect 246211 90051 246277 90052
rect 249155 90116 249221 90117
rect 249155 90052 249156 90116
rect 249220 90052 249221 90116
rect 249155 90051 249221 90052
rect 351643 90116 351709 90117
rect 351643 90052 351644 90116
rect 351708 90052 351709 90116
rect 351643 90051 351709 90052
rect 245843 89164 245909 89165
rect 245843 89100 245844 89164
rect 245908 89100 245909 89164
rect 245843 89099 245909 89100
rect 249158 88893 249218 90051
rect 249155 88892 249221 88893
rect 249155 88842 249156 88892
rect 249220 88842 249221 88892
rect 249155 88484 249221 88485
rect 249155 88420 249156 88484
rect 249220 88420 249221 88484
rect 249155 88419 249221 88420
rect 242531 86036 242597 86037
rect 242531 85972 242532 86036
rect 242596 85972 242597 86036
rect 242531 85971 242597 85972
rect 182550 83725 182610 85206
rect 182547 83724 182613 83725
rect 182547 83660 182548 83724
rect 182612 83660 182613 83724
rect 182547 83659 182613 83660
rect 242715 76516 242781 76517
rect 242715 76452 242716 76516
rect 242780 76452 242781 76516
rect 242715 76451 242781 76452
rect 242718 73882 242778 76451
rect 249158 75565 249218 88419
rect 261667 87532 261733 87533
rect 261667 87468 261668 87532
rect 261732 87468 261733 87532
rect 261667 87467 261733 87468
rect 252651 86172 252717 86173
rect 252651 86108 252652 86172
rect 252716 86108 252717 86172
rect 252651 86107 252717 86108
rect 249155 75564 249221 75565
rect 249155 75500 249156 75564
rect 249220 75500 249221 75564
rect 249155 75499 249221 75500
rect 252654 75429 252714 86107
rect 252651 75428 252717 75429
rect 252651 75364 252652 75428
rect 252716 75364 252717 75428
rect 252651 75363 252717 75364
rect 237382 59602 237442 68886
rect 173902 52445 173962 53246
rect 173899 52444 173965 52445
rect 173899 52380 173900 52444
rect 173964 52380 173965 52444
rect 173899 52379 173965 52380
rect 191379 50404 191445 50405
rect 191379 50340 191380 50404
rect 191444 50340 191445 50404
rect 191379 50339 191445 50340
rect 191382 48722 191442 50339
rect 199659 50268 199725 50269
rect 199659 50204 199660 50268
rect 199724 50204 199725 50268
rect 199659 50203 199725 50204
rect 169302 48574 169730 48634
rect 147836 47894 148018 47954
rect 147836 47892 147837 47894
rect 147771 47891 147837 47892
rect 147958 45781 148018 47894
rect 168747 47956 168813 47957
rect 168747 47892 168748 47956
rect 168812 47892 168813 47956
rect 168747 47891 168813 47892
rect 169670 47821 169730 48574
rect 169667 47820 169733 47821
rect 169667 47756 169668 47820
rect 169732 47756 169733 47820
rect 169667 47755 169733 47756
rect 157526 45917 157586 46446
rect 158998 46053 159058 47126
rect 158995 46052 159061 46053
rect 158995 45988 158996 46052
rect 159060 45988 159061 46052
rect 158995 45987 159061 45988
rect 157523 45916 157589 45917
rect 157523 45852 157524 45916
rect 157588 45852 157589 45916
rect 157523 45851 157589 45852
rect 147955 45780 148021 45781
rect 147955 45716 147956 45780
rect 148020 45716 148021 45780
rect 147955 45715 148021 45716
rect 169670 44829 169730 47755
rect 199662 46682 199722 50203
rect 169667 44828 169733 44829
rect 169667 44764 169668 44828
rect 169732 44764 169733 44828
rect 169667 44763 169733 44764
rect 118147 44692 118213 44693
rect 118147 44628 118148 44692
rect 118212 44628 118213 44692
rect 118147 44627 118213 44628
rect 207758 39117 207818 53246
rect 211987 53124 212053 53125
rect 211987 53060 211988 53124
rect 212052 53060 212053 53124
rect 211987 53059 212053 53060
rect 211990 43469 212050 53059
rect 227998 51765 228058 53246
rect 227995 51764 228061 51765
rect 227995 51700 227996 51764
rect 228060 51700 228061 51764
rect 227995 51699 228061 51700
rect 238302 50762 238362 59366
rect 237566 48093 237626 50526
rect 261670 49314 261730 87467
rect 262771 86988 262837 86989
rect 262771 86924 262772 86988
rect 262836 86924 262837 86988
rect 262771 86923 262837 86924
rect 261851 75428 261917 75429
rect 261851 75364 261852 75428
rect 261916 75364 261917 75428
rect 261851 75363 261917 75364
rect 261486 49254 261730 49314
rect 237563 48092 237629 48093
rect 237563 48028 237564 48092
rect 237628 48028 237629 48092
rect 237563 48027 237629 48028
rect 248606 47957 248666 48486
rect 261486 48042 261546 49254
rect 248603 47956 248669 47957
rect 248603 47892 248604 47956
rect 248668 47892 248669 47956
rect 248603 47891 248669 47892
rect 261854 46682 261914 75363
rect 262774 49314 262834 86923
rect 263507 86852 263573 86853
rect 263507 86788 263508 86852
rect 263572 86788 263573 86852
rect 263507 86787 263573 86788
rect 263139 86716 263205 86717
rect 263139 86652 263140 86716
rect 263204 86652 263205 86716
rect 263139 86651 263205 86652
rect 263142 51354 263202 86651
rect 263142 51294 263386 51354
rect 263326 50082 263386 51294
rect 263510 50674 263570 86787
rect 263510 50614 263754 50674
rect 262554 49254 262834 49314
rect 262406 48093 262466 49166
rect 262403 48092 262469 48093
rect 262403 48028 262404 48092
rect 262468 48028 262469 48092
rect 262403 48027 262469 48028
rect 252654 46053 252714 46446
rect 252651 46052 252717 46053
rect 252651 45988 252652 46052
rect 252716 45988 252717 46052
rect 252651 45987 252717 45988
rect 263326 45781 263386 49846
rect 263694 49314 263754 50614
rect 263878 49994 263938 88606
rect 351646 77877 351706 90051
rect 352014 79234 352074 96174
rect 356795 87396 356861 87397
rect 356795 87332 356796 87396
rect 356860 87332 356861 87396
rect 356795 87331 356861 87332
rect 351830 79174 352074 79234
rect 351830 77877 351890 79174
rect 351643 77876 351709 77877
rect 351643 77812 351644 77876
rect 351708 77812 351709 77876
rect 351643 77811 351709 77812
rect 351827 77876 351893 77877
rect 351827 77812 351828 77876
rect 351892 77812 351893 77876
rect 351827 77811 351893 77812
rect 307115 53396 307181 53397
rect 307115 53332 307116 53396
rect 307180 53332 307181 53396
rect 307115 53331 307181 53332
rect 266638 52445 266698 53246
rect 266635 52444 266701 52445
rect 266635 52380 266636 52444
rect 266700 52380 266701 52444
rect 266635 52379 266701 52380
rect 263878 49934 264490 49994
rect 263510 49254 263754 49314
rect 263510 46053 263570 49254
rect 263878 48093 263938 48486
rect 263875 48092 263941 48093
rect 263875 48028 263876 48092
rect 263940 48028 263941 48092
rect 263875 48027 263941 48028
rect 264430 47413 264490 49934
rect 263875 47412 263941 47413
rect 263875 47362 263876 47412
rect 263940 47362 263941 47412
rect 264427 47412 264493 47413
rect 264427 47348 264428 47412
rect 264492 47348 264493 47412
rect 264427 47347 264493 47348
rect 263507 46052 263573 46053
rect 263507 45988 263508 46052
rect 263572 45988 263573 46052
rect 263507 45987 263573 45988
rect 263323 45780 263389 45781
rect 263323 45716 263324 45780
rect 263388 45716 263389 45780
rect 263323 45715 263389 45716
rect 211987 43468 212053 43469
rect 211987 43404 211988 43468
rect 212052 43404 212053 43468
rect 211987 43403 212053 43404
rect 301598 39117 301658 53246
rect 207755 39116 207821 39117
rect 207755 39052 207756 39116
rect 207820 39052 207821 39116
rect 207755 39051 207821 39052
rect 301595 39116 301661 39117
rect 301595 39052 301596 39116
rect 301660 39052 301661 39116
rect 301595 39051 301661 39052
rect 307118 37757 307178 53331
rect 321838 51765 321898 53246
rect 321835 51764 321901 51765
rect 321835 51700 321836 51764
rect 321900 51700 321901 51764
rect 321835 51699 321901 51700
rect 330851 49996 330917 49997
rect 330851 49932 330852 49996
rect 330916 49994 330917 49996
rect 330916 49934 331466 49994
rect 330916 49932 330917 49934
rect 330851 49931 330917 49932
rect 331406 45373 331466 49934
rect 356798 46053 356858 87331
rect 435740 75720 439740 106120
rect 435740 75484 435862 75720
rect 436098 75484 436182 75720
rect 436418 75484 436502 75720
rect 436738 75484 436822 75720
rect 437058 75484 437142 75720
rect 437378 75484 437462 75720
rect 437698 75484 437782 75720
rect 438018 75484 438102 75720
rect 438338 75484 438422 75720
rect 438658 75484 438742 75720
rect 438978 75484 439062 75720
rect 439298 75484 439382 75720
rect 439618 75484 439740 75720
rect 356795 46052 356861 46053
rect 356795 45988 356796 46052
rect 356860 45988 356861 46052
rect 356795 45987 356861 45988
rect 331403 45372 331469 45373
rect 331403 45308 331404 45372
rect 331468 45308 331469 45372
rect 331403 45307 331469 45308
rect 435740 45084 439740 75484
rect 435740 44848 435862 45084
rect 436098 44848 436182 45084
rect 436418 44848 436502 45084
rect 436738 44848 436822 45084
rect 437058 44848 437142 45084
rect 437378 44848 437462 45084
rect 437698 44848 437782 45084
rect 438018 44848 438102 45084
rect 438338 44848 438422 45084
rect 438658 44848 438742 45084
rect 438978 44848 439062 45084
rect 439298 44848 439382 45084
rect 439618 44848 439740 45084
rect 307115 37756 307181 37757
rect 307115 37692 307116 37756
rect 307180 37692 307181 37756
rect 307115 37691 307181 37692
rect 5000 14212 5122 14448
rect 5358 14212 5442 14448
rect 5678 14212 5762 14448
rect 5998 14212 6082 14448
rect 6318 14212 6402 14448
rect 6638 14212 6722 14448
rect 6958 14212 7042 14448
rect 7278 14212 7362 14448
rect 7598 14212 7682 14448
rect 7918 14212 8002 14448
rect 8238 14212 8322 14448
rect 8558 14212 8642 14448
rect 8878 14212 9000 14448
rect 5000 8878 9000 14212
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 435740 14448 439740 44848
rect 435740 14212 435862 14448
rect 436098 14212 436182 14448
rect 436418 14212 436502 14448
rect 436738 14212 436822 14448
rect 437058 14212 437142 14448
rect 437378 14212 437462 14448
rect 437698 14212 437782 14448
rect 438018 14212 438102 14448
rect 438338 14212 438422 14448
rect 438658 14212 438742 14448
rect 438978 14212 439062 14448
rect 439298 14212 439382 14448
rect 439618 14212 439740 14448
rect 435740 8878 439740 14212
rect 435740 8642 435862 8878
rect 436098 8642 436182 8878
rect 436418 8642 436502 8878
rect 436738 8642 436822 8878
rect 437058 8642 437142 8878
rect 437378 8642 437462 8878
rect 437698 8642 437782 8878
rect 438018 8642 438102 8878
rect 438338 8642 438422 8878
rect 438658 8642 438742 8878
rect 438978 8642 439062 8878
rect 439298 8642 439382 8878
rect 439618 8642 439740 8878
rect 435740 8558 439740 8642
rect 435740 8322 435862 8558
rect 436098 8322 436182 8558
rect 436418 8322 436502 8558
rect 436738 8322 436822 8558
rect 437058 8322 437142 8558
rect 437378 8322 437462 8558
rect 437698 8322 437782 8558
rect 438018 8322 438102 8558
rect 438338 8322 438422 8558
rect 438658 8322 438742 8558
rect 438978 8322 439062 8558
rect 439298 8322 439382 8558
rect 439618 8322 439740 8558
rect 435740 8238 439740 8322
rect 435740 8002 435862 8238
rect 436098 8002 436182 8238
rect 436418 8002 436502 8238
rect 436738 8002 436822 8238
rect 437058 8002 437142 8238
rect 437378 8002 437462 8238
rect 437698 8002 437782 8238
rect 438018 8002 438102 8238
rect 438338 8002 438422 8238
rect 438658 8002 438742 8238
rect 438978 8002 439062 8238
rect 439298 8002 439382 8238
rect 439618 8002 439740 8238
rect 435740 7918 439740 8002
rect 435740 7682 435862 7918
rect 436098 7682 436182 7918
rect 436418 7682 436502 7918
rect 436738 7682 436822 7918
rect 437058 7682 437142 7918
rect 437378 7682 437462 7918
rect 437698 7682 437782 7918
rect 438018 7682 438102 7918
rect 438338 7682 438422 7918
rect 438658 7682 438742 7918
rect 438978 7682 439062 7918
rect 439298 7682 439382 7918
rect 439618 7682 439740 7918
rect 435740 7598 439740 7682
rect 435740 7362 435862 7598
rect 436098 7362 436182 7598
rect 436418 7362 436502 7598
rect 436738 7362 436822 7598
rect 437058 7362 437142 7598
rect 437378 7362 437462 7598
rect 437698 7362 437782 7598
rect 438018 7362 438102 7598
rect 438338 7362 438422 7598
rect 438658 7362 438742 7598
rect 438978 7362 439062 7598
rect 439298 7362 439382 7598
rect 439618 7362 439740 7598
rect 435740 7278 439740 7362
rect 435740 7042 435862 7278
rect 436098 7042 436182 7278
rect 436418 7042 436502 7278
rect 436738 7042 436822 7278
rect 437058 7042 437142 7278
rect 437378 7042 437462 7278
rect 437698 7042 437782 7278
rect 438018 7042 438102 7278
rect 438338 7042 438422 7278
rect 438658 7042 438742 7278
rect 438978 7042 439062 7278
rect 439298 7042 439382 7278
rect 439618 7042 439740 7278
rect 435740 6958 439740 7042
rect 435740 6722 435862 6958
rect 436098 6722 436182 6958
rect 436418 6722 436502 6958
rect 436738 6722 436822 6958
rect 437058 6722 437142 6958
rect 437378 6722 437462 6958
rect 437698 6722 437782 6958
rect 438018 6722 438102 6958
rect 438338 6722 438422 6958
rect 438658 6722 438742 6958
rect 438978 6722 439062 6958
rect 439298 6722 439382 6958
rect 439618 6722 439740 6958
rect 435740 6638 439740 6722
rect 435740 6402 435862 6638
rect 436098 6402 436182 6638
rect 436418 6402 436502 6638
rect 436738 6402 436822 6638
rect 437058 6402 437142 6638
rect 437378 6402 437462 6638
rect 437698 6402 437782 6638
rect 438018 6402 438102 6638
rect 438338 6402 438422 6638
rect 438658 6402 438742 6638
rect 438978 6402 439062 6638
rect 439298 6402 439382 6638
rect 439618 6402 439740 6638
rect 435740 6318 439740 6402
rect 435740 6082 435862 6318
rect 436098 6082 436182 6318
rect 436418 6082 436502 6318
rect 436738 6082 436822 6318
rect 437058 6082 437142 6318
rect 437378 6082 437462 6318
rect 437698 6082 437782 6318
rect 438018 6082 438102 6318
rect 438338 6082 438422 6318
rect 438658 6082 438742 6318
rect 438978 6082 439062 6318
rect 439298 6082 439382 6318
rect 439618 6082 439740 6318
rect 435740 5998 439740 6082
rect 435740 5762 435862 5998
rect 436098 5762 436182 5998
rect 436418 5762 436502 5998
rect 436738 5762 436822 5998
rect 437058 5762 437142 5998
rect 437378 5762 437462 5998
rect 437698 5762 437782 5998
rect 438018 5762 438102 5998
rect 438338 5762 438422 5998
rect 438658 5762 438742 5998
rect 438978 5762 439062 5998
rect 439298 5762 439382 5998
rect 439618 5762 439740 5998
rect 435740 5678 439740 5762
rect 435740 5442 435862 5678
rect 436098 5442 436182 5678
rect 436418 5442 436502 5678
rect 436738 5442 436822 5678
rect 437058 5442 437142 5678
rect 437378 5442 437462 5678
rect 437698 5442 437782 5678
rect 438018 5442 438102 5678
rect 438338 5442 438422 5678
rect 438658 5442 438742 5678
rect 438978 5442 439062 5678
rect 439298 5442 439382 5678
rect 439618 5442 439740 5678
rect 435740 5358 439740 5442
rect 435740 5122 435862 5358
rect 436098 5122 436182 5358
rect 436418 5122 436502 5358
rect 436738 5122 436822 5358
rect 437058 5122 437142 5358
rect 437378 5122 437462 5358
rect 437698 5122 437782 5358
rect 438018 5122 438102 5358
rect 438338 5122 438422 5358
rect 438658 5122 438742 5358
rect 438978 5122 439062 5358
rect 439298 5122 439382 5358
rect 439618 5122 439740 5358
rect 435740 5000 439740 5122
rect 440740 366762 444740 401642
rect 440740 366526 440862 366762
rect 441098 366526 441182 366762
rect 441418 366526 441502 366762
rect 441738 366526 441822 366762
rect 442058 366526 442142 366762
rect 442378 366526 442462 366762
rect 442698 366526 442782 366762
rect 443018 366526 443102 366762
rect 443338 366526 443422 366762
rect 443658 366526 443742 366762
rect 443978 366526 444062 366762
rect 444298 366526 444382 366762
rect 444618 366526 444740 366762
rect 440740 336126 444740 366526
rect 440740 335890 440862 336126
rect 441098 335890 441182 336126
rect 441418 335890 441502 336126
rect 441738 335890 441822 336126
rect 442058 335890 442142 336126
rect 442378 335890 442462 336126
rect 442698 335890 442782 336126
rect 443018 335890 443102 336126
rect 443338 335890 443422 336126
rect 443658 335890 443742 336126
rect 443978 335890 444062 336126
rect 444298 335890 444382 336126
rect 444618 335890 444740 336126
rect 440740 305490 444740 335890
rect 440740 305254 440862 305490
rect 441098 305254 441182 305490
rect 441418 305254 441502 305490
rect 441738 305254 441822 305490
rect 442058 305254 442142 305490
rect 442378 305254 442462 305490
rect 442698 305254 442782 305490
rect 443018 305254 443102 305490
rect 443338 305254 443422 305490
rect 443658 305254 443742 305490
rect 443978 305254 444062 305490
rect 444298 305254 444382 305490
rect 444618 305254 444740 305490
rect 440740 274854 444740 305254
rect 440740 274618 440862 274854
rect 441098 274618 441182 274854
rect 441418 274618 441502 274854
rect 441738 274618 441822 274854
rect 442058 274618 442142 274854
rect 442378 274618 442462 274854
rect 442698 274618 442782 274854
rect 443018 274618 443102 274854
rect 443338 274618 443422 274854
rect 443658 274618 443742 274854
rect 443978 274618 444062 274854
rect 444298 274618 444382 274854
rect 444618 274618 444740 274854
rect 440740 244218 444740 274618
rect 440740 243982 440862 244218
rect 441098 243982 441182 244218
rect 441418 243982 441502 244218
rect 441738 243982 441822 244218
rect 442058 243982 442142 244218
rect 442378 243982 442462 244218
rect 442698 243982 442782 244218
rect 443018 243982 443102 244218
rect 443338 243982 443422 244218
rect 443658 243982 443742 244218
rect 443978 243982 444062 244218
rect 444298 243982 444382 244218
rect 444618 243982 444740 244218
rect 440740 213582 444740 243982
rect 440740 213346 440862 213582
rect 441098 213346 441182 213582
rect 441418 213346 441502 213582
rect 441738 213346 441822 213582
rect 442058 213346 442142 213582
rect 442378 213346 442462 213582
rect 442698 213346 442782 213582
rect 443018 213346 443102 213582
rect 443338 213346 443422 213582
rect 443658 213346 443742 213582
rect 443978 213346 444062 213582
rect 444298 213346 444382 213582
rect 444618 213346 444740 213582
rect 440740 182946 444740 213346
rect 440740 182710 440862 182946
rect 441098 182710 441182 182946
rect 441418 182710 441502 182946
rect 441738 182710 441822 182946
rect 442058 182710 442142 182946
rect 442378 182710 442462 182946
rect 442698 182710 442782 182946
rect 443018 182710 443102 182946
rect 443338 182710 443422 182946
rect 443658 182710 443742 182946
rect 443978 182710 444062 182946
rect 444298 182710 444382 182946
rect 444618 182710 444740 182946
rect 440740 152310 444740 182710
rect 440740 152074 440862 152310
rect 441098 152074 441182 152310
rect 441418 152074 441502 152310
rect 441738 152074 441822 152310
rect 442058 152074 442142 152310
rect 442378 152074 442462 152310
rect 442698 152074 442782 152310
rect 443018 152074 443102 152310
rect 443338 152074 443422 152310
rect 443658 152074 443742 152310
rect 443978 152074 444062 152310
rect 444298 152074 444382 152310
rect 444618 152074 444740 152310
rect 440740 121674 444740 152074
rect 440740 121438 440862 121674
rect 441098 121438 441182 121674
rect 441418 121438 441502 121674
rect 441738 121438 441822 121674
rect 442058 121438 442142 121674
rect 442378 121438 442462 121674
rect 442698 121438 442782 121674
rect 443018 121438 443102 121674
rect 443338 121438 443422 121674
rect 443658 121438 443742 121674
rect 443978 121438 444062 121674
rect 444298 121438 444382 121674
rect 444618 121438 444740 121674
rect 440740 91038 444740 121438
rect 440740 90802 440862 91038
rect 441098 90802 441182 91038
rect 441418 90802 441502 91038
rect 441738 90802 441822 91038
rect 442058 90802 442142 91038
rect 442378 90802 442462 91038
rect 442698 90802 442782 91038
rect 443018 90802 443102 91038
rect 443338 90802 443422 91038
rect 443658 90802 443742 91038
rect 443978 90802 444062 91038
rect 444298 90802 444382 91038
rect 444618 90802 444740 91038
rect 440740 60402 444740 90802
rect 440740 60166 440862 60402
rect 441098 60166 441182 60402
rect 441418 60166 441502 60402
rect 441738 60166 441822 60402
rect 442058 60166 442142 60402
rect 442378 60166 442462 60402
rect 442698 60166 442782 60402
rect 443018 60166 443102 60402
rect 443338 60166 443422 60402
rect 443658 60166 443742 60402
rect 443978 60166 444062 60402
rect 444298 60166 444382 60402
rect 444618 60166 444740 60402
rect 440740 29766 444740 60166
rect 440740 29530 440862 29766
rect 441098 29530 441182 29766
rect 441418 29530 441502 29766
rect 441738 29530 441822 29766
rect 442058 29530 442142 29766
rect 442378 29530 442462 29766
rect 442698 29530 442782 29766
rect 443018 29530 443102 29766
rect 443338 29530 443422 29766
rect 443658 29530 443742 29766
rect 443978 29530 444062 29766
rect 444298 29530 444382 29766
rect 444618 29530 444740 29766
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 440740 3878 444740 29530
rect 440740 3642 440862 3878
rect 441098 3642 441182 3878
rect 441418 3642 441502 3878
rect 441738 3642 441822 3878
rect 442058 3642 442142 3878
rect 442378 3642 442462 3878
rect 442698 3642 442782 3878
rect 443018 3642 443102 3878
rect 443338 3642 443422 3878
rect 443658 3642 443742 3878
rect 443978 3642 444062 3878
rect 444298 3642 444382 3878
rect 444618 3642 444740 3878
rect 440740 3558 444740 3642
rect 440740 3322 440862 3558
rect 441098 3322 441182 3558
rect 441418 3322 441502 3558
rect 441738 3322 441822 3558
rect 442058 3322 442142 3558
rect 442378 3322 442462 3558
rect 442698 3322 442782 3558
rect 443018 3322 443102 3558
rect 443338 3322 443422 3558
rect 443658 3322 443742 3558
rect 443978 3322 444062 3558
rect 444298 3322 444382 3558
rect 444618 3322 444740 3558
rect 440740 3238 444740 3322
rect 440740 3002 440862 3238
rect 441098 3002 441182 3238
rect 441418 3002 441502 3238
rect 441738 3002 441822 3238
rect 442058 3002 442142 3238
rect 442378 3002 442462 3238
rect 442698 3002 442782 3238
rect 443018 3002 443102 3238
rect 443338 3002 443422 3238
rect 443658 3002 443742 3238
rect 443978 3002 444062 3238
rect 444298 3002 444382 3238
rect 444618 3002 444740 3238
rect 440740 2918 444740 3002
rect 440740 2682 440862 2918
rect 441098 2682 441182 2918
rect 441418 2682 441502 2918
rect 441738 2682 441822 2918
rect 442058 2682 442142 2918
rect 442378 2682 442462 2918
rect 442698 2682 442782 2918
rect 443018 2682 443102 2918
rect 443338 2682 443422 2918
rect 443658 2682 443742 2918
rect 443978 2682 444062 2918
rect 444298 2682 444382 2918
rect 444618 2682 444740 2918
rect 440740 2598 444740 2682
rect 440740 2362 440862 2598
rect 441098 2362 441182 2598
rect 441418 2362 441502 2598
rect 441738 2362 441822 2598
rect 442058 2362 442142 2598
rect 442378 2362 442462 2598
rect 442698 2362 442782 2598
rect 443018 2362 443102 2598
rect 443338 2362 443422 2598
rect 443658 2362 443742 2598
rect 443978 2362 444062 2598
rect 444298 2362 444382 2598
rect 444618 2362 444740 2598
rect 440740 2278 444740 2362
rect 440740 2042 440862 2278
rect 441098 2042 441182 2278
rect 441418 2042 441502 2278
rect 441738 2042 441822 2278
rect 442058 2042 442142 2278
rect 442378 2042 442462 2278
rect 442698 2042 442782 2278
rect 443018 2042 443102 2278
rect 443338 2042 443422 2278
rect 443658 2042 443742 2278
rect 443978 2042 444062 2278
rect 444298 2042 444382 2278
rect 444618 2042 444740 2278
rect 440740 1958 444740 2042
rect 440740 1722 440862 1958
rect 441098 1722 441182 1958
rect 441418 1722 441502 1958
rect 441738 1722 441822 1958
rect 442058 1722 442142 1958
rect 442378 1722 442462 1958
rect 442698 1722 442782 1958
rect 443018 1722 443102 1958
rect 443338 1722 443422 1958
rect 443658 1722 443742 1958
rect 443978 1722 444062 1958
rect 444298 1722 444382 1958
rect 444618 1722 444740 1958
rect 440740 1638 444740 1722
rect 440740 1402 440862 1638
rect 441098 1402 441182 1638
rect 441418 1402 441502 1638
rect 441738 1402 441822 1638
rect 442058 1402 442142 1638
rect 442378 1402 442462 1638
rect 442698 1402 442782 1638
rect 443018 1402 443102 1638
rect 443338 1402 443422 1638
rect 443658 1402 443742 1638
rect 443978 1402 444062 1638
rect 444298 1402 444382 1638
rect 444618 1402 444740 1638
rect 440740 1318 444740 1402
rect 440740 1082 440862 1318
rect 441098 1082 441182 1318
rect 441418 1082 441502 1318
rect 441738 1082 441822 1318
rect 442058 1082 442142 1318
rect 442378 1082 442462 1318
rect 442698 1082 442782 1318
rect 443018 1082 443102 1318
rect 443338 1082 443422 1318
rect 443658 1082 443742 1318
rect 443978 1082 444062 1318
rect 444298 1082 444382 1318
rect 444618 1082 444740 1318
rect 440740 998 444740 1082
rect 440740 762 440862 998
rect 441098 762 441182 998
rect 441418 762 441502 998
rect 441738 762 441822 998
rect 442058 762 442142 998
rect 442378 762 442462 998
rect 442698 762 442782 998
rect 443018 762 443102 998
rect 443338 762 443422 998
rect 443658 762 443742 998
rect 443978 762 444062 998
rect 444298 762 444382 998
rect 444618 762 444740 998
rect 440740 678 444740 762
rect 440740 442 440862 678
rect 441098 442 441182 678
rect 441418 442 441502 678
rect 441738 442 441822 678
rect 442058 442 442142 678
rect 442378 442 442462 678
rect 442698 442 442782 678
rect 443018 442 443102 678
rect 443338 442 443422 678
rect 443658 442 443742 678
rect 443978 442 444062 678
rect 444298 442 444382 678
rect 444618 442 444740 678
rect 440740 358 444740 442
rect 440740 122 440862 358
rect 441098 122 441182 358
rect 441418 122 441502 358
rect 441738 122 441822 358
rect 442058 122 442142 358
rect 442378 122 442462 358
rect 442698 122 442782 358
rect 443018 122 443102 358
rect 443338 122 443422 358
rect 443658 122 443742 358
rect 443978 122 444062 358
rect 444298 122 444382 358
rect 444618 122 444740 358
rect 440740 0 444740 122
<< via4 >>
rect 122 405162 358 405398
rect 442 405162 678 405398
rect 762 405162 998 405398
rect 1082 405162 1318 405398
rect 1402 405162 1638 405398
rect 1722 405162 1958 405398
rect 2042 405162 2278 405398
rect 2362 405162 2598 405398
rect 2682 405162 2918 405398
rect 3002 405162 3238 405398
rect 3322 405162 3558 405398
rect 3642 405162 3878 405398
rect 122 404842 358 405078
rect 442 404842 678 405078
rect 762 404842 998 405078
rect 1082 404842 1318 405078
rect 1402 404842 1638 405078
rect 1722 404842 1958 405078
rect 2042 404842 2278 405078
rect 2362 404842 2598 405078
rect 2682 404842 2918 405078
rect 3002 404842 3238 405078
rect 3322 404842 3558 405078
rect 3642 404842 3878 405078
rect 122 404522 358 404758
rect 442 404522 678 404758
rect 762 404522 998 404758
rect 1082 404522 1318 404758
rect 1402 404522 1638 404758
rect 1722 404522 1958 404758
rect 2042 404522 2278 404758
rect 2362 404522 2598 404758
rect 2682 404522 2918 404758
rect 3002 404522 3238 404758
rect 3322 404522 3558 404758
rect 3642 404522 3878 404758
rect 122 404202 358 404438
rect 442 404202 678 404438
rect 762 404202 998 404438
rect 1082 404202 1318 404438
rect 1402 404202 1638 404438
rect 1722 404202 1958 404438
rect 2042 404202 2278 404438
rect 2362 404202 2598 404438
rect 2682 404202 2918 404438
rect 3002 404202 3238 404438
rect 3322 404202 3558 404438
rect 3642 404202 3878 404438
rect 122 403882 358 404118
rect 442 403882 678 404118
rect 762 403882 998 404118
rect 1082 403882 1318 404118
rect 1402 403882 1638 404118
rect 1722 403882 1958 404118
rect 2042 403882 2278 404118
rect 2362 403882 2598 404118
rect 2682 403882 2918 404118
rect 3002 403882 3238 404118
rect 3322 403882 3558 404118
rect 3642 403882 3878 404118
rect 122 403562 358 403798
rect 442 403562 678 403798
rect 762 403562 998 403798
rect 1082 403562 1318 403798
rect 1402 403562 1638 403798
rect 1722 403562 1958 403798
rect 2042 403562 2278 403798
rect 2362 403562 2598 403798
rect 2682 403562 2918 403798
rect 3002 403562 3238 403798
rect 3322 403562 3558 403798
rect 3642 403562 3878 403798
rect 122 403242 358 403478
rect 442 403242 678 403478
rect 762 403242 998 403478
rect 1082 403242 1318 403478
rect 1402 403242 1638 403478
rect 1722 403242 1958 403478
rect 2042 403242 2278 403478
rect 2362 403242 2598 403478
rect 2682 403242 2918 403478
rect 3002 403242 3238 403478
rect 3322 403242 3558 403478
rect 3642 403242 3878 403478
rect 122 402922 358 403158
rect 442 402922 678 403158
rect 762 402922 998 403158
rect 1082 402922 1318 403158
rect 1402 402922 1638 403158
rect 1722 402922 1958 403158
rect 2042 402922 2278 403158
rect 2362 402922 2598 403158
rect 2682 402922 2918 403158
rect 3002 402922 3238 403158
rect 3322 402922 3558 403158
rect 3642 402922 3878 403158
rect 122 402602 358 402838
rect 442 402602 678 402838
rect 762 402602 998 402838
rect 1082 402602 1318 402838
rect 1402 402602 1638 402838
rect 1722 402602 1958 402838
rect 2042 402602 2278 402838
rect 2362 402602 2598 402838
rect 2682 402602 2918 402838
rect 3002 402602 3238 402838
rect 3322 402602 3558 402838
rect 3642 402602 3878 402838
rect 122 402282 358 402518
rect 442 402282 678 402518
rect 762 402282 998 402518
rect 1082 402282 1318 402518
rect 1402 402282 1638 402518
rect 1722 402282 1958 402518
rect 2042 402282 2278 402518
rect 2362 402282 2598 402518
rect 2682 402282 2918 402518
rect 3002 402282 3238 402518
rect 3322 402282 3558 402518
rect 3642 402282 3878 402518
rect 122 401962 358 402198
rect 442 401962 678 402198
rect 762 401962 998 402198
rect 1082 401962 1318 402198
rect 1402 401962 1638 402198
rect 1722 401962 1958 402198
rect 2042 401962 2278 402198
rect 2362 401962 2598 402198
rect 2682 401962 2918 402198
rect 3002 401962 3238 402198
rect 3322 401962 3558 402198
rect 3642 401962 3878 402198
rect 122 401642 358 401878
rect 442 401642 678 401878
rect 762 401642 998 401878
rect 1082 401642 1318 401878
rect 1402 401642 1638 401878
rect 1722 401642 1958 401878
rect 2042 401642 2278 401878
rect 2362 401642 2598 401878
rect 2682 401642 2918 401878
rect 3002 401642 3238 401878
rect 3322 401642 3558 401878
rect 3642 401642 3878 401878
rect 440862 405162 441098 405398
rect 441182 405162 441418 405398
rect 441502 405162 441738 405398
rect 441822 405162 442058 405398
rect 442142 405162 442378 405398
rect 442462 405162 442698 405398
rect 442782 405162 443018 405398
rect 443102 405162 443338 405398
rect 443422 405162 443658 405398
rect 443742 405162 443978 405398
rect 444062 405162 444298 405398
rect 444382 405162 444618 405398
rect 440862 404842 441098 405078
rect 441182 404842 441418 405078
rect 441502 404842 441738 405078
rect 441822 404842 442058 405078
rect 442142 404842 442378 405078
rect 442462 404842 442698 405078
rect 442782 404842 443018 405078
rect 443102 404842 443338 405078
rect 443422 404842 443658 405078
rect 443742 404842 443978 405078
rect 444062 404842 444298 405078
rect 444382 404842 444618 405078
rect 440862 404522 441098 404758
rect 441182 404522 441418 404758
rect 441502 404522 441738 404758
rect 441822 404522 442058 404758
rect 442142 404522 442378 404758
rect 442462 404522 442698 404758
rect 442782 404522 443018 404758
rect 443102 404522 443338 404758
rect 443422 404522 443658 404758
rect 443742 404522 443978 404758
rect 444062 404522 444298 404758
rect 444382 404522 444618 404758
rect 440862 404202 441098 404438
rect 441182 404202 441418 404438
rect 441502 404202 441738 404438
rect 441822 404202 442058 404438
rect 442142 404202 442378 404438
rect 442462 404202 442698 404438
rect 442782 404202 443018 404438
rect 443102 404202 443338 404438
rect 443422 404202 443658 404438
rect 443742 404202 443978 404438
rect 444062 404202 444298 404438
rect 444382 404202 444618 404438
rect 440862 403882 441098 404118
rect 441182 403882 441418 404118
rect 441502 403882 441738 404118
rect 441822 403882 442058 404118
rect 442142 403882 442378 404118
rect 442462 403882 442698 404118
rect 442782 403882 443018 404118
rect 443102 403882 443338 404118
rect 443422 403882 443658 404118
rect 443742 403882 443978 404118
rect 444062 403882 444298 404118
rect 444382 403882 444618 404118
rect 440862 403562 441098 403798
rect 441182 403562 441418 403798
rect 441502 403562 441738 403798
rect 441822 403562 442058 403798
rect 442142 403562 442378 403798
rect 442462 403562 442698 403798
rect 442782 403562 443018 403798
rect 443102 403562 443338 403798
rect 443422 403562 443658 403798
rect 443742 403562 443978 403798
rect 444062 403562 444298 403798
rect 444382 403562 444618 403798
rect 440862 403242 441098 403478
rect 441182 403242 441418 403478
rect 441502 403242 441738 403478
rect 441822 403242 442058 403478
rect 442142 403242 442378 403478
rect 442462 403242 442698 403478
rect 442782 403242 443018 403478
rect 443102 403242 443338 403478
rect 443422 403242 443658 403478
rect 443742 403242 443978 403478
rect 444062 403242 444298 403478
rect 444382 403242 444618 403478
rect 440862 402922 441098 403158
rect 441182 402922 441418 403158
rect 441502 402922 441738 403158
rect 441822 402922 442058 403158
rect 442142 402922 442378 403158
rect 442462 402922 442698 403158
rect 442782 402922 443018 403158
rect 443102 402922 443338 403158
rect 443422 402922 443658 403158
rect 443742 402922 443978 403158
rect 444062 402922 444298 403158
rect 444382 402922 444618 403158
rect 440862 402602 441098 402838
rect 441182 402602 441418 402838
rect 441502 402602 441738 402838
rect 441822 402602 442058 402838
rect 442142 402602 442378 402838
rect 442462 402602 442698 402838
rect 442782 402602 443018 402838
rect 443102 402602 443338 402838
rect 443422 402602 443658 402838
rect 443742 402602 443978 402838
rect 444062 402602 444298 402838
rect 444382 402602 444618 402838
rect 440862 402282 441098 402518
rect 441182 402282 441418 402518
rect 441502 402282 441738 402518
rect 441822 402282 442058 402518
rect 442142 402282 442378 402518
rect 442462 402282 442698 402518
rect 442782 402282 443018 402518
rect 443102 402282 443338 402518
rect 443422 402282 443658 402518
rect 443742 402282 443978 402518
rect 444062 402282 444298 402518
rect 444382 402282 444618 402518
rect 440862 401962 441098 402198
rect 441182 401962 441418 402198
rect 441502 401962 441738 402198
rect 441822 401962 442058 402198
rect 442142 401962 442378 402198
rect 442462 401962 442698 402198
rect 442782 401962 443018 402198
rect 443102 401962 443338 402198
rect 443422 401962 443658 402198
rect 443742 401962 443978 402198
rect 444062 401962 444298 402198
rect 444382 401962 444618 402198
rect 440862 401642 441098 401878
rect 441182 401642 441418 401878
rect 441502 401642 441738 401878
rect 441822 401642 442058 401878
rect 442142 401642 442378 401878
rect 442462 401642 442698 401878
rect 442782 401642 443018 401878
rect 443102 401642 443338 401878
rect 443422 401642 443658 401878
rect 443742 401642 443978 401878
rect 444062 401642 444298 401878
rect 444382 401642 444618 401878
rect 122 366526 358 366762
rect 442 366526 678 366762
rect 762 366526 998 366762
rect 1082 366526 1318 366762
rect 1402 366526 1638 366762
rect 1722 366526 1958 366762
rect 2042 366526 2278 366762
rect 2362 366526 2598 366762
rect 2682 366526 2918 366762
rect 3002 366526 3238 366762
rect 3322 366526 3558 366762
rect 3642 366526 3878 366762
rect 122 335890 358 336126
rect 442 335890 678 336126
rect 762 335890 998 336126
rect 1082 335890 1318 336126
rect 1402 335890 1638 336126
rect 1722 335890 1958 336126
rect 2042 335890 2278 336126
rect 2362 335890 2598 336126
rect 2682 335890 2918 336126
rect 3002 335890 3238 336126
rect 3322 335890 3558 336126
rect 3642 335890 3878 336126
rect 122 305254 358 305490
rect 442 305254 678 305490
rect 762 305254 998 305490
rect 1082 305254 1318 305490
rect 1402 305254 1638 305490
rect 1722 305254 1958 305490
rect 2042 305254 2278 305490
rect 2362 305254 2598 305490
rect 2682 305254 2918 305490
rect 3002 305254 3238 305490
rect 3322 305254 3558 305490
rect 3642 305254 3878 305490
rect 122 274618 358 274854
rect 442 274618 678 274854
rect 762 274618 998 274854
rect 1082 274618 1318 274854
rect 1402 274618 1638 274854
rect 1722 274618 1958 274854
rect 2042 274618 2278 274854
rect 2362 274618 2598 274854
rect 2682 274618 2918 274854
rect 3002 274618 3238 274854
rect 3322 274618 3558 274854
rect 3642 274618 3878 274854
rect 122 243982 358 244218
rect 442 243982 678 244218
rect 762 243982 998 244218
rect 1082 243982 1318 244218
rect 1402 243982 1638 244218
rect 1722 243982 1958 244218
rect 2042 243982 2278 244218
rect 2362 243982 2598 244218
rect 2682 243982 2918 244218
rect 3002 243982 3238 244218
rect 3322 243982 3558 244218
rect 3642 243982 3878 244218
rect 122 213346 358 213582
rect 442 213346 678 213582
rect 762 213346 998 213582
rect 1082 213346 1318 213582
rect 1402 213346 1638 213582
rect 1722 213346 1958 213582
rect 2042 213346 2278 213582
rect 2362 213346 2598 213582
rect 2682 213346 2918 213582
rect 3002 213346 3238 213582
rect 3322 213346 3558 213582
rect 3642 213346 3878 213582
rect 122 182710 358 182946
rect 442 182710 678 182946
rect 762 182710 998 182946
rect 1082 182710 1318 182946
rect 1402 182710 1638 182946
rect 1722 182710 1958 182946
rect 2042 182710 2278 182946
rect 2362 182710 2598 182946
rect 2682 182710 2918 182946
rect 3002 182710 3238 182946
rect 3322 182710 3558 182946
rect 3642 182710 3878 182946
rect 122 152074 358 152310
rect 442 152074 678 152310
rect 762 152074 998 152310
rect 1082 152074 1318 152310
rect 1402 152074 1638 152310
rect 1722 152074 1958 152310
rect 2042 152074 2278 152310
rect 2362 152074 2598 152310
rect 2682 152074 2918 152310
rect 3002 152074 3238 152310
rect 3322 152074 3558 152310
rect 3642 152074 3878 152310
rect 122 121438 358 121674
rect 442 121438 678 121674
rect 762 121438 998 121674
rect 1082 121438 1318 121674
rect 1402 121438 1638 121674
rect 1722 121438 1958 121674
rect 2042 121438 2278 121674
rect 2362 121438 2598 121674
rect 2682 121438 2918 121674
rect 3002 121438 3238 121674
rect 3322 121438 3558 121674
rect 3642 121438 3878 121674
rect 122 90802 358 91038
rect 442 90802 678 91038
rect 762 90802 998 91038
rect 1082 90802 1318 91038
rect 1402 90802 1638 91038
rect 1722 90802 1958 91038
rect 2042 90802 2278 91038
rect 2362 90802 2598 91038
rect 2682 90802 2918 91038
rect 3002 90802 3238 91038
rect 3322 90802 3558 91038
rect 3642 90802 3878 91038
rect 122 60166 358 60402
rect 442 60166 678 60402
rect 762 60166 998 60402
rect 1082 60166 1318 60402
rect 1402 60166 1638 60402
rect 1722 60166 1958 60402
rect 2042 60166 2278 60402
rect 2362 60166 2598 60402
rect 2682 60166 2918 60402
rect 3002 60166 3238 60402
rect 3322 60166 3558 60402
rect 3642 60166 3878 60402
rect 122 29530 358 29766
rect 442 29530 678 29766
rect 762 29530 998 29766
rect 1082 29530 1318 29766
rect 1402 29530 1638 29766
rect 1722 29530 1958 29766
rect 2042 29530 2278 29766
rect 2362 29530 2598 29766
rect 2682 29530 2918 29766
rect 3002 29530 3238 29766
rect 3322 29530 3558 29766
rect 3642 29530 3878 29766
rect 5122 400162 5358 400398
rect 5442 400162 5678 400398
rect 5762 400162 5998 400398
rect 6082 400162 6318 400398
rect 6402 400162 6638 400398
rect 6722 400162 6958 400398
rect 7042 400162 7278 400398
rect 7362 400162 7598 400398
rect 7682 400162 7918 400398
rect 8002 400162 8238 400398
rect 8322 400162 8558 400398
rect 8642 400162 8878 400398
rect 5122 399842 5358 400078
rect 5442 399842 5678 400078
rect 5762 399842 5998 400078
rect 6082 399842 6318 400078
rect 6402 399842 6638 400078
rect 6722 399842 6958 400078
rect 7042 399842 7278 400078
rect 7362 399842 7598 400078
rect 7682 399842 7918 400078
rect 8002 399842 8238 400078
rect 8322 399842 8558 400078
rect 8642 399842 8878 400078
rect 5122 399522 5358 399758
rect 5442 399522 5678 399758
rect 5762 399522 5998 399758
rect 6082 399522 6318 399758
rect 6402 399522 6638 399758
rect 6722 399522 6958 399758
rect 7042 399522 7278 399758
rect 7362 399522 7598 399758
rect 7682 399522 7918 399758
rect 8002 399522 8238 399758
rect 8322 399522 8558 399758
rect 8642 399522 8878 399758
rect 5122 399202 5358 399438
rect 5442 399202 5678 399438
rect 5762 399202 5998 399438
rect 6082 399202 6318 399438
rect 6402 399202 6638 399438
rect 6722 399202 6958 399438
rect 7042 399202 7278 399438
rect 7362 399202 7598 399438
rect 7682 399202 7918 399438
rect 8002 399202 8238 399438
rect 8322 399202 8558 399438
rect 8642 399202 8878 399438
rect 5122 398882 5358 399118
rect 5442 398882 5678 399118
rect 5762 398882 5998 399118
rect 6082 398882 6318 399118
rect 6402 398882 6638 399118
rect 6722 398882 6958 399118
rect 7042 398882 7278 399118
rect 7362 398882 7598 399118
rect 7682 398882 7918 399118
rect 8002 398882 8238 399118
rect 8322 398882 8558 399118
rect 8642 398882 8878 399118
rect 5122 398562 5358 398798
rect 5442 398562 5678 398798
rect 5762 398562 5998 398798
rect 6082 398562 6318 398798
rect 6402 398562 6638 398798
rect 6722 398562 6958 398798
rect 7042 398562 7278 398798
rect 7362 398562 7598 398798
rect 7682 398562 7918 398798
rect 8002 398562 8238 398798
rect 8322 398562 8558 398798
rect 8642 398562 8878 398798
rect 5122 398242 5358 398478
rect 5442 398242 5678 398478
rect 5762 398242 5998 398478
rect 6082 398242 6318 398478
rect 6402 398242 6638 398478
rect 6722 398242 6958 398478
rect 7042 398242 7278 398478
rect 7362 398242 7598 398478
rect 7682 398242 7918 398478
rect 8002 398242 8238 398478
rect 8322 398242 8558 398478
rect 8642 398242 8878 398478
rect 5122 397922 5358 398158
rect 5442 397922 5678 398158
rect 5762 397922 5998 398158
rect 6082 397922 6318 398158
rect 6402 397922 6638 398158
rect 6722 397922 6958 398158
rect 7042 397922 7278 398158
rect 7362 397922 7598 398158
rect 7682 397922 7918 398158
rect 8002 397922 8238 398158
rect 8322 397922 8558 398158
rect 8642 397922 8878 398158
rect 5122 397602 5358 397838
rect 5442 397602 5678 397838
rect 5762 397602 5998 397838
rect 6082 397602 6318 397838
rect 6402 397602 6638 397838
rect 6722 397602 6958 397838
rect 7042 397602 7278 397838
rect 7362 397602 7598 397838
rect 7682 397602 7918 397838
rect 8002 397602 8238 397838
rect 8322 397602 8558 397838
rect 8642 397602 8878 397838
rect 5122 397282 5358 397518
rect 5442 397282 5678 397518
rect 5762 397282 5998 397518
rect 6082 397282 6318 397518
rect 6402 397282 6638 397518
rect 6722 397282 6958 397518
rect 7042 397282 7278 397518
rect 7362 397282 7598 397518
rect 7682 397282 7918 397518
rect 8002 397282 8238 397518
rect 8322 397282 8558 397518
rect 8642 397282 8878 397518
rect 5122 396962 5358 397198
rect 5442 396962 5678 397198
rect 5762 396962 5998 397198
rect 6082 396962 6318 397198
rect 6402 396962 6638 397198
rect 6722 396962 6958 397198
rect 7042 396962 7278 397198
rect 7362 396962 7598 397198
rect 7682 396962 7918 397198
rect 8002 396962 8238 397198
rect 8322 396962 8558 397198
rect 8642 396962 8878 397198
rect 5122 396642 5358 396878
rect 5442 396642 5678 396878
rect 5762 396642 5998 396878
rect 6082 396642 6318 396878
rect 6402 396642 6638 396878
rect 6722 396642 6958 396878
rect 7042 396642 7278 396878
rect 7362 396642 7598 396878
rect 7682 396642 7918 396878
rect 8002 396642 8238 396878
rect 8322 396642 8558 396878
rect 8642 396642 8878 396878
rect 435862 400162 436098 400398
rect 436182 400162 436418 400398
rect 436502 400162 436738 400398
rect 436822 400162 437058 400398
rect 437142 400162 437378 400398
rect 437462 400162 437698 400398
rect 437782 400162 438018 400398
rect 438102 400162 438338 400398
rect 438422 400162 438658 400398
rect 438742 400162 438978 400398
rect 439062 400162 439298 400398
rect 439382 400162 439618 400398
rect 435862 399842 436098 400078
rect 436182 399842 436418 400078
rect 436502 399842 436738 400078
rect 436822 399842 437058 400078
rect 437142 399842 437378 400078
rect 437462 399842 437698 400078
rect 437782 399842 438018 400078
rect 438102 399842 438338 400078
rect 438422 399842 438658 400078
rect 438742 399842 438978 400078
rect 439062 399842 439298 400078
rect 439382 399842 439618 400078
rect 435862 399522 436098 399758
rect 436182 399522 436418 399758
rect 436502 399522 436738 399758
rect 436822 399522 437058 399758
rect 437142 399522 437378 399758
rect 437462 399522 437698 399758
rect 437782 399522 438018 399758
rect 438102 399522 438338 399758
rect 438422 399522 438658 399758
rect 438742 399522 438978 399758
rect 439062 399522 439298 399758
rect 439382 399522 439618 399758
rect 435862 399202 436098 399438
rect 436182 399202 436418 399438
rect 436502 399202 436738 399438
rect 436822 399202 437058 399438
rect 437142 399202 437378 399438
rect 437462 399202 437698 399438
rect 437782 399202 438018 399438
rect 438102 399202 438338 399438
rect 438422 399202 438658 399438
rect 438742 399202 438978 399438
rect 439062 399202 439298 399438
rect 439382 399202 439618 399438
rect 435862 398882 436098 399118
rect 436182 398882 436418 399118
rect 436502 398882 436738 399118
rect 436822 398882 437058 399118
rect 437142 398882 437378 399118
rect 437462 398882 437698 399118
rect 437782 398882 438018 399118
rect 438102 398882 438338 399118
rect 438422 398882 438658 399118
rect 438742 398882 438978 399118
rect 439062 398882 439298 399118
rect 439382 398882 439618 399118
rect 435862 398562 436098 398798
rect 436182 398562 436418 398798
rect 436502 398562 436738 398798
rect 436822 398562 437058 398798
rect 437142 398562 437378 398798
rect 437462 398562 437698 398798
rect 437782 398562 438018 398798
rect 438102 398562 438338 398798
rect 438422 398562 438658 398798
rect 438742 398562 438978 398798
rect 439062 398562 439298 398798
rect 439382 398562 439618 398798
rect 435862 398242 436098 398478
rect 436182 398242 436418 398478
rect 436502 398242 436738 398478
rect 436822 398242 437058 398478
rect 437142 398242 437378 398478
rect 437462 398242 437698 398478
rect 437782 398242 438018 398478
rect 438102 398242 438338 398478
rect 438422 398242 438658 398478
rect 438742 398242 438978 398478
rect 439062 398242 439298 398478
rect 439382 398242 439618 398478
rect 435862 397922 436098 398158
rect 436182 397922 436418 398158
rect 436502 397922 436738 398158
rect 436822 397922 437058 398158
rect 437142 397922 437378 398158
rect 437462 397922 437698 398158
rect 437782 397922 438018 398158
rect 438102 397922 438338 398158
rect 438422 397922 438658 398158
rect 438742 397922 438978 398158
rect 439062 397922 439298 398158
rect 439382 397922 439618 398158
rect 435862 397602 436098 397838
rect 436182 397602 436418 397838
rect 436502 397602 436738 397838
rect 436822 397602 437058 397838
rect 437142 397602 437378 397838
rect 437462 397602 437698 397838
rect 437782 397602 438018 397838
rect 438102 397602 438338 397838
rect 438422 397602 438658 397838
rect 438742 397602 438978 397838
rect 439062 397602 439298 397838
rect 439382 397602 439618 397838
rect 435862 397282 436098 397518
rect 436182 397282 436418 397518
rect 436502 397282 436738 397518
rect 436822 397282 437058 397518
rect 437142 397282 437378 397518
rect 437462 397282 437698 397518
rect 437782 397282 438018 397518
rect 438102 397282 438338 397518
rect 438422 397282 438658 397518
rect 438742 397282 438978 397518
rect 439062 397282 439298 397518
rect 439382 397282 439618 397518
rect 435862 396962 436098 397198
rect 436182 396962 436418 397198
rect 436502 396962 436738 397198
rect 436822 396962 437058 397198
rect 437142 396962 437378 397198
rect 437462 396962 437698 397198
rect 437782 396962 438018 397198
rect 438102 396962 438338 397198
rect 438422 396962 438658 397198
rect 438742 396962 438978 397198
rect 439062 396962 439298 397198
rect 439382 396962 439618 397198
rect 435862 396642 436098 396878
rect 436182 396642 436418 396878
rect 436502 396642 436738 396878
rect 436822 396642 437058 396878
rect 437142 396642 437378 396878
rect 437462 396642 437698 396878
rect 437782 396642 438018 396878
rect 438102 396642 438338 396878
rect 438422 396642 438658 396878
rect 438742 396642 438978 396878
rect 439062 396642 439298 396878
rect 439382 396642 439618 396878
rect 5122 381844 5358 382080
rect 5442 381844 5678 382080
rect 5762 381844 5998 382080
rect 6082 381844 6318 382080
rect 6402 381844 6638 382080
rect 6722 381844 6958 382080
rect 7042 381844 7278 382080
rect 7362 381844 7598 382080
rect 7682 381844 7918 382080
rect 8002 381844 8238 382080
rect 8322 381844 8558 382080
rect 8642 381844 8878 382080
rect 435862 381844 436098 382080
rect 436182 381844 436418 382080
rect 436502 381844 436738 382080
rect 436822 381844 437058 382080
rect 437142 381844 437378 382080
rect 437462 381844 437698 382080
rect 437782 381844 438018 382080
rect 438102 381844 438338 382080
rect 438422 381844 438658 382080
rect 438742 381844 438978 382080
rect 439062 381844 439298 382080
rect 439382 381844 439618 382080
rect 332054 355846 332290 356082
rect 341622 355846 341858 356082
rect 5122 351208 5358 351444
rect 5442 351208 5678 351444
rect 5762 351208 5998 351444
rect 6082 351208 6318 351444
rect 6402 351208 6638 351444
rect 6722 351208 6958 351444
rect 7042 351208 7278 351444
rect 7362 351208 7598 351444
rect 7682 351208 7918 351444
rect 8002 351208 8238 351444
rect 8322 351208 8558 351444
rect 8642 351208 8878 351444
rect 435862 351208 436098 351444
rect 436182 351208 436418 351444
rect 436502 351208 436738 351444
rect 436822 351208 437058 351444
rect 437142 351208 437378 351444
rect 437462 351208 437698 351444
rect 437782 351208 438018 351444
rect 438102 351208 438338 351444
rect 438422 351208 438658 351444
rect 438742 351208 438978 351444
rect 439062 351208 439298 351444
rect 439382 351208 439618 351444
rect 332054 349726 332290 349962
rect 341070 336806 341306 337042
rect 341070 334766 341306 335002
rect 5122 320572 5358 320808
rect 5442 320572 5678 320808
rect 5762 320572 5998 320808
rect 6082 320572 6318 320808
rect 6402 320572 6638 320808
rect 6722 320572 6958 320808
rect 7042 320572 7278 320808
rect 7362 320572 7598 320808
rect 7682 320572 7918 320808
rect 8002 320572 8238 320808
rect 8322 320572 8558 320808
rect 8642 320572 8878 320808
rect 137198 332196 137434 332282
rect 137198 332132 137284 332196
rect 137284 332132 137348 332196
rect 137348 332132 137434 332196
rect 137198 332046 137434 332132
rect 201598 332196 201834 332282
rect 201598 332132 201684 332196
rect 201684 332132 201748 332196
rect 201748 332132 201834 332196
rect 201598 332046 201834 332132
rect 158542 331366 158778 331602
rect 137198 330836 137434 330922
rect 137198 330772 137284 330836
rect 137284 330772 137348 330836
rect 137348 330772 137434 330836
rect 137198 330686 137434 330772
rect 159462 330686 159698 330922
rect 204358 330686 204594 330922
rect 230854 332196 231090 332282
rect 230854 332132 230940 332196
rect 230940 332132 231004 332196
rect 231004 332132 231090 332196
rect 230854 332046 231090 332132
rect 295438 332046 295674 332282
rect 212086 329326 212322 329562
rect 137382 328796 137618 328882
rect 137382 328732 137468 328796
rect 137468 328732 137532 328796
rect 137532 328732 137618 328796
rect 137382 328646 137618 328732
rect 161670 328796 161906 328882
rect 252566 331366 252802 331602
rect 231222 330836 231458 330922
rect 231222 330772 231308 330836
rect 231308 330772 231372 330836
rect 231372 330772 231458 330836
rect 231222 330686 231458 330772
rect 251830 330686 252066 330922
rect 292678 330836 292914 330922
rect 292678 330772 292764 330836
rect 292764 330772 292828 330836
rect 292828 330772 292914 330836
rect 292678 330686 292914 330772
rect 336286 331366 336522 331602
rect 299302 329326 299538 329562
rect 161670 328732 161756 328796
rect 161756 328732 161820 328796
rect 161820 328732 161906 328796
rect 161670 328646 161906 328732
rect 231774 328796 232010 328882
rect 231774 328732 231860 328796
rect 231860 328732 231924 328796
rect 231924 328732 232010 328796
rect 231774 328646 232010 328732
rect 253302 328796 253538 328882
rect 253302 328732 253388 328796
rect 253388 328732 253452 328796
rect 253452 328732 253538 328796
rect 253302 328646 253538 328732
rect 137382 328116 137618 328202
rect 137382 328052 137468 328116
rect 137468 328052 137532 328116
rect 137532 328052 137618 328116
rect 137382 327966 137618 328052
rect 160566 328116 160802 328202
rect 160566 328052 160652 328116
rect 160652 328052 160716 328116
rect 160716 328052 160802 328116
rect 160566 327966 160802 328052
rect 208590 328116 208826 328202
rect 208590 328052 208676 328116
rect 208676 328052 208740 328116
rect 208740 328052 208826 328116
rect 208590 327966 208826 328052
rect 105182 319806 105418 320042
rect 5122 289936 5358 290172
rect 5442 289936 5678 290172
rect 5762 289936 5998 290172
rect 6082 289936 6318 290172
rect 6402 289936 6638 290172
rect 6722 289936 6958 290172
rect 7042 289936 7278 290172
rect 7362 289936 7598 290172
rect 7682 289936 7918 290172
rect 8002 289936 8238 290172
rect 8322 289936 8558 290172
rect 8642 289936 8878 290172
rect 38574 286486 38810 286722
rect 13550 283766 13786 284002
rect 38574 283766 38810 284002
rect 104446 307566 104682 307802
rect 104506 305254 104742 305490
rect 198506 305254 198742 305490
rect 104446 302806 104682 303042
rect 435862 320572 436098 320808
rect 436182 320572 436418 320808
rect 436502 320572 436738 320808
rect 436822 320572 437058 320808
rect 437142 320572 437378 320808
rect 437462 320572 437698 320808
rect 437782 320572 438018 320808
rect 438102 320572 438338 320808
rect 438422 320572 438658 320808
rect 438742 320572 438978 320808
rect 439062 320572 439298 320808
rect 439382 320572 439618 320808
rect 292506 305254 292742 305490
rect 246126 298726 246362 298962
rect 5122 259300 5358 259536
rect 5442 259300 5678 259536
rect 5762 259300 5998 259536
rect 6082 259300 6318 259536
rect 6402 259300 6638 259536
rect 6722 259300 6958 259536
rect 7042 259300 7278 259536
rect 7362 259300 7598 259536
rect 7682 259300 7918 259536
rect 8002 259300 8238 259536
rect 8322 259300 8558 259536
rect 8642 259300 8878 259536
rect 48510 256036 48746 256122
rect 48510 255972 48596 256036
rect 48596 255972 48660 256036
rect 48660 255972 48746 256036
rect 48510 255886 48746 255972
rect 49062 251806 49298 252042
rect 49062 249236 49298 249322
rect 49062 249172 49148 249236
rect 49148 249172 49212 249236
rect 49212 249172 49298 249236
rect 49062 249086 49298 249172
rect 49062 242966 49298 243202
rect 48326 242286 48562 242522
rect 49062 239788 49148 239802
rect 49148 239788 49212 239802
rect 49212 239788 49298 239802
rect 49062 239566 49298 239788
rect 73166 237526 73402 237762
rect 134622 298196 134858 298282
rect 134622 298132 134708 298196
rect 134708 298132 134772 298196
rect 134772 298132 134858 298196
rect 134622 298046 134858 298132
rect 246126 298046 246362 298282
rect 136830 297366 137066 297602
rect 230670 297366 230906 297602
rect 104630 291246 104866 291482
rect 89146 289936 89382 290172
rect 229198 293966 229434 294202
rect 228646 293286 228882 293522
rect 137750 292756 137986 292842
rect 137750 292692 137836 292756
rect 137836 292692 137900 292756
rect 137900 292692 137986 292756
rect 137750 292606 137986 292692
rect 104630 289206 104866 289442
rect 134622 285126 134858 285362
rect 84390 284596 84626 284682
rect 84390 284532 84476 284596
rect 84476 284532 84540 284596
rect 84540 284532 84626 284596
rect 84390 284446 84626 284532
rect 178598 291246 178834 291482
rect 183146 289936 183382 290172
rect 231774 291396 232010 291482
rect 231774 291332 231860 291396
rect 231860 291332 231924 291396
rect 231924 291332 232010 291396
rect 231774 291246 232010 291332
rect 137750 289356 137986 289442
rect 137750 289292 137836 289356
rect 137836 289292 137900 289356
rect 137900 289292 137986 289356
rect 137750 289206 137986 289292
rect 165534 289206 165770 289442
rect 236006 289206 236242 289442
rect 137198 284446 137434 284682
rect 84574 282406 84810 282642
rect 134622 282406 134858 282642
rect 138486 282406 138722 282642
rect 84574 281876 84810 281962
rect 84574 281812 84660 281876
rect 84660 281812 84724 281876
rect 84724 281812 84810 281876
rect 84574 281726 84810 281812
rect 84574 281196 84810 281282
rect 84574 281132 84660 281196
rect 84660 281132 84724 281196
rect 84724 281132 84810 281196
rect 84574 281046 84810 281132
rect 104506 274618 104742 274854
rect 198506 274618 198742 274854
rect 73902 251126 74138 251362
rect 76110 255886 76346 256122
rect 75190 251806 75426 252042
rect 74822 251126 75058 251362
rect 74270 247726 74506 247962
rect 73902 245006 74138 245242
rect 75190 250446 75426 250682
rect 76110 251126 76346 251362
rect 75558 245006 75794 245242
rect 75742 242966 75978 243202
rect 5122 228664 5358 228900
rect 5442 228664 5678 228900
rect 5762 228664 5998 228900
rect 6082 228664 6318 228900
rect 6402 228664 6638 228900
rect 6722 228664 6958 228900
rect 7042 228664 7278 228900
rect 7362 228664 7598 228900
rect 7682 228664 7918 228900
rect 8002 228664 8238 228900
rect 8322 228664 8558 228900
rect 8642 228664 8878 228900
rect 5122 198028 5358 198264
rect 5442 198028 5678 198264
rect 5762 198028 5998 198264
rect 6082 198028 6318 198264
rect 6402 198028 6638 198264
rect 6722 198028 6958 198264
rect 7042 198028 7278 198264
rect 7362 198028 7598 198264
rect 7682 198028 7918 198264
rect 8002 198028 8238 198264
rect 8322 198028 8558 198264
rect 8642 198028 8878 198264
rect 74132 238886 74368 239122
rect 75374 240246 75610 240482
rect 144006 257246 144242 257482
rect 144006 248406 144242 248642
rect 93774 241076 94010 241162
rect 93774 241012 93860 241076
rect 93860 241012 93924 241076
rect 93924 241012 94010 241076
rect 93774 240926 94010 241012
rect 95982 240926 96218 241162
rect 136830 241606 137066 241842
rect 76110 240246 76346 240482
rect 104814 240246 105050 240482
rect 106470 240396 106706 240482
rect 106470 240332 106556 240396
rect 106556 240332 106620 240396
rect 106620 240332 106706 240396
rect 106470 240246 106706 240332
rect 118614 240396 118850 240482
rect 118614 240332 118700 240396
rect 118700 240332 118764 240396
rect 118764 240332 118850 240396
rect 118614 240246 118850 240332
rect 125790 240260 126026 240482
rect 125790 240246 125876 240260
rect 125876 240246 125940 240260
rect 125940 240246 126026 240260
rect 128550 240260 128786 240482
rect 128550 240246 128636 240260
rect 128636 240246 128700 240260
rect 128700 240246 128786 240260
rect 75742 239566 75978 239802
rect 95062 239716 95298 239802
rect 95062 239652 95148 239716
rect 95148 239652 95212 239716
rect 95212 239652 95298 239716
rect 95062 239566 95298 239652
rect 75742 235636 75978 235722
rect 75742 235572 75828 235636
rect 75828 235572 75892 235636
rect 75892 235572 75978 235636
rect 75742 235486 75978 235572
rect 102238 238206 102474 238442
rect 110334 235708 110420 235722
rect 110420 235708 110484 235722
rect 110484 235708 110570 235722
rect 110334 235486 110570 235708
rect 143638 241606 143874 241842
rect 138670 239566 138906 239802
rect 143638 239566 143874 239802
rect 142718 238356 142954 238442
rect 142718 238292 142804 238356
rect 142804 238292 142868 238356
rect 142868 238292 142954 238356
rect 142718 238206 142954 238292
rect 167742 240246 167978 240482
rect 147870 237526 148106 237762
rect 149158 237526 149394 237762
rect 144006 236846 144242 237082
rect 148606 236846 148842 237082
rect 149526 236180 149762 236402
rect 149526 236166 149612 236180
rect 149612 236166 149676 236180
rect 149676 236166 149762 236180
rect 153390 236316 153626 236402
rect 153390 236252 153476 236316
rect 153476 236252 153540 236316
rect 153540 236252 153626 236316
rect 153390 236166 153626 236252
rect 162774 236316 163010 236402
rect 162774 236252 162860 236316
rect 162860 236252 162924 236316
rect 162924 236252 163010 236316
rect 162774 236166 163010 236252
rect 137750 234956 137986 235042
rect 137750 234892 137836 234956
rect 137836 234892 137900 234956
rect 137900 234892 137986 234956
rect 137750 234806 137986 234892
rect 141062 234806 141298 235042
rect 144926 234956 145162 235042
rect 144926 234892 145012 234956
rect 145012 234892 145076 234956
rect 145076 234892 145162 234956
rect 144926 234806 145162 234892
rect 151918 234956 152154 235042
rect 151918 234892 152004 234956
rect 152004 234892 152068 234956
rect 152068 234892 152154 234956
rect 151918 234806 152154 234892
rect 187798 239716 188034 239802
rect 187798 239652 187884 239716
rect 187884 239652 187948 239716
rect 187948 239652 188034 239716
rect 187798 239566 188034 239652
rect 211166 239716 211402 239802
rect 211166 239652 211252 239716
rect 211252 239652 211316 239716
rect 211316 239652 211402 239716
rect 211166 239566 211402 239652
rect 169030 238206 169266 238442
rect 199942 238356 200178 238442
rect 199942 238292 200028 238356
rect 200028 238292 200092 238356
rect 200092 238292 200178 238356
rect 199942 238206 200178 238292
rect 168478 234806 168714 235042
rect 230854 239036 231090 239122
rect 230854 238972 230940 239036
rect 230940 238972 231004 239036
rect 231004 238972 231090 239036
rect 230854 238886 231090 238972
rect 231774 238356 232010 238442
rect 231774 238292 231860 238356
rect 231860 238292 231924 238356
rect 231924 238292 232010 238356
rect 231774 238206 232010 238292
rect 183750 236996 183986 237082
rect 183750 236932 183836 236996
rect 183836 236932 183900 236996
rect 183900 236932 183986 236996
rect 183750 236846 183986 236932
rect 207118 234956 207354 235042
rect 207118 234892 207204 234956
rect 207204 234892 207268 234956
rect 207268 234892 207354 234956
rect 207118 234806 207354 234892
rect 231774 234956 232010 235042
rect 231774 234892 231860 234956
rect 231860 234892 231924 234956
rect 231924 234892 232010 234956
rect 231774 234806 232010 234892
rect 234718 234956 234954 235042
rect 234718 234892 234804 234956
rect 234804 234892 234868 234956
rect 234868 234892 234954 234956
rect 234718 234806 234954 234892
rect 228830 217126 229066 217362
rect 148606 216596 148842 216682
rect 148606 216532 148692 216596
rect 148692 216532 148756 216596
rect 148756 216532 148842 216596
rect 148606 216446 148842 216532
rect 177494 216596 177730 216682
rect 177494 216532 177580 216596
rect 177580 216532 177644 216596
rect 177644 216532 177730 216596
rect 177494 216446 177730 216532
rect 164798 215086 165034 215322
rect 104506 213346 104742 213582
rect 198506 213346 198742 213582
rect 134622 205036 134858 205122
rect 134622 204972 134708 205036
rect 134708 204972 134772 205036
rect 134772 204972 134858 205036
rect 134622 204886 134858 204972
rect 84574 204428 84660 204442
rect 84660 204428 84724 204442
rect 84724 204428 84810 204442
rect 84574 204206 84810 204428
rect 137750 200956 137986 201042
rect 137750 200892 137836 200956
rect 137836 200892 137900 200956
rect 137900 200892 137986 200956
rect 137750 200806 137986 200892
rect 137934 198766 138170 199002
rect 89146 198028 89382 198264
rect 137934 194006 138170 194242
rect 104506 182710 104742 182946
rect 231774 207756 232010 207842
rect 231774 207692 231860 207756
rect 231860 207692 231924 207756
rect 231924 207692 232010 207756
rect 231774 207606 232010 207692
rect 230670 200806 230906 201042
rect 230670 198766 230906 199002
rect 183146 198028 183382 198264
rect 322670 297366 322906 297602
rect 322670 293436 322906 293522
rect 322670 293372 322756 293436
rect 322756 293372 322820 293436
rect 322820 293372 322906 293436
rect 322670 293286 322906 293372
rect 257718 291246 257954 291482
rect 263606 291396 263842 291482
rect 263606 291332 263692 291396
rect 263692 291332 263756 291396
rect 263756 291332 263842 291396
rect 263606 291246 263842 291332
rect 272622 291246 272858 291482
rect 322670 291246 322906 291482
rect 277146 289936 277382 290172
rect 259374 289206 259610 289442
rect 353214 314366 353450 314602
rect 351742 285126 351978 285362
rect 246126 282406 246362 282642
rect 246126 279006 246362 279242
rect 292506 274618 292742 274854
rect 247782 262006 248018 262242
rect 238030 259966 238266 260202
rect 238030 257246 238266 257482
rect 236558 249086 236794 249322
rect 236926 245006 237162 245242
rect 238030 249086 238266 249322
rect 236926 242286 237162 242522
rect 261950 241606 262186 241842
rect 261582 240246 261818 240482
rect 238030 238206 238266 238442
rect 261950 238206 262186 238442
rect 248702 237526 248938 237762
rect 262870 239566 263106 239802
rect 249806 234806 250042 235042
rect 244286 234126 244522 234362
rect 245942 234276 246178 234362
rect 245942 234212 246028 234276
rect 246028 234212 246092 234276
rect 246092 234212 246178 234276
rect 245942 234126 246178 234212
rect 269126 233446 269362 233682
rect 259558 232916 259794 233002
rect 259558 232852 259644 232916
rect 259644 232852 259708 232916
rect 259708 232852 259794 232916
rect 259558 232766 259794 232852
rect 353582 285276 353818 285362
rect 353582 285212 353668 285276
rect 353668 285212 353732 285276
rect 353732 285212 353818 285276
rect 353582 285126 353818 285212
rect 412094 314366 412330 314602
rect 412094 308246 412330 308482
rect 412094 306206 412330 306442
rect 429390 306206 429626 306442
rect 435862 289936 436098 290172
rect 436182 289936 436418 290172
rect 436502 289936 436738 290172
rect 436822 289936 437058 290172
rect 437142 289936 437378 290172
rect 437462 289936 437698 290172
rect 437782 289936 438018 290172
rect 438102 289936 438338 290172
rect 438422 289936 438658 290172
rect 438742 289936 438978 290172
rect 439062 289936 439298 290172
rect 439382 289936 439618 290172
rect 412094 282406 412330 282642
rect 415038 278326 415274 278562
rect 435862 259300 436098 259536
rect 436182 259300 436418 259536
rect 436502 259300 436738 259536
rect 436822 259300 437058 259536
rect 437142 259300 437378 259536
rect 437462 259300 437698 259536
rect 437782 259300 438018 259536
rect 438102 259300 438338 259536
rect 438422 259300 438658 259536
rect 438742 259300 438978 259536
rect 439062 259300 439298 259536
rect 439382 259300 439618 259536
rect 355606 255886 355842 256122
rect 358550 255900 358786 256122
rect 358550 255886 358636 255900
rect 358636 255886 358700 255900
rect 358700 255886 358786 255900
rect 325062 249086 325298 249322
rect 303718 240396 303954 240482
rect 303718 240332 303804 240396
rect 303804 240332 303868 240396
rect 303868 240332 303954 240396
rect 303718 240246 303954 240332
rect 290470 239716 290706 239802
rect 290470 239652 290556 239716
rect 290556 239652 290620 239716
rect 290620 239652 290706 239716
rect 290470 239566 290706 239652
rect 325614 239566 325850 239802
rect 325246 239036 325482 239122
rect 325246 238972 325332 239036
rect 325332 238972 325396 239036
rect 325396 238972 325482 239036
rect 325246 238886 325482 238972
rect 286790 238356 287026 238442
rect 286790 238292 286876 238356
rect 286876 238292 286940 238356
rect 286940 238292 287026 238356
rect 286790 238206 287026 238292
rect 284214 234806 284450 235042
rect 297462 234806 297698 235042
rect 300958 234956 301194 235042
rect 300958 234892 301044 234956
rect 301044 234892 301108 234956
rect 301108 234892 301194 234956
rect 300958 234806 301194 234892
rect 285134 233446 285370 233682
rect 289918 233596 290154 233682
rect 289918 233532 290004 233596
rect 290004 233532 290068 233596
rect 290068 233532 290154 233596
rect 289918 233446 290154 233532
rect 282558 232916 282794 233002
rect 282558 232852 282644 232916
rect 282644 232852 282708 232916
rect 282708 232852 282794 232916
rect 282558 232766 282794 232852
rect 242630 217126 242866 217362
rect 258638 217126 258874 217362
rect 272622 217126 272858 217362
rect 322854 217140 323090 217362
rect 322854 217126 322940 217140
rect 322940 217126 323004 217140
rect 323004 217126 323090 217140
rect 336838 217126 337074 217362
rect 242630 216596 242866 216682
rect 242630 216532 242716 216596
rect 242716 216532 242780 216596
rect 242780 216532 242866 216596
rect 242630 216446 242866 216532
rect 258638 216596 258874 216682
rect 258638 216532 258724 216596
rect 258724 216532 258788 216596
rect 258788 216532 258874 216596
rect 258638 216446 258874 216532
rect 272622 216596 272858 216682
rect 272622 216532 272708 216596
rect 272708 216532 272772 216596
rect 272772 216532 272858 216596
rect 272622 216446 272858 216532
rect 336654 216596 336890 216682
rect 336654 216532 336740 216596
rect 336740 216532 336804 216596
rect 336804 216532 336890 216596
rect 336654 216446 336890 216532
rect 322854 215766 323090 216002
rect 292506 213346 292742 213582
rect 242446 207606 242682 207842
rect 236006 194686 236242 194922
rect 228646 194006 228882 194242
rect 322670 200956 322906 201042
rect 322670 200892 322756 200956
rect 322756 200892 322820 200956
rect 322820 200892 322906 200956
rect 322670 200806 322906 200892
rect 322670 198780 322906 199002
rect 322670 198766 322756 198780
rect 322756 198766 322820 198780
rect 322820 198766 322906 198780
rect 277146 198028 277382 198264
rect 322670 194836 322906 194922
rect 322670 194772 322756 194836
rect 322756 194772 322820 194836
rect 322820 194772 322906 194836
rect 322670 194686 322906 194772
rect 358550 249236 358786 249322
rect 358550 249172 358636 249236
rect 358636 249172 358700 249236
rect 358700 249172 358786 249236
rect 358550 249086 358786 249172
rect 360390 238886 360626 239122
rect 376882 228664 377118 228900
rect 435862 228664 436098 228900
rect 436182 228664 436418 228900
rect 436502 228664 436738 228900
rect 436822 228664 437058 228900
rect 437142 228664 437378 228900
rect 437462 228664 437698 228900
rect 437782 228664 438018 228900
rect 438102 228664 438338 228900
rect 438422 228664 438658 228900
rect 438742 228664 438978 228900
rect 439062 228664 439298 228900
rect 439382 228664 439618 228900
rect 358550 222036 358786 222122
rect 358550 221972 358636 222036
rect 358636 221972 358700 222036
rect 358700 221972 358786 222036
rect 358550 221886 358786 221972
rect 405838 222036 406074 222122
rect 405838 221972 405924 222036
rect 405924 221972 405988 222036
rect 405988 221972 406074 222036
rect 405838 221886 406074 221972
rect 352662 217126 352898 217362
rect 352662 216596 352898 216682
rect 352662 216532 352748 216596
rect 352748 216532 352812 216596
rect 352812 216532 352898 216596
rect 352662 216446 352898 216532
rect 357446 215916 357682 216002
rect 357446 215852 357532 215916
rect 357532 215852 357596 215916
rect 357596 215852 357682 215916
rect 357446 215766 357682 215852
rect 405838 215916 406074 216002
rect 405838 215852 405924 215916
rect 405924 215852 405988 215916
rect 405988 215852 406074 215916
rect 405838 215766 406074 215852
rect 435862 198028 436098 198264
rect 436182 198028 436418 198264
rect 436502 198028 436738 198264
rect 436822 198028 437058 198264
rect 437142 198028 437378 198264
rect 437462 198028 437698 198264
rect 437782 198028 438018 198264
rect 438102 198028 438338 198264
rect 438422 198028 438658 198264
rect 438742 198028 438978 198264
rect 439062 198028 439298 198264
rect 439382 198028 439618 198264
rect 198506 182710 198742 182946
rect 292506 182710 292742 182946
rect 174734 181086 174970 181322
rect 73534 168166 73770 168402
rect 5122 167392 5358 167628
rect 5442 167392 5678 167628
rect 5762 167392 5998 167628
rect 6082 167392 6318 167628
rect 6402 167392 6638 167628
rect 6722 167392 6958 167628
rect 7042 167392 7278 167628
rect 7362 167392 7598 167628
rect 7682 167392 7918 167628
rect 8002 167392 8238 167628
rect 8322 167392 8558 167628
rect 8642 167392 8878 167628
rect 49062 162268 49148 162282
rect 49148 162268 49212 162282
rect 49212 162268 49298 162282
rect 49062 162046 49298 162268
rect 49062 157966 49298 158202
rect 74638 162046 74874 162282
rect 74454 160686 74690 160922
rect 73718 157286 73954 157522
rect 49062 155396 49298 155482
rect 49062 155332 49148 155396
rect 49148 155332 49212 155396
rect 49212 155332 49298 155396
rect 49062 155246 49298 155332
rect 49062 153206 49298 153442
rect 49062 148446 49298 148682
rect 49062 145726 49298 145962
rect 73902 153206 74138 153442
rect 74270 151166 74506 151402
rect 76662 168166 76898 168402
rect 75558 155246 75794 155482
rect 74638 149806 74874 150042
rect 74270 149126 74506 149362
rect 5122 136756 5358 136992
rect 5442 136756 5678 136992
rect 5762 136756 5998 136992
rect 6082 136756 6318 136992
rect 6402 136756 6638 136992
rect 6722 136756 6958 136992
rect 7042 136756 7278 136992
rect 7362 136756 7598 136992
rect 7682 136756 7918 136992
rect 8002 136756 8238 136992
rect 8322 136756 8558 136992
rect 8642 136756 8878 136992
rect 5122 106120 5358 106356
rect 5442 106120 5678 106356
rect 5762 106120 5998 106356
rect 6082 106120 6318 106356
rect 6402 106120 6638 106356
rect 6722 106120 6958 106356
rect 7042 106120 7278 106356
rect 7362 106120 7598 106356
rect 7682 106120 7918 106356
rect 8002 106120 8238 106356
rect 8322 106120 8558 106356
rect 8642 106120 8878 106356
rect 75006 148446 75242 148682
rect 75190 145726 75426 145962
rect 75190 143686 75426 143922
rect 74822 143006 75058 143242
rect 74638 141646 74874 141882
rect 76662 157966 76898 158202
rect 76294 149806 76530 150042
rect 77582 148446 77818 148682
rect 77030 145046 77266 145282
rect 98742 145196 98978 145282
rect 98742 145132 98828 145196
rect 98828 145132 98892 145196
rect 98892 145132 98978 145196
rect 98742 145046 98978 145132
rect 77582 144366 77818 144602
rect 95062 144516 95298 144602
rect 95062 144452 95148 144516
rect 95148 144452 95212 144516
rect 95212 144452 95298 144516
rect 95062 144366 95298 144452
rect 77950 143686 78186 143922
rect 109598 143156 109834 143242
rect 109598 143092 109684 143156
rect 109684 143092 109748 143156
rect 109748 143092 109834 143156
rect 109598 143006 109834 143092
rect 137014 143006 137250 143242
rect 105918 141868 106004 141882
rect 106004 141868 106068 141882
rect 106068 141868 106154 141882
rect 105918 141646 106154 141868
rect 137382 141116 137618 141202
rect 137382 141052 137468 141116
rect 137468 141052 137532 141116
rect 137532 141052 137618 141116
rect 137382 140966 137618 141052
rect 137566 140436 137802 140522
rect 137566 140372 137652 140436
rect 137652 140372 137716 140436
rect 137716 140372 137802 140436
rect 137566 140286 137802 140372
rect 144006 162046 144242 162282
rect 144006 160006 144242 160242
rect 144006 151166 144242 151402
rect 144006 145046 144242 145282
rect 146950 143006 147186 143242
rect 148790 143006 149026 143242
rect 150262 143006 150498 143242
rect 146398 141116 146634 141202
rect 146398 141052 146484 141116
rect 146484 141052 146548 141116
rect 146548 141052 146634 141116
rect 146398 140966 146634 141052
rect 104506 121438 104742 121674
rect 144926 117166 145162 117402
rect 136830 116636 137066 116722
rect 136830 116572 136916 116636
rect 136916 116572 136980 116636
rect 136980 116572 137066 116636
rect 136830 116486 137066 116572
rect 138118 116636 138354 116722
rect 138118 116572 138204 116636
rect 138204 116572 138268 116636
rect 138268 116572 138354 116636
rect 138118 116486 138354 116572
rect 151918 141116 152154 141202
rect 151918 141052 152004 141116
rect 152004 141052 152068 141116
rect 152068 141052 152154 141116
rect 151918 140966 152154 141052
rect 271334 181766 271570 182002
rect 323406 181988 323492 182002
rect 323492 181988 323556 182002
rect 323556 181988 323642 182002
rect 323406 181766 323642 181988
rect 267470 181236 267706 181322
rect 267470 181172 267556 181236
rect 267556 181172 267620 181236
rect 267620 181172 267706 181236
rect 267470 181086 267706 181172
rect 323038 181086 323274 181322
rect 228646 180406 228882 180642
rect 169214 143686 169450 143922
rect 168478 140966 168714 141202
rect 148974 140286 149210 140522
rect 167558 140286 167794 140522
rect 187798 144516 188034 144602
rect 187798 144452 187884 144516
rect 187884 144452 187948 144516
rect 187948 144452 188034 144516
rect 187798 144366 188034 144452
rect 197182 140508 197268 140522
rect 197268 140508 197332 140522
rect 197332 140508 197418 140522
rect 197182 140286 197418 140508
rect 203070 143686 203306 143922
rect 237662 168166 237898 168402
rect 237294 166126 237530 166362
rect 237294 157286 237530 157522
rect 237294 150486 237530 150722
rect 237662 147766 237898 148002
rect 242630 168166 242866 168402
rect 243366 168166 243602 168402
rect 247046 168166 247282 168402
rect 238030 147086 238266 147322
rect 238030 146406 238266 146642
rect 231038 143156 231274 143242
rect 231038 143092 231124 143156
rect 231124 143092 231188 143156
rect 231188 143092 231274 143156
rect 231038 143006 231274 143092
rect 207486 141116 207722 141202
rect 207486 141052 207572 141116
rect 207572 141052 207636 141116
rect 207636 141052 207722 141116
rect 207486 140966 207722 141052
rect 231590 140286 231826 140522
rect 261582 144366 261818 144602
rect 242814 143006 243050 143242
rect 246310 143006 246546 143242
rect 247230 143006 247466 143242
rect 242446 142326 242682 142562
rect 249806 142476 250042 142562
rect 249806 142412 249892 142476
rect 249892 142412 249956 142476
rect 249956 142412 250042 142476
rect 249806 142326 250042 142412
rect 250358 142476 250594 142562
rect 250358 142412 250444 142476
rect 250444 142412 250508 142476
rect 250508 142412 250594 142476
rect 250358 142326 250594 142412
rect 255142 141646 255378 141882
rect 309790 179268 309876 179282
rect 309876 179268 309940 179282
rect 309940 179268 310026 179282
rect 309790 179046 310026 179268
rect 311078 179196 311314 179282
rect 311078 179132 311164 179196
rect 311164 179132 311228 179196
rect 311228 179132 311314 179196
rect 311078 179046 311314 179132
rect 312550 179268 312636 179282
rect 312636 179268 312700 179282
rect 312700 179268 312786 179282
rect 312550 179046 312786 179268
rect 313654 179196 313890 179282
rect 313654 179132 313740 179196
rect 313740 179132 313804 179196
rect 313804 179132 313890 179196
rect 313654 179046 313890 179132
rect 435862 167392 436098 167628
rect 436182 167392 436418 167628
rect 436502 167392 436738 167628
rect 436822 167392 437058 167628
rect 437142 167392 437378 167628
rect 437462 167392 437698 167628
rect 437782 167392 438018 167628
rect 438102 167392 438338 167628
rect 438422 167392 438658 167628
rect 438742 167392 438978 167628
rect 439062 167392 439298 167628
rect 439382 167392 439618 167628
rect 282374 143836 282610 143922
rect 282374 143772 282460 143836
rect 282460 143772 282524 143836
rect 282524 143772 282610 143836
rect 282374 143686 282610 143772
rect 283662 143836 283898 143922
rect 283662 143772 283748 143836
rect 283748 143772 283812 143836
rect 283812 143772 283898 143836
rect 283662 143686 283898 143772
rect 262870 143006 263106 143242
rect 245206 140286 245442 140522
rect 251278 140286 251514 140522
rect 262318 140286 262554 140522
rect 289918 142476 290154 142562
rect 289918 142412 290004 142476
rect 290004 142412 290068 142476
rect 290068 142412 290154 142476
rect 289918 142326 290154 142412
rect 182830 131446 183066 131682
rect 178598 123966 178834 124202
rect 148422 117846 148658 118082
rect 245758 123966 245994 124202
rect 245390 123286 245626 123522
rect 242630 122620 242866 122842
rect 242630 122606 242716 122620
rect 242716 122606 242780 122620
rect 242780 122606 242866 122620
rect 198506 121438 198742 121674
rect 198470 119886 198706 120122
rect 163694 115806 163930 116042
rect 147686 112556 147922 112642
rect 147686 112492 147772 112556
rect 147772 112492 147836 112556
rect 147836 112492 147922 112556
rect 147686 112406 147922 112492
rect 152102 112406 152338 112642
rect 84574 109700 84810 109922
rect 84574 109686 84660 109700
rect 84660 109686 84724 109700
rect 84724 109686 84810 109700
rect 134622 109836 134858 109922
rect 134622 109772 134708 109836
rect 134708 109772 134772 109836
rect 134772 109772 134858 109836
rect 134622 109686 134858 109772
rect 136830 107116 137066 107202
rect 136830 107052 136916 107116
rect 136916 107052 136980 107116
rect 136980 107052 137066 107116
rect 136830 106966 137066 107052
rect 89146 106120 89382 106356
rect 136830 100996 137066 101082
rect 136830 100932 136916 100996
rect 136916 100932 136980 100996
rect 136980 100932 137066 100996
rect 136830 100846 137066 100932
rect 148422 94726 148658 94962
rect 104506 90802 104742 91038
rect 245390 116486 245626 116722
rect 228646 115806 228882 116042
rect 230670 112406 230906 112642
rect 244102 112406 244338 112642
rect 240054 109836 240290 109922
rect 240054 109772 240140 109836
rect 240140 109772 240204 109836
rect 240204 109772 240290 109836
rect 240054 109686 240290 109772
rect 242078 109686 242314 109922
rect 164798 106966 165034 107202
rect 230854 106966 231090 107202
rect 183146 106120 183382 106356
rect 176022 100316 176258 100402
rect 176022 100252 176108 100316
rect 176108 100252 176172 100316
rect 176172 100252 176258 100316
rect 176022 100166 176258 100252
rect 176942 100316 177178 100402
rect 176942 100252 177028 100316
rect 177028 100252 177092 100316
rect 177092 100252 177178 100316
rect 228646 102206 228882 102442
rect 178046 100846 178282 101082
rect 228646 100860 228882 101082
rect 228646 100846 228732 100860
rect 228732 100846 228796 100860
rect 228796 100846 228882 100860
rect 176942 100166 177178 100252
rect 163694 96086 163930 96322
rect 178046 96086 178282 96322
rect 163694 95406 163930 95642
rect 178046 95406 178282 95642
rect 245758 113086 245994 113322
rect 249070 127366 249306 127602
rect 248518 126836 248754 126922
rect 302246 143836 302482 143922
rect 302246 143772 302332 143836
rect 302332 143772 302396 143836
rect 302396 143772 302482 143836
rect 302246 143686 302482 143772
rect 297646 143156 297882 143242
rect 297646 143092 297732 143156
rect 297732 143092 297796 143156
rect 297796 143092 297882 143156
rect 297646 143006 297882 143092
rect 301878 141116 302114 141202
rect 301878 141052 301964 141116
rect 301964 141052 302028 141116
rect 302028 141052 302114 141116
rect 301878 140966 302114 141052
rect 292494 131446 292730 131682
rect 248518 126772 248604 126836
rect 248604 126772 248668 126836
rect 248668 126772 248754 126836
rect 248518 126686 248754 126772
rect 322670 124116 322906 124202
rect 322670 124052 322756 124116
rect 322756 124052 322820 124116
rect 322820 124052 322906 124116
rect 322670 123966 322906 124052
rect 258638 122620 258874 122842
rect 258638 122606 258724 122620
rect 258724 122606 258788 122620
rect 258788 122606 258874 122620
rect 272622 122620 272858 122842
rect 272622 122606 272708 122620
rect 272708 122606 272772 122620
rect 272772 122606 272858 122620
rect 292506 121438 292742 121674
rect 322670 109836 322906 109922
rect 322670 109772 322756 109836
rect 322756 109772 322820 109836
rect 322820 109772 322906 109836
rect 322670 109686 322906 109772
rect 258822 106966 259058 107202
rect 277146 106120 277382 106356
rect 272622 100846 272858 101082
rect 323038 100996 323274 101082
rect 323038 100932 323124 100996
rect 323124 100932 323188 100996
rect 323188 100932 323274 100996
rect 323038 100846 323274 100932
rect 263054 100316 263290 100402
rect 322670 100388 322756 100402
rect 322756 100388 322820 100402
rect 322820 100388 322906 100402
rect 263054 100252 263140 100316
rect 263140 100252 263204 100316
rect 263204 100252 263290 100316
rect 263054 100166 263290 100252
rect 244654 98806 244890 99042
rect 322670 100166 322906 100388
rect 246126 98806 246362 99042
rect 264342 98806 264578 99042
rect 244102 96086 244338 96322
rect 5122 75484 5358 75720
rect 5442 75484 5678 75720
rect 5762 75484 5998 75720
rect 6082 75484 6318 75720
rect 6402 75484 6638 75720
rect 6722 75484 6958 75720
rect 7042 75484 7278 75720
rect 7362 75484 7598 75720
rect 7682 75484 7918 75720
rect 8002 75484 8238 75720
rect 8322 75484 8558 75720
rect 8642 75484 8878 75720
rect 72430 73646 72666 73882
rect 73350 61406 73586 61642
rect 73902 59366 74138 59602
rect 178598 94726 178834 94962
rect 229014 94876 229250 94962
rect 229014 94812 229100 94876
rect 229100 94812 229164 94876
rect 229164 94812 229250 94876
rect 229014 94726 229250 94812
rect 242446 94726 242682 94962
rect 164798 93366 165034 93602
rect 148422 73646 148658 73882
rect 74638 68886 74874 69122
rect 144742 63446 144978 63682
rect 75006 61406 75242 61642
rect 75374 59366 75610 59602
rect 73350 49166 73586 49402
rect 73166 48486 73402 48722
rect 74454 48486 74690 48722
rect 144742 54606 144978 54842
rect 144742 53926 144978 54162
rect 78870 53246 79106 53482
rect 113462 53246 113698 53482
rect 134070 53246 134306 53482
rect 102422 51356 102658 51442
rect 102422 51292 102508 51356
rect 102508 51292 102572 51356
rect 102572 51292 102658 51356
rect 102422 51206 102658 51292
rect 93590 50676 93826 50762
rect 93590 50612 93676 50676
rect 93676 50612 93740 50676
rect 93740 50612 93826 50676
rect 93590 50526 93826 50612
rect 87150 49316 87386 49402
rect 87150 49252 87236 49316
rect 87236 49252 87300 49316
rect 87300 49252 87386 49316
rect 87150 49166 87386 49252
rect 105182 49316 105418 49402
rect 105182 49252 105268 49316
rect 105268 49252 105332 49316
rect 105332 49252 105418 49316
rect 105182 49166 105418 49252
rect 87150 48486 87386 48722
rect 110334 47276 110570 47362
rect 110334 47212 110420 47276
rect 110420 47212 110484 47276
rect 110484 47212 110570 47276
rect 110334 47126 110570 47212
rect 107390 46446 107626 46682
rect 5122 44848 5358 45084
rect 5442 44848 5678 45084
rect 5762 44848 5998 45084
rect 6082 44848 6318 45084
rect 6402 44848 6638 45084
rect 6722 44848 6958 45084
rect 7042 44848 7278 45084
rect 7362 44848 7598 45084
rect 7682 44848 7918 45084
rect 8002 44848 8238 45084
rect 8322 44848 8558 45084
rect 8642 44848 8878 45084
rect 142718 51206 142954 51442
rect 144742 49166 144978 49402
rect 147870 49166 148106 49402
rect 167926 49166 168162 49402
rect 154678 48486 154914 48722
rect 167558 48486 167794 48722
rect 160014 47956 160250 48042
rect 198506 90802 198742 91038
rect 178598 86566 178834 86802
rect 245758 96086 245994 96322
rect 258638 95406 258874 95642
rect 272622 95406 272858 95642
rect 322670 94046 322906 94282
rect 292506 90802 292742 91038
rect 435862 136756 436098 136992
rect 436182 136756 436418 136992
rect 436502 136756 436738 136992
rect 436822 136756 437058 136992
rect 437142 136756 437378 136992
rect 437462 136756 437698 136992
rect 437782 136756 438018 136992
rect 438102 136756 438338 136992
rect 438422 136756 438658 136992
rect 438742 136756 438978 136992
rect 439062 136756 439298 136992
rect 439382 136756 439618 136992
rect 435862 106120 436098 106356
rect 436182 106120 436418 106356
rect 436502 106120 436738 106356
rect 436822 106120 437058 106356
rect 437142 106120 437378 106356
rect 437462 106120 437698 106356
rect 437782 106120 438018 106356
rect 438102 106120 438338 106356
rect 438422 106120 438658 106356
rect 438742 106120 438978 106356
rect 439062 106120 439298 106356
rect 439382 106120 439618 106356
rect 249070 88828 249156 88842
rect 249156 88828 249220 88842
rect 249220 88828 249306 88842
rect 249070 88606 249306 88828
rect 263790 88606 264026 88842
rect 245022 87926 245258 88162
rect 182462 85206 182698 85442
rect 252014 88076 252250 88162
rect 252014 88012 252100 88076
rect 252100 88012 252164 88076
rect 252164 88012 252250 88076
rect 252014 87926 252250 88012
rect 242630 73646 242866 73882
rect 237294 68886 237530 69122
rect 237294 59366 237530 59602
rect 238214 59366 238450 59602
rect 173814 53246 174050 53482
rect 207670 53246 207906 53482
rect 227910 53246 228146 53482
rect 187246 50676 187482 50762
rect 187246 50612 187332 50676
rect 187332 50612 187396 50676
rect 187396 50612 187482 50676
rect 187246 50526 187482 50612
rect 181726 49316 181962 49402
rect 181726 49252 181812 49316
rect 181812 49252 181876 49316
rect 181876 49252 181962 49316
rect 181726 49166 181962 49252
rect 160014 47892 160100 47956
rect 160100 47892 160164 47956
rect 160164 47892 160250 47956
rect 160014 47806 160250 47892
rect 169030 47806 169266 48042
rect 191294 48486 191530 48722
rect 182094 47956 182330 48042
rect 182094 47892 182180 47956
rect 182180 47892 182244 47956
rect 182244 47892 182330 47956
rect 182094 47806 182330 47892
rect 158910 47126 159146 47362
rect 162774 47276 163010 47362
rect 162774 47212 162860 47276
rect 162860 47212 162924 47276
rect 162924 47212 163010 47276
rect 162774 47126 163010 47212
rect 157438 46446 157674 46682
rect 204174 49316 204410 49402
rect 204174 49252 204260 49316
rect 204260 49252 204324 49316
rect 204324 49252 204410 49316
rect 204174 49166 204410 49252
rect 180990 46596 181226 46682
rect 180990 46532 181076 46596
rect 181076 46532 181140 46596
rect 181140 46532 181226 46596
rect 180990 46446 181226 46532
rect 199574 46446 199810 46682
rect 237478 50526 237714 50762
rect 238214 50526 238450 50762
rect 248518 48486 248754 48722
rect 253854 47956 254090 48042
rect 253854 47892 253940 47956
rect 253940 47892 254004 47956
rect 254004 47892 254090 47956
rect 253854 47806 254090 47892
rect 261398 47806 261634 48042
rect 248518 47276 248754 47362
rect 248518 47212 248604 47276
rect 248604 47212 248668 47276
rect 248668 47212 248754 47276
rect 248518 47126 248754 47212
rect 262318 49166 262554 49402
rect 263238 49846 263474 50082
rect 252566 46446 252802 46682
rect 260294 46596 260530 46682
rect 260294 46532 260380 46596
rect 260380 46532 260444 46596
rect 260444 46532 260530 46596
rect 260294 46446 260530 46532
rect 261766 46446 262002 46682
rect 266550 53246 266786 53482
rect 301510 53246 301746 53482
rect 280350 50676 280586 50762
rect 280350 50612 280436 50676
rect 280436 50612 280500 50676
rect 280500 50612 280586 50676
rect 280350 50526 280586 50612
rect 274830 49996 275066 50082
rect 263790 48486 264026 48722
rect 274830 49932 274916 49996
rect 274916 49932 274980 49996
rect 274980 49932 275066 49996
rect 274830 49846 275066 49932
rect 274830 49316 275066 49402
rect 274830 49252 274916 49316
rect 274916 49252 274980 49316
rect 274980 49252 275066 49316
rect 274830 49166 275066 49252
rect 274830 47956 275066 48042
rect 274830 47892 274916 47956
rect 274916 47892 274980 47956
rect 274980 47892 275066 47956
rect 274830 47806 275066 47892
rect 263790 47348 263876 47362
rect 263876 47348 263940 47362
rect 263940 47348 264026 47362
rect 263790 47126 264026 47348
rect 275750 46596 275986 46682
rect 275750 46532 275836 46596
rect 275836 46532 275900 46596
rect 275900 46532 275986 46596
rect 275750 46446 275986 46532
rect 321750 53246 321986 53482
rect 435862 75484 436098 75720
rect 436182 75484 436418 75720
rect 436502 75484 436738 75720
rect 436822 75484 437058 75720
rect 437142 75484 437378 75720
rect 437462 75484 437698 75720
rect 437782 75484 438018 75720
rect 438102 75484 438338 75720
rect 438422 75484 438658 75720
rect 438742 75484 438978 75720
rect 439062 75484 439298 75720
rect 439382 75484 439618 75720
rect 435862 44848 436098 45084
rect 436182 44848 436418 45084
rect 436502 44848 436738 45084
rect 436822 44848 437058 45084
rect 437142 44848 437378 45084
rect 437462 44848 437698 45084
rect 437782 44848 438018 45084
rect 438102 44848 438338 45084
rect 438422 44848 438658 45084
rect 438742 44848 438978 45084
rect 439062 44848 439298 45084
rect 439382 44848 439618 45084
rect 5122 14212 5358 14448
rect 5442 14212 5678 14448
rect 5762 14212 5998 14448
rect 6082 14212 6318 14448
rect 6402 14212 6638 14448
rect 6722 14212 6958 14448
rect 7042 14212 7278 14448
rect 7362 14212 7598 14448
rect 7682 14212 7918 14448
rect 8002 14212 8238 14448
rect 8322 14212 8558 14448
rect 8642 14212 8878 14448
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 435862 14212 436098 14448
rect 436182 14212 436418 14448
rect 436502 14212 436738 14448
rect 436822 14212 437058 14448
rect 437142 14212 437378 14448
rect 437462 14212 437698 14448
rect 437782 14212 438018 14448
rect 438102 14212 438338 14448
rect 438422 14212 438658 14448
rect 438742 14212 438978 14448
rect 439062 14212 439298 14448
rect 439382 14212 439618 14448
rect 435862 8642 436098 8878
rect 436182 8642 436418 8878
rect 436502 8642 436738 8878
rect 436822 8642 437058 8878
rect 437142 8642 437378 8878
rect 437462 8642 437698 8878
rect 437782 8642 438018 8878
rect 438102 8642 438338 8878
rect 438422 8642 438658 8878
rect 438742 8642 438978 8878
rect 439062 8642 439298 8878
rect 439382 8642 439618 8878
rect 435862 8322 436098 8558
rect 436182 8322 436418 8558
rect 436502 8322 436738 8558
rect 436822 8322 437058 8558
rect 437142 8322 437378 8558
rect 437462 8322 437698 8558
rect 437782 8322 438018 8558
rect 438102 8322 438338 8558
rect 438422 8322 438658 8558
rect 438742 8322 438978 8558
rect 439062 8322 439298 8558
rect 439382 8322 439618 8558
rect 435862 8002 436098 8238
rect 436182 8002 436418 8238
rect 436502 8002 436738 8238
rect 436822 8002 437058 8238
rect 437142 8002 437378 8238
rect 437462 8002 437698 8238
rect 437782 8002 438018 8238
rect 438102 8002 438338 8238
rect 438422 8002 438658 8238
rect 438742 8002 438978 8238
rect 439062 8002 439298 8238
rect 439382 8002 439618 8238
rect 435862 7682 436098 7918
rect 436182 7682 436418 7918
rect 436502 7682 436738 7918
rect 436822 7682 437058 7918
rect 437142 7682 437378 7918
rect 437462 7682 437698 7918
rect 437782 7682 438018 7918
rect 438102 7682 438338 7918
rect 438422 7682 438658 7918
rect 438742 7682 438978 7918
rect 439062 7682 439298 7918
rect 439382 7682 439618 7918
rect 435862 7362 436098 7598
rect 436182 7362 436418 7598
rect 436502 7362 436738 7598
rect 436822 7362 437058 7598
rect 437142 7362 437378 7598
rect 437462 7362 437698 7598
rect 437782 7362 438018 7598
rect 438102 7362 438338 7598
rect 438422 7362 438658 7598
rect 438742 7362 438978 7598
rect 439062 7362 439298 7598
rect 439382 7362 439618 7598
rect 435862 7042 436098 7278
rect 436182 7042 436418 7278
rect 436502 7042 436738 7278
rect 436822 7042 437058 7278
rect 437142 7042 437378 7278
rect 437462 7042 437698 7278
rect 437782 7042 438018 7278
rect 438102 7042 438338 7278
rect 438422 7042 438658 7278
rect 438742 7042 438978 7278
rect 439062 7042 439298 7278
rect 439382 7042 439618 7278
rect 435862 6722 436098 6958
rect 436182 6722 436418 6958
rect 436502 6722 436738 6958
rect 436822 6722 437058 6958
rect 437142 6722 437378 6958
rect 437462 6722 437698 6958
rect 437782 6722 438018 6958
rect 438102 6722 438338 6958
rect 438422 6722 438658 6958
rect 438742 6722 438978 6958
rect 439062 6722 439298 6958
rect 439382 6722 439618 6958
rect 435862 6402 436098 6638
rect 436182 6402 436418 6638
rect 436502 6402 436738 6638
rect 436822 6402 437058 6638
rect 437142 6402 437378 6638
rect 437462 6402 437698 6638
rect 437782 6402 438018 6638
rect 438102 6402 438338 6638
rect 438422 6402 438658 6638
rect 438742 6402 438978 6638
rect 439062 6402 439298 6638
rect 439382 6402 439618 6638
rect 435862 6082 436098 6318
rect 436182 6082 436418 6318
rect 436502 6082 436738 6318
rect 436822 6082 437058 6318
rect 437142 6082 437378 6318
rect 437462 6082 437698 6318
rect 437782 6082 438018 6318
rect 438102 6082 438338 6318
rect 438422 6082 438658 6318
rect 438742 6082 438978 6318
rect 439062 6082 439298 6318
rect 439382 6082 439618 6318
rect 435862 5762 436098 5998
rect 436182 5762 436418 5998
rect 436502 5762 436738 5998
rect 436822 5762 437058 5998
rect 437142 5762 437378 5998
rect 437462 5762 437698 5998
rect 437782 5762 438018 5998
rect 438102 5762 438338 5998
rect 438422 5762 438658 5998
rect 438742 5762 438978 5998
rect 439062 5762 439298 5998
rect 439382 5762 439618 5998
rect 435862 5442 436098 5678
rect 436182 5442 436418 5678
rect 436502 5442 436738 5678
rect 436822 5442 437058 5678
rect 437142 5442 437378 5678
rect 437462 5442 437698 5678
rect 437782 5442 438018 5678
rect 438102 5442 438338 5678
rect 438422 5442 438658 5678
rect 438742 5442 438978 5678
rect 439062 5442 439298 5678
rect 439382 5442 439618 5678
rect 435862 5122 436098 5358
rect 436182 5122 436418 5358
rect 436502 5122 436738 5358
rect 436822 5122 437058 5358
rect 437142 5122 437378 5358
rect 437462 5122 437698 5358
rect 437782 5122 438018 5358
rect 438102 5122 438338 5358
rect 438422 5122 438658 5358
rect 438742 5122 438978 5358
rect 439062 5122 439298 5358
rect 439382 5122 439618 5358
rect 440862 366526 441098 366762
rect 441182 366526 441418 366762
rect 441502 366526 441738 366762
rect 441822 366526 442058 366762
rect 442142 366526 442378 366762
rect 442462 366526 442698 366762
rect 442782 366526 443018 366762
rect 443102 366526 443338 366762
rect 443422 366526 443658 366762
rect 443742 366526 443978 366762
rect 444062 366526 444298 366762
rect 444382 366526 444618 366762
rect 440862 335890 441098 336126
rect 441182 335890 441418 336126
rect 441502 335890 441738 336126
rect 441822 335890 442058 336126
rect 442142 335890 442378 336126
rect 442462 335890 442698 336126
rect 442782 335890 443018 336126
rect 443102 335890 443338 336126
rect 443422 335890 443658 336126
rect 443742 335890 443978 336126
rect 444062 335890 444298 336126
rect 444382 335890 444618 336126
rect 440862 305254 441098 305490
rect 441182 305254 441418 305490
rect 441502 305254 441738 305490
rect 441822 305254 442058 305490
rect 442142 305254 442378 305490
rect 442462 305254 442698 305490
rect 442782 305254 443018 305490
rect 443102 305254 443338 305490
rect 443422 305254 443658 305490
rect 443742 305254 443978 305490
rect 444062 305254 444298 305490
rect 444382 305254 444618 305490
rect 440862 274618 441098 274854
rect 441182 274618 441418 274854
rect 441502 274618 441738 274854
rect 441822 274618 442058 274854
rect 442142 274618 442378 274854
rect 442462 274618 442698 274854
rect 442782 274618 443018 274854
rect 443102 274618 443338 274854
rect 443422 274618 443658 274854
rect 443742 274618 443978 274854
rect 444062 274618 444298 274854
rect 444382 274618 444618 274854
rect 440862 243982 441098 244218
rect 441182 243982 441418 244218
rect 441502 243982 441738 244218
rect 441822 243982 442058 244218
rect 442142 243982 442378 244218
rect 442462 243982 442698 244218
rect 442782 243982 443018 244218
rect 443102 243982 443338 244218
rect 443422 243982 443658 244218
rect 443742 243982 443978 244218
rect 444062 243982 444298 244218
rect 444382 243982 444618 244218
rect 440862 213346 441098 213582
rect 441182 213346 441418 213582
rect 441502 213346 441738 213582
rect 441822 213346 442058 213582
rect 442142 213346 442378 213582
rect 442462 213346 442698 213582
rect 442782 213346 443018 213582
rect 443102 213346 443338 213582
rect 443422 213346 443658 213582
rect 443742 213346 443978 213582
rect 444062 213346 444298 213582
rect 444382 213346 444618 213582
rect 440862 182710 441098 182946
rect 441182 182710 441418 182946
rect 441502 182710 441738 182946
rect 441822 182710 442058 182946
rect 442142 182710 442378 182946
rect 442462 182710 442698 182946
rect 442782 182710 443018 182946
rect 443102 182710 443338 182946
rect 443422 182710 443658 182946
rect 443742 182710 443978 182946
rect 444062 182710 444298 182946
rect 444382 182710 444618 182946
rect 440862 152074 441098 152310
rect 441182 152074 441418 152310
rect 441502 152074 441738 152310
rect 441822 152074 442058 152310
rect 442142 152074 442378 152310
rect 442462 152074 442698 152310
rect 442782 152074 443018 152310
rect 443102 152074 443338 152310
rect 443422 152074 443658 152310
rect 443742 152074 443978 152310
rect 444062 152074 444298 152310
rect 444382 152074 444618 152310
rect 440862 121438 441098 121674
rect 441182 121438 441418 121674
rect 441502 121438 441738 121674
rect 441822 121438 442058 121674
rect 442142 121438 442378 121674
rect 442462 121438 442698 121674
rect 442782 121438 443018 121674
rect 443102 121438 443338 121674
rect 443422 121438 443658 121674
rect 443742 121438 443978 121674
rect 444062 121438 444298 121674
rect 444382 121438 444618 121674
rect 440862 90802 441098 91038
rect 441182 90802 441418 91038
rect 441502 90802 441738 91038
rect 441822 90802 442058 91038
rect 442142 90802 442378 91038
rect 442462 90802 442698 91038
rect 442782 90802 443018 91038
rect 443102 90802 443338 91038
rect 443422 90802 443658 91038
rect 443742 90802 443978 91038
rect 444062 90802 444298 91038
rect 444382 90802 444618 91038
rect 440862 60166 441098 60402
rect 441182 60166 441418 60402
rect 441502 60166 441738 60402
rect 441822 60166 442058 60402
rect 442142 60166 442378 60402
rect 442462 60166 442698 60402
rect 442782 60166 443018 60402
rect 443102 60166 443338 60402
rect 443422 60166 443658 60402
rect 443742 60166 443978 60402
rect 444062 60166 444298 60402
rect 444382 60166 444618 60402
rect 440862 29530 441098 29766
rect 441182 29530 441418 29766
rect 441502 29530 441738 29766
rect 441822 29530 442058 29766
rect 442142 29530 442378 29766
rect 442462 29530 442698 29766
rect 442782 29530 443018 29766
rect 443102 29530 443338 29766
rect 443422 29530 443658 29766
rect 443742 29530 443978 29766
rect 444062 29530 444298 29766
rect 444382 29530 444618 29766
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 440862 3642 441098 3878
rect 441182 3642 441418 3878
rect 441502 3642 441738 3878
rect 441822 3642 442058 3878
rect 442142 3642 442378 3878
rect 442462 3642 442698 3878
rect 442782 3642 443018 3878
rect 443102 3642 443338 3878
rect 443422 3642 443658 3878
rect 443742 3642 443978 3878
rect 444062 3642 444298 3878
rect 444382 3642 444618 3878
rect 440862 3322 441098 3558
rect 441182 3322 441418 3558
rect 441502 3322 441738 3558
rect 441822 3322 442058 3558
rect 442142 3322 442378 3558
rect 442462 3322 442698 3558
rect 442782 3322 443018 3558
rect 443102 3322 443338 3558
rect 443422 3322 443658 3558
rect 443742 3322 443978 3558
rect 444062 3322 444298 3558
rect 444382 3322 444618 3558
rect 440862 3002 441098 3238
rect 441182 3002 441418 3238
rect 441502 3002 441738 3238
rect 441822 3002 442058 3238
rect 442142 3002 442378 3238
rect 442462 3002 442698 3238
rect 442782 3002 443018 3238
rect 443102 3002 443338 3238
rect 443422 3002 443658 3238
rect 443742 3002 443978 3238
rect 444062 3002 444298 3238
rect 444382 3002 444618 3238
rect 440862 2682 441098 2918
rect 441182 2682 441418 2918
rect 441502 2682 441738 2918
rect 441822 2682 442058 2918
rect 442142 2682 442378 2918
rect 442462 2682 442698 2918
rect 442782 2682 443018 2918
rect 443102 2682 443338 2918
rect 443422 2682 443658 2918
rect 443742 2682 443978 2918
rect 444062 2682 444298 2918
rect 444382 2682 444618 2918
rect 440862 2362 441098 2598
rect 441182 2362 441418 2598
rect 441502 2362 441738 2598
rect 441822 2362 442058 2598
rect 442142 2362 442378 2598
rect 442462 2362 442698 2598
rect 442782 2362 443018 2598
rect 443102 2362 443338 2598
rect 443422 2362 443658 2598
rect 443742 2362 443978 2598
rect 444062 2362 444298 2598
rect 444382 2362 444618 2598
rect 440862 2042 441098 2278
rect 441182 2042 441418 2278
rect 441502 2042 441738 2278
rect 441822 2042 442058 2278
rect 442142 2042 442378 2278
rect 442462 2042 442698 2278
rect 442782 2042 443018 2278
rect 443102 2042 443338 2278
rect 443422 2042 443658 2278
rect 443742 2042 443978 2278
rect 444062 2042 444298 2278
rect 444382 2042 444618 2278
rect 440862 1722 441098 1958
rect 441182 1722 441418 1958
rect 441502 1722 441738 1958
rect 441822 1722 442058 1958
rect 442142 1722 442378 1958
rect 442462 1722 442698 1958
rect 442782 1722 443018 1958
rect 443102 1722 443338 1958
rect 443422 1722 443658 1958
rect 443742 1722 443978 1958
rect 444062 1722 444298 1958
rect 444382 1722 444618 1958
rect 440862 1402 441098 1638
rect 441182 1402 441418 1638
rect 441502 1402 441738 1638
rect 441822 1402 442058 1638
rect 442142 1402 442378 1638
rect 442462 1402 442698 1638
rect 442782 1402 443018 1638
rect 443102 1402 443338 1638
rect 443422 1402 443658 1638
rect 443742 1402 443978 1638
rect 444062 1402 444298 1638
rect 444382 1402 444618 1638
rect 440862 1082 441098 1318
rect 441182 1082 441418 1318
rect 441502 1082 441738 1318
rect 441822 1082 442058 1318
rect 442142 1082 442378 1318
rect 442462 1082 442698 1318
rect 442782 1082 443018 1318
rect 443102 1082 443338 1318
rect 443422 1082 443658 1318
rect 443742 1082 443978 1318
rect 444062 1082 444298 1318
rect 444382 1082 444618 1318
rect 440862 762 441098 998
rect 441182 762 441418 998
rect 441502 762 441738 998
rect 441822 762 442058 998
rect 442142 762 442378 998
rect 442462 762 442698 998
rect 442782 762 443018 998
rect 443102 762 443338 998
rect 443422 762 443658 998
rect 443742 762 443978 998
rect 444062 762 444298 998
rect 444382 762 444618 998
rect 440862 442 441098 678
rect 441182 442 441418 678
rect 441502 442 441738 678
rect 441822 442 442058 678
rect 442142 442 442378 678
rect 442462 442 442698 678
rect 442782 442 443018 678
rect 443102 442 443338 678
rect 443422 442 443658 678
rect 443742 442 443978 678
rect 444062 442 444298 678
rect 444382 442 444618 678
rect 440862 122 441098 358
rect 441182 122 441418 358
rect 441502 122 441738 358
rect 441822 122 442058 358
rect 442142 122 442378 358
rect 442462 122 442698 358
rect 442782 122 443018 358
rect 443102 122 443338 358
rect 443422 122 443658 358
rect 443742 122 443978 358
rect 444062 122 444298 358
rect 444382 122 444618 358
<< metal5 >>
rect 0 405398 444740 405520
rect 0 405162 122 405398
rect 358 405162 442 405398
rect 678 405162 762 405398
rect 998 405162 1082 405398
rect 1318 405162 1402 405398
rect 1638 405162 1722 405398
rect 1958 405162 2042 405398
rect 2278 405162 2362 405398
rect 2598 405162 2682 405398
rect 2918 405162 3002 405398
rect 3238 405162 3322 405398
rect 3558 405162 3642 405398
rect 3878 405162 440862 405398
rect 441098 405162 441182 405398
rect 441418 405162 441502 405398
rect 441738 405162 441822 405398
rect 442058 405162 442142 405398
rect 442378 405162 442462 405398
rect 442698 405162 442782 405398
rect 443018 405162 443102 405398
rect 443338 405162 443422 405398
rect 443658 405162 443742 405398
rect 443978 405162 444062 405398
rect 444298 405162 444382 405398
rect 444618 405162 444740 405398
rect 0 405078 444740 405162
rect 0 404842 122 405078
rect 358 404842 442 405078
rect 678 404842 762 405078
rect 998 404842 1082 405078
rect 1318 404842 1402 405078
rect 1638 404842 1722 405078
rect 1958 404842 2042 405078
rect 2278 404842 2362 405078
rect 2598 404842 2682 405078
rect 2918 404842 3002 405078
rect 3238 404842 3322 405078
rect 3558 404842 3642 405078
rect 3878 404842 440862 405078
rect 441098 404842 441182 405078
rect 441418 404842 441502 405078
rect 441738 404842 441822 405078
rect 442058 404842 442142 405078
rect 442378 404842 442462 405078
rect 442698 404842 442782 405078
rect 443018 404842 443102 405078
rect 443338 404842 443422 405078
rect 443658 404842 443742 405078
rect 443978 404842 444062 405078
rect 444298 404842 444382 405078
rect 444618 404842 444740 405078
rect 0 404758 444740 404842
rect 0 404522 122 404758
rect 358 404522 442 404758
rect 678 404522 762 404758
rect 998 404522 1082 404758
rect 1318 404522 1402 404758
rect 1638 404522 1722 404758
rect 1958 404522 2042 404758
rect 2278 404522 2362 404758
rect 2598 404522 2682 404758
rect 2918 404522 3002 404758
rect 3238 404522 3322 404758
rect 3558 404522 3642 404758
rect 3878 404522 440862 404758
rect 441098 404522 441182 404758
rect 441418 404522 441502 404758
rect 441738 404522 441822 404758
rect 442058 404522 442142 404758
rect 442378 404522 442462 404758
rect 442698 404522 442782 404758
rect 443018 404522 443102 404758
rect 443338 404522 443422 404758
rect 443658 404522 443742 404758
rect 443978 404522 444062 404758
rect 444298 404522 444382 404758
rect 444618 404522 444740 404758
rect 0 404438 444740 404522
rect 0 404202 122 404438
rect 358 404202 442 404438
rect 678 404202 762 404438
rect 998 404202 1082 404438
rect 1318 404202 1402 404438
rect 1638 404202 1722 404438
rect 1958 404202 2042 404438
rect 2278 404202 2362 404438
rect 2598 404202 2682 404438
rect 2918 404202 3002 404438
rect 3238 404202 3322 404438
rect 3558 404202 3642 404438
rect 3878 404202 440862 404438
rect 441098 404202 441182 404438
rect 441418 404202 441502 404438
rect 441738 404202 441822 404438
rect 442058 404202 442142 404438
rect 442378 404202 442462 404438
rect 442698 404202 442782 404438
rect 443018 404202 443102 404438
rect 443338 404202 443422 404438
rect 443658 404202 443742 404438
rect 443978 404202 444062 404438
rect 444298 404202 444382 404438
rect 444618 404202 444740 404438
rect 0 404118 444740 404202
rect 0 403882 122 404118
rect 358 403882 442 404118
rect 678 403882 762 404118
rect 998 403882 1082 404118
rect 1318 403882 1402 404118
rect 1638 403882 1722 404118
rect 1958 403882 2042 404118
rect 2278 403882 2362 404118
rect 2598 403882 2682 404118
rect 2918 403882 3002 404118
rect 3238 403882 3322 404118
rect 3558 403882 3642 404118
rect 3878 403882 440862 404118
rect 441098 403882 441182 404118
rect 441418 403882 441502 404118
rect 441738 403882 441822 404118
rect 442058 403882 442142 404118
rect 442378 403882 442462 404118
rect 442698 403882 442782 404118
rect 443018 403882 443102 404118
rect 443338 403882 443422 404118
rect 443658 403882 443742 404118
rect 443978 403882 444062 404118
rect 444298 403882 444382 404118
rect 444618 403882 444740 404118
rect 0 403798 444740 403882
rect 0 403562 122 403798
rect 358 403562 442 403798
rect 678 403562 762 403798
rect 998 403562 1082 403798
rect 1318 403562 1402 403798
rect 1638 403562 1722 403798
rect 1958 403562 2042 403798
rect 2278 403562 2362 403798
rect 2598 403562 2682 403798
rect 2918 403562 3002 403798
rect 3238 403562 3322 403798
rect 3558 403562 3642 403798
rect 3878 403562 440862 403798
rect 441098 403562 441182 403798
rect 441418 403562 441502 403798
rect 441738 403562 441822 403798
rect 442058 403562 442142 403798
rect 442378 403562 442462 403798
rect 442698 403562 442782 403798
rect 443018 403562 443102 403798
rect 443338 403562 443422 403798
rect 443658 403562 443742 403798
rect 443978 403562 444062 403798
rect 444298 403562 444382 403798
rect 444618 403562 444740 403798
rect 0 403478 444740 403562
rect 0 403242 122 403478
rect 358 403242 442 403478
rect 678 403242 762 403478
rect 998 403242 1082 403478
rect 1318 403242 1402 403478
rect 1638 403242 1722 403478
rect 1958 403242 2042 403478
rect 2278 403242 2362 403478
rect 2598 403242 2682 403478
rect 2918 403242 3002 403478
rect 3238 403242 3322 403478
rect 3558 403242 3642 403478
rect 3878 403242 440862 403478
rect 441098 403242 441182 403478
rect 441418 403242 441502 403478
rect 441738 403242 441822 403478
rect 442058 403242 442142 403478
rect 442378 403242 442462 403478
rect 442698 403242 442782 403478
rect 443018 403242 443102 403478
rect 443338 403242 443422 403478
rect 443658 403242 443742 403478
rect 443978 403242 444062 403478
rect 444298 403242 444382 403478
rect 444618 403242 444740 403478
rect 0 403158 444740 403242
rect 0 402922 122 403158
rect 358 402922 442 403158
rect 678 402922 762 403158
rect 998 402922 1082 403158
rect 1318 402922 1402 403158
rect 1638 402922 1722 403158
rect 1958 402922 2042 403158
rect 2278 402922 2362 403158
rect 2598 402922 2682 403158
rect 2918 402922 3002 403158
rect 3238 402922 3322 403158
rect 3558 402922 3642 403158
rect 3878 402922 440862 403158
rect 441098 402922 441182 403158
rect 441418 402922 441502 403158
rect 441738 402922 441822 403158
rect 442058 402922 442142 403158
rect 442378 402922 442462 403158
rect 442698 402922 442782 403158
rect 443018 402922 443102 403158
rect 443338 402922 443422 403158
rect 443658 402922 443742 403158
rect 443978 402922 444062 403158
rect 444298 402922 444382 403158
rect 444618 402922 444740 403158
rect 0 402838 444740 402922
rect 0 402602 122 402838
rect 358 402602 442 402838
rect 678 402602 762 402838
rect 998 402602 1082 402838
rect 1318 402602 1402 402838
rect 1638 402602 1722 402838
rect 1958 402602 2042 402838
rect 2278 402602 2362 402838
rect 2598 402602 2682 402838
rect 2918 402602 3002 402838
rect 3238 402602 3322 402838
rect 3558 402602 3642 402838
rect 3878 402602 440862 402838
rect 441098 402602 441182 402838
rect 441418 402602 441502 402838
rect 441738 402602 441822 402838
rect 442058 402602 442142 402838
rect 442378 402602 442462 402838
rect 442698 402602 442782 402838
rect 443018 402602 443102 402838
rect 443338 402602 443422 402838
rect 443658 402602 443742 402838
rect 443978 402602 444062 402838
rect 444298 402602 444382 402838
rect 444618 402602 444740 402838
rect 0 402518 444740 402602
rect 0 402282 122 402518
rect 358 402282 442 402518
rect 678 402282 762 402518
rect 998 402282 1082 402518
rect 1318 402282 1402 402518
rect 1638 402282 1722 402518
rect 1958 402282 2042 402518
rect 2278 402282 2362 402518
rect 2598 402282 2682 402518
rect 2918 402282 3002 402518
rect 3238 402282 3322 402518
rect 3558 402282 3642 402518
rect 3878 402282 440862 402518
rect 441098 402282 441182 402518
rect 441418 402282 441502 402518
rect 441738 402282 441822 402518
rect 442058 402282 442142 402518
rect 442378 402282 442462 402518
rect 442698 402282 442782 402518
rect 443018 402282 443102 402518
rect 443338 402282 443422 402518
rect 443658 402282 443742 402518
rect 443978 402282 444062 402518
rect 444298 402282 444382 402518
rect 444618 402282 444740 402518
rect 0 402198 444740 402282
rect 0 401962 122 402198
rect 358 401962 442 402198
rect 678 401962 762 402198
rect 998 401962 1082 402198
rect 1318 401962 1402 402198
rect 1638 401962 1722 402198
rect 1958 401962 2042 402198
rect 2278 401962 2362 402198
rect 2598 401962 2682 402198
rect 2918 401962 3002 402198
rect 3238 401962 3322 402198
rect 3558 401962 3642 402198
rect 3878 401962 440862 402198
rect 441098 401962 441182 402198
rect 441418 401962 441502 402198
rect 441738 401962 441822 402198
rect 442058 401962 442142 402198
rect 442378 401962 442462 402198
rect 442698 401962 442782 402198
rect 443018 401962 443102 402198
rect 443338 401962 443422 402198
rect 443658 401962 443742 402198
rect 443978 401962 444062 402198
rect 444298 401962 444382 402198
rect 444618 401962 444740 402198
rect 0 401878 444740 401962
rect 0 401642 122 401878
rect 358 401642 442 401878
rect 678 401642 762 401878
rect 998 401642 1082 401878
rect 1318 401642 1402 401878
rect 1638 401642 1722 401878
rect 1958 401642 2042 401878
rect 2278 401642 2362 401878
rect 2598 401642 2682 401878
rect 2918 401642 3002 401878
rect 3238 401642 3322 401878
rect 3558 401642 3642 401878
rect 3878 401642 440862 401878
rect 441098 401642 441182 401878
rect 441418 401642 441502 401878
rect 441738 401642 441822 401878
rect 442058 401642 442142 401878
rect 442378 401642 442462 401878
rect 442698 401642 442782 401878
rect 443018 401642 443102 401878
rect 443338 401642 443422 401878
rect 443658 401642 443742 401878
rect 443978 401642 444062 401878
rect 444298 401642 444382 401878
rect 444618 401642 444740 401878
rect 0 401520 444740 401642
rect 5000 400398 439740 400520
rect 5000 400162 5122 400398
rect 5358 400162 5442 400398
rect 5678 400162 5762 400398
rect 5998 400162 6082 400398
rect 6318 400162 6402 400398
rect 6638 400162 6722 400398
rect 6958 400162 7042 400398
rect 7278 400162 7362 400398
rect 7598 400162 7682 400398
rect 7918 400162 8002 400398
rect 8238 400162 8322 400398
rect 8558 400162 8642 400398
rect 8878 400162 435862 400398
rect 436098 400162 436182 400398
rect 436418 400162 436502 400398
rect 436738 400162 436822 400398
rect 437058 400162 437142 400398
rect 437378 400162 437462 400398
rect 437698 400162 437782 400398
rect 438018 400162 438102 400398
rect 438338 400162 438422 400398
rect 438658 400162 438742 400398
rect 438978 400162 439062 400398
rect 439298 400162 439382 400398
rect 439618 400162 439740 400398
rect 5000 400078 439740 400162
rect 5000 399842 5122 400078
rect 5358 399842 5442 400078
rect 5678 399842 5762 400078
rect 5998 399842 6082 400078
rect 6318 399842 6402 400078
rect 6638 399842 6722 400078
rect 6958 399842 7042 400078
rect 7278 399842 7362 400078
rect 7598 399842 7682 400078
rect 7918 399842 8002 400078
rect 8238 399842 8322 400078
rect 8558 399842 8642 400078
rect 8878 399842 435862 400078
rect 436098 399842 436182 400078
rect 436418 399842 436502 400078
rect 436738 399842 436822 400078
rect 437058 399842 437142 400078
rect 437378 399842 437462 400078
rect 437698 399842 437782 400078
rect 438018 399842 438102 400078
rect 438338 399842 438422 400078
rect 438658 399842 438742 400078
rect 438978 399842 439062 400078
rect 439298 399842 439382 400078
rect 439618 399842 439740 400078
rect 5000 399758 439740 399842
rect 5000 399522 5122 399758
rect 5358 399522 5442 399758
rect 5678 399522 5762 399758
rect 5998 399522 6082 399758
rect 6318 399522 6402 399758
rect 6638 399522 6722 399758
rect 6958 399522 7042 399758
rect 7278 399522 7362 399758
rect 7598 399522 7682 399758
rect 7918 399522 8002 399758
rect 8238 399522 8322 399758
rect 8558 399522 8642 399758
rect 8878 399522 435862 399758
rect 436098 399522 436182 399758
rect 436418 399522 436502 399758
rect 436738 399522 436822 399758
rect 437058 399522 437142 399758
rect 437378 399522 437462 399758
rect 437698 399522 437782 399758
rect 438018 399522 438102 399758
rect 438338 399522 438422 399758
rect 438658 399522 438742 399758
rect 438978 399522 439062 399758
rect 439298 399522 439382 399758
rect 439618 399522 439740 399758
rect 5000 399438 439740 399522
rect 5000 399202 5122 399438
rect 5358 399202 5442 399438
rect 5678 399202 5762 399438
rect 5998 399202 6082 399438
rect 6318 399202 6402 399438
rect 6638 399202 6722 399438
rect 6958 399202 7042 399438
rect 7278 399202 7362 399438
rect 7598 399202 7682 399438
rect 7918 399202 8002 399438
rect 8238 399202 8322 399438
rect 8558 399202 8642 399438
rect 8878 399202 435862 399438
rect 436098 399202 436182 399438
rect 436418 399202 436502 399438
rect 436738 399202 436822 399438
rect 437058 399202 437142 399438
rect 437378 399202 437462 399438
rect 437698 399202 437782 399438
rect 438018 399202 438102 399438
rect 438338 399202 438422 399438
rect 438658 399202 438742 399438
rect 438978 399202 439062 399438
rect 439298 399202 439382 399438
rect 439618 399202 439740 399438
rect 5000 399118 439740 399202
rect 5000 398882 5122 399118
rect 5358 398882 5442 399118
rect 5678 398882 5762 399118
rect 5998 398882 6082 399118
rect 6318 398882 6402 399118
rect 6638 398882 6722 399118
rect 6958 398882 7042 399118
rect 7278 398882 7362 399118
rect 7598 398882 7682 399118
rect 7918 398882 8002 399118
rect 8238 398882 8322 399118
rect 8558 398882 8642 399118
rect 8878 398882 435862 399118
rect 436098 398882 436182 399118
rect 436418 398882 436502 399118
rect 436738 398882 436822 399118
rect 437058 398882 437142 399118
rect 437378 398882 437462 399118
rect 437698 398882 437782 399118
rect 438018 398882 438102 399118
rect 438338 398882 438422 399118
rect 438658 398882 438742 399118
rect 438978 398882 439062 399118
rect 439298 398882 439382 399118
rect 439618 398882 439740 399118
rect 5000 398798 439740 398882
rect 5000 398562 5122 398798
rect 5358 398562 5442 398798
rect 5678 398562 5762 398798
rect 5998 398562 6082 398798
rect 6318 398562 6402 398798
rect 6638 398562 6722 398798
rect 6958 398562 7042 398798
rect 7278 398562 7362 398798
rect 7598 398562 7682 398798
rect 7918 398562 8002 398798
rect 8238 398562 8322 398798
rect 8558 398562 8642 398798
rect 8878 398562 435862 398798
rect 436098 398562 436182 398798
rect 436418 398562 436502 398798
rect 436738 398562 436822 398798
rect 437058 398562 437142 398798
rect 437378 398562 437462 398798
rect 437698 398562 437782 398798
rect 438018 398562 438102 398798
rect 438338 398562 438422 398798
rect 438658 398562 438742 398798
rect 438978 398562 439062 398798
rect 439298 398562 439382 398798
rect 439618 398562 439740 398798
rect 5000 398478 439740 398562
rect 5000 398242 5122 398478
rect 5358 398242 5442 398478
rect 5678 398242 5762 398478
rect 5998 398242 6082 398478
rect 6318 398242 6402 398478
rect 6638 398242 6722 398478
rect 6958 398242 7042 398478
rect 7278 398242 7362 398478
rect 7598 398242 7682 398478
rect 7918 398242 8002 398478
rect 8238 398242 8322 398478
rect 8558 398242 8642 398478
rect 8878 398242 435862 398478
rect 436098 398242 436182 398478
rect 436418 398242 436502 398478
rect 436738 398242 436822 398478
rect 437058 398242 437142 398478
rect 437378 398242 437462 398478
rect 437698 398242 437782 398478
rect 438018 398242 438102 398478
rect 438338 398242 438422 398478
rect 438658 398242 438742 398478
rect 438978 398242 439062 398478
rect 439298 398242 439382 398478
rect 439618 398242 439740 398478
rect 5000 398158 439740 398242
rect 5000 397922 5122 398158
rect 5358 397922 5442 398158
rect 5678 397922 5762 398158
rect 5998 397922 6082 398158
rect 6318 397922 6402 398158
rect 6638 397922 6722 398158
rect 6958 397922 7042 398158
rect 7278 397922 7362 398158
rect 7598 397922 7682 398158
rect 7918 397922 8002 398158
rect 8238 397922 8322 398158
rect 8558 397922 8642 398158
rect 8878 397922 435862 398158
rect 436098 397922 436182 398158
rect 436418 397922 436502 398158
rect 436738 397922 436822 398158
rect 437058 397922 437142 398158
rect 437378 397922 437462 398158
rect 437698 397922 437782 398158
rect 438018 397922 438102 398158
rect 438338 397922 438422 398158
rect 438658 397922 438742 398158
rect 438978 397922 439062 398158
rect 439298 397922 439382 398158
rect 439618 397922 439740 398158
rect 5000 397838 439740 397922
rect 5000 397602 5122 397838
rect 5358 397602 5442 397838
rect 5678 397602 5762 397838
rect 5998 397602 6082 397838
rect 6318 397602 6402 397838
rect 6638 397602 6722 397838
rect 6958 397602 7042 397838
rect 7278 397602 7362 397838
rect 7598 397602 7682 397838
rect 7918 397602 8002 397838
rect 8238 397602 8322 397838
rect 8558 397602 8642 397838
rect 8878 397602 435862 397838
rect 436098 397602 436182 397838
rect 436418 397602 436502 397838
rect 436738 397602 436822 397838
rect 437058 397602 437142 397838
rect 437378 397602 437462 397838
rect 437698 397602 437782 397838
rect 438018 397602 438102 397838
rect 438338 397602 438422 397838
rect 438658 397602 438742 397838
rect 438978 397602 439062 397838
rect 439298 397602 439382 397838
rect 439618 397602 439740 397838
rect 5000 397518 439740 397602
rect 5000 397282 5122 397518
rect 5358 397282 5442 397518
rect 5678 397282 5762 397518
rect 5998 397282 6082 397518
rect 6318 397282 6402 397518
rect 6638 397282 6722 397518
rect 6958 397282 7042 397518
rect 7278 397282 7362 397518
rect 7598 397282 7682 397518
rect 7918 397282 8002 397518
rect 8238 397282 8322 397518
rect 8558 397282 8642 397518
rect 8878 397282 435862 397518
rect 436098 397282 436182 397518
rect 436418 397282 436502 397518
rect 436738 397282 436822 397518
rect 437058 397282 437142 397518
rect 437378 397282 437462 397518
rect 437698 397282 437782 397518
rect 438018 397282 438102 397518
rect 438338 397282 438422 397518
rect 438658 397282 438742 397518
rect 438978 397282 439062 397518
rect 439298 397282 439382 397518
rect 439618 397282 439740 397518
rect 5000 397198 439740 397282
rect 5000 396962 5122 397198
rect 5358 396962 5442 397198
rect 5678 396962 5762 397198
rect 5998 396962 6082 397198
rect 6318 396962 6402 397198
rect 6638 396962 6722 397198
rect 6958 396962 7042 397198
rect 7278 396962 7362 397198
rect 7598 396962 7682 397198
rect 7918 396962 8002 397198
rect 8238 396962 8322 397198
rect 8558 396962 8642 397198
rect 8878 396962 435862 397198
rect 436098 396962 436182 397198
rect 436418 396962 436502 397198
rect 436738 396962 436822 397198
rect 437058 396962 437142 397198
rect 437378 396962 437462 397198
rect 437698 396962 437782 397198
rect 438018 396962 438102 397198
rect 438338 396962 438422 397198
rect 438658 396962 438742 397198
rect 438978 396962 439062 397198
rect 439298 396962 439382 397198
rect 439618 396962 439740 397198
rect 5000 396878 439740 396962
rect 5000 396642 5122 396878
rect 5358 396642 5442 396878
rect 5678 396642 5762 396878
rect 5998 396642 6082 396878
rect 6318 396642 6402 396878
rect 6638 396642 6722 396878
rect 6958 396642 7042 396878
rect 7278 396642 7362 396878
rect 7598 396642 7682 396878
rect 7918 396642 8002 396878
rect 8238 396642 8322 396878
rect 8558 396642 8642 396878
rect 8878 396642 435862 396878
rect 436098 396642 436182 396878
rect 436418 396642 436502 396878
rect 436738 396642 436822 396878
rect 437058 396642 437142 396878
rect 437378 396642 437462 396878
rect 437698 396642 437782 396878
rect 438018 396642 438102 396878
rect 438338 396642 438422 396878
rect 438658 396642 438742 396878
rect 438978 396642 439062 396878
rect 439298 396642 439382 396878
rect 439618 396642 439740 396878
rect 5000 396520 439740 396642
rect 0 382080 444740 382122
rect 0 381844 5122 382080
rect 5358 381844 5442 382080
rect 5678 381844 5762 382080
rect 5998 381844 6082 382080
rect 6318 381844 6402 382080
rect 6638 381844 6722 382080
rect 6958 381844 7042 382080
rect 7278 381844 7362 382080
rect 7598 381844 7682 382080
rect 7918 381844 8002 382080
rect 8238 381844 8322 382080
rect 8558 381844 8642 382080
rect 8878 381844 435862 382080
rect 436098 381844 436182 382080
rect 436418 381844 436502 382080
rect 436738 381844 436822 382080
rect 437058 381844 437142 382080
rect 437378 381844 437462 382080
rect 437698 381844 437782 382080
rect 438018 381844 438102 382080
rect 438338 381844 438422 382080
rect 438658 381844 438742 382080
rect 438978 381844 439062 382080
rect 439298 381844 439382 382080
rect 439618 381844 444740 382080
rect 0 381802 444740 381844
rect 0 366762 444740 366804
rect 0 366526 122 366762
rect 358 366526 442 366762
rect 678 366526 762 366762
rect 998 366526 1082 366762
rect 1318 366526 1402 366762
rect 1638 366526 1722 366762
rect 1958 366526 2042 366762
rect 2278 366526 2362 366762
rect 2598 366526 2682 366762
rect 2918 366526 3002 366762
rect 3238 366526 3322 366762
rect 3558 366526 3642 366762
rect 3878 366526 440862 366762
rect 441098 366526 441182 366762
rect 441418 366526 441502 366762
rect 441738 366526 441822 366762
rect 442058 366526 442142 366762
rect 442378 366526 442462 366762
rect 442698 366526 442782 366762
rect 443018 366526 443102 366762
rect 443338 366526 443422 366762
rect 443658 366526 443742 366762
rect 443978 366526 444062 366762
rect 444298 366526 444382 366762
rect 444618 366526 444740 366762
rect 0 366484 444740 366526
rect 332012 356082 341900 356124
rect 332012 355846 332054 356082
rect 332290 355846 341622 356082
rect 341858 355846 341900 356082
rect 332012 355804 341900 355846
rect 0 351444 444740 351486
rect 0 351208 5122 351444
rect 5358 351208 5442 351444
rect 5678 351208 5762 351444
rect 5998 351208 6082 351444
rect 6318 351208 6402 351444
rect 6638 351208 6722 351444
rect 6958 351208 7042 351444
rect 7278 351208 7362 351444
rect 7598 351208 7682 351444
rect 7918 351208 8002 351444
rect 8238 351208 8322 351444
rect 8558 351208 8642 351444
rect 8878 351208 435862 351444
rect 436098 351208 436182 351444
rect 436418 351208 436502 351444
rect 436738 351208 436822 351444
rect 437058 351208 437142 351444
rect 437378 351208 437462 351444
rect 437698 351208 437782 351444
rect 438018 351208 438102 351444
rect 438338 351208 438422 351444
rect 438658 351208 438742 351444
rect 438978 351208 439062 351444
rect 439298 351208 439382 351444
rect 439618 351208 444740 351444
rect 0 351166 444740 351208
rect 332012 349962 341348 350004
rect 332012 349726 332054 349962
rect 332290 349726 341348 349962
rect 332012 349684 341348 349726
rect 341028 339804 341348 349684
rect 341028 339484 341532 339804
rect 341212 338444 341532 339484
rect 341212 338124 341716 338444
rect 341396 337084 341716 338124
rect 341028 337042 341716 337084
rect 341028 336806 341070 337042
rect 341306 336806 341716 337042
rect 341028 336764 341716 336806
rect 0 336126 444740 336168
rect 0 335890 122 336126
rect 358 335890 442 336126
rect 678 335890 762 336126
rect 998 335890 1082 336126
rect 1318 335890 1402 336126
rect 1638 335890 1722 336126
rect 1958 335890 2042 336126
rect 2278 335890 2362 336126
rect 2598 335890 2682 336126
rect 2918 335890 3002 336126
rect 3238 335890 3322 336126
rect 3558 335890 3642 336126
rect 3878 335890 440862 336126
rect 441098 335890 441182 336126
rect 441418 335890 441502 336126
rect 441738 335890 441822 336126
rect 442058 335890 442142 336126
rect 442378 335890 442462 336126
rect 442698 335890 442782 336126
rect 443018 335890 443102 336126
rect 443338 335890 443422 336126
rect 443658 335890 443742 336126
rect 443978 335890 444062 336126
rect 444298 335890 444382 336126
rect 444618 335890 444740 336126
rect 0 335848 444740 335890
rect 336244 335002 341348 335044
rect 336244 334766 341070 335002
rect 341306 334766 341348 335002
rect 336244 334724 341348 334766
rect 137156 332282 201876 332324
rect 137156 332046 137198 332282
rect 137434 332046 201598 332282
rect 201834 332046 201876 332282
rect 137156 332004 201876 332046
rect 230812 332282 295716 332324
rect 230812 332046 230854 332282
rect 231090 332046 295438 332282
rect 295674 332046 295716 332282
rect 230812 332004 295716 332046
rect 158500 331602 158820 332004
rect 158500 331366 158542 331602
rect 158778 331366 158820 331602
rect 158500 331324 158820 331366
rect 252524 331602 252844 332004
rect 252524 331366 252566 331602
rect 252802 331366 252844 331602
rect 252524 331324 252844 331366
rect 336244 331602 336564 334724
rect 336244 331366 336286 331602
rect 336522 331366 336564 331602
rect 336244 331324 336564 331366
rect 137156 330922 204636 330964
rect 137156 330686 137198 330922
rect 137434 330686 159462 330922
rect 159698 330686 204358 330922
rect 204594 330686 204636 330922
rect 137156 330644 204636 330686
rect 231180 330922 292956 330964
rect 231180 330686 231222 330922
rect 231458 330686 251830 330922
rect 252066 330686 292678 330922
rect 292914 330686 292956 330922
rect 231180 330644 292956 330686
rect 161628 329562 212364 329604
rect 161628 329326 212086 329562
rect 212322 329326 212364 329562
rect 161628 329284 212364 329326
rect 253260 329562 299580 329604
rect 253260 329326 299302 329562
rect 299538 329326 299580 329562
rect 253260 329284 299580 329326
rect 161628 328924 161948 329284
rect 253260 328924 253580 329284
rect 137340 328882 161948 328924
rect 137340 328646 137382 328882
rect 137618 328646 161670 328882
rect 161906 328646 161948 328882
rect 137340 328604 161948 328646
rect 231732 328882 253580 328924
rect 231732 328646 231774 328882
rect 232010 328646 253302 328882
rect 253538 328646 253580 328882
rect 231732 328604 253580 328646
rect 137340 328202 208868 328244
rect 137340 327966 137382 328202
rect 137618 327966 160566 328202
rect 160802 327966 208590 328202
rect 208826 327966 208868 328202
rect 137340 327924 208868 327966
rect 0 320808 444740 320850
rect 0 320572 5122 320808
rect 5358 320572 5442 320808
rect 5678 320572 5762 320808
rect 5998 320572 6082 320808
rect 6318 320572 6402 320808
rect 6638 320572 6722 320808
rect 6958 320572 7042 320808
rect 7278 320572 7362 320808
rect 7598 320572 7682 320808
rect 7918 320572 8002 320808
rect 8238 320572 8322 320808
rect 8558 320572 8642 320808
rect 8878 320572 435862 320808
rect 436098 320572 436182 320808
rect 436418 320572 436502 320808
rect 436738 320572 436822 320808
rect 437058 320572 437142 320808
rect 437378 320572 437462 320808
rect 437698 320572 437782 320808
rect 438018 320572 438102 320808
rect 438338 320572 438422 320808
rect 438658 320572 438742 320808
rect 438978 320572 439062 320808
rect 439298 320572 439382 320808
rect 439618 320572 444740 320808
rect 0 320530 444740 320572
rect 105140 320042 105644 320084
rect 105140 319806 105182 320042
rect 105418 319806 105644 320042
rect 105140 319764 105644 319806
rect 105324 313964 105644 319764
rect 353172 314602 412372 314644
rect 353172 314366 353214 314602
rect 353450 314366 412094 314602
rect 412330 314366 412372 314602
rect 353172 314324 412372 314366
rect 105140 313644 105644 313964
rect 105140 312604 105460 313644
rect 104588 312284 105460 312604
rect 104588 309204 104908 312284
rect 104404 308884 104908 309204
rect 104404 307802 104724 308884
rect 412052 308482 413108 308524
rect 412052 308246 412094 308482
rect 412330 308246 413108 308482
rect 412052 308204 413108 308246
rect 104404 307566 104446 307802
rect 104682 307566 104724 307802
rect 104404 307524 104724 307566
rect 412788 306484 413108 308204
rect 412052 306442 429668 306484
rect 412052 306206 412094 306442
rect 412330 306206 429390 306442
rect 429626 306206 429668 306442
rect 412052 306164 429668 306206
rect 0 305490 444740 305532
rect 0 305254 122 305490
rect 358 305254 442 305490
rect 678 305254 762 305490
rect 998 305254 1082 305490
rect 1318 305254 1402 305490
rect 1638 305254 1722 305490
rect 1958 305254 2042 305490
rect 2278 305254 2362 305490
rect 2598 305254 2682 305490
rect 2918 305254 3002 305490
rect 3238 305254 3322 305490
rect 3558 305254 3642 305490
rect 3878 305254 104506 305490
rect 104742 305254 198506 305490
rect 198742 305254 292506 305490
rect 292742 305254 440862 305490
rect 441098 305254 441182 305490
rect 441418 305254 441502 305490
rect 441738 305254 441822 305490
rect 442058 305254 442142 305490
rect 442378 305254 442462 305490
rect 442698 305254 442782 305490
rect 443018 305254 443102 305490
rect 443338 305254 443422 305490
rect 443658 305254 443742 305490
rect 443978 305254 444062 305490
rect 444298 305254 444382 305490
rect 444618 305254 444740 305490
rect 0 305212 444740 305254
rect 104404 304124 113740 304444
rect 104404 303042 104724 304124
rect 104404 302806 104446 303042
rect 104682 302806 104724 303042
rect 104404 302764 104724 302806
rect 113420 298324 113740 304124
rect 246084 298962 248796 299004
rect 246084 298726 246126 298962
rect 246362 298726 248796 298962
rect 246084 298684 248796 298726
rect 248476 298324 248796 298684
rect 104588 298004 113740 298324
rect 104588 291482 104908 298004
rect 113420 296964 113740 298004
rect 118756 298282 134900 298324
rect 118756 298046 134622 298282
rect 134858 298046 134900 298282
rect 118756 298004 134900 298046
rect 246084 298282 248796 298324
rect 246084 298046 246126 298282
rect 246362 298046 248796 298282
rect 246084 298004 248796 298046
rect 118756 296964 119076 298004
rect 136788 297602 322948 297644
rect 136788 297366 136830 297602
rect 137066 297366 230670 297602
rect 230906 297366 322670 297602
rect 322906 297366 322948 297602
rect 136788 297324 322948 297366
rect 113420 296644 119076 296964
rect 202844 295284 205924 295604
rect 202844 294924 203164 295284
rect 200084 294604 203164 294924
rect 205604 294924 205924 295284
rect 206340 295284 222668 295604
rect 206340 294924 206660 295284
rect 205604 294604 206660 294924
rect 173956 293244 193596 293564
rect 137708 292842 142260 292884
rect 137708 292606 137750 292842
rect 137986 292606 142260 292842
rect 137708 292564 142260 292606
rect 104588 291246 104630 291482
rect 104866 291246 104908 291482
rect 104588 291204 104908 291246
rect 141940 291524 142260 292564
rect 173956 292204 174276 293244
rect 171380 291884 174276 292204
rect 193276 292204 193596 293244
rect 200084 292204 200404 294604
rect 205604 293924 206108 294604
rect 222348 294244 222668 295284
rect 222348 294202 229476 294244
rect 222348 293966 229198 294202
rect 229434 293966 229476 294202
rect 222348 293924 229476 293966
rect 292084 293924 306940 294244
rect 292084 293564 292404 293924
rect 193276 291884 200404 292204
rect 201004 293244 209236 293564
rect 171380 291524 171700 291884
rect 201004 291524 201324 293244
rect 141940 291204 171700 291524
rect 178556 291482 201324 291524
rect 178556 291246 178598 291482
rect 178834 291246 201324 291482
rect 178556 291204 201324 291246
rect 208916 291524 209236 293244
rect 220324 293522 228924 293564
rect 220324 293286 228646 293522
rect 228882 293286 228924 293522
rect 220324 293244 228924 293286
rect 270556 293244 292404 293564
rect 299076 293244 305836 293564
rect 220324 291524 220644 293244
rect 241668 292564 251372 292884
rect 241668 291524 241988 292564
rect 208916 291204 220644 291524
rect 231732 291482 241988 291524
rect 231732 291246 231774 291482
rect 232010 291246 241988 291482
rect 231732 291204 241988 291246
rect 251052 291524 251372 292564
rect 270556 292204 270876 293244
rect 267980 291884 270876 292204
rect 267980 291524 268300 291884
rect 299076 291524 299396 293244
rect 251052 291482 257996 291524
rect 251052 291246 257718 291482
rect 257954 291246 257996 291482
rect 251052 291204 257996 291246
rect 263564 291482 268300 291524
rect 263564 291246 263606 291482
rect 263842 291246 268300 291482
rect 263564 291204 268300 291246
rect 272580 291482 299396 291524
rect 272580 291246 272622 291482
rect 272858 291246 299396 291482
rect 272580 291204 299396 291246
rect 305516 291524 305836 293244
rect 306620 292884 306940 293924
rect 316372 293522 322948 293564
rect 316372 293286 322670 293522
rect 322906 293286 322948 293522
rect 316372 293244 322948 293286
rect 306620 292564 315772 292884
rect 315452 292204 315772 292564
rect 316372 292204 316692 293244
rect 315452 291884 316692 292204
rect 305516 291482 322948 291524
rect 305516 291246 322670 291482
rect 322906 291246 322948 291482
rect 305516 291204 322948 291246
rect 0 290172 444740 290214
rect 0 289936 5122 290172
rect 5358 289936 5442 290172
rect 5678 289936 5762 290172
rect 5998 289936 6082 290172
rect 6318 289936 6402 290172
rect 6638 289936 6722 290172
rect 6958 289936 7042 290172
rect 7278 289936 7362 290172
rect 7598 289936 7682 290172
rect 7918 289936 8002 290172
rect 8238 289936 8322 290172
rect 8558 289936 8642 290172
rect 8878 289936 89146 290172
rect 89382 289936 183146 290172
rect 183382 289936 277146 290172
rect 277382 289936 435862 290172
rect 436098 289936 436182 290172
rect 436418 289936 436502 290172
rect 436738 289936 436822 290172
rect 437058 289936 437142 290172
rect 437378 289936 437462 290172
rect 437698 289936 437782 290172
rect 438018 289936 438102 290172
rect 438338 289936 438422 290172
rect 438658 289936 438742 290172
rect 438978 289936 439062 290172
rect 439298 289936 439382 290172
rect 439618 289936 444740 290172
rect 0 289894 444740 289936
rect 92076 289164 93132 289484
rect 92076 288804 92396 289164
rect 91524 288484 92396 288804
rect 92812 288804 93132 289164
rect 104588 289442 104908 289484
rect 104588 289206 104630 289442
rect 104866 289206 104908 289442
rect 104588 288804 104908 289206
rect 137708 289442 165812 289484
rect 137708 289206 137750 289442
rect 137986 289206 165534 289442
rect 165770 289206 165812 289442
rect 137708 289164 165812 289206
rect 235964 289442 259652 289484
rect 235964 289206 236006 289442
rect 236242 289206 259374 289442
rect 259610 289206 259652 289442
rect 235964 289164 259652 289206
rect 92812 288484 104908 288804
rect 29148 286722 38852 286764
rect 29148 286486 38574 286722
rect 38810 286486 38852 286722
rect 29148 286444 38852 286486
rect 29148 285404 29468 286444
rect 21788 285084 29468 285404
rect 41292 285084 51732 285404
rect 21788 284044 22108 285084
rect 41292 284044 41612 285084
rect 13508 284002 22108 284044
rect 13508 283766 13550 284002
rect 13786 283766 22108 284002
rect 13508 283724 22108 283766
rect 38532 284002 41612 284044
rect 38532 283766 38574 284002
rect 38810 283766 41612 284002
rect 38532 283724 41612 283766
rect 51412 284044 51732 285084
rect 84164 284682 84824 284724
rect 84164 284446 84390 284682
rect 84626 284446 84824 284682
rect 84164 284404 84824 284446
rect 51412 283724 60748 284044
rect 60428 283364 60748 283724
rect 71100 283724 79884 284044
rect 71100 283364 71420 283724
rect 60428 283044 71420 283364
rect 79564 283364 79884 283724
rect 84164 283364 84484 284404
rect 91524 284044 91844 288484
rect 79564 283044 84484 283364
rect 84900 283724 91844 284044
rect 92260 285764 101596 286084
rect 84900 282684 85220 283724
rect 84532 282642 85220 282684
rect 84532 282406 84574 282642
rect 84810 282406 85220 282642
rect 84532 282364 85220 282406
rect 92260 282004 92580 285764
rect 101276 284044 101596 285764
rect 102564 285764 106564 286084
rect 102564 284044 102884 285764
rect 106244 285404 106564 285764
rect 106244 285362 134900 285404
rect 106244 285126 134622 285362
rect 134858 285126 134900 285362
rect 106244 285084 134900 285126
rect 351700 285362 353860 285404
rect 351700 285126 351742 285362
rect 351978 285126 353582 285362
rect 353818 285126 353860 285362
rect 351700 285084 353860 285126
rect 110292 284404 128092 284724
rect 110292 284044 110612 284404
rect 96676 283724 99756 284044
rect 101276 283724 102884 284044
rect 103668 283724 110612 284044
rect 96676 283364 96996 283724
rect 84532 281962 92580 282004
rect 84532 281726 84574 281962
rect 84810 281726 92580 281962
rect 84532 281684 92580 281726
rect 95204 283044 96996 283364
rect 99436 283364 99756 283724
rect 103668 283364 103988 283724
rect 99436 283044 103988 283364
rect 127772 283364 128092 284404
rect 128876 284682 137476 284724
rect 128876 284446 137198 284682
rect 137434 284446 137476 284682
rect 128876 284404 137476 284446
rect 128876 283364 129196 284404
rect 127772 283044 129196 283364
rect 95204 281324 95524 283044
rect 134580 282642 138764 282684
rect 134580 282406 134622 282642
rect 134858 282406 138486 282642
rect 138722 282406 138764 282642
rect 134580 282364 138764 282406
rect 246084 282642 248612 282684
rect 246084 282406 246126 282642
rect 246362 282406 248612 282642
rect 246084 282364 248612 282406
rect 412052 282642 415316 282684
rect 412052 282406 412094 282642
rect 412330 282406 415316 282642
rect 412052 282364 415316 282406
rect 84532 281282 95524 281324
rect 84532 281046 84574 281282
rect 84810 281046 95524 281282
rect 84532 281004 95524 281046
rect 248292 279284 248612 282364
rect 246084 279242 248612 279284
rect 246084 279006 246126 279242
rect 246362 279006 248612 279242
rect 246084 278964 248612 279006
rect 414996 278562 415316 282364
rect 414996 278326 415038 278562
rect 415274 278326 415316 278562
rect 414996 278284 415316 278326
rect 0 274854 444740 274896
rect 0 274618 122 274854
rect 358 274618 442 274854
rect 678 274618 762 274854
rect 998 274618 1082 274854
rect 1318 274618 1402 274854
rect 1638 274618 1722 274854
rect 1958 274618 2042 274854
rect 2278 274618 2362 274854
rect 2598 274618 2682 274854
rect 2918 274618 3002 274854
rect 3238 274618 3322 274854
rect 3558 274618 3642 274854
rect 3878 274618 104506 274854
rect 104742 274618 198506 274854
rect 198742 274618 292506 274854
rect 292742 274618 440862 274854
rect 441098 274618 441182 274854
rect 441418 274618 441502 274854
rect 441738 274618 441822 274854
rect 442058 274618 442142 274854
rect 442378 274618 442462 274854
rect 442698 274618 442782 274854
rect 443018 274618 443102 274854
rect 443338 274618 443422 274854
rect 443658 274618 443742 274854
rect 443978 274618 444062 274854
rect 444298 274618 444382 274854
rect 444618 274618 444740 274854
rect 0 274576 444740 274618
rect 247740 262242 248060 262284
rect 247740 262006 247782 262242
rect 248018 262006 248060 262242
rect 247740 260244 248060 262006
rect 237988 260202 248060 260244
rect 237988 259966 238030 260202
rect 238266 259966 248060 260202
rect 237988 259924 248060 259966
rect 0 259536 444740 259578
rect 0 259300 5122 259536
rect 5358 259300 5442 259536
rect 5678 259300 5762 259536
rect 5998 259300 6082 259536
rect 6318 259300 6402 259536
rect 6638 259300 6722 259536
rect 6958 259300 7042 259536
rect 7278 259300 7362 259536
rect 7598 259300 7682 259536
rect 7918 259300 8002 259536
rect 8238 259300 8322 259536
rect 8558 259300 8642 259536
rect 8878 259300 435862 259536
rect 436098 259300 436182 259536
rect 436418 259300 436502 259536
rect 436738 259300 436822 259536
rect 437058 259300 437142 259536
rect 437378 259300 437462 259536
rect 437698 259300 437782 259536
rect 438018 259300 438102 259536
rect 438338 259300 438422 259536
rect 438658 259300 438742 259536
rect 438978 259300 439062 259536
rect 439298 259300 439382 259536
rect 439618 259300 444740 259536
rect 0 259258 444740 259300
rect 143964 257482 148700 257524
rect 143964 257246 144006 257482
rect 144242 257246 148700 257482
rect 143964 257204 148700 257246
rect 237988 257482 248244 257524
rect 237988 257246 238030 257482
rect 238266 257246 248244 257482
rect 237988 257204 248244 257246
rect 48468 256122 76388 256164
rect 48468 255886 48510 256122
rect 48746 255886 76110 256122
rect 76346 255886 76388 256122
rect 48468 255844 76388 255886
rect 49020 252042 75468 252084
rect 49020 251806 49062 252042
rect 49298 251806 75190 252042
rect 75426 251806 75468 252042
rect 49020 251764 75468 251806
rect 73860 251362 75100 251404
rect 73860 251126 73902 251362
rect 74138 251126 74822 251362
rect 75058 251126 75100 251362
rect 73860 251084 75100 251126
rect 75516 251362 76388 251404
rect 75516 251126 76110 251362
rect 76346 251126 76388 251362
rect 75516 251084 76388 251126
rect 75516 250724 75836 251084
rect 75148 250682 75836 250724
rect 75148 250446 75190 250682
rect 75426 250446 75836 250682
rect 75148 250404 75836 250446
rect 49020 249322 68108 249364
rect 49020 249086 49062 249322
rect 49298 249086 68108 249322
rect 49020 249044 68108 249086
rect 67788 248004 68108 249044
rect 148380 248684 148700 257204
rect 236516 249322 238308 249364
rect 236516 249086 236558 249322
rect 236794 249086 238030 249322
rect 238266 249086 238308 249322
rect 236516 249044 238308 249086
rect 143964 248642 148700 248684
rect 143964 248406 144006 248642
rect 144242 248406 148700 248642
rect 143964 248364 148700 248406
rect 67788 247962 74548 248004
rect 67788 247726 74270 247962
rect 74506 247726 74548 247962
rect 67788 247684 74548 247726
rect 247924 245284 248244 257204
rect 355564 256122 358828 256164
rect 355564 255886 355606 256122
rect 355842 255886 358550 256122
rect 358786 255886 358828 256122
rect 355564 255844 358828 255886
rect 325020 249322 358828 249364
rect 325020 249086 325062 249322
rect 325298 249086 358550 249322
rect 358786 249086 358828 249322
rect 325020 249044 358828 249086
rect 73860 245242 75836 245284
rect 73860 245006 73902 245242
rect 74138 245006 75558 245242
rect 75794 245006 75836 245242
rect 73860 244964 75836 245006
rect 236884 245242 248244 245284
rect 236884 245006 236926 245242
rect 237162 245006 248244 245242
rect 236884 244964 248244 245006
rect 0 244218 444740 244260
rect 0 243982 122 244218
rect 358 243982 442 244218
rect 678 243982 762 244218
rect 998 243982 1082 244218
rect 1318 243982 1402 244218
rect 1638 243982 1722 244218
rect 1958 243982 2042 244218
rect 2278 243982 2362 244218
rect 2598 243982 2682 244218
rect 2918 243982 3002 244218
rect 3238 243982 3322 244218
rect 3558 243982 3642 244218
rect 3878 243982 440862 244218
rect 441098 243982 441182 244218
rect 441418 243982 441502 244218
rect 441738 243982 441822 244218
rect 442058 243982 442142 244218
rect 442378 243982 442462 244218
rect 442698 243982 442782 244218
rect 443018 243982 443102 244218
rect 443338 243982 443422 244218
rect 443658 243982 443742 244218
rect 443978 243982 444062 244218
rect 444298 243982 444382 244218
rect 444618 243982 444740 244218
rect 0 243940 444740 243982
rect 49020 243202 76020 243244
rect 49020 242966 49062 243202
rect 49298 242966 75742 243202
rect 75978 242966 76020 243202
rect 49020 242924 76020 242966
rect 48284 242522 60748 242564
rect 48284 242286 48326 242522
rect 48562 242286 60748 242522
rect 48284 242244 60748 242286
rect 236884 242522 242908 242564
rect 236884 242286 236926 242522
rect 237162 242286 242908 242522
rect 236884 242244 242908 242286
rect 51044 240884 51548 242244
rect 60428 241884 60748 242244
rect 242588 241884 242908 242244
rect 60428 241564 74732 241884
rect 74412 240524 74732 241564
rect 95204 241564 96260 241884
rect 95204 241204 95524 241564
rect 93732 241162 95524 241204
rect 93732 240926 93774 241162
rect 94010 240926 95524 241162
rect 93732 240884 95524 240926
rect 95940 241162 96260 241564
rect 95940 240926 95982 241162
rect 96218 240926 96260 241162
rect 95940 240884 96260 240926
rect 128508 241842 137108 241884
rect 128508 241606 136830 241842
rect 137066 241606 137108 241842
rect 128508 241564 137108 241606
rect 143596 241842 152748 241884
rect 143596 241606 143638 241842
rect 143874 241606 152748 241842
rect 143596 241564 152748 241606
rect 74412 240482 76388 240524
rect 74412 240246 75374 240482
rect 75610 240246 76110 240482
rect 76346 240246 76388 240482
rect 74412 240204 76388 240246
rect 104772 240482 106748 240524
rect 104772 240246 104814 240482
rect 105050 240246 106470 240482
rect 106706 240246 106748 240482
rect 104772 240204 106748 240246
rect 118572 240482 126068 240524
rect 118572 240246 118614 240482
rect 118850 240246 125790 240482
rect 126026 240246 126068 240482
rect 118572 240204 126068 240246
rect 128508 240482 128828 241564
rect 128508 240246 128550 240482
rect 128786 240246 128828 240482
rect 128508 240204 128828 240246
rect 152428 240524 152748 241564
rect 176716 241564 188812 241884
rect 242588 241842 262228 241884
rect 242588 241606 261950 241842
rect 262186 241606 262228 241842
rect 242588 241564 262228 241606
rect 176716 240524 177036 241564
rect 152428 240204 153484 240524
rect 167700 240482 177036 240524
rect 167700 240246 167742 240482
rect 167978 240246 177036 240482
rect 167700 240204 177036 240246
rect 153164 239844 153484 240204
rect 188492 239844 188812 241564
rect 292452 241204 292956 241884
rect 282884 240884 283940 241204
rect 282884 240524 283204 240884
rect 224924 240204 229476 240524
rect 49020 239802 73444 239844
rect 49020 239566 49062 239802
rect 49298 239566 73444 239802
rect 49020 239524 73444 239566
rect 75700 239802 143916 239844
rect 75700 239566 75742 239802
rect 75978 239566 95062 239802
rect 95298 239566 138670 239802
rect 138906 239566 143638 239802
rect 143874 239566 143916 239802
rect 75700 239524 143916 239566
rect 149116 239802 188076 239844
rect 149116 239566 187798 239802
rect 188034 239566 188076 239802
rect 149116 239524 188076 239566
rect 188492 239524 196172 239844
rect 73124 237762 73444 239524
rect 74090 239122 80620 239164
rect 74090 238886 74132 239122
rect 74368 238886 80620 239122
rect 74090 238844 80620 238886
rect 80300 238484 80620 238844
rect 80300 238442 102516 238484
rect 80300 238206 102238 238442
rect 102474 238206 102516 238442
rect 80300 238164 102516 238206
rect 142676 238442 148148 238484
rect 142676 238206 142718 238442
rect 142954 238206 148148 238442
rect 142676 238164 148148 238206
rect 73124 237526 73166 237762
rect 73402 237526 73444 237762
rect 73124 237484 73444 237526
rect 147828 237762 148148 238164
rect 147828 237526 147870 237762
rect 148106 237526 148148 237762
rect 147828 237484 148148 237526
rect 149116 237762 149436 239524
rect 195852 239164 196172 239524
rect 211124 239802 211444 239844
rect 211124 239566 211166 239802
rect 211402 239566 211444 239802
rect 211124 239164 211444 239566
rect 224924 239164 225244 240204
rect 195852 238844 225244 239164
rect 229156 239164 229476 240204
rect 250316 240204 254868 240524
rect 235228 239524 248980 239844
rect 235228 239164 235548 239524
rect 229156 239122 235548 239164
rect 229156 238886 230854 239122
rect 231090 238886 235548 239122
rect 229156 238844 235548 238886
rect 248660 239164 248980 239524
rect 250316 239164 250636 240204
rect 248660 238844 250636 239164
rect 254548 239164 254868 240204
rect 259884 240482 283204 240524
rect 259884 240246 261582 240482
rect 261818 240246 283204 240482
rect 259884 240204 283204 240246
rect 283620 240524 283940 240884
rect 292084 240884 303996 241204
rect 292084 240524 292404 240884
rect 283620 240204 292404 240524
rect 303676 240482 303996 240884
rect 303676 240246 303718 240482
rect 303954 240246 303996 240482
rect 303676 240204 303996 240246
rect 259884 239164 260204 240204
rect 262828 239802 325892 239844
rect 262828 239566 262870 239802
rect 263106 239566 290470 239802
rect 290706 239566 325614 239802
rect 325850 239566 325892 239802
rect 262828 239524 325892 239566
rect 254548 238844 260204 239164
rect 325204 239122 360668 239164
rect 325204 238886 325246 239122
rect 325482 238886 360390 239122
rect 360626 238886 360668 239122
rect 325204 238844 360668 238886
rect 168988 238442 200220 238484
rect 168988 238206 169030 238442
rect 169266 238206 199942 238442
rect 200178 238206 200220 238442
rect 168988 238164 200220 238206
rect 231732 238442 238308 238484
rect 231732 238206 231774 238442
rect 232010 238206 238030 238442
rect 238266 238206 238308 238442
rect 231732 238164 238308 238206
rect 149116 237526 149158 237762
rect 149394 237526 149436 237762
rect 149116 237484 149436 237526
rect 248660 237762 248980 238844
rect 261908 238442 287068 238484
rect 261908 238206 261950 238442
rect 262186 238206 286790 238442
rect 287026 238206 287068 238442
rect 261908 238164 287068 238206
rect 248660 237526 248702 237762
rect 248938 237526 248980 237762
rect 248660 237484 248980 237526
rect 143964 237082 148884 237124
rect 143964 236846 144006 237082
rect 144242 236846 148606 237082
rect 148842 236846 148884 237082
rect 143964 236804 148884 236846
rect 182052 237082 184028 237124
rect 182052 236846 183750 237082
rect 183986 236846 184028 237082
rect 182052 236804 184028 236846
rect 182052 236444 182372 236804
rect 149484 236402 153668 236444
rect 149484 236166 149526 236402
rect 149762 236166 153390 236402
rect 153626 236166 153668 236402
rect 149484 236124 153668 236166
rect 162732 236402 182372 236444
rect 162732 236166 162774 236402
rect 163010 236166 182372 236402
rect 162732 236124 182372 236166
rect 75700 235722 110612 235764
rect 75700 235486 75742 235722
rect 75978 235486 110334 235722
rect 110570 235486 110612 235722
rect 75700 235444 110612 235486
rect 172484 235444 172988 236124
rect 137708 235042 141340 235084
rect 137708 234806 137750 235042
rect 137986 234806 141062 235042
rect 141298 234806 141340 235042
rect 137708 234764 141340 234806
rect 144884 235042 207396 235084
rect 144884 234806 144926 235042
rect 145162 234806 151918 235042
rect 152154 234806 168478 235042
rect 168714 234806 207118 235042
rect 207354 234806 207396 235042
rect 144884 234764 207396 234806
rect 231732 235042 234996 235084
rect 231732 234806 231774 235042
rect 232010 234806 234718 235042
rect 234954 234806 234996 235042
rect 231732 234764 234996 234806
rect 249764 235042 284492 235084
rect 249764 234806 249806 235042
rect 250042 234806 284214 235042
rect 284450 234806 284492 235042
rect 249764 234764 284492 234806
rect 297420 235042 301236 235084
rect 297420 234806 297462 235042
rect 297698 234806 300958 235042
rect 301194 234806 301236 235042
rect 297420 234764 301236 234806
rect 244244 234362 251556 234404
rect 244244 234126 244286 234362
rect 244522 234126 245942 234362
rect 246178 234126 251556 234362
rect 244244 234084 251556 234126
rect 251236 233044 251556 234084
rect 269084 233682 271060 233724
rect 269084 233446 269126 233682
rect 269362 233446 271060 233682
rect 269084 233404 271060 233446
rect 270740 233044 271060 233404
rect 273316 233404 275660 233724
rect 285092 233682 290196 233724
rect 285092 233446 285134 233682
rect 285370 233446 289918 233682
rect 290154 233446 290196 233682
rect 285092 233404 290196 233446
rect 273316 233044 273636 233404
rect 251236 233002 259836 233044
rect 251236 232766 259558 233002
rect 259794 232766 259836 233002
rect 251236 232724 259836 232766
rect 270740 232724 273636 233044
rect 275340 233044 275660 233404
rect 275340 233002 282836 233044
rect 275340 232766 282558 233002
rect 282794 232766 282836 233002
rect 275340 232724 282836 232766
rect 0 228900 444740 228942
rect 0 228664 5122 228900
rect 5358 228664 5442 228900
rect 5678 228664 5762 228900
rect 5998 228664 6082 228900
rect 6318 228664 6402 228900
rect 6638 228664 6722 228900
rect 6958 228664 7042 228900
rect 7278 228664 7362 228900
rect 7598 228664 7682 228900
rect 7918 228664 8002 228900
rect 8238 228664 8322 228900
rect 8558 228664 8642 228900
rect 8878 228664 376882 228900
rect 377118 228664 435862 228900
rect 436098 228664 436182 228900
rect 436418 228664 436502 228900
rect 436738 228664 436822 228900
rect 437058 228664 437142 228900
rect 437378 228664 437462 228900
rect 437698 228664 437782 228900
rect 438018 228664 438102 228900
rect 438338 228664 438422 228900
rect 438658 228664 438742 228900
rect 438978 228664 439062 228900
rect 439298 228664 439382 228900
rect 439618 228664 444740 228900
rect 0 228622 444740 228664
rect 358508 222122 406116 222164
rect 358508 221886 358550 222122
rect 358786 221886 405838 222122
rect 406074 221886 406116 222122
rect 358508 221844 406116 221886
rect 219404 217362 229108 217404
rect 219404 217126 228830 217362
rect 229066 217126 229108 217362
rect 219404 217084 229108 217126
rect 242588 217362 258916 217404
rect 242588 217126 242630 217362
rect 242866 217126 258638 217362
rect 258874 217126 258916 217362
rect 242588 217084 258916 217126
rect 272580 217362 297740 217404
rect 272580 217126 272622 217362
rect 272858 217126 297740 217362
rect 272580 217084 297740 217126
rect 219404 216724 219724 217084
rect 148564 216682 152196 216724
rect 148564 216446 148606 216682
rect 148842 216446 152196 216682
rect 148564 216404 152196 216446
rect 177452 216682 186788 216724
rect 177452 216446 177494 216682
rect 177730 216446 186788 216682
rect 177452 216404 186788 216446
rect 151876 215364 152196 216404
rect 186468 216044 186788 216404
rect 196036 216404 219724 216724
rect 242588 216682 258916 216724
rect 242588 216446 242630 216682
rect 242866 216446 258638 216682
rect 258874 216446 258916 216682
rect 242588 216404 258916 216446
rect 272580 216682 287436 216724
rect 272580 216446 272622 216682
rect 272858 216446 287436 216682
rect 272580 216404 287436 216446
rect 196036 216044 196356 216404
rect 186468 215724 196356 216044
rect 287116 216044 287436 216404
rect 287116 215724 297004 216044
rect 151876 215322 165076 215364
rect 151876 215086 164798 215322
rect 165034 215086 165076 215322
rect 151876 215044 165076 215086
rect 195852 215044 196356 215724
rect 296684 214684 297004 215724
rect 297420 215364 297740 217084
rect 306252 217362 323132 217404
rect 306252 217126 322854 217362
rect 323090 217126 323132 217362
rect 306252 217084 323132 217126
rect 336796 217362 352940 217404
rect 336796 217126 336838 217362
rect 337074 217126 352662 217362
rect 352898 217126 352940 217362
rect 336796 217084 352940 217126
rect 306252 215364 306572 217084
rect 336612 216682 352940 216724
rect 336612 216446 336654 216682
rect 336890 216446 352662 216682
rect 352898 216446 352940 216682
rect 336612 216404 352940 216446
rect 297420 215044 306572 215364
rect 307172 216002 323132 216044
rect 307172 215766 322854 216002
rect 323090 215766 323132 216002
rect 307172 215724 323132 215766
rect 357404 216002 406116 216044
rect 357404 215766 357446 216002
rect 357682 215766 405838 216002
rect 406074 215766 406116 216002
rect 357404 215724 406116 215766
rect 307172 214684 307492 215724
rect 296684 214364 307492 214684
rect 0 213582 444740 213624
rect 0 213346 122 213582
rect 358 213346 442 213582
rect 678 213346 762 213582
rect 998 213346 1082 213582
rect 1318 213346 1402 213582
rect 1638 213346 1722 213582
rect 1958 213346 2042 213582
rect 2278 213346 2362 213582
rect 2598 213346 2682 213582
rect 2918 213346 3002 213582
rect 3238 213346 3322 213582
rect 3558 213346 3642 213582
rect 3878 213346 104506 213582
rect 104742 213346 198506 213582
rect 198742 213346 292506 213582
rect 292742 213346 440862 213582
rect 441098 213346 441182 213582
rect 441418 213346 441502 213582
rect 441738 213346 441822 213582
rect 442058 213346 442142 213582
rect 442378 213346 442462 213582
rect 442698 213346 442782 213582
rect 443018 213346 443102 213582
rect 443338 213346 443422 213582
rect 443658 213346 443742 213582
rect 443978 213346 444062 213582
rect 444298 213346 444382 213582
rect 444618 213346 444740 213582
rect 0 213304 444740 213346
rect 231732 207842 242724 207884
rect 231732 207606 231774 207842
rect 232010 207606 242446 207842
rect 242682 207606 242724 207842
rect 231732 207564 242724 207606
rect 93916 206204 109140 206524
rect 93916 204484 94236 206204
rect 108820 205164 109140 206204
rect 115996 206204 119076 206524
rect 115996 205844 116316 206204
rect 115444 205524 116316 205844
rect 118756 205844 119076 206204
rect 120780 206204 128644 206524
rect 120780 205844 121100 206204
rect 118756 205524 121100 205844
rect 115444 205164 115764 205524
rect 108820 204844 115764 205164
rect 128324 205164 128644 206204
rect 128324 205122 134900 205164
rect 128324 204886 134622 205122
rect 134858 204886 134900 205122
rect 128324 204844 134900 204886
rect 84532 204442 94236 204484
rect 84532 204206 84574 204442
rect 84810 204206 94236 204442
rect 84532 204164 94236 204206
rect 137708 201042 322948 201084
rect 137708 200806 137750 201042
rect 137986 200806 230670 201042
rect 230906 200806 322670 201042
rect 322906 200806 322948 201042
rect 137708 200764 322948 200806
rect 137892 199002 322948 199044
rect 137892 198766 137934 199002
rect 138170 198766 230670 199002
rect 230906 198766 322670 199002
rect 322906 198766 322948 199002
rect 137892 198724 322948 198766
rect 0 198264 444740 198306
rect 0 198028 5122 198264
rect 5358 198028 5442 198264
rect 5678 198028 5762 198264
rect 5998 198028 6082 198264
rect 6318 198028 6402 198264
rect 6638 198028 6722 198264
rect 6958 198028 7042 198264
rect 7278 198028 7362 198264
rect 7598 198028 7682 198264
rect 7918 198028 8002 198264
rect 8238 198028 8322 198264
rect 8558 198028 8642 198264
rect 8878 198028 89146 198264
rect 89382 198028 183146 198264
rect 183382 198028 277146 198264
rect 277382 198028 435862 198264
rect 436098 198028 436182 198264
rect 436418 198028 436502 198264
rect 436738 198028 436822 198264
rect 437058 198028 437142 198264
rect 437378 198028 437462 198264
rect 437698 198028 437782 198264
rect 438018 198028 438102 198264
rect 438338 198028 438422 198264
rect 438658 198028 438742 198264
rect 438978 198028 439062 198264
rect 439298 198028 439382 198264
rect 439618 198028 444740 198264
rect 0 197986 444740 198028
rect 235964 194922 322948 194964
rect 235964 194686 236006 194922
rect 236242 194686 322670 194922
rect 322906 194686 322948 194922
rect 235964 194644 322948 194686
rect 137892 194242 228924 194284
rect 137892 194006 137934 194242
rect 138170 194006 228646 194242
rect 228882 194006 228924 194242
rect 137892 193964 228924 194006
rect 0 182946 444740 182988
rect 0 182710 122 182946
rect 358 182710 442 182946
rect 678 182710 762 182946
rect 998 182710 1082 182946
rect 1318 182710 1402 182946
rect 1638 182710 1722 182946
rect 1958 182710 2042 182946
rect 2278 182710 2362 182946
rect 2598 182710 2682 182946
rect 2918 182710 3002 182946
rect 3238 182710 3322 182946
rect 3558 182710 3642 182946
rect 3878 182710 104506 182946
rect 104742 182710 198506 182946
rect 198742 182710 292506 182946
rect 292742 182710 440862 182946
rect 441098 182710 441182 182946
rect 441418 182710 441502 182946
rect 441738 182710 441822 182946
rect 442058 182710 442142 182946
rect 442378 182710 442462 182946
rect 442698 182710 442782 182946
rect 443018 182710 443102 182946
rect 443338 182710 443422 182946
rect 443658 182710 443742 182946
rect 443978 182710 444062 182946
rect 444298 182710 444382 182946
rect 444618 182710 444740 182946
rect 0 182668 444740 182710
rect 318948 182044 323684 182316
rect 215172 181724 219908 182044
rect 271292 182002 310804 182044
rect 271292 181766 271334 182002
rect 271570 181766 310804 182002
rect 271292 181724 310804 181766
rect 174692 181322 196356 181364
rect 174692 181086 174734 181322
rect 174970 181086 196356 181322
rect 174692 181044 196356 181086
rect 196036 180004 196356 181044
rect 215172 180684 215492 181724
rect 205788 180364 215492 180684
rect 219588 180684 219908 181724
rect 267428 181322 283388 181364
rect 267428 181086 267470 181322
rect 267706 181086 283388 181322
rect 267428 181044 283388 181086
rect 219588 180642 228924 180684
rect 219588 180406 228646 180642
rect 228882 180406 228924 180642
rect 219588 180364 228924 180406
rect 205788 180004 206108 180364
rect 196036 179684 206108 180004
rect 283068 180004 283388 181044
rect 292452 181044 302708 181364
rect 292452 180004 292772 181044
rect 283068 179684 292772 180004
rect 302388 180004 302708 181044
rect 302388 179684 310068 180004
rect 309748 179282 310068 179684
rect 309748 179046 309790 179282
rect 310026 179046 310068 179282
rect 309748 179004 310068 179046
rect 310484 179324 310804 181724
rect 312876 182002 323684 182044
rect 312876 181996 323406 182002
rect 312876 181724 319268 181996
rect 323364 181766 323406 181996
rect 323642 181766 323684 182002
rect 323364 181724 323684 181766
rect 312876 181364 313196 181724
rect 312508 181044 313196 181364
rect 321524 181322 323316 181364
rect 321524 181086 323038 181322
rect 323274 181086 323316 181322
rect 321524 181044 323316 181086
rect 310484 179282 311356 179324
rect 310484 179046 311078 179282
rect 311314 179046 311356 179282
rect 310484 179004 311356 179046
rect 312508 179282 312828 181044
rect 321524 180004 321844 181044
rect 312508 179046 312550 179282
rect 312786 179046 312828 179282
rect 312508 179004 312828 179046
rect 313612 179684 321844 180004
rect 313612 179282 313932 179684
rect 313612 179046 313654 179282
rect 313890 179046 313932 179282
rect 313612 179004 313932 179046
rect 73492 168402 76940 168444
rect 73492 168166 73534 168402
rect 73770 168166 76662 168402
rect 76898 168166 76940 168402
rect 73492 168124 76940 168166
rect 237620 168402 242908 168444
rect 237620 168166 237662 168402
rect 237898 168166 242630 168402
rect 242866 168166 242908 168402
rect 237620 168124 242908 168166
rect 243324 168402 247324 168444
rect 243324 168166 243366 168402
rect 243602 168166 247046 168402
rect 247282 168166 247324 168402
rect 243324 168124 247324 168166
rect 0 167628 444740 167670
rect 0 167392 5122 167628
rect 5358 167392 5442 167628
rect 5678 167392 5762 167628
rect 5998 167392 6082 167628
rect 6318 167392 6402 167628
rect 6638 167392 6722 167628
rect 6958 167392 7042 167628
rect 7278 167392 7362 167628
rect 7598 167392 7682 167628
rect 7918 167392 8002 167628
rect 8238 167392 8322 167628
rect 8558 167392 8642 167628
rect 8878 167392 435862 167628
rect 436098 167392 436182 167628
rect 436418 167392 436502 167628
rect 436738 167392 436822 167628
rect 437058 167392 437142 167628
rect 437378 167392 437462 167628
rect 437698 167392 437782 167628
rect 438018 167392 438102 167628
rect 438338 167392 438422 167628
rect 438658 167392 438742 167628
rect 438978 167392 439062 167628
rect 439298 167392 439382 167628
rect 439618 167392 444740 167628
rect 0 167350 444740 167392
rect 237252 166362 247508 166404
rect 237252 166126 237294 166362
rect 237530 166126 247508 166362
rect 237252 166084 247508 166126
rect 247188 162324 247508 166084
rect 49020 162282 74916 162324
rect 49020 162046 49062 162282
rect 49298 162046 74638 162282
rect 74874 162046 74916 162282
rect 49020 162004 74916 162046
rect 143964 162282 148884 162324
rect 143964 162046 144006 162282
rect 144242 162046 148884 162282
rect 143964 162004 148884 162046
rect 247188 162004 248428 162324
rect 74412 160922 74732 162004
rect 74412 160686 74454 160922
rect 74690 160686 74732 160922
rect 74412 160644 74732 160686
rect 148564 160284 148884 162004
rect 248108 160284 248428 162004
rect 143964 160242 148884 160284
rect 143964 160006 144006 160242
rect 144242 160006 148884 160242
rect 143964 159964 148884 160006
rect 242588 159964 248428 160284
rect 49020 158202 76940 158244
rect 49020 157966 49062 158202
rect 49298 157966 76662 158202
rect 76898 157966 76940 158202
rect 49020 157924 76940 157966
rect 73676 157522 73996 157924
rect 242588 157564 242908 159964
rect 73676 157286 73718 157522
rect 73954 157286 73996 157522
rect 73676 157244 73996 157286
rect 237252 157522 242908 157564
rect 237252 157286 237294 157522
rect 237530 157286 242908 157522
rect 237252 157244 242908 157286
rect 49020 155482 75836 155524
rect 49020 155246 49062 155482
rect 49298 155246 75558 155482
rect 75794 155246 75836 155482
rect 49020 155204 75836 155246
rect 49020 153442 74180 153484
rect 49020 153206 49062 153442
rect 49298 153206 73902 153442
rect 74138 153206 74180 153442
rect 49020 153164 74180 153206
rect 0 152310 444740 152352
rect 0 152074 122 152310
rect 358 152074 442 152310
rect 678 152074 762 152310
rect 998 152074 1082 152310
rect 1318 152074 1402 152310
rect 1638 152074 1722 152310
rect 1958 152074 2042 152310
rect 2278 152074 2362 152310
rect 2598 152074 2682 152310
rect 2918 152074 3002 152310
rect 3238 152074 3322 152310
rect 3558 152074 3642 152310
rect 3878 152074 440862 152310
rect 441098 152074 441182 152310
rect 441418 152074 441502 152310
rect 441738 152074 441822 152310
rect 442058 152074 442142 152310
rect 442378 152074 442462 152310
rect 442698 152074 442782 152310
rect 443018 152074 443102 152310
rect 443338 152074 443422 152310
rect 443658 152074 443742 152310
rect 443978 152074 444062 152310
rect 444298 152074 444382 152310
rect 444618 152074 444740 152310
rect 0 152032 444740 152074
rect 74228 151402 74548 151444
rect 74228 151166 74270 151402
rect 74506 151166 74548 151402
rect 74228 150764 74548 151166
rect 143964 151402 145388 151444
rect 143964 151166 144006 151402
rect 144242 151166 145388 151402
rect 143964 151124 145388 151166
rect 73860 150444 74548 150764
rect 73860 149404 74180 150444
rect 74596 150042 76572 150084
rect 74596 149806 74638 150042
rect 74874 149806 76294 150042
rect 76530 149806 76572 150042
rect 74596 149764 76572 149806
rect 73860 149362 74548 149404
rect 73860 149126 74270 149362
rect 74506 149126 74548 149362
rect 73860 149084 74548 149126
rect 49020 148682 77860 148724
rect 49020 148446 49062 148682
rect 49298 148446 75006 148682
rect 75242 148446 77582 148682
rect 77818 148446 77860 148682
rect 49020 148404 77860 148446
rect 49020 145962 75468 146004
rect 49020 145726 49062 145962
rect 49298 145726 75190 145962
rect 75426 145726 75468 145962
rect 49020 145684 75468 145726
rect 145068 145324 145388 151124
rect 237252 150722 246588 150764
rect 237252 150486 237294 150722
rect 237530 150486 246588 150722
rect 237252 150444 246588 150486
rect 237620 148002 243828 148044
rect 237620 147766 237662 148002
rect 237898 147766 243828 148002
rect 237620 147724 243828 147766
rect 237988 147322 242540 147364
rect 237988 147086 238030 147322
rect 238266 147086 242540 147322
rect 237988 147044 242540 147086
rect 242220 146684 242540 147044
rect 237988 146642 242540 146684
rect 237988 146406 238030 146642
rect 238266 146406 242540 146642
rect 237988 146364 242540 146406
rect 76988 145282 145388 145324
rect 76988 145046 77030 145282
rect 77266 145046 98742 145282
rect 98978 145046 144006 145282
rect 144242 145046 145388 145282
rect 76988 145004 145388 145046
rect 147644 145004 149068 145324
rect 147644 144644 147964 145004
rect 77540 144602 147964 144644
rect 77540 144366 77582 144602
rect 77818 144366 95062 144602
rect 95298 144366 147964 144602
rect 77540 144324 147964 144366
rect 148748 144644 149068 145004
rect 148748 144602 188076 144644
rect 148748 144366 187798 144602
rect 188034 144366 188076 144602
rect 148748 144324 188076 144366
rect 75148 143922 78228 143964
rect 75148 143686 75190 143922
rect 75426 143686 77950 143922
rect 78186 143686 78228 143922
rect 75148 143644 78228 143686
rect 74780 143242 147228 143284
rect 74780 143006 74822 143242
rect 75058 143006 109598 143242
rect 109834 143006 137014 143242
rect 137250 143006 146950 143242
rect 147186 143006 147228 143242
rect 74780 142964 147228 143006
rect 148748 143242 149068 144324
rect 164204 143644 167284 143964
rect 148748 143006 148790 143242
rect 149026 143006 149068 143242
rect 148748 142964 149068 143006
rect 150220 143242 156980 143284
rect 150220 143006 150262 143242
rect 150498 143006 156980 143242
rect 150220 142964 156980 143006
rect 156660 141924 156980 142964
rect 164204 141924 164524 143644
rect 166964 142604 167284 143644
rect 167700 143922 203348 143964
rect 167700 143686 169214 143922
rect 169450 143686 203070 143922
rect 203306 143686 203348 143922
rect 167700 143644 203348 143686
rect 167700 142604 168020 143644
rect 230996 143242 243092 143284
rect 230996 143006 231038 143242
rect 231274 143006 242814 143242
rect 243050 143006 243092 143242
rect 230996 142964 243092 143006
rect 243508 142604 243828 147724
rect 246268 143242 246588 150444
rect 262092 145004 264620 145324
rect 262092 144644 262412 145004
rect 261540 144602 262412 144644
rect 261540 144366 261582 144602
rect 261818 144366 262412 144602
rect 261540 144324 262412 144366
rect 262092 143284 262412 144324
rect 264300 143964 264620 145004
rect 264300 143922 282652 143964
rect 264300 143686 282374 143922
rect 282610 143686 282652 143922
rect 264300 143644 282652 143686
rect 283620 143922 302524 143964
rect 283620 143686 283662 143922
rect 283898 143686 302246 143922
rect 302482 143686 302524 143922
rect 283620 143644 302524 143686
rect 246268 143006 246310 143242
rect 246546 143006 246588 143242
rect 246268 142964 246588 143006
rect 247188 143242 262412 143284
rect 247188 143006 247230 143242
rect 247466 143006 262412 143242
rect 247188 142964 262412 143006
rect 262828 143242 297924 143284
rect 262828 143006 262870 143242
rect 263106 143006 297646 143242
rect 297882 143006 297924 143242
rect 262828 142964 297924 143006
rect 166964 142284 168020 142604
rect 242404 142562 243828 142604
rect 242404 142326 242446 142562
rect 242682 142326 243828 142562
rect 242404 142284 243828 142326
rect 249764 142562 250636 142604
rect 249764 142326 249806 142562
rect 250042 142326 250358 142562
rect 250594 142326 250636 142562
rect 249764 142284 250636 142326
rect 273500 142562 290196 142604
rect 273500 142326 289918 142562
rect 290154 142326 290196 142562
rect 273500 142284 290196 142326
rect 273500 141924 273820 142284
rect 74596 141882 106196 141924
rect 74596 141646 74638 141882
rect 74874 141646 105918 141882
rect 106154 141646 106196 141882
rect 74596 141604 106196 141646
rect 156660 141604 164524 141924
rect 255100 141882 273820 141924
rect 255100 141646 255142 141882
rect 255378 141646 273820 141882
rect 255100 141604 273820 141646
rect 137340 141202 146676 141244
rect 137340 140966 137382 141202
rect 137618 140966 146398 141202
rect 146634 140966 146676 141202
rect 137340 140924 146676 140966
rect 147092 141202 207764 141244
rect 147092 140966 151918 141202
rect 152154 140966 168478 141202
rect 168714 140966 207486 141202
rect 207722 140966 207764 141202
rect 147092 140924 207764 140966
rect 263564 140924 268852 141244
rect 147092 140564 147412 140924
rect 263564 140564 263884 140924
rect 137524 140522 147412 140564
rect 137524 140286 137566 140522
rect 137802 140286 147412 140522
rect 137524 140244 147412 140286
rect 148932 140522 197460 140564
rect 148932 140286 148974 140522
rect 149210 140286 167558 140522
rect 167794 140286 197182 140522
rect 197418 140286 197460 140522
rect 148932 140244 197460 140286
rect 231548 140522 245484 140564
rect 231548 140286 231590 140522
rect 231826 140286 245206 140522
rect 245442 140286 245484 140522
rect 231548 140244 245484 140286
rect 251236 140522 263884 140564
rect 251236 140286 251278 140522
rect 251514 140286 262318 140522
rect 262554 140286 263884 140522
rect 251236 140244 263884 140286
rect 268532 140564 268852 140924
rect 292820 141202 302156 141244
rect 292820 140966 301878 141202
rect 302114 140966 302156 141202
rect 292820 140924 302156 140966
rect 268532 140244 273452 140564
rect 273132 139884 273452 140244
rect 273868 140244 292404 140564
rect 273868 139884 274188 140244
rect 273132 139564 274188 139884
rect 292084 139884 292404 140244
rect 292820 139884 293140 140924
rect 292084 139564 293140 139884
rect 0 136992 444740 137034
rect 0 136756 5122 136992
rect 5358 136756 5442 136992
rect 5678 136756 5762 136992
rect 5998 136756 6082 136992
rect 6318 136756 6402 136992
rect 6638 136756 6722 136992
rect 6958 136756 7042 136992
rect 7278 136756 7362 136992
rect 7598 136756 7682 136992
rect 7918 136756 8002 136992
rect 8238 136756 8322 136992
rect 8558 136756 8642 136992
rect 8878 136756 435862 136992
rect 436098 136756 436182 136992
rect 436418 136756 436502 136992
rect 436738 136756 436822 136992
rect 437058 136756 437142 136992
rect 437378 136756 437462 136992
rect 437698 136756 437782 136992
rect 438018 136756 438102 136992
rect 438338 136756 438422 136992
rect 438658 136756 438742 136992
rect 438978 136756 439062 136992
rect 439298 136756 439382 136992
rect 439618 136756 444740 136992
rect 0 136714 444740 136756
rect 182788 131682 183108 131724
rect 182788 131446 182830 131682
rect 183066 131446 183108 131682
rect 182788 124244 183108 131446
rect 292268 131682 292772 131724
rect 292268 131446 292494 131682
rect 292730 131446 292772 131682
rect 292268 131404 292772 131446
rect 249028 127602 249532 127644
rect 249028 127366 249070 127602
rect 249306 127366 249532 127602
rect 249028 127324 249532 127366
rect 248476 126922 248796 126964
rect 248476 126686 248518 126922
rect 248754 126686 248796 126922
rect 248476 124244 248796 126686
rect 178556 124202 183108 124244
rect 178556 123966 178598 124202
rect 178834 123966 183108 124202
rect 178556 123924 183108 123966
rect 245716 124202 248796 124244
rect 245716 123966 245758 124202
rect 245994 123966 248796 124202
rect 245716 123924 248796 123966
rect 249212 123564 249532 127324
rect 292268 123564 292588 131404
rect 296684 123564 297188 124244
rect 316188 124202 322948 124244
rect 316188 123966 322670 124202
rect 322906 123966 322948 124202
rect 316188 123924 322948 123966
rect 245348 123522 249532 123564
rect 245348 123286 245390 123522
rect 245626 123286 249532 123522
rect 245348 123244 249532 123286
rect 287116 123244 306572 123564
rect 287116 122884 287436 123244
rect 242588 122842 258916 122884
rect 242588 122606 242630 122842
rect 242866 122606 258638 122842
rect 258874 122606 258916 122842
rect 242588 122564 258916 122606
rect 272580 122842 287436 122884
rect 272580 122606 272622 122842
rect 272858 122606 287436 122842
rect 272580 122564 287436 122606
rect 306252 122884 306572 123244
rect 316188 122884 316508 123924
rect 306252 122564 316508 122884
rect 0 121674 444740 121716
rect 0 121438 122 121674
rect 358 121438 442 121674
rect 678 121438 762 121674
rect 998 121438 1082 121674
rect 1318 121438 1402 121674
rect 1638 121438 1722 121674
rect 1958 121438 2042 121674
rect 2278 121438 2362 121674
rect 2598 121438 2682 121674
rect 2918 121438 3002 121674
rect 3238 121438 3322 121674
rect 3558 121438 3642 121674
rect 3878 121438 104506 121674
rect 104742 121438 198506 121674
rect 198742 121438 292506 121674
rect 292742 121438 440862 121674
rect 441098 121438 441182 121674
rect 441418 121438 441502 121674
rect 441738 121438 441822 121674
rect 442058 121438 442142 121674
rect 442378 121438 442462 121674
rect 442698 121438 442782 121674
rect 443018 121438 443102 121674
rect 443338 121438 443422 121674
rect 443658 121438 443742 121674
rect 443978 121438 444062 121674
rect 444298 121438 444382 121674
rect 444618 121438 444740 121674
rect 0 121396 444740 121438
rect 198244 120122 198748 120164
rect 198244 119886 198470 120122
rect 198706 119886 198748 120122
rect 198244 119844 198748 119886
rect 198244 118804 198564 119844
rect 154452 118484 158268 118804
rect 154452 118124 154772 118484
rect 145068 118082 154772 118124
rect 145068 117846 148422 118082
rect 148658 117846 154772 118082
rect 145068 117804 154772 117846
rect 145068 117444 145388 117804
rect 144884 117402 145388 117444
rect 144884 117166 144926 117402
rect 145162 117166 145388 117402
rect 144884 117124 145388 117166
rect 157948 116764 158268 118484
rect 196404 118484 208684 118804
rect 196404 116764 196724 118484
rect 208364 118124 208684 118484
rect 208364 117804 210156 118124
rect 209836 117444 210156 117804
rect 209836 117124 215676 117444
rect 136788 116722 138396 116764
rect 136788 116486 136830 116722
rect 137066 116486 138118 116722
rect 138354 116486 138396 116722
rect 136788 116444 138396 116486
rect 157580 116444 158268 116764
rect 190516 116444 196724 116764
rect 157580 116084 157900 116444
rect 190516 116084 190836 116444
rect 157580 116042 190836 116084
rect 157580 115806 163694 116042
rect 163930 115806 190836 116042
rect 157580 115764 190836 115806
rect 215356 116084 215676 117124
rect 235228 116722 245668 116764
rect 235228 116486 245390 116722
rect 245626 116486 245668 116722
rect 235228 116444 245668 116486
rect 235228 116084 235548 116444
rect 215356 116042 235548 116084
rect 215356 115806 228646 116042
rect 228882 115806 235548 116042
rect 215356 115764 235548 115806
rect 245716 113322 246036 113364
rect 245716 113086 245758 113322
rect 245994 113086 246036 113322
rect 245716 112684 246036 113086
rect 147644 112642 246036 112684
rect 147644 112406 147686 112642
rect 147922 112406 152102 112642
rect 152338 112406 230670 112642
rect 230906 112406 244102 112642
rect 244338 112406 246036 112642
rect 147644 112364 246036 112406
rect 84532 109922 90188 109964
rect 84532 109686 84574 109922
rect 84810 109686 90188 109922
rect 84532 109644 90188 109686
rect 89868 109284 90188 109644
rect 99436 109644 109508 109964
rect 99436 109284 99756 109644
rect 89868 108964 99756 109284
rect 109188 109284 109508 109644
rect 118756 109922 134900 109964
rect 118756 109686 134622 109922
rect 134858 109686 134900 109922
rect 118756 109644 134900 109686
rect 240012 109922 322948 109964
rect 240012 109686 240054 109922
rect 240290 109686 242078 109922
rect 242314 109686 322670 109922
rect 322906 109686 322948 109922
rect 240012 109644 322948 109686
rect 118756 109284 119076 109644
rect 109188 108964 119076 109284
rect 99252 108284 99756 108964
rect 118572 108284 119076 108964
rect 244612 108284 250084 108604
rect 244612 107244 244932 108284
rect 136788 107202 165076 107244
rect 136788 106966 136830 107202
rect 137066 106966 164798 107202
rect 165034 106966 165076 107202
rect 136788 106924 165076 106966
rect 230812 107202 244932 107244
rect 230812 106966 230854 107202
rect 231090 106966 244932 107202
rect 230812 106924 244932 106966
rect 249764 107244 250084 108284
rect 249764 107202 259100 107244
rect 249764 106966 258822 107202
rect 259058 106966 259100 107202
rect 249764 106924 259100 106966
rect 0 106356 444740 106398
rect 0 106120 5122 106356
rect 5358 106120 5442 106356
rect 5678 106120 5762 106356
rect 5998 106120 6082 106356
rect 6318 106120 6402 106356
rect 6638 106120 6722 106356
rect 6958 106120 7042 106356
rect 7278 106120 7362 106356
rect 7598 106120 7682 106356
rect 7918 106120 8002 106356
rect 8238 106120 8322 106356
rect 8558 106120 8642 106356
rect 8878 106120 89146 106356
rect 89382 106120 183146 106356
rect 183382 106120 277146 106356
rect 277382 106120 435862 106356
rect 436098 106120 436182 106356
rect 436418 106120 436502 106356
rect 436738 106120 436822 106356
rect 437058 106120 437142 106356
rect 437378 106120 437462 106356
rect 437698 106120 437782 106356
rect 438018 106120 438102 106356
rect 438338 106120 438422 106356
rect 438658 106120 438742 106356
rect 438978 106120 439062 106356
rect 439298 106120 439382 106356
rect 439618 106120 444740 106356
rect 0 106078 444740 106120
rect 200268 102164 209972 102484
rect 200268 101124 200588 102164
rect 209652 101124 209972 102164
rect 219772 102442 228924 102484
rect 219772 102206 228646 102442
rect 228882 102206 228924 102442
rect 219772 102164 228924 102206
rect 296868 102164 306572 102484
rect 219772 101124 220092 102164
rect 296868 101124 297188 102164
rect 306252 101124 306572 102164
rect 136788 101082 138396 101124
rect 136788 100846 136830 101082
rect 137066 100846 138396 101082
rect 136788 100804 138396 100846
rect 138076 99764 138396 100804
rect 150404 100804 154956 101124
rect 178004 101082 200588 101124
rect 178004 100846 178046 101082
rect 178282 100846 200588 101082
rect 178004 100804 200588 100846
rect 201004 100804 209236 101124
rect 209652 100804 220092 101124
rect 220692 101082 234628 101124
rect 220692 100846 228646 101082
rect 228882 100846 234628 101082
rect 220692 100804 234628 100846
rect 272580 101082 297188 101124
rect 272580 100846 272622 101082
rect 272858 100846 297188 101082
rect 272580 100804 297188 100846
rect 297604 100804 305836 101124
rect 306252 101082 323316 101124
rect 306252 100846 323038 101082
rect 323274 100846 323316 101082
rect 306252 100804 323316 100846
rect 150404 100444 150724 100804
rect 140836 100124 150724 100444
rect 140836 99764 141156 100124
rect 138076 99444 141156 99764
rect 154636 99084 154956 100804
rect 201004 100444 201324 100804
rect 158316 100402 176300 100444
rect 158316 100166 176022 100402
rect 176258 100166 176300 100402
rect 158316 100124 176300 100166
rect 176900 100402 183844 100444
rect 176900 100166 176942 100402
rect 177178 100166 183844 100402
rect 176900 100124 183844 100166
rect 158316 99084 158636 100124
rect 154636 98764 158636 99084
rect 183524 99084 183844 100124
rect 190332 100124 201324 100444
rect 208916 100444 209236 100804
rect 208916 100124 219908 100444
rect 190332 99084 190652 100124
rect 219588 99764 219908 100124
rect 220692 99764 221012 100804
rect 219588 99444 221012 99764
rect 234308 99764 234628 100804
rect 297604 100444 297924 100804
rect 251236 100124 254316 100444
rect 251236 99764 251556 100124
rect 234308 99444 241988 99764
rect 183524 98764 190652 99084
rect 241668 98404 241988 99444
rect 251052 99444 251556 99764
rect 253996 99764 254316 100124
rect 260804 100402 263332 100444
rect 260804 100166 263054 100402
rect 263290 100166 263332 100402
rect 260804 100124 263332 100166
rect 273132 100124 277868 100444
rect 260804 99764 261124 100124
rect 253996 99444 261124 99764
rect 244612 99042 246404 99084
rect 244612 98806 244654 99042
rect 244890 98806 246126 99042
rect 246362 98806 246404 99042
rect 244612 98764 246404 98806
rect 251052 98404 251372 99444
rect 273132 99084 273452 100124
rect 264300 99042 273452 99084
rect 264300 98806 264342 99042
rect 264578 98806 273452 99042
rect 264300 98764 273452 98806
rect 277548 99084 277868 100124
rect 286932 100124 297924 100444
rect 305516 100444 305836 100804
rect 305516 100402 322948 100444
rect 305516 100166 322670 100402
rect 322906 100166 322948 100402
rect 305516 100124 322948 100166
rect 286932 99084 287252 100124
rect 277548 98764 287252 99084
rect 241668 98084 251372 98404
rect 160892 96322 163972 96364
rect 160892 96086 163694 96322
rect 163930 96086 163972 96322
rect 160892 96044 163972 96086
rect 178004 96322 181268 96364
rect 178004 96086 178046 96322
rect 178282 96086 181268 96322
rect 178004 96044 181268 96086
rect 160892 95684 161212 96044
rect 180948 95684 181268 96044
rect 211308 96044 220828 96364
rect 244060 96322 246036 96364
rect 244060 96086 244102 96322
rect 244338 96086 245758 96322
rect 245994 96086 246036 96322
rect 244060 96044 246036 96086
rect 211308 95684 211628 96044
rect 160892 95642 163972 95684
rect 160892 95406 163694 95642
rect 163930 95406 163972 95642
rect 160892 95364 163972 95406
rect 178004 95642 181268 95684
rect 178004 95406 178046 95642
rect 178282 95406 181268 95642
rect 178004 95364 181268 95406
rect 181684 95364 186788 95684
rect 181684 95004 182004 95364
rect 148380 94962 161948 95004
rect 148380 94726 148422 94962
rect 148658 94726 161948 94962
rect 148380 94684 161948 94726
rect 178556 94962 182004 95004
rect 178556 94726 178598 94962
rect 178834 94726 182004 94962
rect 178556 94684 182004 94726
rect 186468 95004 186788 95364
rect 196036 95364 211628 95684
rect 196036 95004 196356 95364
rect 186468 94684 196356 95004
rect 220508 95004 220828 96044
rect 250868 95642 258916 95684
rect 250868 95548 258638 95642
rect 250730 95406 258638 95548
rect 258874 95406 258916 95642
rect 250730 95364 258916 95406
rect 272580 95642 283388 95684
rect 272580 95406 272622 95642
rect 272858 95406 283388 95642
rect 272580 95364 283388 95406
rect 250730 95228 251188 95364
rect 250730 95004 251050 95228
rect 220508 94962 229292 95004
rect 220508 94726 229014 94962
rect 229250 94726 229292 94962
rect 220508 94684 229292 94726
rect 242404 94962 251050 95004
rect 242404 94726 242446 94962
rect 242682 94726 251050 94962
rect 242404 94684 251050 94726
rect 283068 95004 283388 95364
rect 292636 95364 312276 95684
rect 292636 95004 292956 95364
rect 283068 94684 292956 95004
rect 161628 93644 161948 94684
rect 195852 94004 196356 94684
rect 292452 94004 292956 94684
rect 311956 94324 312276 95364
rect 311956 94282 322948 94324
rect 311956 94046 322670 94282
rect 322906 94046 322948 94282
rect 311956 94004 322948 94046
rect 161628 93602 165076 93644
rect 161628 93366 164798 93602
rect 165034 93366 165076 93602
rect 161628 93324 165076 93366
rect 0 91038 444740 91080
rect 0 90802 122 91038
rect 358 90802 442 91038
rect 678 90802 762 91038
rect 998 90802 1082 91038
rect 1318 90802 1402 91038
rect 1638 90802 1722 91038
rect 1958 90802 2042 91038
rect 2278 90802 2362 91038
rect 2598 90802 2682 91038
rect 2918 90802 3002 91038
rect 3238 90802 3322 91038
rect 3558 90802 3642 91038
rect 3878 90802 104506 91038
rect 104742 90802 198506 91038
rect 198742 90802 292506 91038
rect 292742 90802 440862 91038
rect 441098 90802 441182 91038
rect 441418 90802 441502 91038
rect 441738 90802 441822 91038
rect 442058 90802 442142 91038
rect 442378 90802 442462 91038
rect 442698 90802 442782 91038
rect 443018 90802 443102 91038
rect 443338 90802 443422 91038
rect 443658 90802 443742 91038
rect 443978 90802 444062 91038
rect 444298 90802 444382 91038
rect 444618 90802 444740 91038
rect 0 90760 444740 90802
rect 249028 88842 264068 88884
rect 249028 88606 249070 88842
rect 249306 88606 263790 88842
rect 264026 88606 264068 88842
rect 249028 88564 264068 88606
rect 244980 88162 252292 88204
rect 244980 87926 245022 88162
rect 245258 87926 252014 88162
rect 252250 87926 252292 88162
rect 244980 87884 252292 87926
rect 178556 86802 182740 86844
rect 178556 86566 178598 86802
rect 178834 86566 182740 86802
rect 178556 86524 182740 86566
rect 182420 85442 182740 86524
rect 182420 85206 182462 85442
rect 182698 85206 182740 85442
rect 182420 85164 182740 85206
rect 0 75720 444740 75762
rect 0 75484 5122 75720
rect 5358 75484 5442 75720
rect 5678 75484 5762 75720
rect 5998 75484 6082 75720
rect 6318 75484 6402 75720
rect 6638 75484 6722 75720
rect 6958 75484 7042 75720
rect 7278 75484 7362 75720
rect 7598 75484 7682 75720
rect 7918 75484 8002 75720
rect 8238 75484 8322 75720
rect 8558 75484 8642 75720
rect 8878 75484 435862 75720
rect 436098 75484 436182 75720
rect 436418 75484 436502 75720
rect 436738 75484 436822 75720
rect 437058 75484 437142 75720
rect 437378 75484 437462 75720
rect 437698 75484 437782 75720
rect 438018 75484 438102 75720
rect 438338 75484 438422 75720
rect 438658 75484 438742 75720
rect 438978 75484 439062 75720
rect 439298 75484 439382 75720
rect 439618 75484 444740 75720
rect 0 75442 444740 75484
rect 72388 73882 72708 73924
rect 72388 73646 72430 73882
rect 72666 73646 72708 73882
rect 72388 69164 72708 73646
rect 148380 73882 148700 73924
rect 148380 73646 148422 73882
rect 148658 73646 148700 73882
rect 148380 70524 148700 73646
rect 242588 73882 242908 73924
rect 242588 73646 242630 73882
rect 242866 73646 242908 73882
rect 148380 70204 148884 70524
rect 72388 69122 74916 69164
rect 72388 68886 74638 69122
rect 74874 68886 74916 69122
rect 72388 68844 74916 68886
rect 148564 63724 148884 70204
rect 242588 69164 242908 73646
rect 237252 69122 242908 69164
rect 237252 68886 237294 69122
rect 237530 68886 242908 69122
rect 237252 68844 242908 68886
rect 144700 63682 148884 63724
rect 144700 63446 144742 63682
rect 144978 63446 148884 63682
rect 144700 63404 148884 63446
rect 73308 61642 75284 61684
rect 73308 61406 73350 61642
rect 73586 61406 75006 61642
rect 75242 61406 75284 61642
rect 73308 61364 75284 61406
rect 0 60402 444740 60444
rect 0 60166 122 60402
rect 358 60166 442 60402
rect 678 60166 762 60402
rect 998 60166 1082 60402
rect 1318 60166 1402 60402
rect 1638 60166 1722 60402
rect 1958 60166 2042 60402
rect 2278 60166 2362 60402
rect 2598 60166 2682 60402
rect 2918 60166 3002 60402
rect 3238 60166 3322 60402
rect 3558 60166 3642 60402
rect 3878 60166 440862 60402
rect 441098 60166 441182 60402
rect 441418 60166 441502 60402
rect 441738 60166 441822 60402
rect 442058 60166 442142 60402
rect 442378 60166 442462 60402
rect 442698 60166 442782 60402
rect 443018 60166 443102 60402
rect 443338 60166 443422 60402
rect 443658 60166 443742 60402
rect 443978 60166 444062 60402
rect 444298 60166 444382 60402
rect 444618 60166 444740 60402
rect 0 60124 444740 60166
rect 73860 59602 75652 59644
rect 73860 59366 73902 59602
rect 74138 59366 75374 59602
rect 75610 59366 75652 59602
rect 73860 59324 75652 59366
rect 237252 59602 238492 59644
rect 237252 59366 237294 59602
rect 237530 59366 238214 59602
rect 238450 59366 238492 59602
rect 237252 59324 238492 59366
rect 144700 54842 148148 54884
rect 144700 54606 144742 54842
rect 144978 54606 148148 54842
rect 144700 54564 148148 54606
rect 147828 54204 148148 54564
rect 144700 54162 148148 54204
rect 144700 53926 144742 54162
rect 144978 53926 148148 54162
rect 144700 53884 148148 53926
rect 78828 53482 134348 53524
rect 78828 53246 78870 53482
rect 79106 53246 113462 53482
rect 113698 53246 134070 53482
rect 134306 53246 134348 53482
rect 78828 53204 134348 53246
rect 173772 53482 228188 53524
rect 173772 53246 173814 53482
rect 174050 53246 207670 53482
rect 207906 53246 227910 53482
rect 228146 53246 228188 53482
rect 173772 53204 228188 53246
rect 266508 53482 322028 53524
rect 266508 53246 266550 53482
rect 266786 53246 301510 53482
rect 301746 53246 321750 53482
rect 321986 53246 322028 53482
rect 266508 53204 322028 53246
rect 102380 51442 142996 51484
rect 102380 51206 102422 51442
rect 102658 51206 142718 51442
rect 142954 51206 142996 51442
rect 102380 51164 142996 51206
rect 93548 50762 280628 50804
rect 93548 50526 93590 50762
rect 93826 50526 187246 50762
rect 187482 50526 237478 50762
rect 237714 50526 238214 50762
rect 238450 50526 280350 50762
rect 280586 50526 280628 50762
rect 93548 50484 280628 50526
rect 73308 49402 87428 49444
rect 73308 49166 73350 49402
rect 73586 49166 87150 49402
rect 87386 49166 87428 49402
rect 73308 49124 87428 49166
rect 105140 49402 145020 49444
rect 105140 49166 105182 49402
rect 105418 49166 144742 49402
rect 144978 49166 145020 49402
rect 105140 49124 145020 49166
rect 147828 49402 148148 50484
rect 263196 50082 275108 50124
rect 263196 49846 263238 50082
rect 263474 49846 274830 50082
rect 275066 49846 275108 50082
rect 263196 49804 275108 49846
rect 147828 49166 147870 49402
rect 148106 49166 148148 49402
rect 147828 49124 148148 49166
rect 167884 49402 182004 49444
rect 167884 49166 167926 49402
rect 168162 49166 181726 49402
rect 181962 49166 182004 49402
rect 167884 49124 182004 49166
rect 204132 49402 275108 49444
rect 204132 49166 204174 49402
rect 204410 49166 262318 49402
rect 262554 49166 274830 49402
rect 275066 49166 275108 49402
rect 204132 49124 275108 49166
rect 73124 48722 87428 48764
rect 73124 48486 73166 48722
rect 73402 48486 74454 48722
rect 74690 48486 87150 48722
rect 87386 48486 87428 48722
rect 73124 48444 87428 48486
rect 154636 48722 191572 48764
rect 154636 48486 154678 48722
rect 154914 48486 167558 48722
rect 167794 48486 191294 48722
rect 191530 48486 191572 48722
rect 154636 48444 191572 48486
rect 248476 48722 264068 48764
rect 248476 48486 248518 48722
rect 248754 48486 263790 48722
rect 264026 48486 264068 48722
rect 248476 48444 264068 48486
rect 159972 48042 182372 48084
rect 159972 47806 160014 48042
rect 160250 47806 169030 48042
rect 169266 47806 182094 48042
rect 182330 47806 182372 48042
rect 159972 47764 182372 47806
rect 253812 48042 275108 48084
rect 253812 47806 253854 48042
rect 254090 47806 261398 48042
rect 261634 47806 274830 48042
rect 275066 47806 275108 48042
rect 253812 47764 275108 47806
rect 110292 47362 159188 47404
rect 110292 47126 110334 47362
rect 110570 47126 158910 47362
rect 159146 47126 159188 47362
rect 110292 47084 159188 47126
rect 162732 47362 181222 47404
rect 162732 47126 162774 47362
rect 163010 47126 181222 47362
rect 162732 47084 181222 47126
rect 180902 46724 181222 47084
rect 190332 47084 199852 47404
rect 248476 47362 264068 47404
rect 248476 47126 248518 47362
rect 248754 47126 263790 47362
rect 264026 47126 264068 47362
rect 248476 47084 264068 47126
rect 107348 46682 157716 46724
rect 107348 46446 107390 46682
rect 107626 46446 157438 46682
rect 157674 46446 157716 46682
rect 107348 46404 157716 46446
rect 180902 46682 181562 46724
rect 180902 46446 180990 46682
rect 181226 46446 181562 46682
rect 180902 46404 181562 46446
rect 180902 46044 181222 46404
rect 190332 46044 190652 47084
rect 199532 46724 199852 47084
rect 199532 46682 252844 46724
rect 199532 46446 199574 46682
rect 199810 46446 252566 46682
rect 252802 46446 252844 46682
rect 199532 46404 252844 46446
rect 260252 46682 276028 46724
rect 260252 46446 260294 46682
rect 260530 46446 261766 46682
rect 262002 46446 275750 46682
rect 275986 46446 276028 46682
rect 260252 46404 276028 46446
rect 180902 45724 190652 46044
rect 0 45084 444740 45126
rect 0 44848 5122 45084
rect 5358 44848 5442 45084
rect 5678 44848 5762 45084
rect 5998 44848 6082 45084
rect 6318 44848 6402 45084
rect 6638 44848 6722 45084
rect 6958 44848 7042 45084
rect 7278 44848 7362 45084
rect 7598 44848 7682 45084
rect 7918 44848 8002 45084
rect 8238 44848 8322 45084
rect 8558 44848 8642 45084
rect 8878 44848 435862 45084
rect 436098 44848 436182 45084
rect 436418 44848 436502 45084
rect 436738 44848 436822 45084
rect 437058 44848 437142 45084
rect 437378 44848 437462 45084
rect 437698 44848 437782 45084
rect 438018 44848 438102 45084
rect 438338 44848 438422 45084
rect 438658 44848 438742 45084
rect 438978 44848 439062 45084
rect 439298 44848 439382 45084
rect 439618 44848 444740 45084
rect 0 44806 444740 44848
rect 0 29766 444740 29808
rect 0 29530 122 29766
rect 358 29530 442 29766
rect 678 29530 762 29766
rect 998 29530 1082 29766
rect 1318 29530 1402 29766
rect 1638 29530 1722 29766
rect 1958 29530 2042 29766
rect 2278 29530 2362 29766
rect 2598 29530 2682 29766
rect 2918 29530 3002 29766
rect 3238 29530 3322 29766
rect 3558 29530 3642 29766
rect 3878 29530 440862 29766
rect 441098 29530 441182 29766
rect 441418 29530 441502 29766
rect 441738 29530 441822 29766
rect 442058 29530 442142 29766
rect 442378 29530 442462 29766
rect 442698 29530 442782 29766
rect 443018 29530 443102 29766
rect 443338 29530 443422 29766
rect 443658 29530 443742 29766
rect 443978 29530 444062 29766
rect 444298 29530 444382 29766
rect 444618 29530 444740 29766
rect 0 29488 444740 29530
rect 0 14448 444740 14490
rect 0 14212 5122 14448
rect 5358 14212 5442 14448
rect 5678 14212 5762 14448
rect 5998 14212 6082 14448
rect 6318 14212 6402 14448
rect 6638 14212 6722 14448
rect 6958 14212 7042 14448
rect 7278 14212 7362 14448
rect 7598 14212 7682 14448
rect 7918 14212 8002 14448
rect 8238 14212 8322 14448
rect 8558 14212 8642 14448
rect 8878 14212 435862 14448
rect 436098 14212 436182 14448
rect 436418 14212 436502 14448
rect 436738 14212 436822 14448
rect 437058 14212 437142 14448
rect 437378 14212 437462 14448
rect 437698 14212 437782 14448
rect 438018 14212 438102 14448
rect 438338 14212 438422 14448
rect 438658 14212 438742 14448
rect 438978 14212 439062 14448
rect 439298 14212 439382 14448
rect 439618 14212 444740 14448
rect 0 14170 444740 14212
rect 5000 8878 439740 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 435862 8878
rect 436098 8642 436182 8878
rect 436418 8642 436502 8878
rect 436738 8642 436822 8878
rect 437058 8642 437142 8878
rect 437378 8642 437462 8878
rect 437698 8642 437782 8878
rect 438018 8642 438102 8878
rect 438338 8642 438422 8878
rect 438658 8642 438742 8878
rect 438978 8642 439062 8878
rect 439298 8642 439382 8878
rect 439618 8642 439740 8878
rect 5000 8558 439740 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 435862 8558
rect 436098 8322 436182 8558
rect 436418 8322 436502 8558
rect 436738 8322 436822 8558
rect 437058 8322 437142 8558
rect 437378 8322 437462 8558
rect 437698 8322 437782 8558
rect 438018 8322 438102 8558
rect 438338 8322 438422 8558
rect 438658 8322 438742 8558
rect 438978 8322 439062 8558
rect 439298 8322 439382 8558
rect 439618 8322 439740 8558
rect 5000 8238 439740 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 435862 8238
rect 436098 8002 436182 8238
rect 436418 8002 436502 8238
rect 436738 8002 436822 8238
rect 437058 8002 437142 8238
rect 437378 8002 437462 8238
rect 437698 8002 437782 8238
rect 438018 8002 438102 8238
rect 438338 8002 438422 8238
rect 438658 8002 438742 8238
rect 438978 8002 439062 8238
rect 439298 8002 439382 8238
rect 439618 8002 439740 8238
rect 5000 7918 439740 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 435862 7918
rect 436098 7682 436182 7918
rect 436418 7682 436502 7918
rect 436738 7682 436822 7918
rect 437058 7682 437142 7918
rect 437378 7682 437462 7918
rect 437698 7682 437782 7918
rect 438018 7682 438102 7918
rect 438338 7682 438422 7918
rect 438658 7682 438742 7918
rect 438978 7682 439062 7918
rect 439298 7682 439382 7918
rect 439618 7682 439740 7918
rect 5000 7598 439740 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 435862 7598
rect 436098 7362 436182 7598
rect 436418 7362 436502 7598
rect 436738 7362 436822 7598
rect 437058 7362 437142 7598
rect 437378 7362 437462 7598
rect 437698 7362 437782 7598
rect 438018 7362 438102 7598
rect 438338 7362 438422 7598
rect 438658 7362 438742 7598
rect 438978 7362 439062 7598
rect 439298 7362 439382 7598
rect 439618 7362 439740 7598
rect 5000 7278 439740 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 435862 7278
rect 436098 7042 436182 7278
rect 436418 7042 436502 7278
rect 436738 7042 436822 7278
rect 437058 7042 437142 7278
rect 437378 7042 437462 7278
rect 437698 7042 437782 7278
rect 438018 7042 438102 7278
rect 438338 7042 438422 7278
rect 438658 7042 438742 7278
rect 438978 7042 439062 7278
rect 439298 7042 439382 7278
rect 439618 7042 439740 7278
rect 5000 6958 439740 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 435862 6958
rect 436098 6722 436182 6958
rect 436418 6722 436502 6958
rect 436738 6722 436822 6958
rect 437058 6722 437142 6958
rect 437378 6722 437462 6958
rect 437698 6722 437782 6958
rect 438018 6722 438102 6958
rect 438338 6722 438422 6958
rect 438658 6722 438742 6958
rect 438978 6722 439062 6958
rect 439298 6722 439382 6958
rect 439618 6722 439740 6958
rect 5000 6638 439740 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 435862 6638
rect 436098 6402 436182 6638
rect 436418 6402 436502 6638
rect 436738 6402 436822 6638
rect 437058 6402 437142 6638
rect 437378 6402 437462 6638
rect 437698 6402 437782 6638
rect 438018 6402 438102 6638
rect 438338 6402 438422 6638
rect 438658 6402 438742 6638
rect 438978 6402 439062 6638
rect 439298 6402 439382 6638
rect 439618 6402 439740 6638
rect 5000 6318 439740 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 435862 6318
rect 436098 6082 436182 6318
rect 436418 6082 436502 6318
rect 436738 6082 436822 6318
rect 437058 6082 437142 6318
rect 437378 6082 437462 6318
rect 437698 6082 437782 6318
rect 438018 6082 438102 6318
rect 438338 6082 438422 6318
rect 438658 6082 438742 6318
rect 438978 6082 439062 6318
rect 439298 6082 439382 6318
rect 439618 6082 439740 6318
rect 5000 5998 439740 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 435862 5998
rect 436098 5762 436182 5998
rect 436418 5762 436502 5998
rect 436738 5762 436822 5998
rect 437058 5762 437142 5998
rect 437378 5762 437462 5998
rect 437698 5762 437782 5998
rect 438018 5762 438102 5998
rect 438338 5762 438422 5998
rect 438658 5762 438742 5998
rect 438978 5762 439062 5998
rect 439298 5762 439382 5998
rect 439618 5762 439740 5998
rect 5000 5678 439740 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 435862 5678
rect 436098 5442 436182 5678
rect 436418 5442 436502 5678
rect 436738 5442 436822 5678
rect 437058 5442 437142 5678
rect 437378 5442 437462 5678
rect 437698 5442 437782 5678
rect 438018 5442 438102 5678
rect 438338 5442 438422 5678
rect 438658 5442 438742 5678
rect 438978 5442 439062 5678
rect 439298 5442 439382 5678
rect 439618 5442 439740 5678
rect 5000 5358 439740 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 435862 5358
rect 436098 5122 436182 5358
rect 436418 5122 436502 5358
rect 436738 5122 436822 5358
rect 437058 5122 437142 5358
rect 437378 5122 437462 5358
rect 437698 5122 437782 5358
rect 438018 5122 438102 5358
rect 438338 5122 438422 5358
rect 438658 5122 438742 5358
rect 438978 5122 439062 5358
rect 439298 5122 439382 5358
rect 439618 5122 439740 5358
rect 5000 5000 439740 5122
rect 0 3878 444740 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 440862 3878
rect 441098 3642 441182 3878
rect 441418 3642 441502 3878
rect 441738 3642 441822 3878
rect 442058 3642 442142 3878
rect 442378 3642 442462 3878
rect 442698 3642 442782 3878
rect 443018 3642 443102 3878
rect 443338 3642 443422 3878
rect 443658 3642 443742 3878
rect 443978 3642 444062 3878
rect 444298 3642 444382 3878
rect 444618 3642 444740 3878
rect 0 3558 444740 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 440862 3558
rect 441098 3322 441182 3558
rect 441418 3322 441502 3558
rect 441738 3322 441822 3558
rect 442058 3322 442142 3558
rect 442378 3322 442462 3558
rect 442698 3322 442782 3558
rect 443018 3322 443102 3558
rect 443338 3322 443422 3558
rect 443658 3322 443742 3558
rect 443978 3322 444062 3558
rect 444298 3322 444382 3558
rect 444618 3322 444740 3558
rect 0 3238 444740 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 440862 3238
rect 441098 3002 441182 3238
rect 441418 3002 441502 3238
rect 441738 3002 441822 3238
rect 442058 3002 442142 3238
rect 442378 3002 442462 3238
rect 442698 3002 442782 3238
rect 443018 3002 443102 3238
rect 443338 3002 443422 3238
rect 443658 3002 443742 3238
rect 443978 3002 444062 3238
rect 444298 3002 444382 3238
rect 444618 3002 444740 3238
rect 0 2918 444740 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 440862 2918
rect 441098 2682 441182 2918
rect 441418 2682 441502 2918
rect 441738 2682 441822 2918
rect 442058 2682 442142 2918
rect 442378 2682 442462 2918
rect 442698 2682 442782 2918
rect 443018 2682 443102 2918
rect 443338 2682 443422 2918
rect 443658 2682 443742 2918
rect 443978 2682 444062 2918
rect 444298 2682 444382 2918
rect 444618 2682 444740 2918
rect 0 2598 444740 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 440862 2598
rect 441098 2362 441182 2598
rect 441418 2362 441502 2598
rect 441738 2362 441822 2598
rect 442058 2362 442142 2598
rect 442378 2362 442462 2598
rect 442698 2362 442782 2598
rect 443018 2362 443102 2598
rect 443338 2362 443422 2598
rect 443658 2362 443742 2598
rect 443978 2362 444062 2598
rect 444298 2362 444382 2598
rect 444618 2362 444740 2598
rect 0 2278 444740 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 440862 2278
rect 441098 2042 441182 2278
rect 441418 2042 441502 2278
rect 441738 2042 441822 2278
rect 442058 2042 442142 2278
rect 442378 2042 442462 2278
rect 442698 2042 442782 2278
rect 443018 2042 443102 2278
rect 443338 2042 443422 2278
rect 443658 2042 443742 2278
rect 443978 2042 444062 2278
rect 444298 2042 444382 2278
rect 444618 2042 444740 2278
rect 0 1958 444740 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 440862 1958
rect 441098 1722 441182 1958
rect 441418 1722 441502 1958
rect 441738 1722 441822 1958
rect 442058 1722 442142 1958
rect 442378 1722 442462 1958
rect 442698 1722 442782 1958
rect 443018 1722 443102 1958
rect 443338 1722 443422 1958
rect 443658 1722 443742 1958
rect 443978 1722 444062 1958
rect 444298 1722 444382 1958
rect 444618 1722 444740 1958
rect 0 1638 444740 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 440862 1638
rect 441098 1402 441182 1638
rect 441418 1402 441502 1638
rect 441738 1402 441822 1638
rect 442058 1402 442142 1638
rect 442378 1402 442462 1638
rect 442698 1402 442782 1638
rect 443018 1402 443102 1638
rect 443338 1402 443422 1638
rect 443658 1402 443742 1638
rect 443978 1402 444062 1638
rect 444298 1402 444382 1638
rect 444618 1402 444740 1638
rect 0 1318 444740 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 440862 1318
rect 441098 1082 441182 1318
rect 441418 1082 441502 1318
rect 441738 1082 441822 1318
rect 442058 1082 442142 1318
rect 442378 1082 442462 1318
rect 442698 1082 442782 1318
rect 443018 1082 443102 1318
rect 443338 1082 443422 1318
rect 443658 1082 443742 1318
rect 443978 1082 444062 1318
rect 444298 1082 444382 1318
rect 444618 1082 444740 1318
rect 0 998 444740 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 440862 998
rect 441098 762 441182 998
rect 441418 762 441502 998
rect 441738 762 441822 998
rect 442058 762 442142 998
rect 442378 762 442462 998
rect 442698 762 442782 998
rect 443018 762 443102 998
rect 443338 762 443422 998
rect 443658 762 443742 998
rect 443978 762 444062 998
rect 444298 762 444382 998
rect 444618 762 444740 998
rect 0 678 444740 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 440862 678
rect 441098 442 441182 678
rect 441418 442 441502 678
rect 441738 442 441822 678
rect 442058 442 442142 678
rect 442378 442 442462 678
rect 442698 442 442782 678
rect 443018 442 443102 678
rect 443338 442 443422 678
rect 443658 442 443742 678
rect 443978 442 444062 678
rect 444298 442 444382 678
rect 444618 442 444740 678
rect 0 358 444740 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 440862 358
rect 441098 122 441182 358
rect 441418 122 441502 358
rect 441738 122 441822 358
rect 442058 122 442142 358
rect 442378 122 442462 358
rect 442698 122 442782 358
rect 443018 122 443102 358
rect 443338 122 443422 358
rect 443658 122 443742 358
rect 443978 122 444062 358
rect 444298 122 444382 358
rect 444618 122 444740 358
rect 0 0 444740 122
use sb_0__0_  sb_0__0_
timestamp 1603804930
transform 1 0 48895 0 1 47824
box 1 0 27528 28000
use grid_io_bottom  grid_io_bottom_1__0_
timestamp 1603804930
transform 1 0 89896 0 1 18824
box 0 0 38862 16000
use cbx_1__0_  cbx_1__0_
timestamp 1603804930
transform 1 0 89896 0 1 53824
box 0 0 40000 16000
use sb_1__0_  sb_1__0_
timestamp 1603804930
transform 1 0 142896 0 1 47824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_2__0_
timestamp 1603804930
transform 1 0 183896 0 1 18824
box 0 0 38862 16000
use cbx_1__0_  cbx_2__0_
timestamp 1603804930
transform 1 0 183896 0 1 53824
box 0 0 40000 16000
use sb_1__0_  sb_2__0_
timestamp 1603804930
transform 1 0 236896 0 1 47824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_3__0_
timestamp 1603804930
transform 1 0 277896 0 1 18824
box 0 0 38862 16000
use cbx_1__0_  cbx_3__0_
timestamp 1603804930
transform 1 0 277896 0 1 53824
box 0 0 40000 16000
use sb_3__0_  sb_3__0_
timestamp 1603804930
transform 1 0 330896 0 1 47824
box 0 0 27403 28000
use grid_io_left  grid_io_left_0__1_
timestamp 1603804930
transform 1 0 19896 0 1 88824
box 0 0 16000 38752
use cby_0__1_  cby_0__1_
timestamp 1603804930
transform 1 0 54896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_1__1_
timestamp 1603804930
transform 1 0 84896 0 1 83824
box 0 0 50000 50000
use cby_1__1_  cby_1__1_
timestamp 1603804930
transform 1 0 148896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_2__1_
timestamp 1603804930
transform 1 0 178896 0 1 83824
box 0 0 50000 50000
use cby_1__1_  cby_2__1_
timestamp 1603804930
transform 1 0 242896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_3__1_
timestamp 1603804930
transform 1 0 272896 0 1 83824
box 0 0 50000 50000
use cby_3__1_  cby_3__1_
timestamp 1603804930
transform 1 0 336896 0 1 88824
box 0 0 16000 40000
use grid_io_right  grid_io_right_4__1_
timestamp 1603804930
transform 1 0 408896 0 1 88824
box 0 0 16000 38752
use grid_io_left  grid_io_left_0__2_
timestamp 1603804930
transform 1 0 19896 0 1 182824
box 0 0 16000 38752
use sb_0__1_  sb_0__1_
timestamp 1603804930
transform 1 0 48896 0 1 141824
box 0 0 28000 28000
use cby_0__1_  cby_0__2_
timestamp 1603804930
transform 1 0 54896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_1__2_
timestamp 1603804930
transform 1 0 84896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_1__1_
timestamp 1603804930
transform 1 0 89896 0 1 147824
box 0 0 40000 16000
use sb_1__1_  sb_1__1_
timestamp 1603804930
transform 1 0 142896 0 1 141824
box 0 0 28000 28000
use cby_1__1_  cby_1__2_
timestamp 1603804930
transform 1 0 148896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1603804930
transform 1 0 178896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_2__1_
timestamp 1603804930
transform 1 0 183896 0 1 147824
box 0 0 40000 16000
use sb_1__1_  sb_2__1_
timestamp 1603804930
transform 1 0 236896 0 1 141824
box 0 0 28000 28000
use cby_1__1_  cby_2__2_
timestamp 1603804930
transform 1 0 242896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_3__2_
timestamp 1603804930
transform 1 0 272896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_3__1_
timestamp 1603804930
transform 1 0 277896 0 1 147824
box 0 0 40000 16000
use sb_3__1_  sb_3__1_
timestamp 1603804930
transform 1 0 330896 0 1 141824
box 0 0 28000 28000
use cby_3__1_  cby_3__2_
timestamp 1603804930
transform 1 0 336896 0 1 182824
box 0 0 16000 40000
use grid_io_right  grid_io_right_4__2_
timestamp 1603804930
transform 1 0 408896 0 1 182824
box 0 0 16000 38752
use sb_0__1_  sb_0__2_
timestamp 1603804930
transform 1 0 48896 0 1 235824
box 0 0 28000 28000
use cbx_1__1_  cbx_1__2_
timestamp 1603804930
transform 1 0 89896 0 1 241824
box 0 0 40000 16000
use sb_1__1_  sb_1__2_
timestamp 1603804930
transform 1 0 142896 0 1 235824
box 0 0 28000 28000
use cbx_1__1_  cbx_2__2_
timestamp 1603804930
transform 1 0 183896 0 1 241824
box 0 0 40000 16000
use sb_1__1_  sb_2__2_
timestamp 1603804930
transform 1 0 236896 0 1 235824
box 0 0 28000 28000
use cbx_1__1_  cbx_3__2_
timestamp 1603804930
transform 1 0 277896 0 1 241824
box 0 0 40000 16000
use sb_3__1_  sb_3__2_
timestamp 1603804930
transform 1 0 330896 0 1 235824
box 0 0 28000 28000
use decoder6to61  decoder6to61_0_
timestamp 1603804930
transform 1 0 371896 0 1 212824
box 0 0 22854 24000
use grid_io_left  grid_io_left_0__3_
timestamp 1603804930
transform 1 0 19896 0 1 276824
box 0 0 16000 38752
use cby_0__1_  cby_0__3_
timestamp 1603804930
transform 1 0 54896 0 1 276824
box 0 0 16000 40000
use grid_clb  grid_clb_1__3_
timestamp 1603804930
transform 1 0 84896 0 1 271824
box 0 0 50000 50000
use cby_1__1_  cby_1__3_
timestamp 1603804930
transform 1 0 148896 0 1 276824
box 0 0 16000 40000
use grid_clb  grid_clb_2__3_
timestamp 1603804930
transform 1 0 178896 0 1 271824
box 0 0 50000 50000
use cby_1__1_  cby_2__3_
timestamp 1603804930
transform 1 0 242896 0 1 276824
box 0 0 16000 40000
use grid_clb  grid_clb_3__3_
timestamp 1603804930
transform 1 0 272896 0 1 271824
box 0 0 50000 50000
use cby_3__1_  cby_3__3_
timestamp 1603804930
transform 1 0 336896 0 1 276824
box 0 0 16000 40000
use grid_io_right  grid_io_right_4__3_
timestamp 1603804930
transform 1 0 408896 0 1 276824
box 0 0 16000 38752
use sb_0__3_  sb_0__3_
timestamp 1603804930
transform 1 0 48895 0 1 329824
box 1 0 27528 28000
use grid_io_top  grid_io_top_1__4_
timestamp 1603804930
transform 1 0 89896 0 1 370824
box 0 0 38934 16000
use cbx_1__3_  cbx_1__3_
timestamp 1603804930
transform 1 0 89896 0 1 335824
box 0 0 40000 16000
use sb_1__3_  sb_1__3_
timestamp 1603804930
transform 1 0 142896 0 1 329824
box 0 0 28000 27464
use grid_io_top  grid_io_top_2__4_
timestamp 1603804930
transform 1 0 183896 0 1 370824
box 0 0 38934 16000
use cbx_1__3_  cbx_2__3_
timestamp 1603804930
transform 1 0 183896 0 1 335824
box 0 0 40000 16000
use sb_1__3_  sb_2__3_
timestamp 1603804930
transform 1 0 236896 0 1 329824
box 0 0 28000 27464
use grid_io_top  grid_io_top_3__4_
timestamp 1603804930
transform 1 0 277896 0 1 370824
box 0 0 38934 16000
use cbx_1__3_  cbx_3__3_
timestamp 1603804930
transform 1 0 277896 0 1 335824
box 0 0 40000 16000
use sb_3__3_  sb_3__3_
timestamp 1603804930
transform 1 0 330896 0 1 329824
box 0 0 27587 27464
<< labels >>
rlabel metal3 s 9896 272808 10376 272928 6 address[0]
port 0 nsew default input
rlabel metal3 s 434416 342168 434896 342288 6 address[10]
port 1 nsew default input
rlabel metal3 s 434416 354272 434896 354392 6 address[11]
port 2 nsew default input
rlabel metal3 s 9896 294296 10376 294416 6 address[12]
port 3 nsew default input
rlabel metal3 s 9896 305040 10376 305160 6 address[13]
port 4 nsew default input
rlabel metal2 s 368438 396344 368494 396824 6 address[14]
port 5 nsew default input
rlabel metal3 s 9896 315920 10376 316040 6 address[15]
port 6 nsew default input
rlabel metal2 s 325474 8824 325530 9304 6 address[1]
port 7 nsew default input
rlabel metal3 s 434416 305720 434896 305840 6 address[2]
port 8 nsew default input
rlabel metal2 s 338354 8824 338410 9304 6 address[3]
port 9 nsew default input
rlabel metal2 s 351234 8824 351290 9304 6 address[4]
port 10 nsew default input
rlabel metal2 s 341942 396344 341998 396824 6 address[5]
port 11 nsew default input
rlabel metal3 s 434416 317824 434896 317944 6 address[6]
port 12 nsew default input
rlabel metal3 s 9896 283552 10376 283672 6 address[7]
port 13 nsew default input
rlabel metal3 s 434416 330064 434896 330184 6 address[8]
port 14 nsew default input
rlabel metal2 s 364114 8824 364170 9304 6 address[9]
port 15 nsew default input
rlabel metal2 s 395026 396344 395082 396824 6 clk
port 16 nsew default input
rlabel metal3 s 9896 326664 10376 326784 6 data_in
port 17 nsew default input
rlabel metal2 s 376994 8824 377050 9304 6 enable
port 18 nsew default input
rlabel metal2 s 23162 396344 23218 396824 6 gfpga_pad_GPIO_PAD[0]
port 19 nsew default bidirectional
rlabel metal2 s 129422 396344 129478 396824 6 gfpga_pad_GPIO_PAD[10]
port 20 nsew default bidirectional
rlabel metal2 s 155918 396344 155974 396824 6 gfpga_pad_GPIO_PAD[11]
port 21 nsew default bidirectional
rlabel metal2 s 182506 396344 182562 396824 6 gfpga_pad_GPIO_PAD[12]
port 22 nsew default bidirectional
rlabel metal2 s 209094 396344 209150 396824 6 gfpga_pad_GPIO_PAD[13]
port 23 nsew default bidirectional
rlabel metal3 s 434416 366376 434896 366496 6 gfpga_pad_GPIO_PAD[14]
port 24 nsew default bidirectional
rlabel metal3 s 9896 380520 10376 380640 6 gfpga_pad_GPIO_PAD[15]
port 25 nsew default bidirectional
rlabel metal2 s 421614 396344 421670 396824 6 gfpga_pad_GPIO_PAD[16]
port 26 nsew default bidirectional
rlabel metal3 s 434416 378480 434896 378600 6 gfpga_pad_GPIO_PAD[17]
port 27 nsew default bidirectional
rlabel metal2 s 415634 8824 415690 9304 6 gfpga_pad_GPIO_PAD[18]
port 28 nsew default bidirectional
rlabel metal3 s 434416 390584 434896 390704 6 gfpga_pad_GPIO_PAD[19]
port 29 nsew default bidirectional
rlabel metal2 s 49658 396344 49714 396824 6 gfpga_pad_GPIO_PAD[1]
port 30 nsew default bidirectional
rlabel metal2 s 235682 396344 235738 396824 6 gfpga_pad_GPIO_PAD[20]
port 31 nsew default bidirectional
rlabel metal2 s 262178 396344 262234 396824 6 gfpga_pad_GPIO_PAD[21]
port 32 nsew default bidirectional
rlabel metal2 s 288766 396344 288822 396824 6 gfpga_pad_GPIO_PAD[22]
port 33 nsew default bidirectional
rlabel metal2 s 315354 396344 315410 396824 6 gfpga_pad_GPIO_PAD[23]
port 34 nsew default bidirectional
rlabel metal3 s 434416 14816 434896 14936 6 gfpga_pad_GPIO_PAD[24]
port 35 nsew default bidirectional
rlabel metal3 s 434416 26920 434896 27040 6 gfpga_pad_GPIO_PAD[25]
port 36 nsew default bidirectional
rlabel metal3 s 434416 39024 434896 39144 6 gfpga_pad_GPIO_PAD[26]
port 37 nsew default bidirectional
rlabel metal3 s 434416 51128 434896 51248 6 gfpga_pad_GPIO_PAD[27]
port 38 nsew default bidirectional
rlabel metal3 s 434416 63232 434896 63352 6 gfpga_pad_GPIO_PAD[28]
port 39 nsew default bidirectional
rlabel metal3 s 434416 75336 434896 75456 6 gfpga_pad_GPIO_PAD[29]
port 40 nsew default bidirectional
rlabel metal2 s 76246 396344 76302 396824 6 gfpga_pad_GPIO_PAD[2]
port 41 nsew default bidirectional
rlabel metal3 s 434416 87440 434896 87560 6 gfpga_pad_GPIO_PAD[30]
port 42 nsew default bidirectional
rlabel metal3 s 434416 99680 434896 99800 6 gfpga_pad_GPIO_PAD[31]
port 43 nsew default bidirectional
rlabel metal3 s 434416 111784 434896 111904 6 gfpga_pad_GPIO_PAD[32]
port 44 nsew default bidirectional
rlabel metal3 s 434416 123888 434896 124008 6 gfpga_pad_GPIO_PAD[33]
port 45 nsew default bidirectional
rlabel metal3 s 434416 135992 434896 136112 6 gfpga_pad_GPIO_PAD[34]
port 46 nsew default bidirectional
rlabel metal3 s 434416 148096 434896 148216 6 gfpga_pad_GPIO_PAD[35]
port 47 nsew default bidirectional
rlabel metal3 s 434416 160200 434896 160320 6 gfpga_pad_GPIO_PAD[36]
port 48 nsew default bidirectional
rlabel metal3 s 434416 172440 434896 172560 6 gfpga_pad_GPIO_PAD[37]
port 49 nsew default bidirectional
rlabel metal3 s 434416 184544 434896 184664 6 gfpga_pad_GPIO_PAD[38]
port 50 nsew default bidirectional
rlabel metal3 s 434416 196648 434896 196768 6 gfpga_pad_GPIO_PAD[39]
port 51 nsew default bidirectional
rlabel metal2 s 102834 396344 102890 396824 6 gfpga_pad_GPIO_PAD[3]
port 52 nsew default bidirectional
rlabel metal3 s 434416 208752 434896 208872 6 gfpga_pad_GPIO_PAD[40]
port 53 nsew default bidirectional
rlabel metal3 s 434416 220856 434896 220976 6 gfpga_pad_GPIO_PAD[41]
port 54 nsew default bidirectional
rlabel metal3 s 434416 232960 434896 233080 6 gfpga_pad_GPIO_PAD[42]
port 55 nsew default bidirectional
rlabel metal3 s 434416 245064 434896 245184 6 gfpga_pad_GPIO_PAD[43]
port 56 nsew default bidirectional
rlabel metal3 s 434416 257304 434896 257424 6 gfpga_pad_GPIO_PAD[44]
port 57 nsew default bidirectional
rlabel metal3 s 434416 269408 434896 269528 6 gfpga_pad_GPIO_PAD[45]
port 58 nsew default bidirectional
rlabel metal3 s 434416 281512 434896 281632 6 gfpga_pad_GPIO_PAD[46]
port 59 nsew default bidirectional
rlabel metal3 s 434416 293616 434896 293736 6 gfpga_pad_GPIO_PAD[47]
port 60 nsew default bidirectional
rlabel metal2 s 16354 8824 16410 9304 6 gfpga_pad_GPIO_PAD[48]
port 61 nsew default bidirectional
rlabel metal2 s 29234 8824 29290 9304 6 gfpga_pad_GPIO_PAD[49]
port 62 nsew default bidirectional
rlabel metal3 s 9896 337408 10376 337528 6 gfpga_pad_GPIO_PAD[4]
port 63 nsew default bidirectional
rlabel metal2 s 42114 8824 42170 9304 6 gfpga_pad_GPIO_PAD[50]
port 64 nsew default bidirectional
rlabel metal2 s 54994 8824 55050 9304 6 gfpga_pad_GPIO_PAD[51]
port 65 nsew default bidirectional
rlabel metal2 s 67874 8824 67930 9304 6 gfpga_pad_GPIO_PAD[52]
port 66 nsew default bidirectional
rlabel metal2 s 80754 8824 80810 9304 6 gfpga_pad_GPIO_PAD[53]
port 67 nsew default bidirectional
rlabel metal2 s 93634 8824 93690 9304 6 gfpga_pad_GPIO_PAD[54]
port 68 nsew default bidirectional
rlabel metal2 s 106514 8824 106570 9304 6 gfpga_pad_GPIO_PAD[55]
port 69 nsew default bidirectional
rlabel metal2 s 119394 8824 119450 9304 6 gfpga_pad_GPIO_PAD[56]
port 70 nsew default bidirectional
rlabel metal2 s 132274 8824 132330 9304 6 gfpga_pad_GPIO_PAD[57]
port 71 nsew default bidirectional
rlabel metal2 s 145154 8824 145210 9304 6 gfpga_pad_GPIO_PAD[58]
port 72 nsew default bidirectional
rlabel metal2 s 158034 8824 158090 9304 6 gfpga_pad_GPIO_PAD[59]
port 73 nsew default bidirectional
rlabel metal3 s 9896 348152 10376 348272 6 gfpga_pad_GPIO_PAD[5]
port 74 nsew default bidirectional
rlabel metal2 s 170914 8824 170970 9304 6 gfpga_pad_GPIO_PAD[60]
port 75 nsew default bidirectional
rlabel metal2 s 183794 8824 183850 9304 6 gfpga_pad_GPIO_PAD[61]
port 76 nsew default bidirectional
rlabel metal2 s 196674 8824 196730 9304 6 gfpga_pad_GPIO_PAD[62]
port 77 nsew default bidirectional
rlabel metal2 s 209554 8824 209610 9304 6 gfpga_pad_GPIO_PAD[63]
port 78 nsew default bidirectional
rlabel metal2 s 222434 8824 222490 9304 6 gfpga_pad_GPIO_PAD[64]
port 79 nsew default bidirectional
rlabel metal2 s 235314 8824 235370 9304 6 gfpga_pad_GPIO_PAD[65]
port 80 nsew default bidirectional
rlabel metal2 s 248194 8824 248250 9304 6 gfpga_pad_GPIO_PAD[66]
port 81 nsew default bidirectional
rlabel metal2 s 261074 8824 261130 9304 6 gfpga_pad_GPIO_PAD[67]
port 82 nsew default bidirectional
rlabel metal2 s 273954 8824 274010 9304 6 gfpga_pad_GPIO_PAD[68]
port 83 nsew default bidirectional
rlabel metal2 s 286834 8824 286890 9304 6 gfpga_pad_GPIO_PAD[69]
port 84 nsew default bidirectional
rlabel metal3 s 9896 359032 10376 359152 6 gfpga_pad_GPIO_PAD[6]
port 85 nsew default bidirectional
rlabel metal2 s 299714 8824 299770 9304 6 gfpga_pad_GPIO_PAD[70]
port 86 nsew default bidirectional
rlabel metal2 s 312594 8824 312650 9304 6 gfpga_pad_GPIO_PAD[71]
port 87 nsew default bidirectional
rlabel metal3 s 9896 14136 10376 14256 6 gfpga_pad_GPIO_PAD[72]
port 88 nsew default bidirectional
rlabel metal3 s 9896 24880 10376 25000 6 gfpga_pad_GPIO_PAD[73]
port 89 nsew default bidirectional
rlabel metal3 s 9896 35624 10376 35744 6 gfpga_pad_GPIO_PAD[74]
port 90 nsew default bidirectional
rlabel metal3 s 9896 46368 10376 46488 6 gfpga_pad_GPIO_PAD[75]
port 91 nsew default bidirectional
rlabel metal3 s 9896 57248 10376 57368 6 gfpga_pad_GPIO_PAD[76]
port 92 nsew default bidirectional
rlabel metal3 s 9896 67992 10376 68112 6 gfpga_pad_GPIO_PAD[77]
port 93 nsew default bidirectional
rlabel metal3 s 9896 78736 10376 78856 6 gfpga_pad_GPIO_PAD[78]
port 94 nsew default bidirectional
rlabel metal3 s 9896 89480 10376 89600 6 gfpga_pad_GPIO_PAD[79]
port 95 nsew default bidirectional
rlabel metal2 s 389874 8824 389930 9304 6 gfpga_pad_GPIO_PAD[7]
port 96 nsew default bidirectional
rlabel metal3 s 9896 100360 10376 100480 6 gfpga_pad_GPIO_PAD[80]
port 97 nsew default bidirectional
rlabel metal3 s 9896 111104 10376 111224 6 gfpga_pad_GPIO_PAD[81]
port 98 nsew default bidirectional
rlabel metal3 s 9896 121848 10376 121968 6 gfpga_pad_GPIO_PAD[82]
port 99 nsew default bidirectional
rlabel metal3 s 9896 132592 10376 132712 6 gfpga_pad_GPIO_PAD[83]
port 100 nsew default bidirectional
rlabel metal3 s 9896 143472 10376 143592 6 gfpga_pad_GPIO_PAD[84]
port 101 nsew default bidirectional
rlabel metal3 s 9896 154216 10376 154336 6 gfpga_pad_GPIO_PAD[85]
port 102 nsew default bidirectional
rlabel metal3 s 9896 164960 10376 165080 6 gfpga_pad_GPIO_PAD[86]
port 103 nsew default bidirectional
rlabel metal3 s 9896 175704 10376 175824 6 gfpga_pad_GPIO_PAD[87]
port 104 nsew default bidirectional
rlabel metal3 s 9896 186584 10376 186704 6 gfpga_pad_GPIO_PAD[88]
port 105 nsew default bidirectional
rlabel metal3 s 9896 197328 10376 197448 6 gfpga_pad_GPIO_PAD[89]
port 106 nsew default bidirectional
rlabel metal2 s 402754 8824 402810 9304 6 gfpga_pad_GPIO_PAD[8]
port 107 nsew default bidirectional
rlabel metal3 s 9896 208072 10376 208192 6 gfpga_pad_GPIO_PAD[90]
port 108 nsew default bidirectional
rlabel metal3 s 9896 218816 10376 218936 6 gfpga_pad_GPIO_PAD[91]
port 109 nsew default bidirectional
rlabel metal3 s 9896 229696 10376 229816 6 gfpga_pad_GPIO_PAD[92]
port 110 nsew default bidirectional
rlabel metal3 s 9896 240440 10376 240560 6 gfpga_pad_GPIO_PAD[93]
port 111 nsew default bidirectional
rlabel metal3 s 9896 251184 10376 251304 6 gfpga_pad_GPIO_PAD[94]
port 112 nsew default bidirectional
rlabel metal3 s 9896 261928 10376 262048 6 gfpga_pad_GPIO_PAD[95]
port 113 nsew default bidirectional
rlabel metal3 s 9896 369776 10376 369896 6 gfpga_pad_GPIO_PAD[9]
port 114 nsew default bidirectional
rlabel metal2 s 428514 8824 428570 9304 6 reset
port 115 nsew default input
rlabel metal3 s 9896 391264 10376 391384 6 set
port 116 nsew default input
rlabel metal5 s 5000 5000 439740 9000 8 vpwr
port 117 nsew default input
rlabel metal5 s 0 0 444740 4000 8 vgnd
port 118 nsew default input
<< properties >>
string FIXED_BBOX 0 0 444740 405520
<< end >>
