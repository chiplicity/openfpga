VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_bottom
  CLASS BLOCK ;
  FOREIGN grid_io_bottom ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 80.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 40.160 200.000 40.760 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.910 77.600 100.190 80.000 ;
    END
  END ccff_tail
  PIN gfpga_pad_GPIO_A
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.430 77.600 128.710 80.000 ;
    END
  END gfpga_pad_GPIO_A
  PIN gfpga_pad_GPIO_IE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 2.400 ;
    END
  END gfpga_pad_GPIO_IE
  PIN gfpga_pad_GPIO_OE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.950 77.600 157.230 80.000 ;
    END
  END gfpga_pad_GPIO_OE
  PIN gfpga_pad_GPIO_Y
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END gfpga_pad_GPIO_Y
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.470 77.600 185.750 80.000 ;
    END
  END prog_clk
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 77.600 14.630 80.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.870 77.600 43.150 80.000 ;
    END
  END top_width_0_height_0__pin_1_lower
  PIN top_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 77.600 71.670 80.000 ;
    END
  END top_width_0_height_0__pin_1_upper
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 38.055 10.640 39.655 68.240 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 71.385 10.640 72.985 68.240 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 68.085 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 68.240 ;
      LAYER met2 ;
        RECT 14.910 77.320 42.590 77.600 ;
        RECT 43.430 77.320 71.110 77.600 ;
        RECT 71.950 77.320 99.630 77.600 ;
        RECT 100.470 77.320 128.150 77.600 ;
        RECT 128.990 77.320 156.670 77.600 ;
        RECT 157.510 77.320 185.190 77.600 ;
        RECT 14.350 2.680 185.750 77.320 ;
        RECT 14.350 2.400 99.630 2.680 ;
        RECT 100.470 2.400 185.750 2.680 ;
      LAYER met3 ;
        RECT 2.400 41.160 197.600 68.165 ;
        RECT 2.800 39.760 197.200 41.160 ;
        RECT 2.400 10.715 197.600 39.760 ;
      LAYER met4 ;
        RECT 40.055 10.640 70.985 68.240 ;
        RECT 73.385 10.640 172.985 68.240 ;
  END
END grid_io_bottom
END LIBRARY

