magic
tech sky130A
magscale 1 2
timestamp 1606223963
<< locali >>
rect 9413 12087 9447 12189
rect 4077 11611 4111 11781
rect 12173 11679 12207 11849
rect 6377 10455 6411 10693
rect 10885 10115 10919 10217
rect 11989 9911 12023 10149
rect 14013 9979 14047 10081
rect 12817 9367 12851 9469
rect 3341 8959 3375 9129
rect 9413 8823 9447 9129
rect 6285 6239 6319 6409
rect 10057 6171 10091 6409
rect 12541 6171 12575 6341
rect 11529 5695 11563 5865
rect 14105 5151 14139 5321
rect 6469 4675 6503 4777
rect 3617 3927 3651 4233
rect 15301 2499 15335 2601
rect 13921 2363 13955 2465
<< viali >>
rect 8953 14569 8987 14603
rect 8033 14501 8067 14535
rect 6193 14433 6227 14467
rect 7941 14433 7975 14467
rect 9045 14433 9079 14467
rect 15945 14433 15979 14467
rect 6285 14365 6319 14399
rect 6469 14365 6503 14399
rect 8125 14365 8159 14399
rect 9229 14365 9263 14399
rect 5825 14229 5859 14263
rect 7573 14229 7607 14263
rect 8585 14229 8619 14263
rect 16129 14229 16163 14263
rect 2697 13889 2731 13923
rect 2881 13889 2915 13923
rect 5273 13889 5307 13923
rect 6193 13889 6227 13923
rect 6377 13889 6411 13923
rect 7665 13889 7699 13923
rect 7849 13889 7883 13923
rect 9229 13889 9263 13923
rect 10701 13889 10735 13923
rect 15669 13889 15703 13923
rect 9137 13821 9171 13855
rect 10609 13821 10643 13855
rect 15577 13821 15611 13855
rect 5089 13753 5123 13787
rect 9045 13753 9079 13787
rect 2237 13685 2271 13719
rect 2605 13685 2639 13719
rect 4721 13685 4755 13719
rect 5181 13685 5215 13719
rect 5733 13685 5767 13719
rect 6101 13685 6135 13719
rect 7205 13685 7239 13719
rect 7573 13685 7607 13719
rect 8677 13685 8711 13719
rect 10149 13685 10183 13719
rect 10517 13685 10551 13719
rect 15117 13685 15151 13719
rect 15485 13685 15519 13719
rect 16129 13685 16163 13719
rect 4905 13481 4939 13515
rect 8585 13481 8619 13515
rect 10149 13481 10183 13515
rect 15577 13481 15611 13515
rect 5825 13413 5859 13447
rect 5917 13413 5951 13447
rect 7481 13413 7515 13447
rect 11713 13413 11747 13447
rect 12725 13413 12759 13447
rect 16037 13413 16071 13447
rect 2513 13345 2547 13379
rect 4813 13345 4847 13379
rect 7389 13345 7423 13379
rect 8677 13345 8711 13379
rect 10057 13345 10091 13379
rect 13369 13345 13403 13379
rect 13636 13345 13670 13379
rect 15945 13345 15979 13379
rect 2605 13277 2639 13311
rect 2697 13277 2731 13311
rect 5089 13277 5123 13311
rect 6009 13277 6043 13311
rect 7573 13277 7607 13311
rect 8769 13277 8803 13311
rect 10333 13277 10367 13311
rect 11805 13277 11839 13311
rect 11989 13277 12023 13311
rect 12817 13277 12851 13311
rect 12909 13277 12943 13311
rect 16129 13277 16163 13311
rect 2145 13141 2179 13175
rect 4445 13141 4479 13175
rect 5457 13141 5491 13175
rect 7021 13141 7055 13175
rect 8217 13141 8251 13175
rect 9689 13141 9723 13175
rect 11345 13141 11379 13175
rect 12357 13141 12391 13175
rect 14749 13141 14783 13175
rect 3801 12937 3835 12971
rect 13829 12869 13863 12903
rect 2421 12801 2455 12835
rect 3433 12801 3467 12835
rect 4353 12801 4387 12835
rect 5457 12801 5491 12835
rect 7389 12801 7423 12835
rect 7573 12801 7607 12835
rect 8493 12801 8527 12835
rect 9597 12801 9631 12835
rect 11897 12801 11931 12835
rect 12449 12801 12483 12835
rect 2145 12733 2179 12767
rect 5181 12733 5215 12767
rect 7297 12733 7331 12767
rect 8309 12733 8343 12767
rect 9413 12733 9447 12767
rect 10057 12733 10091 12767
rect 10324 12733 10358 12767
rect 14105 12733 14139 12767
rect 15945 12733 15979 12767
rect 3157 12665 3191 12699
rect 4169 12665 4203 12699
rect 8401 12665 8435 12699
rect 9505 12665 9539 12699
rect 12694 12665 12728 12699
rect 14372 12665 14406 12699
rect 1777 12597 1811 12631
rect 2237 12597 2271 12631
rect 2789 12597 2823 12631
rect 3249 12597 3283 12631
rect 4261 12597 4295 12631
rect 4813 12597 4847 12631
rect 5273 12597 5307 12631
rect 6929 12597 6963 12631
rect 7941 12597 7975 12631
rect 9045 12597 9079 12631
rect 11437 12597 11471 12631
rect 15485 12597 15519 12631
rect 16129 12597 16163 12631
rect 1961 12393 1995 12427
rect 2053 12393 2087 12427
rect 2605 12393 2639 12427
rect 5825 12393 5859 12427
rect 7941 12393 7975 12427
rect 9045 12393 9079 12427
rect 9689 12393 9723 12427
rect 11897 12393 11931 12427
rect 15485 12393 15519 12427
rect 10784 12325 10818 12359
rect 2973 12257 3007 12291
rect 3065 12257 3099 12291
rect 4344 12257 4378 12291
rect 6828 12257 6862 12291
rect 8953 12257 8987 12291
rect 10517 12257 10551 12291
rect 12633 12257 12667 12291
rect 13820 12257 13854 12291
rect 15853 12257 15887 12291
rect 2237 12189 2271 12223
rect 3157 12189 3191 12223
rect 4077 12189 4111 12223
rect 6561 12189 6595 12223
rect 9229 12189 9263 12223
rect 9413 12189 9447 12223
rect 12725 12189 12759 12223
rect 12817 12189 12851 12223
rect 13553 12189 13587 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 1593 12053 1627 12087
rect 5457 12053 5491 12087
rect 8585 12053 8619 12087
rect 9413 12053 9447 12087
rect 12265 12053 12299 12087
rect 14933 12053 14967 12087
rect 3893 11849 3927 11883
rect 4169 11849 4203 11883
rect 5365 11849 5399 11883
rect 8401 11849 8435 11883
rect 10057 11849 10091 11883
rect 10333 11849 10367 11883
rect 11345 11849 11379 11883
rect 12173 11849 12207 11883
rect 13461 11849 13495 11883
rect 4077 11781 4111 11815
rect 1961 11713 1995 11747
rect 2145 11713 2179 11747
rect 2513 11645 2547 11679
rect 2780 11645 2814 11679
rect 4813 11713 4847 11747
rect 5917 11713 5951 11747
rect 10885 11713 10919 11747
rect 11989 11713 12023 11747
rect 13001 11713 13035 11747
rect 13921 11713 13955 11747
rect 14013 11713 14047 11747
rect 16129 11713 16163 11747
rect 5733 11645 5767 11679
rect 7021 11645 7055 11679
rect 7288 11645 7322 11679
rect 8677 11645 8711 11679
rect 8933 11645 8967 11679
rect 12173 11645 12207 11679
rect 13829 11645 13863 11679
rect 14473 11645 14507 11679
rect 4077 11577 4111 11611
rect 4537 11577 4571 11611
rect 10701 11577 10735 11611
rect 11713 11577 11747 11611
rect 14740 11577 14774 11611
rect 1501 11509 1535 11543
rect 1869 11509 1903 11543
rect 4629 11509 4663 11543
rect 5825 11509 5859 11543
rect 10793 11509 10827 11543
rect 11805 11509 11839 11543
rect 12449 11509 12483 11543
rect 12817 11509 12851 11543
rect 12909 11509 12943 11543
rect 15853 11509 15887 11543
rect 4169 11305 4203 11339
rect 7297 11305 7331 11339
rect 9045 11305 9079 11339
rect 11345 11305 11379 11339
rect 12265 11305 12299 11339
rect 2412 11237 2446 11271
rect 4537 11237 4571 11271
rect 7849 11237 7883 11271
rect 8953 11237 8987 11271
rect 10210 11237 10244 11271
rect 1593 11169 1627 11203
rect 2145 11169 2179 11203
rect 5448 11169 5482 11203
rect 7205 11169 7239 11203
rect 8493 11169 8527 11203
rect 11713 11169 11747 11203
rect 12633 11169 12667 11203
rect 13461 11169 13495 11203
rect 13921 11169 13955 11203
rect 14657 11169 14691 11203
rect 15761 11169 15795 11203
rect 15853 11169 15887 11203
rect 4629 11101 4663 11135
rect 4813 11101 4847 11135
rect 5181 11101 5215 11135
rect 7389 11101 7423 11135
rect 9229 11101 9263 11135
rect 9965 11101 9999 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 14013 11101 14047 11135
rect 14105 11101 14139 11135
rect 16037 11101 16071 11135
rect 6561 11033 6595 11067
rect 6837 11033 6871 11067
rect 8309 11033 8343 11067
rect 8585 11033 8619 11067
rect 11897 11033 11931 11067
rect 13277 11033 13311 11067
rect 13553 11033 13587 11067
rect 14841 11033 14875 11067
rect 1777 10965 1811 10999
rect 3525 10965 3559 10999
rect 15393 10965 15427 10999
rect 2789 10761 2823 10795
rect 6837 10761 6871 10795
rect 9229 10761 9263 10795
rect 9597 10761 9631 10795
rect 11345 10761 11379 10795
rect 6377 10693 6411 10727
rect 10333 10693 10367 10727
rect 1409 10625 1443 10659
rect 3617 10625 3651 10659
rect 5641 10625 5675 10659
rect 1676 10557 1710 10591
rect 3433 10557 3467 10591
rect 4077 10557 4111 10591
rect 4905 10557 4939 10591
rect 5365 10557 5399 10591
rect 7389 10625 7423 10659
rect 10885 10625 10919 10659
rect 11989 10625 12023 10659
rect 14933 10625 14967 10659
rect 6653 10557 6687 10591
rect 7205 10557 7239 10591
rect 7849 10557 7883 10591
rect 8116 10557 8150 10591
rect 9781 10557 9815 10591
rect 10701 10557 10735 10591
rect 12449 10557 12483 10591
rect 14381 10557 14415 10591
rect 7297 10489 7331 10523
rect 10793 10489 10827 10523
rect 11713 10489 11747 10523
rect 12694 10489 12728 10523
rect 15200 10489 15234 10523
rect 3065 10421 3099 10455
rect 3525 10421 3559 10455
rect 4261 10421 4295 10455
rect 4721 10421 4755 10455
rect 4997 10421 5031 10455
rect 5457 10421 5491 10455
rect 6377 10421 6411 10455
rect 6469 10421 6503 10455
rect 9873 10421 9907 10455
rect 11805 10421 11839 10455
rect 13829 10421 13863 10455
rect 14565 10421 14599 10455
rect 16313 10421 16347 10455
rect 1961 10217 1995 10251
rect 2973 10217 3007 10251
rect 5733 10217 5767 10251
rect 8217 10217 8251 10251
rect 10425 10217 10459 10251
rect 10517 10217 10551 10251
rect 10885 10217 10919 10251
rect 12081 10217 12115 10251
rect 12541 10217 12575 10251
rect 13093 10217 13127 10251
rect 13553 10217 13587 10251
rect 14565 10217 14599 10251
rect 15669 10217 15703 10251
rect 2329 10149 2363 10183
rect 2421 10149 2455 10183
rect 3433 10149 3467 10183
rect 4598 10149 4632 10183
rect 9045 10149 9079 10183
rect 11989 10149 12023 10183
rect 15761 10149 15795 10183
rect 1409 10081 1443 10115
rect 3341 10081 3375 10115
rect 4353 10081 4387 10115
rect 7104 10081 7138 10115
rect 8953 10081 8987 10115
rect 10885 10081 10919 10115
rect 11437 10081 11471 10115
rect 2605 10013 2639 10047
rect 3617 10013 3651 10047
rect 6837 10013 6871 10047
rect 9229 10013 9263 10047
rect 10609 10013 10643 10047
rect 11529 10013 11563 10047
rect 11713 10013 11747 10047
rect 1593 9945 1627 9979
rect 12449 10081 12483 10115
rect 13461 10081 13495 10115
rect 14013 10081 14047 10115
rect 14473 10081 14507 10115
rect 12633 10013 12667 10047
rect 13645 10013 13679 10047
rect 14749 10013 14783 10047
rect 15853 10013 15887 10047
rect 14013 9945 14047 9979
rect 14105 9945 14139 9979
rect 8585 9877 8619 9911
rect 10057 9877 10091 9911
rect 11069 9877 11103 9911
rect 11989 9877 12023 9911
rect 15301 9877 15335 9911
rect 8217 9673 8251 9707
rect 2789 9605 2823 9639
rect 3065 9605 3099 9639
rect 4997 9605 5031 9639
rect 8585 9605 8619 9639
rect 3617 9537 3651 9571
rect 5549 9537 5583 9571
rect 9229 9537 9263 9571
rect 11989 9537 12023 9571
rect 15209 9537 15243 9571
rect 15301 9537 15335 9571
rect 1409 9469 1443 9503
rect 1676 9469 1710 9503
rect 4077 9469 4111 9503
rect 5457 9469 5491 9503
rect 6009 9469 6043 9503
rect 6837 9469 6871 9503
rect 9597 9469 9631 9503
rect 11805 9469 11839 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 15117 9469 15151 9503
rect 15853 9469 15887 9503
rect 3433 9401 3467 9435
rect 7104 9401 7138 9435
rect 8953 9401 8987 9435
rect 9864 9401 9898 9435
rect 12449 9401 12483 9435
rect 13176 9401 13210 9435
rect 16129 9401 16163 9435
rect 3525 9333 3559 9367
rect 4261 9333 4295 9367
rect 5365 9333 5399 9367
rect 6193 9333 6227 9367
rect 9045 9333 9079 9367
rect 10977 9333 11011 9367
rect 11345 9333 11379 9367
rect 11713 9333 11747 9367
rect 12817 9333 12851 9367
rect 14289 9333 14323 9367
rect 14749 9333 14783 9367
rect 1593 9129 1627 9163
rect 3341 9129 3375 9163
rect 2136 9061 2170 9095
rect 1777 8993 1811 9027
rect 1869 8993 1903 9027
rect 9413 9129 9447 9163
rect 9689 9129 9723 9163
rect 12081 9129 12115 9163
rect 14013 9129 14047 9163
rect 14381 9129 14415 9163
rect 15301 9129 15335 9163
rect 4506 9061 4540 9095
rect 3525 8993 3559 9027
rect 4261 8993 4295 9027
rect 5917 8993 5951 9027
rect 6173 8993 6207 9027
rect 7757 8993 7791 9027
rect 7941 8993 7975 9027
rect 8208 8993 8242 9027
rect 3341 8925 3375 8959
rect 3249 8857 3283 8891
rect 7573 8857 7607 8891
rect 15761 9061 15795 9095
rect 10057 8993 10091 9027
rect 10968 8993 11002 9027
rect 12613 8993 12647 9027
rect 15669 8993 15703 9027
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 10701 8925 10735 8959
rect 12357 8925 12391 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 15853 8925 15887 8959
rect 13737 8857 13771 8891
rect 5641 8789 5675 8823
rect 7297 8789 7331 8823
rect 9321 8789 9355 8823
rect 9413 8789 9447 8823
rect 2145 8585 2179 8619
rect 4537 8585 4571 8619
rect 12633 8585 12667 8619
rect 1777 8517 1811 8551
rect 9505 8517 9539 8551
rect 11437 8517 11471 8551
rect 11529 8517 11563 8551
rect 14197 8517 14231 8551
rect 14473 8517 14507 8551
rect 2697 8449 2731 8483
rect 5825 8449 5859 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 10057 8449 10091 8483
rect 12081 8449 12115 8483
rect 12817 8449 12851 8483
rect 15025 8449 15059 8483
rect 16037 8449 16071 8483
rect 1593 8381 1627 8415
rect 3157 8381 3191 8415
rect 8217 8381 8251 8415
rect 11989 8381 12023 8415
rect 12474 8381 12508 8415
rect 13084 8381 13118 8415
rect 14841 8381 14875 8415
rect 15945 8381 15979 8415
rect 3424 8313 3458 8347
rect 4813 8313 4847 8347
rect 6285 8313 6319 8347
rect 7205 8313 7239 8347
rect 10302 8313 10336 8347
rect 11897 8313 11931 8347
rect 15853 8313 15887 8347
rect 2513 8245 2547 8279
rect 2605 8245 2639 8279
rect 5273 8245 5307 8279
rect 5641 8245 5675 8279
rect 5733 8245 5767 8279
rect 6837 8245 6871 8279
rect 14933 8245 14967 8279
rect 15485 8245 15519 8279
rect 2973 8041 3007 8075
rect 3341 8041 3375 8075
rect 6745 8041 6779 8075
rect 7113 8041 7147 8075
rect 7849 8041 7883 8075
rect 9045 8041 9079 8075
rect 11805 8041 11839 8075
rect 12081 8041 12115 8075
rect 13461 8041 13495 8075
rect 14105 8041 14139 8075
rect 15761 8041 15795 8075
rect 4344 7973 4378 8007
rect 6101 7973 6135 8007
rect 7205 7973 7239 8007
rect 9137 7973 9171 8007
rect 12541 7973 12575 8007
rect 14473 7973 14507 8007
rect 1409 7905 1443 7939
rect 2329 7905 2363 7939
rect 3433 7905 3467 7939
rect 8217 7905 8251 7939
rect 9873 7905 9907 7939
rect 10692 7905 10726 7939
rect 12449 7905 12483 7939
rect 15669 7905 15703 7939
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 3617 7837 3651 7871
rect 4077 7837 4111 7871
rect 6193 7837 6227 7871
rect 6285 7837 6319 7871
rect 7297 7837 7331 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 9321 7837 9355 7871
rect 10425 7837 10459 7871
rect 12633 7837 12667 7871
rect 13553 7837 13587 7871
rect 13645 7837 13679 7871
rect 14565 7837 14599 7871
rect 14749 7837 14783 7871
rect 15853 7837 15887 7871
rect 1593 7769 1627 7803
rect 13093 7769 13127 7803
rect 1961 7701 1995 7735
rect 5457 7701 5491 7735
rect 5733 7701 5767 7735
rect 8677 7701 8711 7735
rect 10057 7701 10091 7735
rect 15301 7701 15335 7735
rect 2237 7497 2271 7531
rect 4629 7497 4663 7531
rect 6837 7497 6871 7531
rect 8309 7497 8343 7531
rect 12449 7497 12483 7531
rect 14013 7497 14047 7531
rect 16221 7497 16255 7531
rect 7941 7429 7975 7463
rect 10057 7429 10091 7463
rect 11713 7429 11747 7463
rect 2789 7361 2823 7395
rect 5641 7361 5675 7395
rect 7389 7361 7423 7395
rect 12909 7361 12943 7395
rect 13093 7361 13127 7395
rect 14381 7361 14415 7395
rect 1593 7293 1627 7327
rect 3249 7293 3283 7327
rect 3516 7293 3550 7327
rect 5549 7293 5583 7327
rect 6101 7293 6135 7327
rect 7205 7293 7239 7327
rect 7757 7293 7791 7327
rect 8125 7293 8159 7327
rect 8677 7293 8711 7327
rect 10333 7293 10367 7327
rect 12173 7293 12207 7327
rect 13829 7293 13863 7327
rect 14648 7293 14682 7327
rect 16037 7293 16071 7327
rect 2697 7225 2731 7259
rect 8944 7225 8978 7259
rect 10600 7225 10634 7259
rect 1777 7157 1811 7191
rect 2605 7157 2639 7191
rect 5089 7157 5123 7191
rect 5457 7157 5491 7191
rect 6285 7157 6319 7191
rect 7297 7157 7331 7191
rect 11989 7157 12023 7191
rect 12817 7157 12851 7191
rect 15761 7157 15795 7191
rect 1961 6953 1995 6987
rect 3341 6953 3375 6987
rect 3433 6953 3467 6987
rect 4353 6953 4387 6987
rect 4721 6953 4755 6987
rect 4813 6953 4847 6987
rect 6745 6953 6779 6987
rect 10517 6953 10551 6987
rect 11529 6953 11563 6987
rect 15669 6953 15703 6987
rect 5632 6885 5666 6919
rect 1409 6817 1443 6851
rect 2329 6817 2363 6851
rect 2421 6817 2455 6851
rect 5365 6817 5399 6851
rect 7021 6817 7055 6851
rect 7288 6817 7322 6851
rect 8861 6817 8895 6851
rect 9045 6817 9079 6851
rect 11621 6817 11655 6851
rect 12541 6817 12575 6851
rect 13277 6817 13311 6851
rect 14197 6817 14231 6851
rect 15761 6817 15795 6851
rect 2513 6749 2547 6783
rect 3617 6749 3651 6783
rect 4905 6749 4939 6783
rect 9689 6749 9723 6783
rect 10609 6749 10643 6783
rect 10793 6749 10827 6783
rect 11713 6749 11747 6783
rect 12633 6749 12667 6783
rect 12817 6749 12851 6783
rect 14289 6749 14323 6783
rect 14473 6749 14507 6783
rect 15853 6749 15887 6783
rect 1593 6681 1627 6715
rect 8677 6681 8711 6715
rect 11161 6681 11195 6715
rect 12173 6681 12207 6715
rect 13829 6681 13863 6715
rect 2973 6613 3007 6647
rect 8401 6613 8435 6647
rect 9229 6613 9263 6647
rect 10149 6613 10183 6647
rect 13461 6613 13495 6647
rect 15301 6613 15335 6647
rect 5457 6409 5491 6443
rect 6285 6409 6319 6443
rect 8769 6409 8803 6443
rect 10057 6409 10091 6443
rect 10149 6409 10183 6443
rect 5917 6273 5951 6307
rect 6009 6273 6043 6307
rect 6469 6341 6503 6375
rect 6929 6273 6963 6307
rect 9689 6273 9723 6307
rect 1501 6205 1535 6239
rect 3157 6205 3191 6239
rect 3801 6205 3835 6239
rect 6285 6205 6319 6239
rect 6653 6205 6687 6239
rect 7196 6205 7230 6239
rect 8585 6205 8619 6239
rect 12541 6341 12575 6375
rect 10793 6273 10827 6307
rect 11713 6273 11747 6307
rect 11529 6205 11563 6239
rect 1768 6137 1802 6171
rect 4046 6137 4080 6171
rect 5825 6137 5859 6171
rect 10057 6137 10091 6171
rect 14289 6273 14323 6307
rect 12633 6205 12667 6239
rect 14556 6205 14590 6239
rect 15945 6205 15979 6239
rect 12541 6137 12575 6171
rect 12900 6137 12934 6171
rect 2881 6069 2915 6103
rect 3341 6069 3375 6103
rect 5181 6069 5215 6103
rect 8309 6069 8343 6103
rect 9137 6069 9171 6103
rect 9505 6069 9539 6103
rect 9597 6069 9631 6103
rect 10517 6069 10551 6103
rect 10609 6069 10643 6103
rect 11161 6069 11195 6103
rect 11621 6069 11655 6103
rect 14013 6069 14047 6103
rect 15669 6069 15703 6103
rect 16129 6069 16163 6103
rect 7297 5865 7331 5899
rect 10609 5865 10643 5899
rect 11069 5865 11103 5899
rect 11529 5865 11563 5899
rect 14197 5865 14231 5899
rect 15761 5865 15795 5899
rect 15853 5865 15887 5899
rect 4813 5797 4847 5831
rect 1593 5729 1627 5763
rect 2329 5729 2363 5763
rect 2596 5729 2630 5763
rect 5724 5729 5758 5763
rect 7113 5729 7147 5763
rect 8033 5729 8067 5763
rect 8677 5729 8711 5763
rect 10057 5729 10091 5763
rect 10977 5729 11011 5763
rect 13277 5797 13311 5831
rect 11877 5729 11911 5763
rect 14105 5729 14139 5763
rect 14749 5729 14783 5763
rect 4905 5661 4939 5695
rect 4997 5661 5031 5695
rect 5457 5661 5491 5695
rect 8125 5661 8159 5695
rect 8217 5661 8251 5695
rect 8953 5661 8987 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 14381 5661 14415 5695
rect 15945 5661 15979 5695
rect 13001 5593 13035 5627
rect 1777 5525 1811 5559
rect 3709 5525 3743 5559
rect 4445 5525 4479 5559
rect 6837 5525 6871 5559
rect 7665 5525 7699 5559
rect 10241 5525 10275 5559
rect 13737 5525 13771 5559
rect 15393 5525 15427 5559
rect 1685 5321 1719 5355
rect 5641 5321 5675 5355
rect 6837 5321 6871 5355
rect 11713 5321 11747 5355
rect 14105 5321 14139 5355
rect 2329 5185 2363 5219
rect 3249 5185 3283 5219
rect 4261 5185 4295 5219
rect 7389 5185 7423 5219
rect 7849 5185 7883 5219
rect 10333 5185 10367 5219
rect 13737 5185 13771 5219
rect 2053 5117 2087 5151
rect 3065 5117 3099 5151
rect 3709 5117 3743 5151
rect 5917 5117 5951 5151
rect 7205 5117 7239 5151
rect 9505 5117 9539 5151
rect 12173 5117 12207 5151
rect 12449 5117 12483 5151
rect 13553 5117 13587 5151
rect 14105 5117 14139 5151
rect 14197 5117 14231 5151
rect 14464 5117 14498 5151
rect 15853 5117 15887 5151
rect 3157 5049 3191 5083
rect 4528 5049 4562 5083
rect 6193 5049 6227 5083
rect 7297 5049 7331 5083
rect 8116 5049 8150 5083
rect 9781 5049 9815 5083
rect 10600 5049 10634 5083
rect 12725 5049 12759 5083
rect 2145 4981 2179 5015
rect 2697 4981 2731 5015
rect 3893 4981 3927 5015
rect 9229 4981 9263 5015
rect 11989 4981 12023 5015
rect 13185 4981 13219 5015
rect 13645 4981 13679 5015
rect 15577 4981 15611 5015
rect 16037 4981 16071 5015
rect 3065 4777 3099 4811
rect 6469 4777 6503 4811
rect 8953 4777 8987 4811
rect 13093 4777 13127 4811
rect 13369 4777 13403 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15669 4777 15703 4811
rect 15761 4777 15795 4811
rect 1952 4709 1986 4743
rect 6101 4709 6135 4743
rect 9045 4709 9079 4743
rect 9934 4709 9968 4743
rect 1685 4641 1719 4675
rect 3341 4641 3375 4675
rect 4344 4641 4378 4675
rect 5825 4641 5859 4675
rect 6469 4641 6503 4675
rect 6561 4641 6595 4675
rect 6828 4641 6862 4675
rect 8401 4641 8435 4675
rect 9689 4641 9723 4675
rect 11529 4641 11563 4675
rect 11980 4641 12014 4675
rect 13553 4641 13587 4675
rect 14657 4641 14691 4675
rect 4077 4573 4111 4607
rect 9229 4573 9263 4607
rect 11713 4573 11747 4607
rect 14105 4573 14139 4607
rect 14289 4573 14323 4607
rect 15853 4573 15887 4607
rect 8217 4505 8251 4539
rect 3525 4437 3559 4471
rect 5457 4437 5491 4471
rect 7941 4437 7975 4471
rect 8585 4437 8619 4471
rect 11069 4437 11103 4471
rect 11345 4437 11379 4471
rect 14841 4437 14875 4471
rect 15301 4437 15335 4471
rect 3617 4233 3651 4267
rect 2329 4097 2363 4131
rect 3341 4097 3375 4131
rect 2145 3961 2179 3995
rect 3157 3961 3191 3995
rect 10609 4165 10643 4199
rect 4353 4097 4387 4131
rect 6377 4097 6411 4131
rect 7757 4097 7791 4131
rect 8861 4097 8895 4131
rect 11437 4097 11471 4131
rect 11897 4097 11931 4131
rect 13001 4097 13035 4131
rect 13921 4097 13955 4131
rect 14105 4097 14139 4131
rect 15025 4097 15059 4131
rect 15945 4097 15979 4131
rect 16037 4097 16071 4131
rect 4813 4029 4847 4063
rect 6101 4029 6135 4063
rect 8585 4029 8619 4063
rect 9229 4029 9263 4063
rect 11253 4029 11287 4063
rect 14841 4029 14875 4063
rect 14933 4029 14967 4063
rect 15853 4029 15887 4063
rect 4261 3961 4295 3995
rect 5089 3961 5123 3995
rect 6193 3961 6227 3995
rect 9474 3961 9508 3995
rect 12817 3961 12851 3995
rect 1777 3893 1811 3927
rect 2237 3893 2271 3927
rect 2789 3893 2823 3927
rect 3249 3893 3283 3927
rect 3617 3893 3651 3927
rect 3801 3893 3835 3927
rect 4169 3893 4203 3927
rect 5733 3893 5767 3927
rect 7205 3893 7239 3927
rect 7573 3893 7607 3927
rect 7665 3893 7699 3927
rect 8217 3893 8251 3927
rect 8677 3893 8711 3927
rect 10885 3893 10919 3927
rect 11345 3893 11379 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 13461 3893 13495 3927
rect 13829 3893 13863 3927
rect 14473 3893 14507 3927
rect 15485 3893 15519 3927
rect 2145 3689 2179 3723
rect 2789 3689 2823 3723
rect 3249 3689 3283 3723
rect 4905 3689 4939 3723
rect 5917 3689 5951 3723
rect 6561 3689 6595 3723
rect 6929 3689 6963 3723
rect 7573 3689 7607 3723
rect 9045 3689 9079 3723
rect 10609 3689 10643 3723
rect 10977 3689 11011 3723
rect 12633 3689 12667 3723
rect 14565 3689 14599 3723
rect 15669 3689 15703 3723
rect 15761 3689 15795 3723
rect 7941 3621 7975 3655
rect 8033 3621 8067 3655
rect 12541 3621 12575 3655
rect 13452 3621 13486 3655
rect 2237 3553 2271 3587
rect 3157 3553 3191 3587
rect 6009 3553 6043 3587
rect 7021 3553 7055 3587
rect 8953 3553 8987 3587
rect 9689 3553 9723 3587
rect 9965 3553 9999 3587
rect 11621 3553 11655 3587
rect 2421 3485 2455 3519
rect 3341 3485 3375 3519
rect 4077 3485 4111 3519
rect 4997 3485 5031 3519
rect 5181 3485 5215 3519
rect 6193 3485 6227 3519
rect 7205 3485 7239 3519
rect 8125 3485 8159 3519
rect 9229 3485 9263 3519
rect 11069 3485 11103 3519
rect 11253 3485 11287 3519
rect 12725 3485 12759 3519
rect 13185 3485 13219 3519
rect 15853 3485 15887 3519
rect 1777 3349 1811 3383
rect 4537 3349 4571 3383
rect 5549 3349 5583 3383
rect 8585 3349 8619 3383
rect 11805 3349 11839 3383
rect 12173 3349 12207 3383
rect 15301 3349 15335 3383
rect 2789 3145 2823 3179
rect 4169 3145 4203 3179
rect 7113 3145 7147 3179
rect 8309 3145 8343 3179
rect 11713 3145 11747 3179
rect 13829 3145 13863 3179
rect 6377 3077 6411 3111
rect 9321 3077 9355 3111
rect 14105 3077 14139 3111
rect 1409 3009 1443 3043
rect 3801 3009 3835 3043
rect 4813 3009 4847 3043
rect 5733 3009 5767 3043
rect 7757 3009 7791 3043
rect 8953 3009 8987 3043
rect 9965 3009 9999 3043
rect 14565 3009 14599 3043
rect 14657 3009 14691 3043
rect 15393 3009 15427 3043
rect 3525 2941 3559 2975
rect 3617 2941 3651 2975
rect 5641 2941 5675 2975
rect 6193 2941 6227 2975
rect 8677 2941 8711 2975
rect 9689 2941 9723 2975
rect 10333 2941 10367 2975
rect 10600 2941 10634 2975
rect 12449 2941 12483 2975
rect 12705 2941 12739 2975
rect 14473 2941 14507 2975
rect 15117 2941 15151 2975
rect 15853 2941 15887 2975
rect 1654 2873 1688 2907
rect 4629 2873 4663 2907
rect 5549 2873 5583 2907
rect 7573 2873 7607 2907
rect 16129 2873 16163 2907
rect 3157 2805 3191 2839
rect 4537 2805 4571 2839
rect 5181 2805 5215 2839
rect 7481 2805 7515 2839
rect 8769 2805 8803 2839
rect 9781 2805 9815 2839
rect 3341 2601 3375 2635
rect 4997 2601 5031 2635
rect 5457 2601 5491 2635
rect 7021 2601 7055 2635
rect 7389 2601 7423 2635
rect 8677 2601 8711 2635
rect 9045 2601 9079 2635
rect 9137 2601 9171 2635
rect 10425 2601 10459 2635
rect 10885 2601 10919 2635
rect 11437 2601 11471 2635
rect 11897 2601 11931 2635
rect 15301 2601 15335 2635
rect 5365 2533 5399 2567
rect 7481 2533 7515 2567
rect 10793 2533 10827 2567
rect 11805 2533 11839 2567
rect 15761 2533 15795 2567
rect 1685 2465 1719 2499
rect 2237 2465 2271 2499
rect 3433 2465 3467 2499
rect 4261 2465 4295 2499
rect 6101 2465 6135 2499
rect 8033 2465 8067 2499
rect 9781 2465 9815 2499
rect 12633 2465 12667 2499
rect 13461 2465 13495 2499
rect 13921 2465 13955 2499
rect 14013 2465 14047 2499
rect 14841 2465 14875 2499
rect 15301 2465 15335 2499
rect 15485 2465 15519 2499
rect 2513 2397 2547 2431
rect 3617 2397 3651 2431
rect 4537 2397 4571 2431
rect 5549 2397 5583 2431
rect 6377 2397 6411 2431
rect 7573 2397 7607 2431
rect 9229 2397 9263 2431
rect 10977 2397 11011 2431
rect 12081 2397 12115 2431
rect 12817 2397 12851 2431
rect 14289 2397 14323 2431
rect 13921 2329 13955 2363
rect 1869 2261 1903 2295
rect 2973 2261 3007 2295
rect 8217 2261 8251 2295
rect 9965 2261 9999 2295
rect 13645 2261 13679 2295
rect 15025 2261 15059 2295
<< metal1 >>
rect 4062 15172 4068 15224
rect 4120 15212 4126 15224
rect 8938 15212 8944 15224
rect 4120 15184 8944 15212
rect 4120 15172 4126 15184
rect 8938 15172 8944 15184
rect 8996 15172 9002 15224
rect 9306 15172 9312 15224
rect 9364 15212 9370 15224
rect 14918 15212 14924 15224
rect 9364 15184 14924 15212
rect 9364 15172 9370 15184
rect 14918 15172 14924 15184
rect 14976 15172 14982 15224
rect 1104 14714 16836 14736
rect 1104 14662 6246 14714
rect 6298 14662 6310 14714
rect 6362 14662 6374 14714
rect 6426 14662 6438 14714
rect 6490 14662 11510 14714
rect 11562 14662 11574 14714
rect 11626 14662 11638 14714
rect 11690 14662 11702 14714
rect 11754 14662 16836 14714
rect 1104 14640 16836 14662
rect 8938 14600 8944 14612
rect 8899 14572 8944 14600
rect 8938 14560 8944 14572
rect 8996 14600 9002 14612
rect 10318 14600 10324 14612
rect 8996 14572 10324 14600
rect 8996 14560 9002 14572
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 8021 14535 8079 14541
rect 8021 14501 8033 14535
rect 8067 14532 8079 14535
rect 11054 14532 11060 14544
rect 8067 14504 11060 14532
rect 8067 14501 8079 14504
rect 8021 14495 8079 14501
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6638 14464 6644 14476
rect 6227 14436 6644 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14464 7987 14467
rect 8754 14464 8760 14476
rect 7975 14436 8760 14464
rect 7975 14433 7987 14436
rect 7929 14427 7987 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 9033 14467 9091 14473
rect 9033 14433 9045 14467
rect 9079 14464 9091 14467
rect 10410 14464 10416 14476
rect 9079 14436 10416 14464
rect 9079 14433 9091 14436
rect 9033 14427 9091 14433
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 10744 14436 15945 14464
rect 10744 14424 10750 14436
rect 15933 14433 15945 14436
rect 15979 14433 15991 14467
rect 15933 14427 15991 14433
rect 6086 14356 6092 14408
rect 6144 14396 6150 14408
rect 6273 14399 6331 14405
rect 6273 14396 6285 14399
rect 6144 14368 6285 14396
rect 6144 14356 6150 14368
rect 6273 14365 6285 14368
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14396 6515 14399
rect 7098 14396 7104 14408
rect 6503 14368 7104 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 8110 14396 8116 14408
rect 8071 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 9214 14396 9220 14408
rect 9175 14368 9220 14396
rect 9214 14356 9220 14368
rect 9272 14356 9278 14408
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 5534 14260 5540 14272
rect 4120 14232 5540 14260
rect 4120 14220 4126 14232
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5813 14263 5871 14269
rect 5813 14229 5825 14263
rect 5859 14260 5871 14263
rect 6178 14260 6184 14272
rect 5859 14232 6184 14260
rect 5859 14229 5871 14232
rect 5813 14223 5871 14229
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 7561 14263 7619 14269
rect 7561 14229 7573 14263
rect 7607 14260 7619 14263
rect 7650 14260 7656 14272
rect 7607 14232 7656 14260
rect 7607 14229 7619 14232
rect 7561 14223 7619 14229
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 8570 14260 8576 14272
rect 8531 14232 8576 14260
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 16117 14263 16175 14269
rect 16117 14229 16129 14263
rect 16163 14260 16175 14263
rect 16298 14260 16304 14272
rect 16163 14232 16304 14260
rect 16163 14229 16175 14232
rect 16117 14223 16175 14229
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 1104 14170 16836 14192
rect 1104 14118 3614 14170
rect 3666 14118 3678 14170
rect 3730 14118 3742 14170
rect 3794 14118 3806 14170
rect 3858 14118 8878 14170
rect 8930 14118 8942 14170
rect 8994 14118 9006 14170
rect 9058 14118 9070 14170
rect 9122 14118 14142 14170
rect 14194 14118 14206 14170
rect 14258 14118 14270 14170
rect 14322 14118 14334 14170
rect 14386 14118 16836 14170
rect 1104 14096 16836 14118
rect 9490 14056 9496 14068
rect 2700 14028 9496 14056
rect 2700 13929 2728 14028
rect 9490 14016 9496 14028
rect 9548 14056 9554 14068
rect 14826 14056 14832 14068
rect 9548 14028 14832 14056
rect 9548 14016 9554 14028
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 5534 13948 5540 14000
rect 5592 13988 5598 14000
rect 13538 13988 13544 14000
rect 5592 13960 13544 13988
rect 5592 13948 5598 13960
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2869 13923 2927 13929
rect 2869 13889 2881 13923
rect 2915 13920 2927 13923
rect 3142 13920 3148 13932
rect 2915 13892 3148 13920
rect 2915 13889 2927 13892
rect 2869 13883 2927 13889
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5132 13892 5273 13920
rect 5132 13880 5138 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 6178 13920 6184 13932
rect 6139 13892 6184 13920
rect 5261 13883 5319 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13920 6423 13923
rect 6914 13920 6920 13932
rect 6411 13892 6920 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 7650 13920 7656 13932
rect 7611 13892 7656 13920
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 7834 13920 7840 13932
rect 7795 13892 7840 13920
rect 7834 13880 7840 13892
rect 7892 13920 7898 13932
rect 9214 13920 9220 13932
rect 7892 13892 9220 13920
rect 7892 13880 7898 13892
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 9916 13892 10701 13920
rect 9916 13880 9922 13892
rect 10689 13889 10701 13892
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 15252 13892 15669 13920
rect 15252 13880 15258 13892
rect 15657 13889 15669 13892
rect 15703 13889 15715 13923
rect 15657 13883 15715 13889
rect 3970 13812 3976 13864
rect 4028 13852 4034 13864
rect 8386 13852 8392 13864
rect 4028 13824 8392 13852
rect 4028 13812 4034 13824
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 9306 13852 9312 13864
rect 9171 13824 9312 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 10594 13852 10600 13864
rect 10555 13824 10600 13852
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 15562 13852 15568 13864
rect 15523 13824 15568 13852
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 4890 13744 4896 13796
rect 4948 13784 4954 13796
rect 5077 13787 5135 13793
rect 5077 13784 5089 13787
rect 4948 13756 5089 13784
rect 4948 13744 4954 13756
rect 5077 13753 5089 13756
rect 5123 13784 5135 13787
rect 7374 13784 7380 13796
rect 5123 13756 7380 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 9033 13787 9091 13793
rect 9033 13753 9045 13787
rect 9079 13784 9091 13787
rect 9674 13784 9680 13796
rect 9079 13756 9680 13784
rect 9079 13753 9091 13756
rect 9033 13747 9091 13753
rect 9674 13744 9680 13756
rect 9732 13744 9738 13796
rect 9784 13756 12480 13784
rect 2222 13716 2228 13728
rect 2183 13688 2228 13716
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 2593 13719 2651 13725
rect 2593 13685 2605 13719
rect 2639 13716 2651 13719
rect 3326 13716 3332 13728
rect 2639 13688 3332 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 3326 13676 3332 13688
rect 3384 13676 3390 13728
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4709 13719 4767 13725
rect 4709 13716 4721 13719
rect 4580 13688 4721 13716
rect 4580 13676 4586 13688
rect 4709 13685 4721 13688
rect 4755 13685 4767 13719
rect 5166 13716 5172 13728
rect 5127 13688 5172 13716
rect 4709 13679 4767 13685
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 6089 13719 6147 13725
rect 6089 13685 6101 13719
rect 6135 13716 6147 13719
rect 7006 13716 7012 13728
rect 6135 13688 7012 13716
rect 6135 13685 6147 13688
rect 6089 13679 6147 13685
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 7190 13716 7196 13728
rect 7151 13688 7196 13716
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7561 13719 7619 13725
rect 7561 13685 7573 13719
rect 7607 13716 7619 13719
rect 7742 13716 7748 13728
rect 7607 13688 7748 13716
rect 7607 13685 7619 13688
rect 7561 13679 7619 13685
rect 7742 13676 7748 13688
rect 7800 13676 7806 13728
rect 8662 13716 8668 13728
rect 8623 13688 8668 13716
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 9784 13716 9812 13756
rect 10134 13716 10140 13728
rect 8904 13688 9812 13716
rect 10095 13688 10140 13716
rect 8904 13676 8910 13688
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10502 13716 10508 13728
rect 10463 13688 10508 13716
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 12452 13716 12480 13756
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 13354 13784 13360 13796
rect 12584 13756 13360 13784
rect 12584 13744 12590 13756
rect 13354 13744 13360 13756
rect 13412 13744 13418 13796
rect 14918 13716 14924 13728
rect 12452 13688 14924 13716
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 15102 13716 15108 13728
rect 15063 13688 15108 13716
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 15470 13716 15476 13728
rect 15431 13688 15476 13716
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 15712 13688 16129 13716
rect 15712 13676 15718 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 1104 13626 16836 13648
rect 1104 13574 6246 13626
rect 6298 13574 6310 13626
rect 6362 13574 6374 13626
rect 6426 13574 6438 13626
rect 6490 13574 11510 13626
rect 11562 13574 11574 13626
rect 11626 13574 11638 13626
rect 11690 13574 11702 13626
rect 11754 13574 16836 13626
rect 1104 13552 16836 13574
rect 4893 13515 4951 13521
rect 4893 13481 4905 13515
rect 4939 13512 4951 13515
rect 8573 13515 8631 13521
rect 4939 13484 8064 13512
rect 4939 13481 4951 13484
rect 4893 13475 4951 13481
rect 8036 13456 8064 13484
rect 8573 13481 8585 13515
rect 8619 13512 8631 13515
rect 8662 13512 8668 13524
rect 8619 13484 8668 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 10134 13512 10140 13524
rect 10095 13484 10140 13512
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10244 13484 15056 13512
rect 5813 13447 5871 13453
rect 5813 13413 5825 13447
rect 5859 13413 5871 13447
rect 5813 13407 5871 13413
rect 5905 13447 5963 13453
rect 5905 13413 5917 13447
rect 5951 13444 5963 13447
rect 7469 13447 7527 13453
rect 5951 13416 6040 13444
rect 5951 13413 5963 13416
rect 5905 13407 5963 13413
rect 2498 13376 2504 13388
rect 2459 13348 2504 13376
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13376 4859 13379
rect 5626 13376 5632 13388
rect 4847 13348 5632 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 5828 13376 5856 13407
rect 5736 13348 5856 13376
rect 6012 13376 6040 13416
rect 7469 13413 7481 13447
rect 7515 13444 7527 13447
rect 7558 13444 7564 13456
rect 7515 13416 7564 13444
rect 7515 13413 7527 13416
rect 7469 13407 7527 13413
rect 7558 13404 7564 13416
rect 7616 13404 7622 13456
rect 8018 13404 8024 13456
rect 8076 13444 8082 13456
rect 10244 13444 10272 13484
rect 15028 13456 15056 13484
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15565 13515 15623 13521
rect 15565 13512 15577 13515
rect 15528 13484 15577 13512
rect 15528 13472 15534 13484
rect 15565 13481 15577 13484
rect 15611 13481 15623 13515
rect 15565 13475 15623 13481
rect 8076 13416 10272 13444
rect 11701 13447 11759 13453
rect 8076 13404 8082 13416
rect 11701 13413 11713 13447
rect 11747 13444 11759 13447
rect 12526 13444 12532 13456
rect 11747 13416 12532 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 12713 13447 12771 13453
rect 12713 13444 12725 13447
rect 12636 13416 12725 13444
rect 6012 13348 6224 13376
rect 2590 13308 2596 13320
rect 2551 13280 2596 13308
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 5074 13308 5080 13320
rect 2740 13280 2785 13308
rect 5035 13280 5080 13308
rect 2740 13268 2746 13280
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 5736 13240 5764 13348
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 6052 13280 6097 13308
rect 6052 13268 6058 13280
rect 5810 13240 5816 13252
rect 5736 13212 5816 13240
rect 5810 13200 5816 13212
rect 5868 13200 5874 13252
rect 5902 13200 5908 13252
rect 5960 13240 5966 13252
rect 6196 13240 6224 13348
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 7377 13379 7435 13385
rect 7377 13376 7389 13379
rect 6880 13348 7389 13376
rect 6880 13336 6886 13348
rect 7377 13345 7389 13348
rect 7423 13345 7435 13379
rect 7834 13376 7840 13388
rect 7377 13339 7435 13345
rect 7576 13348 7840 13376
rect 7576 13317 7604 13348
rect 7834 13336 7840 13348
rect 7892 13376 7898 13388
rect 8202 13376 8208 13388
rect 7892 13348 8208 13376
rect 7892 13336 7898 13348
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 8665 13379 8723 13385
rect 8665 13376 8677 13379
rect 8628 13348 8677 13376
rect 8628 13336 8634 13348
rect 8665 13345 8677 13348
rect 8711 13345 8723 13379
rect 8665 13339 8723 13345
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 8904 13348 10057 13376
rect 8904 13336 8910 13348
rect 10045 13345 10057 13348
rect 10091 13376 10103 13379
rect 10686 13376 10692 13388
rect 10091 13348 10692 13376
rect 10091 13345 10103 13348
rect 10045 13339 10103 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 11882 13336 11888 13388
rect 11940 13376 11946 13388
rect 12636 13376 12664 13416
rect 12713 13413 12725 13416
rect 12759 13413 12771 13447
rect 12713 13407 12771 13413
rect 12820 13416 14412 13444
rect 12820 13376 12848 13416
rect 11940 13348 12664 13376
rect 12728 13348 12848 13376
rect 13357 13379 13415 13385
rect 11940 13336 11946 13348
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 7708 13280 8769 13308
rect 7708 13268 7714 13280
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10870 13308 10876 13320
rect 10367 13280 10876 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 11974 13308 11980 13320
rect 11935 13280 11980 13308
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12728 13240 12756 13348
rect 13357 13345 13369 13379
rect 13403 13376 13415 13379
rect 13446 13376 13452 13388
rect 13403 13348 13452 13376
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 13630 13385 13636 13388
rect 13624 13339 13636 13385
rect 13688 13376 13694 13388
rect 13688 13348 13724 13376
rect 13630 13336 13636 13339
rect 13688 13336 13694 13348
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 5960 13212 12756 13240
rect 12820 13240 12848 13271
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 14384 13308 14412 13416
rect 15010 13404 15016 13456
rect 15068 13444 15074 13456
rect 16025 13447 16083 13453
rect 16025 13444 16037 13447
rect 15068 13416 16037 13444
rect 15068 13404 15074 13416
rect 16025 13413 16037 13416
rect 16071 13413 16083 13447
rect 16025 13407 16083 13413
rect 15930 13376 15936 13388
rect 15891 13348 15936 13376
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 16390 13376 16396 13388
rect 16040 13348 16396 13376
rect 16040 13308 16068 13348
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 12952 13280 12997 13308
rect 14384 13280 16068 13308
rect 16117 13311 16175 13317
rect 12952 13268 12958 13280
rect 16117 13277 16129 13311
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 13078 13240 13084 13252
rect 12820 13212 13084 13240
rect 5960 13200 5966 13212
rect 13078 13200 13084 13212
rect 13136 13240 13142 13252
rect 13136 13212 13308 13240
rect 13136 13200 13142 13212
rect 2130 13172 2136 13184
rect 2091 13144 2136 13172
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 4430 13172 4436 13184
rect 4391 13144 4436 13172
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 5166 13132 5172 13184
rect 5224 13172 5230 13184
rect 5445 13175 5503 13181
rect 5445 13172 5457 13175
rect 5224 13144 5457 13172
rect 5224 13132 5230 13144
rect 5445 13141 5457 13144
rect 5491 13141 5503 13175
rect 5445 13135 5503 13141
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13172 7067 13175
rect 7282 13172 7288 13184
rect 7055 13144 7288 13172
rect 7055 13141 7067 13144
rect 7009 13135 7067 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8205 13175 8263 13181
rect 8205 13141 8217 13175
rect 8251 13172 8263 13175
rect 8294 13172 8300 13184
rect 8251 13144 8300 13172
rect 8251 13141 8263 13144
rect 8205 13135 8263 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 9490 13172 9496 13184
rect 9272 13144 9496 13172
rect 9272 13132 9278 13144
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 9766 13172 9772 13184
rect 9723 13144 9772 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 12250 13172 12256 13184
rect 11379 13144 12256 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 13170 13172 13176 13184
rect 12391 13144 13176 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 13280 13172 13308 13212
rect 16022 13200 16028 13252
rect 16080 13240 16086 13252
rect 16132 13240 16160 13271
rect 16080 13212 16160 13240
rect 16080 13200 16086 13212
rect 14458 13172 14464 13184
rect 13280 13144 14464 13172
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 14737 13175 14795 13181
rect 14737 13141 14749 13175
rect 14783 13172 14795 13175
rect 14826 13172 14832 13184
rect 14783 13144 14832 13172
rect 14783 13141 14795 13144
rect 14737 13135 14795 13141
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 1104 13082 16836 13104
rect 1104 13030 3614 13082
rect 3666 13030 3678 13082
rect 3730 13030 3742 13082
rect 3794 13030 3806 13082
rect 3858 13030 8878 13082
rect 8930 13030 8942 13082
rect 8994 13030 9006 13082
rect 9058 13030 9070 13082
rect 9122 13030 14142 13082
rect 14194 13030 14206 13082
rect 14258 13030 14270 13082
rect 14322 13030 14334 13082
rect 14386 13030 16836 13082
rect 1104 13008 16836 13030
rect 3789 12971 3847 12977
rect 3789 12937 3801 12971
rect 3835 12968 3847 12971
rect 4706 12968 4712 12980
rect 3835 12940 4712 12968
rect 3835 12937 3847 12940
rect 3789 12931 3847 12937
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 13446 12968 13452 12980
rect 6880 12940 10088 12968
rect 6880 12928 6886 12940
rect 4154 12900 4160 12912
rect 3436 12872 4160 12900
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 2682 12832 2688 12844
rect 2455 12804 2688 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 3436 12841 3464 12872
rect 4154 12860 4160 12872
rect 4212 12860 4218 12912
rect 5350 12860 5356 12912
rect 5408 12900 5414 12912
rect 5408 12872 9444 12900
rect 5408 12860 5414 12872
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3970 12792 3976 12844
rect 4028 12832 4034 12844
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4028 12804 4353 12832
rect 4028 12792 4034 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 5442 12832 5448 12844
rect 5403 12804 5448 12832
rect 4341 12795 4399 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 7190 12792 7196 12844
rect 7248 12832 7254 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7248 12804 7389 12832
rect 7248 12792 7254 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 7650 12832 7656 12844
rect 7607 12804 7656 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 8478 12832 8484 12844
rect 8439 12804 8484 12832
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 2133 12767 2191 12773
rect 2133 12733 2145 12767
rect 2179 12764 2191 12767
rect 2222 12764 2228 12776
rect 2179 12736 2228 12764
rect 2179 12733 2191 12736
rect 2133 12727 2191 12733
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 5166 12764 5172 12776
rect 5127 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 7282 12764 7288 12776
rect 7243 12736 7288 12764
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7668 12764 7696 12792
rect 7926 12764 7932 12776
rect 7668 12736 7932 12764
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8294 12764 8300 12776
rect 8255 12736 8300 12764
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 9416 12773 9444 12872
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9858 12832 9864 12844
rect 9631 12804 9864 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 10060 12832 10088 12940
rect 12452 12940 13452 12968
rect 11882 12832 11888 12844
rect 10060 12804 10180 12832
rect 11843 12804 11888 12832
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12733 9459 12767
rect 9401 12727 9459 12733
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 10008 12736 10057 12764
rect 10008 12724 10014 12736
rect 10045 12733 10057 12736
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 3145 12699 3203 12705
rect 3145 12665 3157 12699
rect 3191 12696 3203 12699
rect 3418 12696 3424 12708
rect 3191 12668 3424 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 4157 12699 4215 12705
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 4203 12668 4844 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 1762 12628 1768 12640
rect 1723 12600 1768 12628
rect 1762 12588 1768 12600
rect 1820 12588 1826 12640
rect 2222 12628 2228 12640
rect 2183 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12588 2286 12640
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3237 12631 3295 12637
rect 2832 12600 2877 12628
rect 2832 12588 2838 12600
rect 3237 12597 3249 12631
rect 3283 12628 3295 12631
rect 4062 12628 4068 12640
rect 3283 12600 4068 12628
rect 3283 12597 3295 12600
rect 3237 12591 3295 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4246 12628 4252 12640
rect 4207 12600 4252 12628
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4816 12637 4844 12668
rect 6932 12668 8401 12696
rect 4801 12631 4859 12637
rect 4801 12597 4813 12631
rect 4847 12597 4859 12631
rect 4801 12591 4859 12597
rect 5258 12588 5264 12640
rect 5316 12628 5322 12640
rect 6932 12637 6960 12668
rect 8389 12665 8401 12668
rect 8435 12665 8447 12699
rect 9490 12696 9496 12708
rect 9451 12668 9496 12696
rect 8389 12659 8447 12665
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 10152 12696 10180 12804
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 12452 12841 12480 12940
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13630 12860 13636 12912
rect 13688 12900 13694 12912
rect 13817 12903 13875 12909
rect 13817 12900 13829 12903
rect 13688 12872 13829 12900
rect 13688 12860 13694 12872
rect 13817 12869 13829 12872
rect 13863 12869 13875 12903
rect 13817 12863 13875 12869
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 10312 12767 10370 12773
rect 10312 12733 10324 12767
rect 10358 12764 10370 12767
rect 12066 12764 12072 12776
rect 10358 12736 12072 12764
rect 10358 12733 10370 12736
rect 10312 12727 10370 12733
rect 12066 12724 12072 12736
rect 12124 12764 12130 12776
rect 12124 12736 12848 12764
rect 12124 12724 12130 12736
rect 12820 12708 12848 12736
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 13504 12736 14105 12764
rect 13504 12724 13510 12736
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 15933 12767 15991 12773
rect 15933 12764 15945 12767
rect 14093 12727 14151 12733
rect 14200 12736 15945 12764
rect 10410 12696 10416 12708
rect 10152 12668 10416 12696
rect 10410 12656 10416 12668
rect 10468 12656 10474 12708
rect 11256 12668 11560 12696
rect 6917 12631 6975 12637
rect 5316 12600 5361 12628
rect 5316 12588 5322 12600
rect 6917 12597 6929 12631
rect 6963 12597 6975 12631
rect 7926 12628 7932 12640
rect 7887 12600 7932 12628
rect 6917 12591 6975 12597
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 9030 12628 9036 12640
rect 8991 12600 9036 12628
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 11256 12628 11284 12668
rect 9180 12600 11284 12628
rect 9180 12588 9186 12600
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11425 12631 11483 12637
rect 11425 12628 11437 12631
rect 11388 12600 11437 12628
rect 11388 12588 11394 12600
rect 11425 12597 11437 12600
rect 11471 12597 11483 12631
rect 11532 12628 11560 12668
rect 11974 12656 11980 12708
rect 12032 12696 12038 12708
rect 12682 12699 12740 12705
rect 12682 12696 12694 12699
rect 12032 12668 12694 12696
rect 12032 12656 12038 12668
rect 12682 12665 12694 12668
rect 12728 12665 12740 12699
rect 12682 12659 12740 12665
rect 12802 12656 12808 12708
rect 12860 12656 12866 12708
rect 14200 12628 14228 12736
rect 15933 12733 15945 12736
rect 15979 12733 15991 12767
rect 15933 12727 15991 12733
rect 14360 12699 14418 12705
rect 14360 12665 14372 12699
rect 14406 12696 14418 12699
rect 15194 12696 15200 12708
rect 14406 12668 15200 12696
rect 14406 12665 14418 12668
rect 14360 12659 14418 12665
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 11532 12600 14228 12628
rect 11425 12591 11483 12597
rect 14734 12588 14740 12640
rect 14792 12628 14798 12640
rect 15473 12631 15531 12637
rect 15473 12628 15485 12631
rect 14792 12600 15485 12628
rect 14792 12588 14798 12600
rect 15473 12597 15485 12600
rect 15519 12597 15531 12631
rect 16114 12628 16120 12640
rect 16075 12600 16120 12628
rect 15473 12591 15531 12597
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 1104 12538 16836 12560
rect 1104 12486 6246 12538
rect 6298 12486 6310 12538
rect 6362 12486 6374 12538
rect 6426 12486 6438 12538
rect 6490 12486 11510 12538
rect 11562 12486 11574 12538
rect 11626 12486 11638 12538
rect 11690 12486 11702 12538
rect 11754 12486 16836 12538
rect 1104 12464 16836 12486
rect 1762 12384 1768 12436
rect 1820 12424 1826 12436
rect 1949 12427 2007 12433
rect 1949 12424 1961 12427
rect 1820 12396 1961 12424
rect 1820 12384 1826 12396
rect 1949 12393 1961 12396
rect 1995 12393 2007 12427
rect 1949 12387 2007 12393
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2590 12424 2596 12436
rect 2551 12396 2596 12424
rect 2590 12384 2596 12396
rect 2648 12384 2654 12436
rect 5810 12424 5816 12436
rect 5771 12396 5816 12424
rect 5810 12384 5816 12396
rect 5868 12384 5874 12436
rect 7834 12384 7840 12436
rect 7892 12424 7898 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7892 12396 7941 12424
rect 7892 12384 7898 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 7929 12387 7987 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10502 12384 10508 12436
rect 10560 12384 10566 12436
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 11974 12424 11980 12436
rect 11931 12396 11980 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 14458 12424 14464 12436
rect 12308 12396 14464 12424
rect 12308 12384 12314 12396
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 15473 12427 15531 12433
rect 15473 12393 15485 12427
rect 15519 12424 15531 12427
rect 15562 12424 15568 12436
rect 15519 12396 15568 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 4614 12316 4620 12368
rect 4672 12356 4678 12368
rect 10520 12356 10548 12384
rect 4672 12328 10548 12356
rect 10772 12359 10830 12365
rect 4672 12316 4678 12328
rect 10772 12325 10784 12359
rect 10818 12356 10830 12359
rect 11330 12356 11336 12368
rect 10818 12328 11336 12356
rect 10818 12325 10830 12328
rect 10772 12319 10830 12325
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 12526 12316 12532 12368
rect 12584 12356 12590 12368
rect 14642 12356 14648 12368
rect 12584 12328 14648 12356
rect 12584 12316 12590 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 15212 12328 16068 12356
rect 2958 12288 2964 12300
rect 2919 12260 2964 12288
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 4332 12291 4390 12297
rect 3108 12260 3153 12288
rect 3108 12248 3114 12260
rect 4332 12257 4344 12291
rect 4378 12288 4390 12291
rect 5810 12288 5816 12300
rect 4378 12260 5816 12288
rect 4378 12257 4390 12260
rect 4332 12251 4390 12257
rect 5810 12248 5816 12260
rect 5868 12288 5874 12300
rect 5994 12288 6000 12300
rect 5868 12260 6000 12288
rect 5868 12248 5874 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6816 12291 6874 12297
rect 6816 12257 6828 12291
rect 6862 12288 6874 12291
rect 8202 12288 8208 12300
rect 6862 12260 8208 12288
rect 6862 12257 6874 12260
rect 6816 12251 6874 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12288 8999 12291
rect 10318 12288 10324 12300
rect 8987 12260 10324 12288
rect 8987 12257 8999 12260
rect 8941 12251 8999 12257
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10428 12260 10517 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2866 12220 2872 12232
rect 2271 12192 2872 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 2590 12112 2596 12164
rect 2648 12152 2654 12164
rect 4080 12152 4108 12183
rect 2648 12124 4108 12152
rect 2648 12112 2654 12124
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 4080 12084 4108 12124
rect 4338 12084 4344 12096
rect 4080 12056 4344 12084
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5442 12084 5448 12096
rect 4856 12056 5448 12084
rect 4856 12044 4862 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 6178 12084 6184 12096
rect 5684 12056 6184 12084
rect 5684 12044 5690 12056
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 6564 12084 6592 12183
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 9122 12220 9128 12232
rect 7800 12192 9128 12220
rect 7800 12180 7806 12192
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12220 9275 12223
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 9263 12192 9413 12220
rect 9263 12189 9275 12192
rect 9217 12183 9275 12189
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10428 12220 10456 12260
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 12342 12288 12348 12300
rect 10505 12251 10563 12257
rect 10612 12260 12348 12288
rect 10612 12220 10640 12260
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 12618 12288 12624 12300
rect 12579 12260 12624 12288
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 13808 12291 13866 12297
rect 13808 12257 13820 12291
rect 13854 12288 13866 12291
rect 14826 12288 14832 12300
rect 13854 12260 14832 12288
rect 13854 12257 13866 12260
rect 13808 12251 13866 12257
rect 14826 12248 14832 12260
rect 14884 12288 14890 12300
rect 15212 12288 15240 12328
rect 14884 12260 15240 12288
rect 14884 12248 14890 12260
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15841 12291 15899 12297
rect 15841 12288 15853 12291
rect 15528 12260 15853 12288
rect 15528 12248 15534 12260
rect 15841 12257 15853 12260
rect 15887 12257 15899 12291
rect 15841 12251 15899 12257
rect 16040 12232 16068 12328
rect 10008 12192 10456 12220
rect 10520 12192 10640 12220
rect 10008 12180 10014 12192
rect 7558 12112 7564 12164
rect 7616 12152 7622 12164
rect 10520 12152 10548 12192
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 12492 12192 12725 12220
rect 12492 12180 12498 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 7616 12124 10548 12152
rect 12728 12152 12756 12183
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 12860 12192 12905 12220
rect 12860 12180 12866 12192
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 13504 12192 13553 12220
rect 13504 12180 13510 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 14976 12192 15945 12220
rect 14976 12180 14982 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16080 12192 16125 12220
rect 16080 12180 16086 12192
rect 13078 12152 13084 12164
rect 12728 12124 13084 12152
rect 7616 12112 7622 12124
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 6730 12084 6736 12096
rect 6564 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 9306 12084 9312 12096
rect 8619 12056 9312 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 10042 12084 10048 12096
rect 9447 12056 10048 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 10042 12044 10048 12056
rect 10100 12084 10106 12096
rect 10870 12084 10876 12096
rect 10100 12056 10876 12084
rect 10100 12044 10106 12056
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 12253 12087 12311 12093
rect 12253 12053 12265 12087
rect 12299 12084 12311 12087
rect 13906 12084 13912 12096
rect 12299 12056 13912 12084
rect 12299 12053 12311 12056
rect 12253 12047 12311 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12084 14979 12087
rect 15194 12084 15200 12096
rect 14967 12056 15200 12084
rect 14967 12053 14979 12056
rect 14921 12047 14979 12053
rect 15194 12044 15200 12056
rect 15252 12084 15258 12096
rect 15838 12084 15844 12096
rect 15252 12056 15844 12084
rect 15252 12044 15258 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 1104 11994 16836 12016
rect 1104 11942 3614 11994
rect 3666 11942 3678 11994
rect 3730 11942 3742 11994
rect 3794 11942 3806 11994
rect 3858 11942 8878 11994
rect 8930 11942 8942 11994
rect 8994 11942 9006 11994
rect 9058 11942 9070 11994
rect 9122 11942 14142 11994
rect 14194 11942 14206 11994
rect 14258 11942 14270 11994
rect 14322 11942 14334 11994
rect 14386 11942 16836 11994
rect 1104 11920 16836 11942
rect 2774 11880 2780 11892
rect 2056 11852 2780 11880
rect 2056 11812 2084 11852
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 3881 11883 3939 11889
rect 3881 11849 3893 11883
rect 3927 11880 3939 11883
rect 3970 11880 3976 11892
rect 3927 11852 3976 11880
rect 3927 11849 3939 11852
rect 3881 11843 3939 11849
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4246 11880 4252 11892
rect 4203 11852 4252 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4798 11880 4804 11892
rect 4488 11852 4804 11880
rect 4488 11840 4494 11852
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5353 11883 5411 11889
rect 5353 11880 5365 11883
rect 5316 11852 5365 11880
rect 5316 11840 5322 11852
rect 5353 11849 5365 11852
rect 5399 11849 5411 11883
rect 5353 11843 5411 11849
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 8389 11883 8447 11889
rect 5592 11852 7972 11880
rect 5592 11840 5598 11852
rect 1964 11784 2084 11812
rect 4065 11815 4123 11821
rect 1964 11753 1992 11784
rect 4065 11781 4077 11815
rect 4111 11812 4123 11815
rect 6086 11812 6092 11824
rect 4111 11784 6092 11812
rect 4111 11781 4123 11784
rect 4065 11775 4123 11781
rect 6086 11772 6092 11784
rect 6144 11772 6150 11824
rect 7944 11812 7972 11852
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 8478 11880 8484 11892
rect 8435 11852 8484 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8588 11852 9628 11880
rect 8588 11812 8616 11852
rect 7944 11784 8616 11812
rect 9600 11812 9628 11852
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 9916 11852 10057 11880
rect 9916 11840 9922 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10318 11880 10324 11892
rect 10279 11852 10324 11880
rect 10045 11843 10103 11849
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 11333 11883 11391 11889
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 11790 11880 11796 11892
rect 11379 11852 11796 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 13078 11880 13084 11892
rect 12207 11852 13084 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13412 11852 13461 11880
rect 13412 11840 13418 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13449 11843 13507 11849
rect 10594 11812 10600 11824
rect 9600 11784 10600 11812
rect 10594 11772 10600 11784
rect 10652 11812 10658 11824
rect 10962 11812 10968 11824
rect 10652 11784 10968 11812
rect 10652 11772 10658 11784
rect 10962 11772 10968 11784
rect 11020 11772 11026 11824
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 12584 11784 14044 11812
rect 12584 11772 12590 11784
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11713 2007 11747
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 1949 11707 2007 11713
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 4798 11744 4804 11756
rect 3568 11716 4568 11744
rect 4759 11716 4804 11744
rect 3568 11704 3574 11716
rect 2501 11679 2559 11685
rect 1504 11648 2452 11676
rect 1504 11549 1532 11648
rect 2424 11608 2452 11648
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 2590 11676 2596 11688
rect 2547 11648 2596 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 2590 11636 2596 11648
rect 2648 11636 2654 11688
rect 2768 11679 2826 11685
rect 2768 11645 2780 11679
rect 2814 11676 2826 11679
rect 4430 11676 4436 11688
rect 2814 11648 4436 11676
rect 2814 11645 2826 11648
rect 2768 11639 2826 11645
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 4540 11676 4568 11716
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5868 11716 5917 11744
rect 5868 11704 5874 11716
rect 5905 11713 5917 11716
rect 5951 11744 5963 11747
rect 6546 11744 6552 11756
rect 5951 11716 6552 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 6656 11716 7144 11744
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 4540 11648 5733 11676
rect 5721 11645 5733 11648
rect 5767 11676 5779 11679
rect 6656 11676 6684 11716
rect 5767 11648 6684 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6788 11648 7021 11676
rect 6788 11636 6794 11648
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7116 11676 7144 11716
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8536 11716 8800 11744
rect 8536 11704 8542 11716
rect 7276 11679 7334 11685
rect 7116 11648 7236 11676
rect 7009 11639 7067 11645
rect 4065 11611 4123 11617
rect 4065 11608 4077 11611
rect 2424 11580 4077 11608
rect 4065 11577 4077 11580
rect 4111 11577 4123 11611
rect 4065 11571 4123 11577
rect 4525 11611 4583 11617
rect 4525 11577 4537 11611
rect 4571 11608 4583 11611
rect 6822 11608 6828 11620
rect 4571 11580 6828 11608
rect 4571 11577 4583 11580
rect 4525 11571 4583 11577
rect 6822 11568 6828 11580
rect 6880 11568 6886 11620
rect 7208 11608 7236 11648
rect 7276 11645 7288 11679
rect 7322 11676 7334 11679
rect 7834 11676 7840 11688
rect 7322 11648 7840 11676
rect 7322 11645 7334 11648
rect 7276 11639 7334 11645
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 8662 11676 8668 11688
rect 8623 11648 8668 11676
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 8772 11676 8800 11716
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10873 11747 10931 11753
rect 10873 11744 10885 11747
rect 9916 11716 10885 11744
rect 9916 11704 9922 11716
rect 10873 11713 10885 11716
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11388 11716 11989 11744
rect 11388 11704 11394 11716
rect 11977 11713 11989 11716
rect 12023 11744 12035 11747
rect 12023 11716 12296 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 8921 11679 8979 11685
rect 8921 11676 8933 11679
rect 8772 11648 8933 11676
rect 8921 11645 8933 11648
rect 8967 11645 8979 11679
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 8921 11639 8979 11645
rect 9048 11648 12173 11676
rect 9048 11608 9076 11648
rect 12161 11645 12173 11648
rect 12207 11645 12219 11679
rect 12268 11676 12296 11716
rect 12802 11704 12808 11756
rect 12860 11744 12866 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12860 11716 13001 11744
rect 12860 11704 12866 11716
rect 12989 11713 13001 11716
rect 13035 11744 13047 11747
rect 13262 11744 13268 11756
rect 13035 11716 13268 11744
rect 13035 11713 13047 11716
rect 12989 11707 13047 11713
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 13906 11744 13912 11756
rect 13867 11716 13912 11744
rect 13906 11704 13912 11716
rect 13964 11704 13970 11756
rect 14016 11753 14044 11784
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15988 11716 16129 11744
rect 15988 11704 15994 11716
rect 16117 11713 16129 11716
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 12526 11676 12532 11688
rect 12268 11648 12532 11676
rect 12161 11639 12219 11645
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 13228 11648 13829 11676
rect 13228 11636 13234 11648
rect 13817 11645 13829 11648
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 7208 11580 9076 11608
rect 10689 11611 10747 11617
rect 10689 11577 10701 11611
rect 10735 11608 10747 11611
rect 11238 11608 11244 11620
rect 10735 11580 11244 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 11701 11611 11759 11617
rect 11701 11577 11713 11611
rect 11747 11608 11759 11611
rect 11747 11580 12480 11608
rect 11747 11577 11759 11580
rect 11701 11571 11759 11577
rect 1489 11543 1547 11549
rect 1489 11509 1501 11543
rect 1535 11509 1547 11543
rect 1854 11540 1860 11552
rect 1815 11512 1860 11540
rect 1489 11503 1547 11509
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 5626 11540 5632 11552
rect 4663 11512 5632 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 7558 11540 7564 11552
rect 5859 11512 7564 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 10594 11540 10600 11552
rect 8444 11512 10600 11540
rect 8444 11500 8450 11512
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 10778 11540 10784 11552
rect 10739 11512 10784 11540
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 12452 11549 12480 11580
rect 13446 11568 13452 11620
rect 13504 11608 13510 11620
rect 14476 11608 14504 11639
rect 14734 11617 14740 11620
rect 14728 11608 14740 11617
rect 13504 11580 14504 11608
rect 14695 11580 14740 11608
rect 13504 11568 13510 11580
rect 14728 11571 14740 11580
rect 14734 11568 14740 11571
rect 14792 11568 14798 11620
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11388 11512 11805 11540
rect 11388 11500 11394 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11509 12495 11543
rect 12437 11503 12495 11509
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12584 11512 12817 11540
rect 12584 11500 12590 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 12952 11512 12997 11540
rect 12952 11500 12958 11512
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15841 11543 15899 11549
rect 15841 11540 15853 11543
rect 15252 11512 15853 11540
rect 15252 11500 15258 11512
rect 15841 11509 15853 11512
rect 15887 11509 15899 11543
rect 15841 11503 15899 11509
rect 1104 11450 16836 11472
rect 1104 11398 6246 11450
rect 6298 11398 6310 11450
rect 6362 11398 6374 11450
rect 6426 11398 6438 11450
rect 6490 11398 11510 11450
rect 11562 11398 11574 11450
rect 11626 11398 11638 11450
rect 11690 11398 11702 11450
rect 11754 11398 16836 11450
rect 1104 11376 16836 11398
rect 2590 11336 2596 11348
rect 2148 11308 2596 11336
rect 1394 11228 1400 11280
rect 1452 11268 1458 11280
rect 2148 11268 2176 11308
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 4203 11308 7297 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 7285 11299 7343 11305
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9306 11336 9312 11348
rect 9079 11308 9312 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 10928 11308 11345 11336
rect 10928 11296 10934 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 12894 11336 12900 11348
rect 12299 11308 12900 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 13688 11308 14228 11336
rect 13688 11296 13694 11308
rect 1452 11240 2176 11268
rect 1452 11228 1458 11240
rect 2148 11209 2176 11240
rect 2400 11271 2458 11277
rect 2400 11237 2412 11271
rect 2446 11268 2458 11271
rect 3970 11268 3976 11280
rect 2446 11240 3976 11268
rect 2446 11237 2458 11240
rect 2400 11231 2458 11237
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11268 4583 11271
rect 4614 11268 4620 11280
rect 4571 11240 4620 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11169 1639 11203
rect 1581 11163 1639 11169
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11169 2191 11203
rect 4540 11200 4568 11231
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 5534 11268 5540 11280
rect 4724 11240 5540 11268
rect 2133 11163 2191 11169
rect 2240 11172 4568 11200
rect 1596 11132 1624 11163
rect 2240 11132 2268 11172
rect 1596 11104 2268 11132
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 3936 11104 4629 11132
rect 3936 11092 3942 11104
rect 4617 11101 4629 11104
rect 4663 11132 4675 11135
rect 4724 11132 4752 11240
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 6086 11228 6092 11280
rect 6144 11268 6150 11280
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 6144 11240 7849 11268
rect 6144 11228 6150 11240
rect 7837 11237 7849 11240
rect 7883 11237 7895 11271
rect 7837 11231 7895 11237
rect 8941 11271 8999 11277
rect 8941 11237 8953 11271
rect 8987 11268 8999 11271
rect 9766 11268 9772 11280
rect 8987 11240 9772 11268
rect 8987 11237 8999 11240
rect 8941 11231 8999 11237
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 9858 11228 9864 11280
rect 9916 11268 9922 11280
rect 10198 11271 10256 11277
rect 10198 11268 10210 11271
rect 9916 11240 10210 11268
rect 9916 11228 9922 11240
rect 10198 11237 10210 11240
rect 10244 11237 10256 11271
rect 10198 11231 10256 11237
rect 10327 11240 13492 11268
rect 5442 11209 5448 11212
rect 5436 11200 5448 11209
rect 4816 11172 5448 11200
rect 4816 11141 4844 11172
rect 5436 11163 5448 11172
rect 5442 11160 5448 11163
rect 5500 11160 5506 11212
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 6604 11172 6868 11200
rect 6604 11160 6610 11172
rect 4663 11104 4752 11132
rect 4801 11135 4859 11141
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4801 11101 4813 11135
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 6730 11132 6736 11144
rect 5169 11095 5227 11101
rect 6196 11104 6736 11132
rect 5074 11064 5080 11076
rect 3068 11036 5080 11064
rect 1765 10999 1823 11005
rect 1765 10965 1777 10999
rect 1811 10996 1823 10999
rect 2038 10996 2044 11008
rect 1811 10968 2044 10996
rect 1811 10965 1823 10968
rect 1765 10959 1823 10965
rect 2038 10956 2044 10968
rect 2096 10956 2102 11008
rect 2130 10956 2136 11008
rect 2188 10996 2194 11008
rect 3068 10996 3096 11036
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 3510 10996 3516 11008
rect 2188 10968 3096 10996
rect 3471 10968 3516 10996
rect 2188 10956 2194 10968
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 5184 10996 5212 11095
rect 6196 10996 6224 11104
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6840 11132 6868 11172
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 7156 11172 7205 11200
rect 7156 11160 7162 11172
rect 7193 11169 7205 11172
rect 7239 11200 7251 11203
rect 7742 11200 7748 11212
rect 7239 11172 7748 11200
rect 7239 11169 7251 11172
rect 7193 11163 7251 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 9582 11200 9588 11212
rect 8527 11172 9588 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 9582 11160 9588 11172
rect 9640 11200 9646 11212
rect 10327 11200 10355 11240
rect 9640 11172 10355 11200
rect 9640 11160 9646 11172
rect 10594 11160 10600 11212
rect 10652 11200 10658 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 10652 11172 11713 11200
rect 10652 11160 10658 11172
rect 11701 11169 11713 11172
rect 11747 11200 11759 11203
rect 12526 11200 12532 11212
rect 11747 11172 12532 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 13170 11200 13176 11212
rect 12667 11172 13176 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 13464 11209 13492 11240
rect 13722 11228 13728 11280
rect 13780 11268 13786 11280
rect 13780 11240 14136 11268
rect 13780 11228 13786 11240
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11169 13507 11203
rect 13906 11200 13912 11212
rect 13867 11172 13912 11200
rect 13449 11163 13507 11169
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 7374 11132 7380 11144
rect 6840 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 8662 11132 8668 11144
rect 8312 11104 8668 11132
rect 6546 11064 6552 11076
rect 6507 11036 6552 11064
rect 6546 11024 6552 11036
rect 6604 11024 6610 11076
rect 6822 11064 6828 11076
rect 6783 11036 6828 11064
rect 6822 11024 6828 11036
rect 6880 11024 6886 11076
rect 8312 11073 8340 11104
rect 8662 11092 8668 11104
rect 8720 11132 8726 11144
rect 9214 11132 9220 11144
rect 8720 11104 9076 11132
rect 9175 11104 9220 11132
rect 8720 11092 8726 11104
rect 8297 11067 8355 11073
rect 8297 11033 8309 11067
rect 8343 11033 8355 11067
rect 8297 11027 8355 11033
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 8754 11064 8760 11076
rect 8619 11036 8760 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 8846 11024 8852 11076
rect 8904 11024 8910 11076
rect 9048 11064 9076 11104
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9950 11132 9956 11144
rect 9863 11104 9956 11132
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 9766 11064 9772 11076
rect 9048 11036 9772 11064
rect 9766 11024 9772 11036
rect 9824 11064 9830 11076
rect 9968 11064 9996 11092
rect 9824 11036 9996 11064
rect 11885 11067 11943 11073
rect 9824 11024 9830 11036
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 12250 11064 12256 11076
rect 11931 11036 12256 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 12820 11064 12848 11095
rect 13078 11092 13084 11144
rect 13136 11132 13142 11144
rect 13722 11132 13728 11144
rect 13136 11104 13728 11132
rect 13136 11092 13142 11104
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13998 11132 14004 11144
rect 13959 11104 14004 11132
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 14108 11141 14136 11240
rect 14200 11200 14228 11308
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 14200 11172 14657 11200
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 15749 11203 15807 11209
rect 15749 11200 15761 11203
rect 15344 11172 15761 11200
rect 15344 11160 15350 11172
rect 15749 11169 15761 11172
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 15930 11200 15936 11212
rect 15887 11172 15936 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11101 14151 11135
rect 16022 11132 16028 11144
rect 15983 11104 16028 11132
rect 14093 11095 14151 11101
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 12584 11036 12848 11064
rect 13265 11067 13323 11073
rect 12584 11024 12590 11036
rect 13265 11033 13277 11067
rect 13311 11064 13323 11067
rect 13446 11064 13452 11076
rect 13311 11036 13452 11064
rect 13311 11033 13323 11036
rect 13265 11027 13323 11033
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 14550 11064 14556 11076
rect 13587 11036 14556 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 14642 11024 14648 11076
rect 14700 11064 14706 11076
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 14700 11036 14841 11064
rect 14700 11024 14706 11036
rect 14829 11033 14841 11036
rect 14875 11033 14887 11067
rect 15470 11064 15476 11076
rect 14829 11027 14887 11033
rect 14936 11036 15476 11064
rect 5184 10968 6224 10996
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 8864 10996 8892 11024
rect 8720 10968 8892 10996
rect 8720 10956 8726 10968
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 12894 10996 12900 11008
rect 10652 10968 12900 10996
rect 10652 10956 10658 10968
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 14936 10996 14964 11036
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 15378 10996 15384 11008
rect 13412 10968 14964 10996
rect 15339 10968 15384 10996
rect 13412 10956 13418 10968
rect 15378 10956 15384 10968
rect 15436 10956 15442 11008
rect 1104 10906 16836 10928
rect 1104 10854 3614 10906
rect 3666 10854 3678 10906
rect 3730 10854 3742 10906
rect 3794 10854 3806 10906
rect 3858 10854 8878 10906
rect 8930 10854 8942 10906
rect 8994 10854 9006 10906
rect 9058 10854 9070 10906
rect 9122 10854 14142 10906
rect 14194 10854 14206 10906
rect 14258 10854 14270 10906
rect 14322 10854 14334 10906
rect 14386 10854 16836 10906
rect 1104 10832 16836 10854
rect 2590 10752 2596 10804
rect 2648 10792 2654 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2648 10764 2789 10792
rect 2648 10752 2654 10764
rect 2777 10761 2789 10764
rect 2823 10792 2835 10795
rect 3142 10792 3148 10804
rect 2823 10764 3148 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 5534 10792 5540 10804
rect 3988 10764 5540 10792
rect 2406 10684 2412 10736
rect 2464 10724 2470 10736
rect 3988 10724 4016 10764
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 5684 10764 6837 10792
rect 5684 10752 5690 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 8260 10764 9229 10792
rect 8260 10752 8266 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 9582 10792 9588 10804
rect 9543 10764 9588 10792
rect 9217 10755 9275 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 11146 10792 11152 10804
rect 9784 10764 11152 10792
rect 2464 10696 4016 10724
rect 2464 10684 2470 10696
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 4120 10696 4384 10724
rect 4120 10684 4126 10696
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 3510 10656 3516 10668
rect 3160 10628 3516 10656
rect 1664 10591 1722 10597
rect 1664 10557 1676 10591
rect 1710 10588 1722 10591
rect 3160 10588 3188 10628
rect 3510 10616 3516 10628
rect 3568 10656 3574 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3568 10628 3617 10656
rect 3568 10616 3574 10628
rect 3605 10625 3617 10628
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 1710 10560 3188 10588
rect 1710 10557 1722 10560
rect 1664 10551 1722 10557
rect 3234 10548 3240 10600
rect 3292 10588 3298 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3292 10560 3433 10588
rect 3292 10548 3298 10560
rect 3421 10557 3433 10560
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4246 10588 4252 10600
rect 4111 10560 4252 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 2774 10480 2780 10532
rect 2832 10520 2838 10532
rect 4356 10520 4384 10696
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 6365 10727 6423 10733
rect 4672 10696 6224 10724
rect 4672 10684 4678 10696
rect 5626 10656 5632 10668
rect 4908 10628 5488 10656
rect 5587 10628 5632 10656
rect 4908 10597 4936 10628
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 4982 10548 4988 10600
rect 5040 10588 5046 10600
rect 5350 10588 5356 10600
rect 5040 10560 5212 10588
rect 5311 10560 5356 10588
rect 5040 10548 5046 10560
rect 5184 10520 5212 10560
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 5460 10588 5488 10628
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 6086 10588 6092 10600
rect 5460 10560 6092 10588
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6196 10588 6224 10696
rect 6365 10693 6377 10727
rect 6411 10724 6423 10727
rect 6411 10696 7604 10724
rect 6411 10693 6423 10696
rect 6365 10687 6423 10693
rect 6822 10616 6828 10668
rect 6880 10656 6886 10668
rect 6880 10628 7328 10656
rect 6880 10616 6886 10628
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6196 10560 6653 10588
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 6788 10560 7205 10588
rect 6788 10548 6794 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7300 10588 7328 10628
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 7576 10656 7604 10696
rect 7432 10628 7477 10656
rect 7576 10628 7972 10656
rect 7432 10616 7438 10628
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 7300 10560 7849 10588
rect 7193 10551 7251 10557
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 2832 10492 5120 10520
rect 5184 10492 7297 10520
rect 2832 10480 2838 10492
rect 2406 10412 2412 10464
rect 2464 10452 2470 10464
rect 3053 10455 3111 10461
rect 3053 10452 3065 10455
rect 2464 10424 3065 10452
rect 2464 10412 2470 10424
rect 3053 10421 3065 10424
rect 3099 10421 3111 10455
rect 3510 10452 3516 10464
rect 3471 10424 3516 10452
rect 3053 10415 3111 10421
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 3936 10424 4261 10452
rect 3936 10412 3942 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 4614 10412 4620 10464
rect 4672 10452 4678 10464
rect 4709 10455 4767 10461
rect 4709 10452 4721 10455
rect 4672 10424 4721 10452
rect 4672 10412 4678 10424
rect 4709 10421 4721 10424
rect 4755 10421 4767 10455
rect 4982 10452 4988 10464
rect 4943 10424 4988 10452
rect 4709 10415 4767 10421
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 5092 10452 5120 10492
rect 7285 10489 7297 10492
rect 7331 10489 7343 10523
rect 7944 10520 7972 10628
rect 8110 10597 8116 10600
rect 8104 10588 8116 10597
rect 8071 10560 8116 10588
rect 8104 10551 8116 10560
rect 8110 10548 8116 10551
rect 8168 10548 8174 10600
rect 9490 10588 9496 10600
rect 9140 10560 9496 10588
rect 9140 10532 9168 10560
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9784 10597 9812 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11330 10792 11336 10804
rect 11291 10764 11336 10792
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 15654 10792 15660 10804
rect 11440 10764 15660 10792
rect 10321 10727 10379 10733
rect 10321 10693 10333 10727
rect 10367 10724 10379 10727
rect 10594 10724 10600 10736
rect 10367 10696 10600 10724
rect 10367 10693 10379 10696
rect 10321 10687 10379 10693
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 11440 10724 11468 10764
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 10796 10696 11468 10724
rect 9769 10591 9827 10597
rect 9769 10557 9781 10591
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 10796 10588 10824 10696
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12066 10656 12072 10668
rect 12023 10628 12072 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 10735 10560 10824 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 9122 10520 9128 10532
rect 7944 10492 9128 10520
rect 7285 10483 7343 10489
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 9456 10492 10793 10520
rect 9456 10480 9462 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 10781 10483 10839 10489
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 5092 10424 5457 10452
rect 5445 10421 5457 10424
rect 5491 10452 5503 10455
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 5491 10424 6377 10452
rect 5491 10421 5503 10424
rect 5445 10415 5503 10421
rect 6365 10421 6377 10424
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 6457 10455 6515 10461
rect 6457 10421 6469 10455
rect 6503 10452 6515 10455
rect 6822 10452 6828 10464
rect 6503 10424 6828 10452
rect 6503 10421 6515 10424
rect 6457 10415 6515 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7098 10452 7104 10464
rect 6972 10424 7104 10452
rect 6972 10412 6978 10424
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 9582 10452 9588 10464
rect 7524 10424 9588 10452
rect 7524 10412 7530 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10594 10412 10600 10464
rect 10652 10452 10658 10464
rect 10888 10452 10916 10619
rect 12066 10616 12072 10628
rect 12124 10616 12130 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 13464 10628 14933 10656
rect 13464 10600 13492 10628
rect 14921 10625 14933 10628
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 13446 10588 13452 10600
rect 12483 10560 13452 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14369 10591 14427 10597
rect 14369 10588 14381 10591
rect 13872 10560 14381 10588
rect 13872 10548 13878 10560
rect 14369 10557 14381 10560
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 11701 10523 11759 10529
rect 11701 10489 11713 10523
rect 11747 10520 11759 10523
rect 11747 10492 12572 10520
rect 11747 10489 11759 10492
rect 11701 10483 11759 10489
rect 10652 10424 10916 10452
rect 11793 10455 11851 10461
rect 10652 10412 10658 10424
rect 11793 10421 11805 10455
rect 11839 10452 11851 10455
rect 12066 10452 12072 10464
rect 11839 10424 12072 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 12544 10452 12572 10492
rect 12618 10480 12624 10532
rect 12676 10529 12682 10532
rect 12676 10523 12740 10529
rect 12676 10489 12694 10523
rect 12728 10489 12740 10523
rect 12676 10483 12740 10489
rect 12676 10480 12682 10483
rect 13170 10480 13176 10532
rect 13228 10520 13234 10532
rect 15194 10529 15200 10532
rect 15188 10520 15200 10529
rect 13228 10492 14964 10520
rect 15155 10492 15200 10520
rect 13228 10480 13234 10492
rect 12802 10452 12808 10464
rect 12544 10424 12808 10452
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13262 10412 13268 10464
rect 13320 10452 13326 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13320 10424 13829 10452
rect 13320 10412 13326 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14553 10455 14611 10461
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 14826 10452 14832 10464
rect 14599 10424 14832 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 14936 10452 14964 10492
rect 15188 10483 15200 10492
rect 15194 10480 15200 10483
rect 15252 10480 15258 10532
rect 16301 10455 16359 10461
rect 16301 10452 16313 10455
rect 14936 10424 16313 10452
rect 16301 10421 16313 10424
rect 16347 10421 16359 10455
rect 16301 10415 16359 10421
rect 1104 10362 16836 10384
rect 1104 10310 6246 10362
rect 6298 10310 6310 10362
rect 6362 10310 6374 10362
rect 6426 10310 6438 10362
rect 6490 10310 11510 10362
rect 11562 10310 11574 10362
rect 11626 10310 11638 10362
rect 11690 10310 11702 10362
rect 11754 10310 16836 10362
rect 1104 10288 16836 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 2498 10248 2504 10260
rect 1995 10220 2504 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 2958 10248 2964 10260
rect 2919 10220 2964 10248
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 3292 10220 5396 10248
rect 3292 10208 3298 10220
rect 2314 10180 2320 10192
rect 2275 10152 2320 10180
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 2406 10140 2412 10192
rect 2464 10180 2470 10192
rect 3421 10183 3479 10189
rect 3421 10180 3433 10183
rect 2464 10152 2509 10180
rect 2608 10152 3433 10180
rect 2464 10140 2470 10152
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2498 10072 2504 10124
rect 2556 10112 2562 10124
rect 2608 10112 2636 10152
rect 3421 10149 3433 10152
rect 3467 10180 3479 10183
rect 4062 10180 4068 10192
rect 3467 10152 4068 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 4430 10140 4436 10192
rect 4488 10180 4494 10192
rect 4586 10183 4644 10189
rect 4586 10180 4598 10183
rect 4488 10152 4598 10180
rect 4488 10140 4494 10152
rect 4586 10149 4598 10152
rect 4632 10149 4644 10183
rect 5368 10180 5396 10220
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5626 10248 5632 10260
rect 5500 10220 5632 10248
rect 5500 10208 5506 10220
rect 5626 10208 5632 10220
rect 5684 10248 5690 10260
rect 5721 10251 5779 10257
rect 5721 10248 5733 10251
rect 5684 10220 5733 10248
rect 5684 10208 5690 10220
rect 5721 10217 5733 10220
rect 5767 10217 5779 10251
rect 5721 10211 5779 10217
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 7466 10248 7472 10260
rect 6052 10220 7472 10248
rect 6052 10208 6058 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 8168 10220 8217 10248
rect 8168 10208 8174 10220
rect 8205 10217 8217 10220
rect 8251 10217 8263 10251
rect 10410 10248 10416 10260
rect 10371 10220 10416 10248
rect 8205 10211 8263 10217
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10248 10563 10251
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10551 10220 10885 10248
rect 10551 10217 10563 10220
rect 10505 10211 10563 10217
rect 10873 10217 10885 10220
rect 10919 10248 10931 10251
rect 11882 10248 11888 10260
rect 10919 10220 11888 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 12066 10248 12072 10260
rect 12027 10220 12072 10248
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12529 10251 12587 10257
rect 12529 10248 12541 10251
rect 12176 10220 12541 10248
rect 5368 10152 7880 10180
rect 4586 10143 4644 10149
rect 2556 10084 2636 10112
rect 3329 10115 3387 10121
rect 2556 10072 2562 10084
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 4338 10112 4344 10124
rect 3375 10084 4016 10112
rect 4299 10084 4344 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 3988 10044 4016 10084
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 5994 10112 6000 10124
rect 4448 10084 6000 10112
rect 4448 10044 4476 10084
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 7098 10121 7104 10124
rect 7092 10112 7104 10121
rect 7059 10084 7104 10112
rect 7092 10075 7104 10084
rect 7098 10072 7104 10075
rect 7156 10072 7162 10124
rect 6822 10044 6828 10056
rect 3660 10016 3705 10044
rect 3988 10016 4476 10044
rect 6783 10016 6828 10044
rect 3660 10004 3666 10016
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7852 10044 7880 10152
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 8536 10152 9045 10180
rect 8536 10140 8542 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 11977 10183 12035 10189
rect 11977 10180 11989 10183
rect 9033 10143 9091 10149
rect 9140 10152 11989 10180
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 8352 10084 8953 10112
rect 8352 10072 8358 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 9140 10112 9168 10152
rect 11977 10149 11989 10152
rect 12023 10149 12035 10183
rect 11977 10143 12035 10149
rect 8941 10075 8999 10081
rect 9048 10084 9168 10112
rect 9048 10044 9076 10084
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 10873 10115 10931 10121
rect 10873 10112 10885 10115
rect 9640 10084 10885 10112
rect 9640 10072 9646 10084
rect 10873 10081 10885 10084
rect 10919 10081 10931 10115
rect 11422 10112 11428 10124
rect 10873 10075 10931 10081
rect 10971 10084 11428 10112
rect 9214 10044 9220 10056
rect 7852 10016 9076 10044
rect 9127 10016 9220 10044
rect 9214 10004 9220 10016
rect 9272 10044 9278 10056
rect 10226 10044 10232 10056
rect 9272 10016 10232 10044
rect 9272 10004 9278 10016
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10594 10044 10600 10056
rect 10555 10016 10600 10044
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10971 10044 10999 10084
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 12176 10112 12204 10220
rect 12529 10217 12541 10220
rect 12575 10217 12587 10251
rect 12529 10211 12587 10217
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12860 10220 13093 10248
rect 12860 10208 12866 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 13081 10211 13139 10217
rect 13541 10251 13599 10257
rect 13541 10217 13553 10251
rect 13587 10248 13599 10251
rect 13722 10248 13728 10260
rect 13587 10220 13728 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14550 10248 14556 10260
rect 14511 10220 14556 10248
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 15657 10251 15715 10257
rect 15657 10248 15669 10251
rect 15436 10220 15669 10248
rect 15436 10208 15442 10220
rect 15657 10217 15669 10220
rect 15703 10217 15715 10251
rect 15657 10211 15715 10217
rect 15194 10180 15200 10192
rect 11532 10084 12204 10112
rect 12268 10152 15200 10180
rect 10704 10016 10999 10044
rect 1578 9976 1584 9988
rect 1539 9948 1584 9976
rect 1578 9936 1584 9948
rect 1636 9936 1642 9988
rect 2038 9936 2044 9988
rect 2096 9976 2102 9988
rect 3234 9976 3240 9988
rect 2096 9948 3240 9976
rect 2096 9936 2102 9948
rect 3234 9936 3240 9948
rect 3292 9936 3298 9988
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 3384 9948 3464 9976
rect 3384 9936 3390 9948
rect 3436 9920 3464 9948
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 6730 9976 6736 9988
rect 5684 9948 6736 9976
rect 5684 9936 5690 9948
rect 6730 9936 6736 9948
rect 6788 9936 6794 9988
rect 9398 9976 9404 9988
rect 7760 9948 9404 9976
rect 3418 9868 3424 9920
rect 3476 9868 3482 9920
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 4982 9908 4988 9920
rect 4304 9880 4988 9908
rect 4304 9868 4310 9880
rect 4982 9868 4988 9880
rect 5040 9908 5046 9920
rect 7760 9908 7788 9948
rect 9398 9936 9404 9948
rect 9456 9936 9462 9988
rect 10704 9976 10732 10016
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11532 10053 11560 10084
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11112 10016 11529 10044
rect 11112 10004 11118 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10044 11759 10047
rect 12268 10044 12296 10152
rect 15194 10140 15200 10152
rect 15252 10140 15258 10192
rect 15746 10180 15752 10192
rect 15707 10152 15752 10180
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 12526 10112 12532 10124
rect 12483 10084 12532 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 14001 10115 14059 10121
rect 13495 10084 13768 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 12618 10044 12624 10056
rect 11747 10016 12296 10044
rect 12579 10016 12624 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 12618 10004 12624 10016
rect 12676 10044 12682 10056
rect 13633 10047 13691 10053
rect 13633 10044 13645 10047
rect 12676 10016 13645 10044
rect 12676 10004 12682 10016
rect 13633 10013 13645 10016
rect 13679 10013 13691 10047
rect 13740 10044 13768 10084
rect 14001 10081 14013 10115
rect 14047 10112 14059 10115
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 14047 10084 14473 10112
rect 14047 10081 14059 10084
rect 14001 10075 14059 10081
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 16022 10112 16028 10124
rect 14461 10075 14519 10081
rect 15212 10084 16028 10112
rect 14182 10044 14188 10056
rect 13740 10016 14188 10044
rect 13633 10007 13691 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14274 10004 14280 10056
rect 14332 10044 14338 10056
rect 14550 10044 14556 10056
rect 14332 10016 14556 10044
rect 14332 10004 14338 10016
rect 14550 10004 14556 10016
rect 14608 10004 14614 10056
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 15212 10044 15240 10084
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 15838 10044 15844 10056
rect 14783 10016 15240 10044
rect 15799 10016 15844 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 9600 9948 10732 9976
rect 8570 9908 8576 9920
rect 5040 9880 7788 9908
rect 8531 9880 8576 9908
rect 5040 9868 5046 9880
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 9600 9908 9628 9948
rect 10778 9936 10784 9988
rect 10836 9976 10842 9988
rect 14001 9979 14059 9985
rect 14001 9976 14013 9979
rect 10836 9948 14013 9976
rect 10836 9936 10842 9948
rect 14001 9945 14013 9948
rect 14047 9945 14059 9979
rect 14001 9939 14059 9945
rect 14093 9979 14151 9985
rect 14093 9945 14105 9979
rect 14139 9976 14151 9979
rect 15746 9976 15752 9988
rect 14139 9948 15752 9976
rect 14139 9945 14151 9948
rect 14093 9939 14151 9945
rect 15746 9936 15752 9948
rect 15804 9936 15810 9988
rect 8720 9880 9628 9908
rect 8720 9868 8726 9880
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10045 9911 10103 9917
rect 10045 9908 10057 9911
rect 9732 9880 10057 9908
rect 9732 9868 9738 9880
rect 10045 9877 10057 9880
rect 10091 9877 10103 9911
rect 11054 9908 11060 9920
rect 11015 9880 11060 9908
rect 10045 9871 10103 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9908 12035 9911
rect 14918 9908 14924 9920
rect 12023 9880 14924 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 14918 9868 14924 9880
rect 14976 9868 14982 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15289 9911 15347 9917
rect 15289 9908 15301 9911
rect 15252 9880 15301 9908
rect 15252 9868 15258 9880
rect 15289 9877 15301 9880
rect 15335 9877 15347 9911
rect 15289 9871 15347 9877
rect 1104 9818 16836 9840
rect 1104 9766 3614 9818
rect 3666 9766 3678 9818
rect 3730 9766 3742 9818
rect 3794 9766 3806 9818
rect 3858 9766 8878 9818
rect 8930 9766 8942 9818
rect 8994 9766 9006 9818
rect 9058 9766 9070 9818
rect 9122 9766 14142 9818
rect 14194 9766 14206 9818
rect 14258 9766 14270 9818
rect 14322 9766 14334 9818
rect 14386 9766 16836 9818
rect 1104 9744 16836 9766
rect 5166 9704 5172 9716
rect 3896 9676 5172 9704
rect 2682 9596 2688 9648
rect 2740 9636 2746 9648
rect 2777 9639 2835 9645
rect 2777 9636 2789 9639
rect 2740 9608 2789 9636
rect 2740 9596 2746 9608
rect 2777 9605 2789 9608
rect 2823 9605 2835 9639
rect 3050 9636 3056 9648
rect 3011 9608 3056 9636
rect 2777 9599 2835 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 3234 9596 3240 9648
rect 3292 9596 3298 9648
rect 3252 9568 3280 9596
rect 3068 9540 3280 9568
rect 3068 9512 3096 9540
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3568 9540 3617 9568
rect 3568 9528 3574 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1486 9500 1492 9512
rect 1443 9472 1492 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 1664 9503 1722 9509
rect 1664 9469 1676 9503
rect 1710 9500 1722 9503
rect 2590 9500 2596 9512
rect 1710 9472 2596 9500
rect 1710 9469 1722 9472
rect 1664 9463 1722 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 3050 9460 3056 9512
rect 3108 9460 3114 9512
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3896 9500 3924 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5592 9676 6868 9704
rect 5592 9664 5598 9676
rect 4522 9636 4528 9648
rect 4172 9608 4528 9636
rect 4062 9500 4068 9512
rect 3292 9472 3924 9500
rect 4023 9472 4068 9500
rect 3292 9460 3298 9472
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9432 3479 9435
rect 3786 9432 3792 9444
rect 3467 9404 3792 9432
rect 3467 9401 3479 9404
rect 3421 9395 3479 9401
rect 3786 9392 3792 9404
rect 3844 9392 3850 9444
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 2188 9336 3525 9364
rect 2188 9324 2194 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3513 9327 3571 9333
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 4172 9364 4200 9608
rect 4522 9596 4528 9608
rect 4580 9596 4586 9648
rect 4706 9596 4712 9648
rect 4764 9596 4770 9648
rect 4985 9639 5043 9645
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 5626 9636 5632 9648
rect 5031 9608 5632 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 6840 9636 6868 9676
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 8205 9707 8263 9713
rect 8205 9704 8217 9707
rect 7156 9676 8217 9704
rect 7156 9664 7162 9676
rect 8205 9673 8217 9676
rect 8251 9673 8263 9707
rect 8205 9667 8263 9673
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 10652 9676 11928 9704
rect 10652 9664 10658 9676
rect 6788 9608 6868 9636
rect 8573 9639 8631 9645
rect 6788 9596 6794 9608
rect 8573 9605 8585 9639
rect 8619 9636 8631 9639
rect 9398 9636 9404 9648
rect 8619 9608 9404 9636
rect 8619 9605 8631 9608
rect 8573 9599 8631 9605
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 11900 9636 11928 9676
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 14550 9704 14556 9716
rect 12584 9676 13860 9704
rect 12584 9664 12590 9676
rect 13832 9636 13860 9676
rect 14384 9676 14556 9704
rect 14384 9648 14412 9676
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 14090 9636 14096 9648
rect 11900 9608 12020 9636
rect 13832 9608 14096 9636
rect 4246 9528 4252 9580
rect 4304 9568 4310 9580
rect 4614 9568 4620 9580
rect 4304 9540 4620 9568
rect 4304 9528 4310 9540
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 3936 9336 4200 9364
rect 4249 9367 4307 9373
rect 3936 9324 3942 9336
rect 4249 9333 4261 9367
rect 4295 9364 4307 9367
rect 4522 9364 4528 9376
rect 4295 9336 4528 9364
rect 4295 9333 4307 9336
rect 4249 9327 4307 9333
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 4724 9364 4752 9596
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 11992 9577 12020 9608
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14366 9596 14372 9648
rect 14424 9596 14430 9648
rect 14734 9596 14740 9648
rect 14792 9636 14798 9648
rect 14792 9608 15332 9636
rect 14792 9596 14798 9608
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9568 9275 9571
rect 11977 9571 12035 9577
rect 9263 9540 9720 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 5074 9460 5080 9512
rect 5132 9460 5138 9512
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5408 9472 5457 9500
rect 5408 9460 5414 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5960 9472 6009 9500
rect 5960 9460 5966 9472
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 5997 9463 6055 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 9582 9500 9588 9512
rect 7892 9472 9588 9500
rect 7892 9460 7898 9472
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 9692 9500 9720 9540
rect 10888 9540 11284 9568
rect 10888 9500 10916 9540
rect 11256 9500 11284 9540
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 11606 9500 11612 9512
rect 9692 9472 10916 9500
rect 10971 9472 11100 9500
rect 11256 9472 11612 9500
rect 5092 9376 5120 9460
rect 7092 9435 7150 9441
rect 7092 9401 7104 9435
rect 7138 9432 7150 9435
rect 7190 9432 7196 9444
rect 7138 9404 7196 9432
rect 7138 9401 7150 9404
rect 7092 9395 7150 9401
rect 7190 9392 7196 9404
rect 7248 9432 7254 9444
rect 7466 9432 7472 9444
rect 7248 9404 7472 9432
rect 7248 9392 7254 9404
rect 7466 9392 7472 9404
rect 7524 9392 7530 9444
rect 8941 9435 8999 9441
rect 8941 9401 8953 9435
rect 8987 9432 8999 9435
rect 9674 9432 9680 9444
rect 8987 9404 9680 9432
rect 8987 9401 8999 9404
rect 8941 9395 8999 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9858 9441 9864 9444
rect 9852 9395 9864 9441
rect 9916 9432 9922 9444
rect 10042 9432 10048 9444
rect 9916 9404 10048 9432
rect 9858 9392 9864 9395
rect 9916 9392 9922 9404
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10971 9432 10999 9472
rect 10152 9404 10999 9432
rect 11072 9432 11100 9472
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 11698 9460 11704 9512
rect 11756 9500 11762 9512
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 11756 9472 11805 9500
rect 11756 9460 11762 9472
rect 11793 9469 11805 9472
rect 11839 9469 11851 9503
rect 11992 9500 12020 9531
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 15010 9568 15016 9580
rect 14700 9540 15016 9568
rect 14700 9528 14706 9540
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 15194 9568 15200 9580
rect 15155 9540 15200 9568
rect 15194 9528 15200 9540
rect 15252 9528 15258 9580
rect 15304 9577 15332 9608
rect 15289 9571 15347 9577
rect 15289 9537 15301 9571
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 12805 9503 12863 9509
rect 11992 9472 12664 9500
rect 11793 9463 11851 9469
rect 11072 9404 11376 9432
rect 4672 9336 4752 9364
rect 4672 9324 4678 9336
rect 5074 9324 5080 9376
rect 5132 9324 5138 9376
rect 5353 9367 5411 9373
rect 5353 9333 5365 9367
rect 5399 9364 5411 9367
rect 5442 9364 5448 9376
rect 5399 9336 5448 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6181 9367 6239 9373
rect 6181 9364 6193 9367
rect 5960 9336 6193 9364
rect 5960 9324 5966 9336
rect 6181 9333 6193 9336
rect 6227 9333 6239 9367
rect 6181 9327 6239 9333
rect 9033 9367 9091 9373
rect 9033 9333 9045 9367
rect 9079 9364 9091 9367
rect 10152 9364 10180 9404
rect 9079 9336 10180 9364
rect 9079 9333 9091 9336
rect 9033 9327 9091 9333
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 11348 9373 11376 9404
rect 11422 9392 11428 9444
rect 11480 9392 11486 9444
rect 12437 9435 12495 9441
rect 12437 9401 12449 9435
rect 12483 9432 12495 9435
rect 12526 9432 12532 9444
rect 12483 9404 12532 9432
rect 12483 9401 12495 9404
rect 12437 9395 12495 9401
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12636 9432 12664 9472
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12851 9472 12909 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 15102 9500 15108 9512
rect 15063 9472 15108 9500
rect 12897 9463 12955 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 15841 9503 15899 9509
rect 15841 9469 15853 9503
rect 15887 9469 15899 9503
rect 15841 9463 15899 9469
rect 13170 9441 13176 9444
rect 13164 9432 13176 9441
rect 12636 9404 13176 9432
rect 13164 9395 13176 9404
rect 13170 9392 13176 9395
rect 13228 9392 13234 9444
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 15856 9432 15884 9463
rect 14056 9404 15884 9432
rect 16117 9435 16175 9441
rect 14056 9392 14062 9404
rect 16117 9401 16129 9435
rect 16163 9432 16175 9435
rect 16574 9432 16580 9444
rect 16163 9404 16580 9432
rect 16163 9401 16175 9404
rect 16117 9395 16175 9401
rect 16574 9392 16580 9404
rect 16632 9392 16638 9444
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10284 9336 10977 9364
rect 10284 9324 10290 9336
rect 10965 9333 10977 9336
rect 11011 9333 11023 9367
rect 10965 9327 11023 9333
rect 11333 9367 11391 9373
rect 11333 9333 11345 9367
rect 11379 9333 11391 9367
rect 11440 9364 11468 9392
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11440 9336 11713 9364
rect 11333 9327 11391 9333
rect 11701 9333 11713 9336
rect 11747 9364 11759 9367
rect 12066 9364 12072 9376
rect 11747 9336 12072 9364
rect 11747 9333 11759 9336
rect 11701 9327 11759 9333
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 12710 9364 12716 9376
rect 12400 9336 12716 9364
rect 12400 9324 12406 9336
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 13446 9364 13452 9376
rect 12860 9336 13452 9364
rect 12860 9324 12866 9336
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 14274 9364 14280 9376
rect 14235 9336 14280 9364
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 14792 9336 14837 9364
rect 14792 9324 14798 9336
rect 1104 9274 16836 9296
rect 1104 9222 6246 9274
rect 6298 9222 6310 9274
rect 6362 9222 6374 9274
rect 6426 9222 6438 9274
rect 6490 9222 11510 9274
rect 11562 9222 11574 9274
rect 11626 9222 11638 9274
rect 11690 9222 11702 9274
rect 11754 9222 16836 9274
rect 1104 9200 16836 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1544 9132 1593 9160
rect 1544 9120 1550 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 1596 9092 1624 9123
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2406 9160 2412 9172
rect 2004 9132 2412 9160
rect 2004 9120 2010 9132
rect 2406 9120 2412 9132
rect 2464 9160 2470 9172
rect 3329 9163 3387 9169
rect 2464 9132 2912 9160
rect 2464 9120 2470 9132
rect 2124 9095 2182 9101
rect 1596 9064 1900 9092
rect 1872 9033 1900 9064
rect 2124 9061 2136 9095
rect 2170 9092 2182 9095
rect 2682 9092 2688 9104
rect 2170 9064 2688 9092
rect 2170 9061 2182 9064
rect 2124 9055 2182 9061
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 2884 9092 2912 9132
rect 3329 9129 3341 9163
rect 3375 9160 3387 9163
rect 4062 9160 4068 9172
rect 3375 9132 4068 9160
rect 3375 9129 3387 9132
rect 3329 9123 3387 9129
rect 4062 9120 4068 9132
rect 4120 9160 4126 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 4120 9132 9413 9160
rect 4120 9120 4126 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 12069 9163 12127 9169
rect 12069 9129 12081 9163
rect 12115 9160 12127 9163
rect 12618 9160 12624 9172
rect 12115 9132 12624 9160
rect 12115 9129 12127 9132
rect 12069 9123 12127 9129
rect 2884 9064 4108 9092
rect 4080 9036 4108 9064
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 4338 9092 4344 9104
rect 4212 9064 4344 9092
rect 4212 9052 4218 9064
rect 4338 9052 4344 9064
rect 4396 9092 4402 9104
rect 4494 9095 4552 9101
rect 4494 9092 4506 9095
rect 4396 9064 4506 9092
rect 4396 9052 4402 9064
rect 4494 9061 4506 9064
rect 4540 9061 4552 9095
rect 4494 9055 4552 9061
rect 4706 9052 4712 9104
rect 4764 9052 4770 9104
rect 6822 9092 6828 9104
rect 5920 9064 6828 9092
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 8993 1823 9027
rect 1765 8987 1823 8993
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 1946 9024 1952 9036
rect 1903 8996 1952 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 1780 8820 1808 8987
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 3513 9027 3571 9033
rect 3513 9024 3525 9027
rect 2556 8996 3525 9024
rect 2556 8984 2562 8996
rect 3513 8993 3525 8996
rect 3559 8993 3571 9027
rect 3513 8987 3571 8993
rect 4062 8984 4068 9036
rect 4120 8984 4126 9036
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4724 9024 4752 9052
rect 4295 8996 4752 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 5810 9024 5816 9036
rect 5684 8996 5816 9024
rect 5684 8984 5690 8996
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 5920 9033 5948 9064
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 8662 9092 8668 9104
rect 7760 9064 8668 9092
rect 7760 9033 7788 9064
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 9692 9092 9720 9123
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 13998 9160 14004 9172
rect 13959 9132 14004 9160
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14369 9163 14427 9169
rect 14369 9129 14381 9163
rect 14415 9160 14427 9163
rect 15289 9163 15347 9169
rect 15289 9160 15301 9163
rect 14415 9132 15301 9160
rect 14415 9129 14427 9132
rect 14369 9123 14427 9129
rect 15289 9129 15301 9132
rect 15335 9129 15347 9163
rect 15289 9123 15347 9129
rect 15749 9095 15807 9101
rect 15749 9092 15761 9095
rect 9692 9064 15761 9092
rect 15749 9061 15761 9064
rect 15795 9061 15807 9095
rect 15749 9055 15807 9061
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 8993 5963 9027
rect 6161 9027 6219 9033
rect 6161 9024 6173 9027
rect 5905 8987 5963 8993
rect 6012 8996 6173 9024
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3329 8959 3387 8965
rect 3329 8956 3341 8959
rect 3108 8928 3341 8956
rect 3108 8916 3114 8928
rect 3329 8925 3341 8928
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 6012 8956 6040 8996
rect 6161 8993 6173 8996
rect 6207 8993 6219 9027
rect 6161 8987 6219 8993
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 8993 7803 9027
rect 7745 8987 7803 8993
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 7892 8996 7941 9024
rect 7892 8984 7898 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 8196 9027 8254 9033
rect 8196 8993 8208 9027
rect 8242 9024 8254 9027
rect 9214 9024 9220 9036
rect 8242 8996 9220 9024
rect 8242 8993 8254 8996
rect 8196 8987 8254 8993
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 9024 10106 9036
rect 10226 9024 10232 9036
rect 10100 8996 10232 9024
rect 10100 8984 10106 8996
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10956 9027 11014 9033
rect 10956 8993 10968 9027
rect 11002 9024 11014 9027
rect 12066 9024 12072 9036
rect 11002 8996 12072 9024
rect 11002 8993 11014 8996
rect 10956 8987 11014 8993
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12601 9027 12659 9033
rect 12601 9024 12613 9027
rect 12492 8996 12613 9024
rect 12492 8984 12498 8996
rect 12601 8993 12613 8996
rect 12647 9024 12659 9027
rect 14274 9024 14280 9036
rect 12647 8996 14280 9024
rect 12647 8993 12659 8996
rect 12601 8987 12659 8993
rect 14274 8984 14280 8996
rect 14332 9024 14338 9036
rect 15657 9027 15715 9033
rect 14332 8996 14679 9024
rect 14332 8984 14338 8996
rect 9858 8956 9864 8968
rect 5316 8928 6040 8956
rect 8956 8928 9864 8956
rect 5316 8916 5322 8928
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 3237 8891 3295 8897
rect 3237 8888 3249 8891
rect 2924 8860 3249 8888
rect 2924 8848 2930 8860
rect 3237 8857 3249 8860
rect 3283 8888 3295 8891
rect 3418 8888 3424 8900
rect 3283 8860 3424 8888
rect 3283 8857 3295 8860
rect 3237 8851 3295 8857
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 4246 8820 4252 8832
rect 1780 8792 4252 8820
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 5644 8829 5672 8928
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7561 8891 7619 8897
rect 7561 8888 7573 8891
rect 7248 8860 7573 8888
rect 7248 8848 7254 8860
rect 7561 8857 7573 8860
rect 7607 8857 7619 8891
rect 7561 8851 7619 8857
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 5592 8792 5641 8820
rect 5592 8780 5598 8792
rect 5629 8789 5641 8792
rect 5675 8789 5687 8823
rect 5629 8783 5687 8789
rect 7285 8823 7343 8829
rect 7285 8789 7297 8823
rect 7331 8820 7343 8823
rect 7466 8820 7472 8832
rect 7331 8792 7472 8820
rect 7331 8789 7343 8792
rect 7285 8783 7343 8789
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8956 8820 8984 8928
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 10134 8956 10140 8968
rect 10008 8928 10140 8956
rect 10008 8916 10014 8928
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10594 8956 10600 8968
rect 10367 8928 10600 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 10689 8919 10747 8925
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 10704 8888 10732 8919
rect 9732 8860 10732 8888
rect 9732 8848 9738 8860
rect 9306 8820 9312 8832
rect 8260 8792 8984 8820
rect 9267 8792 9312 8820
rect 8260 8780 8266 8792
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 9401 8823 9459 8829
rect 9401 8789 9413 8823
rect 9447 8820 9459 8823
rect 12158 8820 12164 8832
rect 9447 8792 12164 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12360 8820 12388 8919
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 13998 8956 14004 8968
rect 13872 8928 14004 8956
rect 13872 8916 13878 8928
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 14458 8956 14464 8968
rect 14419 8928 14464 8956
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14651 8956 14679 8996
rect 15657 8993 15669 9027
rect 15703 9024 15715 9027
rect 15703 8996 15976 9024
rect 15703 8993 15715 8996
rect 15657 8987 15715 8993
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 14651 8928 15853 8956
rect 14553 8919 14611 8925
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 13446 8848 13452 8900
rect 13504 8888 13510 8900
rect 13725 8891 13783 8897
rect 13725 8888 13737 8891
rect 13504 8860 13737 8888
rect 13504 8848 13510 8860
rect 13725 8857 13737 8860
rect 13771 8888 13783 8891
rect 14568 8888 14596 8919
rect 13771 8860 14596 8888
rect 13771 8857 13783 8860
rect 13725 8851 13783 8857
rect 12710 8820 12716 8832
rect 12360 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 12986 8780 12992 8832
rect 13044 8820 13050 8832
rect 15948 8820 15976 8996
rect 13044 8792 15976 8820
rect 13044 8780 13050 8792
rect 1104 8730 16836 8752
rect 1104 8678 3614 8730
rect 3666 8678 3678 8730
rect 3730 8678 3742 8730
rect 3794 8678 3806 8730
rect 3858 8678 8878 8730
rect 8930 8678 8942 8730
rect 8994 8678 9006 8730
rect 9058 8678 9070 8730
rect 9122 8678 14142 8730
rect 14194 8678 14206 8730
rect 14258 8678 14270 8730
rect 14322 8678 14334 8730
rect 14386 8678 16836 8730
rect 1104 8656 16836 8678
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2222 8616 2228 8628
rect 2179 8588 2228 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2222 8576 2228 8588
rect 2280 8576 2286 8628
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 4525 8619 4583 8625
rect 4525 8616 4537 8619
rect 4396 8588 4537 8616
rect 4396 8576 4402 8588
rect 4525 8585 4537 8588
rect 4571 8585 4583 8619
rect 4525 8579 4583 8585
rect 4890 8576 4896 8628
rect 4948 8576 4954 8628
rect 11882 8616 11888 8628
rect 7300 8588 11888 8616
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 2866 8548 2872 8560
rect 1811 8520 2872 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 4908 8548 4936 8576
rect 4212 8520 4936 8548
rect 4212 8508 4218 8520
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 5316 8520 6960 8548
rect 5316 8508 5322 8520
rect 6932 8492 6960 8520
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2648 8452 2697 8480
rect 2648 8440 2654 8452
rect 2685 8449 2697 8452
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3050 8480 3056 8492
rect 2832 8452 3056 8480
rect 2832 8440 2838 8452
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 4396 8452 5825 8480
rect 4396 8440 4402 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7300 8489 7328 8588
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 12621 8619 12679 8625
rect 12621 8585 12633 8619
rect 12667 8616 12679 8619
rect 13814 8616 13820 8628
rect 12667 8588 13820 8616
rect 12667 8585 12679 8588
rect 12621 8579 12679 8585
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14056 8588 15700 8616
rect 14056 8576 14062 8588
rect 9493 8551 9551 8557
rect 9493 8517 9505 8551
rect 9539 8548 9551 8551
rect 9582 8548 9588 8560
rect 9539 8520 9588 8548
rect 9539 8517 9551 8520
rect 9493 8511 9551 8517
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 11425 8551 11483 8557
rect 11425 8517 11437 8551
rect 11471 8517 11483 8551
rect 11425 8511 11483 8517
rect 11517 8551 11575 8557
rect 11517 8517 11529 8551
rect 11563 8548 11575 8551
rect 12526 8548 12532 8560
rect 11563 8520 12532 8548
rect 11563 8517 11575 8520
rect 11517 8511 11575 8517
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 8110 8480 8116 8492
rect 7515 8452 8116 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 1596 8344 1624 8375
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 2004 8384 3157 8412
rect 2004 8372 2010 8384
rect 3145 8381 3157 8384
rect 3191 8381 3203 8415
rect 7300 8412 7328 8443
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9732 8452 10057 8480
rect 9732 8440 9738 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 3145 8375 3203 8381
rect 3344 8384 7328 8412
rect 3344 8344 3372 8384
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 7800 8384 8217 8412
rect 7800 8372 7806 8384
rect 8205 8381 8217 8384
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 11440 8412 11468 8511
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 14185 8551 14243 8557
rect 14185 8517 14197 8551
rect 14231 8517 14243 8551
rect 14185 8511 14243 8517
rect 14461 8551 14519 8557
rect 14461 8517 14473 8551
rect 14507 8548 14519 8551
rect 15562 8548 15568 8560
rect 14507 8520 15568 8548
rect 14507 8517 14519 8520
rect 14461 8511 14519 8517
rect 12066 8480 12072 8492
rect 12027 8452 12072 8480
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12710 8440 12716 8492
rect 12768 8480 12774 8492
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 12768 8452 12817 8480
rect 12768 8440 12774 8452
rect 12805 8449 12817 8452
rect 12851 8449 12863 8483
rect 14200 8480 14228 8511
rect 15562 8508 15568 8520
rect 15620 8508 15626 8560
rect 15010 8480 15016 8492
rect 14200 8452 15016 8480
rect 12805 8443 12863 8449
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 9272 8384 11468 8412
rect 11977 8415 12035 8421
rect 9272 8372 9278 8384
rect 11977 8381 11989 8415
rect 12023 8412 12035 8415
rect 12158 8412 12164 8424
rect 12023 8384 12164 8412
rect 12023 8381 12035 8384
rect 11977 8375 12035 8381
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 12462 8415 12520 8421
rect 12462 8381 12474 8415
rect 12508 8412 12520 8415
rect 12618 8412 12624 8424
rect 12508 8384 12624 8412
rect 12508 8381 12520 8384
rect 12462 8375 12520 8381
rect 12618 8372 12624 8384
rect 12676 8412 12682 8424
rect 13072 8415 13130 8421
rect 12676 8384 13032 8412
rect 12676 8372 12682 8384
rect 3418 8353 3424 8356
rect 1596 8316 3372 8344
rect 3412 8307 3424 8353
rect 3476 8344 3482 8356
rect 3476 8316 3512 8344
rect 3418 8304 3424 8307
rect 3476 8304 3482 8316
rect 3602 8304 3608 8356
rect 3660 8344 3666 8356
rect 4801 8347 4859 8353
rect 4801 8344 4813 8347
rect 3660 8316 4813 8344
rect 3660 8304 3666 8316
rect 4801 8313 4813 8316
rect 4847 8313 4859 8347
rect 4801 8307 4859 8313
rect 6273 8347 6331 8353
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 7098 8344 7104 8356
rect 6319 8316 7104 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 7098 8304 7104 8316
rect 7156 8304 7162 8356
rect 7193 8347 7251 8353
rect 7193 8313 7205 8347
rect 7239 8344 7251 8347
rect 7282 8344 7288 8356
rect 7239 8316 7288 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 7282 8304 7288 8316
rect 7340 8344 7346 8356
rect 7340 8316 7604 8344
rect 7340 8304 7346 8316
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 2501 8279 2559 8285
rect 2501 8276 2513 8279
rect 2464 8248 2513 8276
rect 2464 8236 2470 8248
rect 2501 8245 2513 8248
rect 2547 8245 2559 8279
rect 2501 8239 2559 8245
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 2648 8248 2693 8276
rect 2648 8236 2654 8248
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 5074 8276 5080 8288
rect 3108 8248 5080 8276
rect 3108 8236 3114 8248
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5258 8276 5264 8288
rect 5219 8248 5264 8276
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 5626 8276 5632 8288
rect 5587 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8236 5690 8288
rect 5721 8279 5779 8285
rect 5721 8245 5733 8279
rect 5767 8276 5779 8279
rect 6730 8276 6736 8288
rect 5767 8248 6736 8276
rect 5767 8245 5779 8248
rect 5721 8239 5779 8245
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 6825 8279 6883 8285
rect 6825 8245 6837 8279
rect 6871 8276 6883 8279
rect 7374 8276 7380 8288
rect 6871 8248 7380 8276
rect 6871 8245 6883 8248
rect 6825 8239 6883 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7576 8276 7604 8316
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 9122 8344 9128 8356
rect 8996 8316 9128 8344
rect 8996 8304 9002 8316
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 10290 8347 10348 8353
rect 10290 8344 10302 8347
rect 9364 8316 10302 8344
rect 9364 8304 9370 8316
rect 10290 8313 10302 8316
rect 10336 8313 10348 8347
rect 10290 8307 10348 8313
rect 11885 8347 11943 8353
rect 11885 8313 11897 8347
rect 11931 8344 11943 8347
rect 12894 8344 12900 8356
rect 11931 8316 12900 8344
rect 11931 8313 11943 8316
rect 11885 8307 11943 8313
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 13004 8344 13032 8384
rect 13072 8381 13084 8415
rect 13118 8412 13130 8415
rect 13446 8412 13452 8424
rect 13118 8384 13452 8412
rect 13118 8381 13130 8384
rect 13072 8375 13130 8381
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8412 14887 8415
rect 14918 8412 14924 8424
rect 14875 8384 14924 8412
rect 14875 8381 14887 8384
rect 14829 8375 14887 8381
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 15672 8412 15700 8588
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 16025 8483 16083 8489
rect 16025 8480 16037 8483
rect 15896 8452 16037 8480
rect 15896 8440 15902 8452
rect 16025 8449 16037 8452
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 15933 8415 15991 8421
rect 15672 8384 15884 8412
rect 13354 8344 13360 8356
rect 13004 8316 13360 8344
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 15286 8344 15292 8356
rect 14936 8316 15292 8344
rect 12066 8276 12072 8288
rect 7576 8248 12072 8276
rect 12066 8236 12072 8248
rect 12124 8236 12130 8288
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 13262 8276 13268 8288
rect 12768 8248 13268 8276
rect 12768 8236 12774 8248
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 14936 8285 14964 8316
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15856 8353 15884 8384
rect 15933 8381 15945 8415
rect 15979 8412 15991 8415
rect 16206 8412 16212 8424
rect 15979 8384 16212 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 15841 8347 15899 8353
rect 15841 8313 15853 8347
rect 15887 8313 15899 8347
rect 15841 8307 15899 8313
rect 14921 8279 14979 8285
rect 14921 8245 14933 8279
rect 14967 8245 14979 8279
rect 15470 8276 15476 8288
rect 15431 8248 15476 8276
rect 14921 8239 14979 8245
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 1104 8186 16836 8208
rect 1104 8134 6246 8186
rect 6298 8134 6310 8186
rect 6362 8134 6374 8186
rect 6426 8134 6438 8186
rect 6490 8134 11510 8186
rect 11562 8134 11574 8186
rect 11626 8134 11638 8186
rect 11690 8134 11702 8186
rect 11754 8134 16836 8186
rect 1104 8112 16836 8134
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 3329 8075 3387 8081
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 5258 8072 5264 8084
rect 3375 8044 5264 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 2976 8004 3004 8035
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 5684 8044 6745 8072
rect 5684 8032 5690 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 6733 8035 6791 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 8294 8072 8300 8084
rect 7883 8044 8300 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8628 8044 9045 8072
rect 8628 8032 8634 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9582 8072 9588 8084
rect 9456 8044 9588 8072
rect 9456 8032 9462 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10502 8072 10508 8084
rect 9876 8044 10508 8072
rect 4338 8013 4344 8016
rect 4332 8004 4344 8013
rect 2976 7976 4200 8004
rect 4299 7976 4344 8004
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2314 7936 2320 7948
rect 2275 7908 2320 7936
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 3421 7939 3479 7945
rect 3421 7905 3433 7939
rect 3467 7936 3479 7939
rect 3510 7936 3516 7948
rect 3467 7908 3516 7936
rect 3467 7905 3479 7908
rect 3421 7899 3479 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 4172 7936 4200 7976
rect 4332 7967 4344 7976
rect 4338 7964 4344 7967
rect 4396 7964 4402 8016
rect 5718 7964 5724 8016
rect 5776 8004 5782 8016
rect 6089 8007 6147 8013
rect 6089 8004 6101 8007
rect 5776 7976 6101 8004
rect 5776 7964 5782 7976
rect 6089 7973 6101 7976
rect 6135 7973 6147 8007
rect 6089 7967 6147 7973
rect 7193 8007 7251 8013
rect 7193 7973 7205 8007
rect 7239 8004 7251 8007
rect 8386 8004 8392 8016
rect 7239 7976 8392 8004
rect 7239 7973 7251 7976
rect 7193 7967 7251 7973
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 9125 8007 9183 8013
rect 9125 8004 9137 8007
rect 8812 7976 9137 8004
rect 8812 7964 8818 7976
rect 9125 7973 9137 7976
rect 9171 7973 9183 8007
rect 9125 7967 9183 7973
rect 5902 7936 5908 7948
rect 4172 7908 5908 7936
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 8205 7939 8263 7945
rect 6288 7908 7328 7936
rect 6288 7880 6316 7908
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 2280 7840 2421 7868
rect 2280 7828 2286 7840
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2590 7868 2596 7880
rect 2551 7840 2596 7868
rect 2409 7831 2467 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 4062 7868 4068 7880
rect 3651 7840 3924 7868
rect 4023 7840 4068 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 2774 7800 2780 7812
rect 1627 7772 2780 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 2774 7760 2780 7772
rect 2832 7760 2838 7812
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 3896 7732 3924 7840
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6178 7868 6184 7880
rect 6052 7840 6184 7868
rect 6052 7828 6058 7840
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6270 7828 6276 7880
rect 6328 7868 6334 7880
rect 7300 7877 7328 7908
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 9766 7936 9772 7948
rect 8251 7908 9772 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 9876 7945 9904 8044
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10962 8072 10968 8084
rect 10836 8044 10968 8072
rect 10836 8032 10842 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11793 8075 11851 8081
rect 11793 8041 11805 8075
rect 11839 8072 11851 8075
rect 11974 8072 11980 8084
rect 11839 8044 11980 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 13449 8075 13507 8081
rect 13449 8072 13461 8075
rect 12115 8044 13461 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 13449 8041 13461 8044
rect 13495 8041 13507 8075
rect 13449 8035 13507 8041
rect 14093 8075 14151 8081
rect 14093 8041 14105 8075
rect 14139 8072 14151 8075
rect 15749 8075 15807 8081
rect 15749 8072 15761 8075
rect 14139 8044 15761 8072
rect 14139 8041 14151 8044
rect 14093 8035 14151 8041
rect 15749 8041 15761 8044
rect 15795 8041 15807 8075
rect 15749 8035 15807 8041
rect 12529 8007 12587 8013
rect 10244 7976 11836 8004
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 7285 7871 7343 7877
rect 6328 7840 6373 7868
rect 6328 7828 6334 7840
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 8076 7840 8309 7868
rect 8076 7828 8082 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 8110 7800 8116 7812
rect 5132 7772 8116 7800
rect 5132 7760 5138 7772
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8202 7760 8208 7812
rect 8260 7800 8266 7812
rect 8404 7800 8432 7831
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8938 7868 8944 7880
rect 8536 7840 8944 7868
rect 8536 7828 8542 7840
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9306 7868 9312 7880
rect 9267 7840 9312 7868
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 10244 7800 10272 7976
rect 11808 7948 11836 7976
rect 12529 7973 12541 8007
rect 12575 8004 12587 8007
rect 12618 8004 12624 8016
rect 12575 7976 12624 8004
rect 12575 7973 12587 7976
rect 12529 7967 12587 7973
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 14461 8007 14519 8013
rect 14461 8004 14473 8007
rect 12768 7976 14473 8004
rect 12768 7964 12774 7976
rect 14461 7973 14473 7976
rect 14507 8004 14519 8007
rect 14642 8004 14648 8016
rect 14507 7976 14648 8004
rect 14507 7973 14519 7976
rect 14461 7967 14519 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 10680 7939 10738 7945
rect 10680 7905 10692 7939
rect 10726 7936 10738 7939
rect 11698 7936 11704 7948
rect 10726 7908 11704 7936
rect 10726 7905 10738 7908
rect 10680 7899 10738 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 11790 7896 11796 7948
rect 11848 7896 11854 7948
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 13262 7936 13268 7948
rect 12483 7908 13268 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 13262 7896 13268 7908
rect 13320 7896 13326 7948
rect 15654 7936 15660 7948
rect 15615 7908 15660 7936
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10376 7840 10425 7868
rect 10376 7828 10382 7840
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7868 12679 7871
rect 13354 7868 13360 7880
rect 12667 7840 13360 7868
rect 12667 7837 12679 7840
rect 12621 7831 12679 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 8260 7772 8432 7800
rect 8496 7772 10272 7800
rect 11716 7772 12204 7800
rect 8260 7760 8266 7772
rect 4430 7732 4436 7744
rect 3896 7704 4436 7732
rect 4430 7692 4436 7704
rect 4488 7732 4494 7744
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 4488 7704 5457 7732
rect 4488 7692 4494 7704
rect 5445 7701 5457 7704
rect 5491 7701 5503 7735
rect 5718 7732 5724 7744
rect 5679 7704 5724 7732
rect 5445 7695 5503 7701
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 8496 7732 8524 7772
rect 6236 7704 8524 7732
rect 8665 7735 8723 7741
rect 6236 7692 6242 7704
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 9490 7732 9496 7744
rect 8711 7704 9496 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10045 7735 10103 7741
rect 10045 7701 10057 7735
rect 10091 7732 10103 7735
rect 11716 7732 11744 7772
rect 10091 7704 11744 7732
rect 12176 7732 12204 7772
rect 12894 7760 12900 7812
rect 12952 7800 12958 7812
rect 13081 7803 13139 7809
rect 13081 7800 13093 7803
rect 12952 7772 13093 7800
rect 12952 7760 12958 7772
rect 13081 7769 13093 7772
rect 13127 7769 13139 7803
rect 13081 7763 13139 7769
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 13648 7800 13676 7831
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 14516 7840 14565 7868
rect 14516 7828 14522 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7868 14795 7871
rect 15010 7868 15016 7880
rect 14783 7840 15016 7868
rect 14783 7837 14795 7840
rect 14737 7831 14795 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15838 7868 15844 7880
rect 15799 7840 15844 7868
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 13228 7772 13676 7800
rect 13228 7760 13234 7772
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14826 7800 14832 7812
rect 13780 7772 14832 7800
rect 13780 7760 13786 7772
rect 14826 7760 14832 7772
rect 14884 7760 14890 7812
rect 14918 7732 14924 7744
rect 12176 7704 14924 7732
rect 10091 7701 10103 7704
rect 10045 7695 10103 7701
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15289 7735 15347 7741
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 15746 7732 15752 7744
rect 15335 7704 15752 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 1104 7642 16836 7664
rect 1104 7590 3614 7642
rect 3666 7590 3678 7642
rect 3730 7590 3742 7642
rect 3794 7590 3806 7642
rect 3858 7590 8878 7642
rect 8930 7590 8942 7642
rect 8994 7590 9006 7642
rect 9058 7590 9070 7642
rect 9122 7590 14142 7642
rect 14194 7590 14206 7642
rect 14258 7590 14270 7642
rect 14322 7590 14334 7642
rect 14386 7590 16836 7642
rect 1104 7568 16836 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 3568 7500 4200 7528
rect 3568 7488 3574 7500
rect 4172 7460 4200 7500
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4396 7500 4629 7528
rect 4396 7488 4402 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 4617 7491 4675 7497
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6788 7500 6837 7528
rect 6788 7488 6794 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 12342 7528 12348 7540
rect 8343 7500 12348 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 13538 7528 13544 7540
rect 12483 7500 13544 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 14001 7531 14059 7537
rect 14001 7497 14013 7531
rect 14047 7528 14059 7531
rect 14642 7528 14648 7540
rect 14047 7500 14648 7528
rect 14047 7497 14059 7500
rect 14001 7491 14059 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 16206 7528 16212 7540
rect 16167 7500 16212 7528
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 7929 7463 7987 7469
rect 7929 7460 7941 7463
rect 4172 7432 7941 7460
rect 7929 7429 7941 7432
rect 7975 7429 7987 7463
rect 10042 7460 10048 7472
rect 10003 7432 10048 7460
rect 7929 7423 7987 7429
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 11698 7460 11704 7472
rect 11659 7432 11704 7460
rect 11698 7420 11704 7432
rect 11756 7460 11762 7472
rect 13170 7460 13176 7472
rect 11756 7432 13176 7460
rect 11756 7420 11762 7432
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 13722 7420 13728 7472
rect 13780 7460 13786 7472
rect 13780 7432 14412 7460
rect 13780 7420 13786 7432
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2464 7364 2789 7392
rect 2464 7352 2470 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 2777 7355 2835 7361
rect 5368 7364 5641 7392
rect 1578 7324 1584 7336
rect 1539 7296 1584 7324
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 2222 7284 2228 7336
rect 2280 7324 2286 7336
rect 3237 7327 3295 7333
rect 3237 7324 3249 7327
rect 2280 7296 3249 7324
rect 2280 7284 2286 7296
rect 3237 7293 3249 7296
rect 3283 7293 3295 7327
rect 3237 7287 3295 7293
rect 3504 7327 3562 7333
rect 3504 7293 3516 7327
rect 3550 7324 3562 7327
rect 5368 7324 5396 7364
rect 5629 7361 5641 7364
rect 5675 7392 5687 7395
rect 6270 7392 6276 7404
rect 5675 7364 6276 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6270 7352 6276 7364
rect 6328 7392 6334 7404
rect 6730 7392 6736 7404
rect 6328 7364 6736 7392
rect 6328 7352 6334 7364
rect 6730 7352 6736 7364
rect 6788 7392 6794 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6788 7364 7389 7392
rect 6788 7352 6794 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12860 7364 12909 7392
rect 12860 7352 12866 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13354 7392 13360 7404
rect 13127 7364 13360 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13354 7352 13360 7364
rect 13412 7392 13418 7404
rect 13538 7392 13544 7404
rect 13412 7364 13544 7392
rect 13412 7352 13418 7364
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 14384 7401 14412 7432
rect 14369 7395 14427 7401
rect 14369 7361 14381 7395
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 3550 7296 5396 7324
rect 3550 7293 3562 7296
rect 3504 7287 3562 7293
rect 1394 7216 1400 7268
rect 1452 7256 1458 7268
rect 2685 7259 2743 7265
rect 2685 7256 2697 7259
rect 1452 7228 2697 7256
rect 1452 7216 1458 7228
rect 2685 7225 2697 7228
rect 2731 7256 2743 7259
rect 3050 7256 3056 7268
rect 2731 7228 3056 7256
rect 2731 7225 2743 7228
rect 2685 7219 2743 7225
rect 3050 7216 3056 7228
rect 3108 7216 3114 7268
rect 3252 7256 3280 7287
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 5500 7296 5549 7324
rect 5500 7284 5506 7296
rect 5537 7293 5549 7296
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7324 6147 7327
rect 6178 7324 6184 7336
rect 6135 7296 6184 7324
rect 6135 7293 6147 7296
rect 6089 7287 6147 7293
rect 4062 7256 4068 7268
rect 3252 7228 4068 7256
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 4246 7216 4252 7268
rect 4304 7256 4310 7268
rect 6104 7256 6132 7287
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 6972 7296 7205 7324
rect 6972 7284 6978 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 7193 7287 7251 7293
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7324 7803 7327
rect 8018 7324 8024 7336
rect 7791 7296 8024 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 4304 7228 6132 7256
rect 7208 7256 7236 7287
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7324 8723 7327
rect 10318 7324 10324 7336
rect 8711 7296 10324 7324
rect 8711 7293 8723 7296
rect 8665 7287 8723 7293
rect 8128 7256 8156 7287
rect 10318 7284 10324 7296
rect 10376 7284 10382 7336
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 10428 7296 12173 7324
rect 7208 7228 8156 7256
rect 4304 7216 4310 7228
rect 750 7148 756 7200
rect 808 7188 814 7200
rect 1765 7191 1823 7197
rect 1765 7188 1777 7191
rect 808 7160 1777 7188
rect 808 7148 814 7160
rect 1765 7157 1777 7160
rect 1811 7157 1823 7191
rect 1765 7151 1823 7157
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7188 2651 7191
rect 3234 7188 3240 7200
rect 2639 7160 3240 7188
rect 2639 7157 2651 7160
rect 2593 7151 2651 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 4522 7188 4528 7200
rect 3568 7160 4528 7188
rect 3568 7148 3574 7160
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 5074 7188 5080 7200
rect 5035 7160 5080 7188
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 5316 7160 5457 7188
rect 5316 7148 5322 7160
rect 5445 7157 5457 7160
rect 5491 7157 5503 7191
rect 5445 7151 5503 7157
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 6273 7191 6331 7197
rect 6273 7188 6285 7191
rect 6052 7160 6285 7188
rect 6052 7148 6058 7160
rect 6273 7157 6285 7160
rect 6319 7157 6331 7191
rect 6273 7151 6331 7157
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7374 7188 7380 7200
rect 7331 7160 7380 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7374 7148 7380 7160
rect 7432 7188 7438 7200
rect 7558 7188 7564 7200
rect 7432 7160 7564 7188
rect 7432 7148 7438 7160
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 8128 7188 8156 7228
rect 8932 7259 8990 7265
rect 8932 7225 8944 7259
rect 8978 7256 8990 7259
rect 9214 7256 9220 7268
rect 8978 7228 9220 7256
rect 8978 7225 8990 7228
rect 8932 7219 8990 7225
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 10428 7256 10456 7296
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 13814 7324 13820 7336
rect 13775 7296 13820 7324
rect 12161 7287 12219 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 14636 7327 14694 7333
rect 14636 7324 14648 7327
rect 14516 7296 14648 7324
rect 14516 7284 14522 7296
rect 14636 7293 14648 7296
rect 14682 7324 14694 7327
rect 15010 7324 15016 7336
rect 14682 7296 15016 7324
rect 14682 7293 14694 7296
rect 14636 7287 14694 7293
rect 15010 7284 15016 7296
rect 15068 7284 15074 7336
rect 16022 7324 16028 7336
rect 15983 7296 16028 7324
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 9456 7228 10456 7256
rect 10588 7259 10646 7265
rect 9456 7216 9462 7228
rect 10588 7225 10600 7259
rect 10634 7256 10646 7259
rect 10778 7256 10784 7268
rect 10634 7228 10784 7256
rect 10634 7225 10646 7228
rect 10588 7219 10646 7225
rect 10778 7216 10784 7228
rect 10836 7216 10842 7268
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 13998 7256 14004 7268
rect 11020 7228 14004 7256
rect 11020 7216 11026 7228
rect 13998 7216 14004 7228
rect 14056 7216 14062 7268
rect 10502 7188 10508 7200
rect 8128 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11977 7191 12035 7197
rect 11977 7188 11989 7191
rect 11204 7160 11989 7188
rect 11204 7148 11210 7160
rect 11977 7157 11989 7160
rect 12023 7188 12035 7191
rect 12066 7188 12072 7200
rect 12023 7160 12072 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 13630 7188 13636 7200
rect 12851 7160 13636 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13630 7148 13636 7160
rect 13688 7188 13694 7200
rect 14274 7188 14280 7200
rect 13688 7160 14280 7188
rect 13688 7148 13694 7160
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 15838 7188 15844 7200
rect 15795 7160 15844 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 1104 7098 16836 7120
rect 1104 7046 6246 7098
rect 6298 7046 6310 7098
rect 6362 7046 6374 7098
rect 6426 7046 6438 7098
rect 6490 7046 11510 7098
rect 11562 7046 11574 7098
rect 11626 7046 11638 7098
rect 11690 7046 11702 7098
rect 11754 7046 16836 7098
rect 1104 7024 16836 7046
rect 1949 6987 2007 6993
rect 1949 6953 1961 6987
rect 1995 6984 2007 6987
rect 2314 6984 2320 6996
rect 1995 6956 2320 6984
rect 1995 6953 2007 6956
rect 1949 6947 2007 6953
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 3329 6987 3387 6993
rect 3329 6984 3341 6987
rect 3292 6956 3341 6984
rect 3292 6944 3298 6956
rect 3329 6953 3341 6956
rect 3375 6953 3387 6987
rect 3329 6947 3387 6953
rect 3421 6987 3479 6993
rect 3421 6953 3433 6987
rect 3467 6984 3479 6987
rect 3467 6956 3740 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 2498 6916 2504 6928
rect 2332 6888 2504 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1762 6848 1768 6860
rect 1443 6820 1768 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2332 6857 2360 6888
rect 2498 6876 2504 6888
rect 2556 6876 2562 6928
rect 3712 6916 3740 6956
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 4341 6987 4399 6993
rect 4341 6984 4353 6987
rect 4212 6956 4353 6984
rect 4212 6944 4218 6956
rect 4341 6953 4353 6956
rect 4387 6953 4399 6987
rect 4706 6984 4712 6996
rect 4667 6956 4712 6984
rect 4341 6947 4399 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 4801 6987 4859 6993
rect 4801 6953 4813 6987
rect 4847 6984 4859 6987
rect 5074 6984 5080 6996
rect 4847 6956 5080 6984
rect 4847 6953 4859 6956
rect 4801 6947 4859 6953
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 6730 6984 6736 6996
rect 6691 6956 6736 6984
rect 6730 6944 6736 6956
rect 6788 6944 6794 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 8110 6984 8116 6996
rect 7340 6956 8116 6984
rect 7340 6944 7346 6956
rect 8110 6944 8116 6956
rect 8168 6984 8174 6996
rect 10042 6984 10048 6996
rect 8168 6956 10048 6984
rect 8168 6944 8174 6956
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10505 6987 10563 6993
rect 10505 6953 10517 6987
rect 10551 6984 10563 6987
rect 10686 6984 10692 6996
rect 10551 6956 10692 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 11517 6987 11575 6993
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 11882 6984 11888 6996
rect 11563 6956 11888 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 11882 6944 11888 6956
rect 11940 6984 11946 6996
rect 13906 6984 13912 6996
rect 11940 6956 13912 6984
rect 11940 6944 11946 6956
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 14274 6944 14280 6996
rect 14332 6984 14338 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 14332 6956 15669 6984
rect 14332 6944 14338 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 15657 6947 15715 6953
rect 4246 6916 4252 6928
rect 3712 6888 4252 6916
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 5626 6925 5632 6928
rect 5620 6916 5632 6925
rect 5587 6888 5632 6916
rect 5620 6879 5632 6888
rect 5626 6876 5632 6879
rect 5684 6876 5690 6928
rect 6822 6876 6828 6928
rect 6880 6916 6886 6928
rect 6880 6888 7420 6916
rect 6880 6876 6886 6888
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2682 6848 2688 6860
rect 2455 6820 2688 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6848 5411 6851
rect 6914 6848 6920 6860
rect 5399 6820 6920 6848
rect 5399 6817 5411 6820
rect 5353 6811 5411 6817
rect 6914 6808 6920 6820
rect 6972 6848 6978 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 6972 6820 7021 6848
rect 6972 6808 6978 6820
rect 7009 6817 7021 6820
rect 7055 6848 7067 6851
rect 7098 6848 7104 6860
rect 7055 6820 7104 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 7282 6857 7288 6860
rect 7276 6848 7288 6857
rect 7243 6820 7288 6848
rect 7276 6811 7288 6820
rect 7282 6808 7288 6811
rect 7340 6808 7346 6860
rect 7392 6848 7420 6888
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 10594 6916 10600 6928
rect 7616 6888 10600 6916
rect 7616 6876 7622 6888
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 11974 6876 11980 6928
rect 12032 6916 12038 6928
rect 16022 6916 16028 6928
rect 12032 6888 16028 6916
rect 12032 6876 12038 6888
rect 16022 6876 16028 6888
rect 16080 6876 16086 6928
rect 8849 6851 8907 6857
rect 8849 6848 8861 6851
rect 7392 6820 8861 6848
rect 8849 6817 8861 6820
rect 8895 6817 8907 6851
rect 8849 6811 8907 6817
rect 9033 6851 9091 6857
rect 9033 6817 9045 6851
rect 9079 6848 9091 6851
rect 9582 6848 9588 6860
rect 9079 6820 9588 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 9916 6820 11621 6848
rect 9916 6808 9922 6820
rect 11609 6817 11621 6820
rect 11655 6848 11667 6851
rect 11790 6848 11796 6860
rect 11655 6820 11796 6848
rect 11655 6817 11667 6820
rect 11609 6811 11667 6817
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 12529 6851 12587 6857
rect 12529 6817 12541 6851
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 2498 6780 2504 6792
rect 2459 6752 2504 6780
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 4246 6780 4252 6792
rect 3651 6752 4252 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4396 6752 4905 6780
rect 4396 6740 4402 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 9674 6780 9680 6792
rect 9635 6752 9680 6780
rect 4893 6743 4951 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10778 6780 10784 6792
rect 10739 6752 10784 6780
rect 10597 6743 10655 6749
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 3050 6712 3056 6724
rect 1627 6684 2176 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2148 6644 2176 6684
rect 2884 6684 3056 6712
rect 2884 6644 2912 6684
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 8662 6712 8668 6724
rect 8623 6684 8668 6712
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 10612 6712 10640 6743
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 12544 6780 12572 6811
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 12952 6820 13277 6848
rect 12952 6808 12958 6820
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 13412 6820 14197 6848
rect 13412 6808 13418 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 14366 6808 14372 6860
rect 14424 6848 14430 6860
rect 14918 6848 14924 6860
rect 14424 6820 14924 6848
rect 14424 6808 14430 6820
rect 14918 6808 14924 6820
rect 14976 6808 14982 6860
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15749 6851 15807 6857
rect 15749 6848 15761 6851
rect 15620 6820 15761 6848
rect 15620 6808 15626 6820
rect 15749 6817 15761 6820
rect 15795 6817 15807 6851
rect 15749 6811 15807 6817
rect 11808 6752 12572 6780
rect 12621 6783 12679 6789
rect 11149 6715 11207 6721
rect 11149 6712 11161 6715
rect 10612 6684 11161 6712
rect 11149 6681 11161 6684
rect 11195 6681 11207 6715
rect 11149 6675 11207 6681
rect 2148 6616 2912 6644
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 6546 6644 6552 6656
rect 3007 6616 6552 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 7248 6616 8401 6644
rect 7248 6604 7254 6616
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 9214 6644 9220 6656
rect 9175 6616 9220 6644
rect 8389 6607 8447 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 10137 6647 10195 6653
rect 10137 6613 10149 6647
rect 10183 6644 10195 6647
rect 11808 6644 11836 6752
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6780 12863 6783
rect 13170 6780 13176 6792
rect 12851 6752 13176 6780
rect 12851 6749 12863 6752
rect 12805 6743 12863 6749
rect 12158 6712 12164 6724
rect 12119 6684 12164 6712
rect 12158 6672 12164 6684
rect 12216 6672 12222 6724
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 12636 6712 12664 6743
rect 13170 6740 13176 6752
rect 13228 6740 13234 6792
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 14056 6752 14289 6780
rect 14056 6740 14062 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14458 6780 14464 6792
rect 14419 6752 14464 6780
rect 14277 6743 14335 6749
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 15838 6780 15844 6792
rect 15799 6752 15844 6780
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 12400 6684 12664 6712
rect 13817 6715 13875 6721
rect 12400 6672 12406 6684
rect 13817 6681 13829 6715
rect 13863 6712 13875 6715
rect 15654 6712 15660 6724
rect 13863 6684 15660 6712
rect 13863 6681 13875 6684
rect 13817 6675 13875 6681
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 10183 6616 11836 6644
rect 13449 6647 13507 6653
rect 10183 6613 10195 6616
rect 10137 6607 10195 6613
rect 13449 6613 13461 6647
rect 13495 6644 13507 6647
rect 15010 6644 15016 6656
rect 13495 6616 15016 6644
rect 13495 6613 13507 6616
rect 13449 6607 13507 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 15286 6644 15292 6656
rect 15247 6616 15292 6644
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 1104 6554 16836 6576
rect 1104 6502 3614 6554
rect 3666 6502 3678 6554
rect 3730 6502 3742 6554
rect 3794 6502 3806 6554
rect 3858 6502 8878 6554
rect 8930 6502 8942 6554
rect 8994 6502 9006 6554
rect 9058 6502 9070 6554
rect 9122 6502 14142 6554
rect 14194 6502 14206 6554
rect 14258 6502 14270 6554
rect 14322 6502 14334 6554
rect 14386 6502 16836 6554
rect 1104 6480 16836 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3142 6440 3148 6452
rect 2556 6412 3148 6440
rect 2556 6400 2562 6412
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 4522 6440 4528 6452
rect 4028 6412 4528 6440
rect 4028 6400 4034 6412
rect 4522 6400 4528 6412
rect 4580 6440 4586 6452
rect 5442 6440 5448 6452
rect 4580 6412 4844 6440
rect 5403 6412 5448 6440
rect 4580 6400 4586 6412
rect 4816 6304 4844 6412
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 6273 6443 6331 6449
rect 6273 6409 6285 6443
rect 6319 6440 6331 6443
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 6319 6412 8769 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 8757 6403 8815 6409
rect 8864 6412 10057 6440
rect 5626 6332 5632 6384
rect 5684 6372 5690 6384
rect 5684 6344 6040 6372
rect 5684 6332 5690 6344
rect 5718 6304 5724 6316
rect 4816 6276 5724 6304
rect 5718 6264 5724 6276
rect 5776 6304 5782 6316
rect 6012 6313 6040 6344
rect 6086 6332 6092 6384
rect 6144 6372 6150 6384
rect 6457 6375 6515 6381
rect 6457 6372 6469 6375
rect 6144 6344 6469 6372
rect 6144 6332 6150 6344
rect 6457 6341 6469 6344
rect 6503 6372 6515 6375
rect 6822 6372 6828 6384
rect 6503 6344 6828 6372
rect 6503 6341 6515 6344
rect 6457 6335 6515 6341
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 8386 6372 8392 6384
rect 8299 6344 8392 6372
rect 8386 6332 8392 6344
rect 8444 6372 8450 6384
rect 8864 6372 8892 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 10137 6443 10195 6449
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 12342 6440 12348 6452
rect 10183 6412 12348 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 12492 6412 15976 6440
rect 12492 6400 12498 6412
rect 8444 6344 8892 6372
rect 8444 6332 8450 6344
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 12529 6375 12587 6381
rect 12529 6372 12541 6375
rect 9272 6344 12541 6372
rect 9272 6332 9278 6344
rect 12529 6341 12541 6344
rect 12575 6341 12587 6375
rect 12529 6335 12587 6341
rect 12618 6332 12624 6384
rect 12676 6332 12682 6384
rect 5905 6307 5963 6313
rect 5905 6304 5917 6307
rect 5776 6276 5917 6304
rect 5776 6264 5782 6276
rect 5905 6273 5917 6276
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 6914 6304 6920 6316
rect 6875 6276 6920 6304
rect 5997 6267 6055 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6236 1547 6239
rect 2314 6236 2320 6248
rect 1535 6208 2320 6236
rect 1535 6205 1547 6208
rect 1489 6199 1547 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 3142 6236 3148 6248
rect 3103 6208 3148 6236
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 1756 6171 1814 6177
rect 1756 6137 1768 6171
rect 1802 6168 1814 6171
rect 2406 6168 2412 6180
rect 1802 6140 2412 6168
rect 1802 6137 1814 6140
rect 1756 6131 1814 6137
rect 2406 6128 2412 6140
rect 2464 6128 2470 6180
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2648 6072 2881 6100
rect 2648 6060 2654 6072
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 2869 6063 2927 6069
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3329 6103 3387 6109
rect 3329 6100 3341 6103
rect 3016 6072 3341 6100
rect 3016 6060 3022 6072
rect 3329 6069 3341 6072
rect 3375 6069 3387 6103
rect 3804 6100 3832 6199
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 7190 6245 7196 6248
rect 6273 6239 6331 6245
rect 6273 6236 6285 6239
rect 3936 6208 6285 6236
rect 3936 6196 3942 6208
rect 6273 6205 6285 6208
rect 6319 6205 6331 6239
rect 6273 6199 6331 6205
rect 6641 6239 6699 6245
rect 6641 6205 6653 6239
rect 6687 6205 6699 6239
rect 7184 6236 7196 6245
rect 7151 6208 7196 6236
rect 6641 6199 6699 6205
rect 7184 6199 7196 6208
rect 3970 6128 3976 6180
rect 4028 6177 4034 6180
rect 4028 6171 4092 6177
rect 4028 6137 4046 6171
rect 4080 6137 4092 6171
rect 4028 6131 4092 6137
rect 4028 6128 4034 6131
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 5813 6171 5871 6177
rect 5813 6168 5825 6171
rect 4764 6140 5825 6168
rect 4764 6128 4770 6140
rect 5813 6137 5825 6140
rect 5859 6168 5871 6171
rect 6454 6168 6460 6180
rect 5859 6140 6460 6168
rect 5859 6137 5871 6140
rect 5813 6131 5871 6137
rect 6454 6128 6460 6140
rect 6512 6128 6518 6180
rect 6656 6168 6684 6199
rect 7190 6196 7196 6199
rect 7248 6196 7254 6248
rect 8404 6236 8432 6332
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 9306 6304 9312 6316
rect 8536 6276 9312 6304
rect 8536 6264 8542 6276
rect 9306 6264 9312 6276
rect 9364 6304 9370 6316
rect 9677 6307 9735 6313
rect 9677 6304 9689 6307
rect 9364 6276 9689 6304
rect 9364 6264 9370 6276
rect 9677 6273 9689 6276
rect 9723 6273 9735 6307
rect 10778 6304 10784 6316
rect 10739 6276 10784 6304
rect 9677 6267 9735 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11330 6304 11336 6316
rect 11204 6276 11336 6304
rect 11204 6264 11210 6276
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 12636 6304 12664 6332
rect 12360 6276 12664 6304
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8404 6208 8585 6236
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 8812 6208 11529 6236
rect 8812 6196 8818 6208
rect 11517 6205 11529 6208
rect 11563 6236 11575 6239
rect 12360 6236 12388 6276
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14277 6307 14335 6313
rect 14277 6304 14289 6307
rect 13780 6276 14289 6304
rect 13780 6264 13786 6276
rect 14277 6273 14289 6276
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 11563 6208 12388 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12492 6208 12633 6236
rect 12492 6196 12498 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 13814 6236 13820 6248
rect 12768 6208 13820 6236
rect 12768 6196 12774 6208
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 14544 6239 14602 6245
rect 14544 6205 14556 6239
rect 14590 6236 14602 6239
rect 15838 6236 15844 6248
rect 14590 6208 15844 6236
rect 14590 6205 14602 6208
rect 14544 6199 14602 6205
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 15948 6245 15976 6412
rect 15933 6239 15991 6245
rect 15933 6205 15945 6239
rect 15979 6205 15991 6239
rect 15933 6199 15991 6205
rect 6730 6168 6736 6180
rect 6656 6140 6736 6168
rect 6730 6128 6736 6140
rect 6788 6128 6794 6180
rect 10045 6171 10103 6177
rect 10045 6137 10057 6171
rect 10091 6168 10103 6171
rect 12529 6171 12587 6177
rect 10091 6140 12296 6168
rect 10091 6137 10103 6140
rect 10045 6131 10103 6137
rect 4338 6100 4344 6112
rect 3804 6072 4344 6100
rect 3329 6063 3387 6069
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5718 6100 5724 6112
rect 5215 6072 5724 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8297 6103 8355 6109
rect 8297 6100 8309 6103
rect 8260 6072 8309 6100
rect 8260 6060 8266 6072
rect 8297 6069 8309 6072
rect 8343 6069 8355 6103
rect 8297 6063 8355 6069
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 9125 6103 9183 6109
rect 9125 6100 9137 6103
rect 8444 6072 9137 6100
rect 8444 6060 8450 6072
rect 9125 6069 9137 6072
rect 9171 6069 9183 6103
rect 9125 6063 9183 6069
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 9493 6103 9551 6109
rect 9493 6100 9505 6103
rect 9364 6072 9505 6100
rect 9364 6060 9370 6072
rect 9493 6069 9505 6072
rect 9539 6069 9551 6103
rect 9493 6063 9551 6069
rect 9585 6103 9643 6109
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 9766 6100 9772 6112
rect 9631 6072 9772 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10502 6100 10508 6112
rect 10463 6072 10508 6100
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 10643 6072 11161 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 11330 6060 11336 6112
rect 11388 6100 11394 6112
rect 11609 6103 11667 6109
rect 11609 6100 11621 6103
rect 11388 6072 11621 6100
rect 11388 6060 11394 6072
rect 11609 6069 11621 6072
rect 11655 6069 11667 6103
rect 12268 6100 12296 6140
rect 12529 6137 12541 6171
rect 12575 6168 12587 6171
rect 12888 6171 12946 6177
rect 12575 6140 12756 6168
rect 12575 6137 12587 6140
rect 12529 6131 12587 6137
rect 12618 6100 12624 6112
rect 12268 6072 12624 6100
rect 11609 6063 11667 6069
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 12728 6100 12756 6140
rect 12888 6137 12900 6171
rect 12934 6168 12946 6171
rect 12934 6140 15700 6168
rect 12934 6137 12946 6140
rect 12888 6131 12946 6137
rect 13446 6100 13452 6112
rect 12728 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 15672 6109 15700 6140
rect 14001 6103 14059 6109
rect 14001 6100 14013 6103
rect 13964 6072 14013 6100
rect 13964 6060 13970 6072
rect 14001 6069 14013 6072
rect 14047 6069 14059 6103
rect 14001 6063 14059 6069
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 15838 6100 15844 6112
rect 15703 6072 15844 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 16114 6100 16120 6112
rect 16075 6072 16120 6100
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 1104 6010 16836 6032
rect 1104 5958 6246 6010
rect 6298 5958 6310 6010
rect 6362 5958 6374 6010
rect 6426 5958 6438 6010
rect 6490 5958 11510 6010
rect 11562 5958 11574 6010
rect 11626 5958 11638 6010
rect 11690 5958 11702 6010
rect 11754 5958 16836 6010
rect 1104 5936 16836 5958
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 4120 5868 7297 5896
rect 4120 5856 4126 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 7285 5859 7343 5865
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 9766 5896 9772 5908
rect 7616 5868 9772 5896
rect 7616 5856 7622 5868
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 10597 5899 10655 5905
rect 10597 5896 10609 5899
rect 10560 5868 10609 5896
rect 10560 5856 10566 5868
rect 10597 5865 10609 5868
rect 10643 5865 10655 5899
rect 10597 5859 10655 5865
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 10962 5896 10968 5908
rect 10744 5868 10968 5896
rect 10744 5856 10750 5868
rect 10962 5856 10968 5868
rect 11020 5896 11026 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 11020 5868 11069 5896
rect 11020 5856 11026 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 11146 5856 11152 5908
rect 11204 5856 11210 5908
rect 11517 5899 11575 5905
rect 11517 5865 11529 5899
rect 11563 5896 11575 5899
rect 12434 5896 12440 5908
rect 11563 5868 12440 5896
rect 11563 5865 11575 5868
rect 11517 5859 11575 5865
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 14185 5899 14243 5905
rect 14185 5896 14197 5899
rect 12676 5868 14197 5896
rect 12676 5856 12682 5868
rect 14185 5865 14197 5868
rect 14231 5865 14243 5899
rect 14185 5859 14243 5865
rect 15378 5856 15384 5908
rect 15436 5896 15442 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15436 5868 15761 5896
rect 15436 5856 15442 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 15749 5859 15807 5865
rect 15841 5899 15899 5905
rect 15841 5865 15853 5899
rect 15887 5896 15899 5899
rect 16390 5896 16396 5908
rect 15887 5868 16396 5896
rect 15887 5865 15899 5868
rect 15841 5859 15899 5865
rect 16390 5856 16396 5868
rect 16448 5856 16454 5908
rect 4338 5828 4344 5840
rect 2332 5800 4344 5828
rect 2332 5772 2360 5800
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 4801 5831 4859 5837
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 9674 5828 9680 5840
rect 4847 5800 9680 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 9784 5828 9812 5856
rect 11164 5828 11192 5856
rect 13262 5828 13268 5840
rect 9784 5800 11100 5828
rect 11072 5772 11100 5800
rect 11164 5800 12011 5828
rect 13223 5800 13268 5828
rect 1581 5763 1639 5769
rect 1581 5729 1593 5763
rect 1627 5760 1639 5763
rect 1670 5760 1676 5772
rect 1627 5732 1676 5760
rect 1627 5729 1639 5732
rect 1581 5723 1639 5729
rect 1670 5720 1676 5732
rect 1728 5720 1734 5772
rect 2314 5760 2320 5772
rect 2227 5732 2320 5760
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 2590 5769 2596 5772
rect 2584 5760 2596 5769
rect 2551 5732 2596 5760
rect 2584 5723 2596 5732
rect 2590 5720 2596 5723
rect 2648 5720 2654 5772
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 5718 5769 5724 5772
rect 4304 5732 5028 5760
rect 4304 5720 4310 5732
rect 4890 5692 4896 5704
rect 4851 5664 4896 5692
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 5000 5701 5028 5732
rect 5712 5723 5724 5769
rect 5776 5760 5782 5772
rect 7101 5763 7159 5769
rect 5776 5732 5812 5760
rect 5718 5720 5724 5723
rect 5776 5720 5782 5732
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 7650 5760 7656 5772
rect 7147 5732 7656 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 5442 5692 5448 5704
rect 5403 5664 5448 5692
rect 4985 5655 5043 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 7116 5568 7144 5723
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 8018 5760 8024 5772
rect 7979 5732 8024 5760
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 8665 5763 8723 5769
rect 8665 5729 8677 5763
rect 8711 5729 8723 5763
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 8665 5723 8723 5729
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7248 5664 8125 5692
rect 7248 5652 7254 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8260 5664 8305 5692
rect 8260 5652 8266 5664
rect 7926 5584 7932 5636
rect 7984 5624 7990 5636
rect 8680 5624 8708 5723
rect 10042 5720 10048 5732
rect 10100 5760 10106 5772
rect 10410 5760 10416 5772
rect 10100 5732 10416 5760
rect 10100 5720 10106 5732
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9306 5692 9312 5704
rect 8987 5664 9312 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 10134 5652 10140 5704
rect 10192 5692 10198 5704
rect 10980 5692 11008 5723
rect 11054 5720 11060 5772
rect 11112 5720 11118 5772
rect 11164 5692 11192 5800
rect 11698 5760 11704 5772
rect 11256 5732 11704 5760
rect 11256 5701 11284 5732
rect 11698 5720 11704 5732
rect 11756 5760 11762 5772
rect 11865 5763 11923 5769
rect 11865 5760 11877 5763
rect 11756 5732 11877 5760
rect 11756 5720 11762 5732
rect 11865 5729 11877 5732
rect 11911 5729 11923 5763
rect 11983 5760 12011 5800
rect 13262 5788 13268 5800
rect 13320 5788 13326 5840
rect 13354 5760 13360 5772
rect 11983 5732 13360 5760
rect 11865 5723 11923 5729
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5760 14151 5763
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14139 5732 14749 5760
rect 14139 5729 14151 5732
rect 14093 5723 14151 5729
rect 14737 5729 14749 5732
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 10192 5664 11192 5692
rect 11241 5695 11299 5701
rect 10192 5652 10198 5664
rect 11241 5661 11253 5695
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11388 5664 11529 5692
rect 11388 5652 11394 5664
rect 11517 5661 11529 5664
rect 11563 5692 11575 5695
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11563 5664 11621 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 14458 5692 14464 5704
rect 14415 5664 14464 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 15930 5652 15936 5704
rect 15988 5692 15994 5704
rect 15988 5664 16033 5692
rect 15988 5652 15994 5664
rect 7984 5596 8708 5624
rect 7984 5584 7990 5596
rect 9214 5584 9220 5636
rect 9272 5624 9278 5636
rect 11422 5624 11428 5636
rect 9272 5596 11428 5624
rect 9272 5584 9278 5596
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 12989 5627 13047 5633
rect 12989 5593 13001 5627
rect 13035 5624 13047 5627
rect 13556 5624 13584 5652
rect 13035 5596 13584 5624
rect 13035 5593 13047 5596
rect 12989 5587 13047 5593
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 3234 5516 3240 5568
rect 3292 5556 3298 5568
rect 3697 5559 3755 5565
rect 3697 5556 3709 5559
rect 3292 5528 3709 5556
rect 3292 5516 3298 5528
rect 3697 5525 3709 5528
rect 3743 5556 3755 5559
rect 3970 5556 3976 5568
rect 3743 5528 3976 5556
rect 3743 5525 3755 5528
rect 3697 5519 3755 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 6730 5556 6736 5568
rect 4479 5528 6736 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 6880 5528 6925 5556
rect 6880 5516 6886 5528
rect 7098 5516 7104 5568
rect 7156 5516 7162 5568
rect 7653 5559 7711 5565
rect 7653 5525 7665 5559
rect 7699 5556 7711 5559
rect 9674 5556 9680 5568
rect 7699 5528 9680 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 10229 5559 10287 5565
rect 10229 5525 10241 5559
rect 10275 5556 10287 5559
rect 12342 5556 12348 5568
rect 10275 5528 12348 5556
rect 10275 5525 10287 5528
rect 10229 5519 10287 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 13596 5528 13737 5556
rect 13596 5516 13602 5528
rect 13725 5525 13737 5528
rect 13771 5525 13783 5559
rect 15378 5556 15384 5568
rect 15339 5528 15384 5556
rect 13725 5519 13783 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 1104 5466 16836 5488
rect 1104 5414 3614 5466
rect 3666 5414 3678 5466
rect 3730 5414 3742 5466
rect 3794 5414 3806 5466
rect 3858 5414 8878 5466
rect 8930 5414 8942 5466
rect 8994 5414 9006 5466
rect 9058 5414 9070 5466
rect 9122 5414 14142 5466
rect 14194 5414 14206 5466
rect 14258 5414 14270 5466
rect 14322 5414 14334 5466
rect 14386 5414 16836 5466
rect 1104 5392 16836 5414
rect 1673 5355 1731 5361
rect 1673 5321 1685 5355
rect 1719 5352 1731 5355
rect 4154 5352 4160 5364
rect 1719 5324 4160 5352
rect 1719 5321 1731 5324
rect 1673 5315 1731 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 5626 5352 5632 5364
rect 4264 5324 5488 5352
rect 5587 5324 5632 5352
rect 4264 5284 4292 5324
rect 2056 5256 4292 5284
rect 2056 5157 2084 5256
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2406 5216 2412 5228
rect 2363 5188 2412 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 4246 5216 4252 5228
rect 4207 5188 4252 5216
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 5460 5216 5488 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 8018 5352 8024 5364
rect 6871 5324 8024 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 11698 5352 11704 5364
rect 11659 5324 11704 5352
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 13354 5352 13360 5364
rect 12492 5324 13360 5352
rect 12492 5312 12498 5324
rect 13354 5312 13360 5324
rect 13412 5352 13418 5364
rect 13722 5352 13728 5364
rect 13412 5324 13728 5352
rect 13412 5312 13418 5324
rect 13722 5312 13728 5324
rect 13780 5352 13786 5364
rect 14093 5355 14151 5361
rect 14093 5352 14105 5355
rect 13780 5324 14105 5352
rect 13780 5312 13786 5324
rect 14093 5321 14105 5324
rect 14139 5321 14151 5355
rect 14918 5352 14924 5364
rect 14093 5315 14151 5321
rect 14200 5324 14924 5352
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6914 5284 6920 5296
rect 5592 5256 6920 5284
rect 5592 5244 5598 5256
rect 6914 5244 6920 5256
rect 6972 5284 6978 5296
rect 6972 5256 7880 5284
rect 6972 5244 6978 5256
rect 5460 5188 6500 5216
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3326 5148 3332 5160
rect 3099 5120 3332 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5117 3755 5151
rect 5626 5148 5632 5160
rect 3697 5111 3755 5117
rect 4448 5120 5632 5148
rect 2498 5040 2504 5092
rect 2556 5080 2562 5092
rect 3145 5083 3203 5089
rect 3145 5080 3157 5083
rect 2556 5052 3157 5080
rect 2556 5040 2562 5052
rect 3145 5049 3157 5052
rect 3191 5049 3203 5083
rect 3712 5080 3740 5111
rect 4448 5080 4476 5120
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 5902 5148 5908 5160
rect 5863 5120 5908 5148
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 3712 5052 4476 5080
rect 4516 5083 4574 5089
rect 3145 5043 3203 5049
rect 4516 5049 4528 5083
rect 4562 5080 4574 5083
rect 4798 5080 4804 5092
rect 4562 5052 4804 5080
rect 4562 5049 4574 5052
rect 4516 5043 4574 5049
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 6181 5083 6239 5089
rect 6181 5080 6193 5083
rect 5500 5052 6193 5080
rect 5500 5040 5506 5052
rect 6181 5049 6193 5052
rect 6227 5049 6239 5083
rect 6181 5043 6239 5049
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 2685 5015 2743 5021
rect 2685 5012 2697 5015
rect 2179 4984 2697 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 2685 4981 2697 4984
rect 2731 4981 2743 5015
rect 2685 4975 2743 4981
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 3881 5015 3939 5021
rect 3881 5012 3893 5015
rect 3476 4984 3893 5012
rect 3476 4972 3482 4984
rect 3881 4981 3893 4984
rect 3927 4981 3939 5015
rect 3881 4975 3939 4981
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 5994 5012 6000 5024
rect 4120 4984 6000 5012
rect 4120 4972 4126 4984
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6472 5012 6500 5188
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 7852 5225 7880 5256
rect 11422 5244 11428 5296
rect 11480 5284 11486 5296
rect 14200 5284 14228 5324
rect 14918 5312 14924 5324
rect 14976 5352 14982 5364
rect 14976 5324 15884 5352
rect 14976 5312 14982 5324
rect 11480 5256 14228 5284
rect 11480 5244 11486 5256
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 7340 5188 7389 5216
rect 7340 5176 7346 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 10318 5216 10324 5228
rect 10279 5188 10324 5216
rect 7837 5179 7895 5185
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 13725 5219 13783 5225
rect 13725 5216 13737 5219
rect 12952 5188 13737 5216
rect 12952 5176 12958 5188
rect 13725 5185 13737 5188
rect 13771 5216 13783 5219
rect 13771 5188 13952 5216
rect 13771 5185 13783 5188
rect 13725 5179 13783 5185
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 6788 5120 7205 5148
rect 6788 5108 6794 5120
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 9490 5148 9496 5160
rect 9451 5120 9496 5148
rect 7193 5111 7251 5117
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 10042 5148 10048 5160
rect 9692 5120 10048 5148
rect 6546 5040 6552 5092
rect 6604 5080 6610 5092
rect 7285 5083 7343 5089
rect 7285 5080 7297 5083
rect 6604 5052 7297 5080
rect 6604 5040 6610 5052
rect 7285 5049 7297 5052
rect 7331 5049 7343 5083
rect 7285 5043 7343 5049
rect 8104 5083 8162 5089
rect 8104 5049 8116 5083
rect 8150 5080 8162 5083
rect 8202 5080 8208 5092
rect 8150 5052 8208 5080
rect 8150 5049 8162 5052
rect 8104 5043 8162 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 9692 5080 9720 5120
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 12161 5151 12219 5157
rect 12161 5148 12173 5151
rect 12124 5120 12173 5148
rect 12124 5108 12130 5120
rect 12161 5117 12173 5120
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5148 12495 5151
rect 12526 5148 12532 5160
rect 12483 5120 12532 5148
rect 12483 5117 12495 5120
rect 12437 5111 12495 5117
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 13538 5148 13544 5160
rect 13499 5120 13544 5148
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 8312 5052 9720 5080
rect 9769 5083 9827 5089
rect 8312 5012 8340 5052
rect 9769 5049 9781 5083
rect 9815 5080 9827 5083
rect 9950 5080 9956 5092
rect 9815 5052 9956 5080
rect 9815 5049 9827 5052
rect 9769 5043 9827 5049
rect 9950 5040 9956 5052
rect 10008 5040 10014 5092
rect 10588 5083 10646 5089
rect 10588 5049 10600 5083
rect 10634 5080 10646 5083
rect 12618 5080 12624 5092
rect 10634 5052 12624 5080
rect 10634 5049 10646 5052
rect 10588 5043 10646 5049
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 12713 5083 12771 5089
rect 12713 5049 12725 5083
rect 12759 5080 12771 5083
rect 13722 5080 13728 5092
rect 12759 5052 13728 5080
rect 12759 5049 12771 5052
rect 12713 5043 12771 5049
rect 13722 5040 13728 5052
rect 13780 5040 13786 5092
rect 9214 5012 9220 5024
rect 6472 4984 8340 5012
rect 9175 4984 9220 5012
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 11974 5012 11980 5024
rect 11935 4984 11980 5012
rect 11974 4972 11980 4984
rect 12032 4972 12038 5024
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 13173 5015 13231 5021
rect 13173 5012 13185 5015
rect 12584 4984 13185 5012
rect 12584 4972 12590 4984
rect 13173 4981 13185 4984
rect 13219 4981 13231 5015
rect 13630 5012 13636 5024
rect 13591 4984 13636 5012
rect 13173 4975 13231 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13924 5012 13952 5188
rect 14458 5157 14464 5160
rect 14093 5151 14151 5157
rect 14093 5117 14105 5151
rect 14139 5148 14151 5151
rect 14185 5151 14243 5157
rect 14185 5148 14197 5151
rect 14139 5120 14197 5148
rect 14139 5117 14151 5120
rect 14093 5111 14151 5117
rect 14185 5117 14197 5120
rect 14231 5117 14243 5151
rect 14452 5148 14464 5157
rect 14419 5120 14464 5148
rect 14185 5111 14243 5117
rect 14452 5111 14464 5120
rect 14458 5108 14464 5111
rect 14516 5108 14522 5160
rect 15856 5157 15884 5324
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5117 15899 5151
rect 15841 5111 15899 5117
rect 15010 5040 15016 5092
rect 15068 5080 15074 5092
rect 15068 5052 16068 5080
rect 15068 5040 15074 5052
rect 16040 5021 16068 5052
rect 15565 5015 15623 5021
rect 15565 5012 15577 5015
rect 13924 4984 15577 5012
rect 15565 4981 15577 4984
rect 15611 4981 15623 5015
rect 15565 4975 15623 4981
rect 16025 5015 16083 5021
rect 16025 4981 16037 5015
rect 16071 4981 16083 5015
rect 16025 4975 16083 4981
rect 1104 4922 16836 4944
rect 1104 4870 6246 4922
rect 6298 4870 6310 4922
rect 6362 4870 6374 4922
rect 6426 4870 6438 4922
rect 6490 4870 11510 4922
rect 11562 4870 11574 4922
rect 11626 4870 11638 4922
rect 11690 4870 11702 4922
rect 11754 4870 16836 4922
rect 1104 4848 16836 4870
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 3053 4811 3111 4817
rect 3053 4808 3065 4811
rect 2464 4780 3065 4808
rect 2464 4768 2470 4780
rect 3053 4777 3065 4780
rect 3099 4777 3111 4811
rect 3234 4808 3240 4820
rect 3053 4771 3111 4777
rect 3160 4780 3240 4808
rect 1940 4743 1998 4749
rect 1940 4709 1952 4743
rect 1986 4740 1998 4743
rect 2682 4740 2688 4752
rect 1986 4712 2688 4740
rect 1986 4709 1998 4712
rect 1940 4703 1998 4709
rect 2682 4700 2688 4712
rect 2740 4740 2746 4752
rect 3160 4740 3188 4780
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 6914 4808 6920 4820
rect 6503 4780 6920 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 8941 4811 8999 4817
rect 8941 4777 8953 4811
rect 8987 4808 8999 4811
rect 11882 4808 11888 4820
rect 8987 4780 11888 4808
rect 8987 4777 8999 4780
rect 8941 4771 8999 4777
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 11974 4768 11980 4820
rect 12032 4768 12038 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12676 4780 13093 4808
rect 12676 4768 12682 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 13081 4771 13139 4777
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15344 4780 15669 4808
rect 15344 4768 15350 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 15746 4768 15752 4820
rect 15804 4808 15810 4820
rect 15804 4780 15849 4808
rect 15804 4768 15810 4780
rect 2740 4712 3188 4740
rect 6089 4743 6147 4749
rect 2740 4700 2746 4712
rect 6089 4709 6101 4743
rect 6135 4740 6147 4743
rect 8018 4740 8024 4752
rect 6135 4712 8024 4740
rect 6135 4709 6147 4712
rect 6089 4703 6147 4709
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 8119 4712 9045 4740
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 1673 4675 1731 4681
rect 1673 4672 1685 4675
rect 1452 4644 1685 4672
rect 1452 4632 1458 4644
rect 1673 4641 1685 4644
rect 1719 4672 1731 4675
rect 2314 4672 2320 4684
rect 1719 4644 2320 4672
rect 1719 4641 1731 4644
rect 1673 4635 1731 4641
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2866 4632 2872 4684
rect 2924 4672 2930 4684
rect 3050 4672 3056 4684
rect 2924 4644 3056 4672
rect 2924 4632 2930 4644
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3326 4672 3332 4684
rect 3287 4644 3332 4672
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 4338 4681 4344 4684
rect 4332 4672 4344 4681
rect 4251 4644 4344 4672
rect 4332 4635 4344 4644
rect 4396 4672 4402 4684
rect 5810 4672 5816 4684
rect 4396 4644 5580 4672
rect 5771 4644 5816 4672
rect 4338 4632 4344 4635
rect 4396 4632 4402 4644
rect 4062 4604 4068 4616
rect 4023 4576 4068 4604
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 5552 4604 5580 4644
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 6822 4681 6828 4684
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 6503 4644 6561 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 6549 4641 6561 4644
rect 6595 4641 6607 4675
rect 6816 4672 6828 4681
rect 6549 4635 6607 4641
rect 6656 4644 6828 4672
rect 6656 4604 6684 4644
rect 6816 4635 6828 4644
rect 6822 4632 6828 4635
rect 6880 4632 6886 4684
rect 7098 4632 7104 4684
rect 7156 4672 7162 4684
rect 8119 4672 8147 4712
rect 9033 4709 9045 4712
rect 9079 4709 9091 4743
rect 9033 4703 9091 4709
rect 9214 4700 9220 4752
rect 9272 4740 9278 4752
rect 9922 4743 9980 4749
rect 9922 4740 9934 4743
rect 9272 4712 9934 4740
rect 9272 4700 9278 4712
rect 9922 4709 9934 4712
rect 9968 4709 9980 4743
rect 11992 4740 12020 4768
rect 9922 4703 9980 4709
rect 11532 4712 13584 4740
rect 7156 4644 8147 4672
rect 8389 4675 8447 4681
rect 7156 4632 7162 4644
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 8662 4672 8668 4684
rect 8435 4644 8668 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4672 9735 4675
rect 9766 4672 9772 4684
rect 9723 4644 9772 4672
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 9766 4632 9772 4644
rect 9824 4672 9830 4684
rect 10318 4672 10324 4684
rect 9824 4644 10324 4672
rect 9824 4632 9830 4644
rect 10318 4632 10324 4644
rect 10376 4672 10382 4684
rect 11532 4681 11560 4712
rect 11517 4675 11575 4681
rect 10376 4644 10732 4672
rect 10376 4632 10382 4644
rect 5552 4576 6500 4604
rect 6472 4480 6500 4576
rect 6564 4576 6684 4604
rect 6564 4548 6592 4576
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 9122 4604 9128 4616
rect 8352 4576 9128 4604
rect 8352 4564 8358 4576
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9398 4604 9404 4616
rect 9263 4576 9404 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 6546 4496 6552 4548
rect 6604 4496 6610 4548
rect 8202 4536 8208 4548
rect 8163 4508 8208 4536
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 10704 4536 10732 4644
rect 11517 4641 11529 4675
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 11968 4675 12026 4681
rect 11968 4641 11980 4675
rect 12014 4672 12026 4675
rect 12894 4672 12900 4684
rect 12014 4644 12900 4672
rect 12014 4641 12026 4644
rect 11968 4635 12026 4641
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 13556 4681 13584 4712
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4641 13599 4675
rect 13541 4635 13599 4641
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 14056 4644 14657 4672
rect 14056 4632 14062 4644
rect 14645 4641 14657 4644
rect 14691 4672 14703 4675
rect 14826 4672 14832 4684
rect 14691 4644 14832 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 11330 4564 11336 4616
rect 11388 4604 11394 4616
rect 11701 4607 11759 4613
rect 11701 4604 11713 4607
rect 11388 4576 11713 4604
rect 11388 4564 11394 4576
rect 11701 4573 11713 4576
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13136 4576 14105 4604
rect 13136 4564 13142 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14458 4604 14464 4616
rect 14323 4576 14464 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15838 4604 15844 4616
rect 15799 4576 15844 4604
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 14918 4536 14924 4548
rect 10704 4508 11376 4536
rect 3510 4468 3516 4480
rect 3471 4440 3516 4468
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 4798 4428 4804 4480
rect 4856 4468 4862 4480
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 4856 4440 5457 4468
rect 4856 4428 4862 4440
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 7929 4471 7987 4477
rect 7929 4468 7941 4471
rect 6512 4440 7941 4468
rect 6512 4428 6518 4440
rect 7929 4437 7941 4440
rect 7975 4437 7987 4471
rect 7929 4431 7987 4437
rect 8573 4471 8631 4477
rect 8573 4437 8585 4471
rect 8619 4468 8631 4471
rect 10870 4468 10876 4480
rect 8619 4440 10876 4468
rect 8619 4437 8631 4440
rect 8573 4431 8631 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11348 4477 11376 4508
rect 13004 4508 14924 4536
rect 11333 4471 11391 4477
rect 11333 4437 11345 4471
rect 11379 4437 11391 4471
rect 11333 4431 11391 4437
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 13004 4468 13032 4508
rect 14918 4496 14924 4508
rect 14976 4496 14982 4548
rect 14826 4468 14832 4480
rect 12400 4440 13032 4468
rect 14787 4440 14832 4468
rect 12400 4428 12406 4440
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15289 4471 15347 4477
rect 15289 4437 15301 4471
rect 15335 4468 15347 4471
rect 15746 4468 15752 4480
rect 15335 4440 15752 4468
rect 15335 4437 15347 4440
rect 15289 4431 15347 4437
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 1104 4378 16836 4400
rect 1104 4326 3614 4378
rect 3666 4326 3678 4378
rect 3730 4326 3742 4378
rect 3794 4326 3806 4378
rect 3858 4326 8878 4378
rect 8930 4326 8942 4378
rect 8994 4326 9006 4378
rect 9058 4326 9070 4378
rect 9122 4326 14142 4378
rect 14194 4326 14206 4378
rect 14258 4326 14270 4378
rect 14322 4326 14334 4378
rect 14386 4326 16836 4378
rect 1104 4304 16836 4326
rect 3605 4267 3663 4273
rect 3605 4233 3617 4267
rect 3651 4264 3663 4267
rect 6730 4264 6736 4276
rect 3651 4236 6736 4264
rect 3651 4233 3663 4236
rect 3605 4227 3663 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 2406 4196 2412 4208
rect 2332 4168 2412 4196
rect 2332 4137 2360 4168
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 2590 4156 2596 4208
rect 2648 4196 2654 4208
rect 6454 4196 6460 4208
rect 2648 4168 4384 4196
rect 2648 4156 2654 4168
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2682 4088 2688 4140
rect 2740 4128 2746 4140
rect 3326 4128 3332 4140
rect 2740 4100 3332 4128
rect 2740 4088 2746 4100
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 4356 4137 4384 4168
rect 6380 4168 6460 4196
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 6380 4137 6408 4168
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 7098 4196 7104 4208
rect 6972 4168 7104 4196
rect 6972 4156 6978 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 9214 4196 9220 4208
rect 8864 4168 9220 4196
rect 6365 4131 6423 4137
rect 5040 4100 6204 4128
rect 5040 4088 5046 4100
rect 1780 4032 3556 4060
rect 1780 3933 1808 4032
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 3145 3995 3203 4001
rect 2179 3964 2820 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3893 1823 3927
rect 1765 3887 1823 3893
rect 2222 3884 2228 3936
rect 2280 3924 2286 3936
rect 2792 3933 2820 3964
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 3528 3992 3556 4032
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4801 4063 4859 4069
rect 4801 4060 4813 4063
rect 4212 4032 4813 4060
rect 4212 4020 4218 4032
rect 4801 4029 4813 4032
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 4948 4032 6101 4060
rect 4948 4020 4954 4032
rect 6089 4029 6101 4032
rect 6135 4029 6147 4063
rect 6176 4060 6204 4100
rect 6365 4097 6377 4131
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 8864 4137 8892 4168
rect 9214 4156 9220 4168
rect 9272 4156 9278 4208
rect 10594 4196 10600 4208
rect 10507 4168 10600 4196
rect 10594 4156 10600 4168
rect 10652 4196 10658 4208
rect 10652 4168 11468 4196
rect 10652 4156 10658 4168
rect 11440 4137 11468 4168
rect 12820 4168 13124 4196
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7340 4100 7757 4128
rect 7340 4088 7346 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 11425 4131 11483 4137
rect 11425 4097 11437 4131
rect 11471 4097 11483 4131
rect 11882 4128 11888 4140
rect 11843 4100 11888 4128
rect 11425 4091 11483 4097
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12820 4128 12848 4168
rect 12124 4100 12848 4128
rect 12124 4088 12130 4100
rect 12894 4088 12900 4140
rect 12952 4128 12958 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12952 4100 13001 4128
rect 12952 4088 12958 4100
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 13096 4128 13124 4168
rect 15838 4156 15844 4208
rect 15896 4196 15902 4208
rect 15896 4168 16068 4196
rect 15896 4156 15902 4168
rect 13262 4128 13268 4140
rect 13096 4100 13268 4128
rect 12989 4091 13047 4097
rect 13262 4088 13268 4100
rect 13320 4128 13326 4140
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13320 4100 13921 4128
rect 13320 4088 13326 4100
rect 13909 4097 13921 4100
rect 13955 4097 13967 4131
rect 14090 4128 14096 4140
rect 14051 4100 14096 4128
rect 13909 4091 13967 4097
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14516 4100 15025 4128
rect 14516 4088 14522 4100
rect 15013 4097 15025 4100
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16040 4137 16068 4168
rect 15933 4131 15991 4137
rect 15933 4128 15945 4131
rect 15528 4100 15945 4128
rect 15528 4088 15534 4100
rect 15933 4097 15945 4100
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16025 4131 16083 4137
rect 16025 4097 16037 4131
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 6176 4032 8585 4060
rect 6089 4023 6147 4029
rect 8573 4029 8585 4032
rect 8619 4060 8631 4063
rect 8754 4060 8760 4072
rect 8619 4032 8760 4060
rect 8619 4029 8631 4032
rect 8573 4023 8631 4029
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9766 4060 9772 4072
rect 9263 4032 9772 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9766 4020 9772 4032
rect 9824 4060 9830 4072
rect 10226 4060 10232 4072
rect 9824 4032 10232 4060
rect 9824 4020 9830 4032
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 11241 4063 11299 4069
rect 11241 4060 11253 4063
rect 10928 4032 11253 4060
rect 10928 4020 10934 4032
rect 11241 4029 11253 4032
rect 11287 4029 11299 4063
rect 11241 4023 11299 4029
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 11974 4060 11980 4072
rect 11388 4032 11980 4060
rect 11388 4020 11394 4032
rect 11974 4020 11980 4032
rect 12032 4060 12038 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 12032 4032 14841 4060
rect 12032 4020 12038 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4060 14979 4063
rect 15194 4060 15200 4072
rect 14967 4032 15200 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 15378 4020 15384 4072
rect 15436 4060 15442 4072
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15436 4032 15853 4060
rect 15436 4020 15442 4032
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 4249 3995 4307 4001
rect 4249 3992 4261 3995
rect 3191 3964 3464 3992
rect 3528 3964 4261 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 2777 3927 2835 3933
rect 2280 3896 2325 3924
rect 2280 3884 2286 3896
rect 2777 3893 2789 3927
rect 2823 3893 2835 3927
rect 2777 3887 2835 3893
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3237 3927 3295 3933
rect 3237 3924 3249 3927
rect 3108 3896 3249 3924
rect 3108 3884 3114 3896
rect 3237 3893 3249 3896
rect 3283 3893 3295 3927
rect 3436 3924 3464 3964
rect 4249 3961 4261 3964
rect 4295 3961 4307 3995
rect 4249 3955 4307 3961
rect 4338 3952 4344 4004
rect 4396 3992 4402 4004
rect 5077 3995 5135 4001
rect 5077 3992 5089 3995
rect 4396 3964 5089 3992
rect 4396 3952 4402 3964
rect 5077 3961 5089 3964
rect 5123 3961 5135 3995
rect 5077 3955 5135 3961
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 6181 3995 6239 4001
rect 6181 3992 6193 3995
rect 5592 3964 6193 3992
rect 5592 3952 5598 3964
rect 6181 3961 6193 3964
rect 6227 3961 6239 3995
rect 6181 3955 6239 3961
rect 7024 3964 8800 3992
rect 3605 3927 3663 3933
rect 3605 3924 3617 3927
rect 3436 3896 3617 3924
rect 3237 3887 3295 3893
rect 3605 3893 3617 3896
rect 3651 3893 3663 3927
rect 3786 3924 3792 3936
rect 3747 3896 3792 3924
rect 3605 3887 3663 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4120 3896 4169 3924
rect 4120 3884 4126 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4157 3887 4215 3893
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 5721 3927 5779 3933
rect 5721 3924 5733 3927
rect 4580 3896 5733 3924
rect 4580 3884 4586 3896
rect 5721 3893 5733 3896
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 7024 3924 7052 3964
rect 7190 3924 7196 3936
rect 5868 3896 7052 3924
rect 7151 3896 7196 3924
rect 5868 3884 5874 3896
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7558 3924 7564 3936
rect 7519 3896 7564 3924
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 8202 3924 8208 3936
rect 7708 3896 7753 3924
rect 8163 3896 8208 3924
rect 7708 3884 7714 3896
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 8352 3896 8677 3924
rect 8352 3884 8358 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 8772 3924 8800 3964
rect 9398 3952 9404 4004
rect 9456 4001 9462 4004
rect 9456 3995 9520 4001
rect 9456 3961 9474 3995
rect 9508 3961 9520 3995
rect 9456 3955 9520 3961
rect 9456 3952 9462 3955
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 12066 3992 12072 4004
rect 11204 3964 12072 3992
rect 11204 3952 11210 3964
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 12805 3995 12863 4001
rect 12805 3961 12817 3995
rect 12851 3992 12863 3995
rect 12851 3964 14504 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 9766 3924 9772 3936
rect 8772 3896 9772 3924
rect 8665 3887 8723 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10873 3927 10931 3933
rect 10873 3893 10885 3927
rect 10919 3924 10931 3927
rect 10962 3924 10968 3936
rect 10919 3896 10968 3924
rect 10919 3893 10931 3896
rect 10873 3887 10931 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 12437 3927 12495 3933
rect 11388 3896 11433 3924
rect 11388 3884 11394 3896
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12618 3924 12624 3936
rect 12483 3896 12624 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13354 3924 13360 3936
rect 12943 3896 13360 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 13814 3924 13820 3936
rect 13504 3896 13549 3924
rect 13775 3896 13820 3924
rect 13504 3884 13510 3896
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14476 3933 14504 3964
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3893 14519 3927
rect 14461 3887 14519 3893
rect 15473 3927 15531 3933
rect 15473 3893 15485 3927
rect 15519 3924 15531 3927
rect 15654 3924 15660 3936
rect 15519 3896 15660 3924
rect 15519 3893 15531 3896
rect 15473 3887 15531 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 1104 3834 16836 3856
rect 1104 3782 6246 3834
rect 6298 3782 6310 3834
rect 6362 3782 6374 3834
rect 6426 3782 6438 3834
rect 6490 3782 11510 3834
rect 11562 3782 11574 3834
rect 11626 3782 11638 3834
rect 11690 3782 11702 3834
rect 11754 3782 16836 3834
rect 1104 3760 16836 3782
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2133 3723 2191 3729
rect 2133 3720 2145 3723
rect 2004 3692 2145 3720
rect 2004 3680 2010 3692
rect 2133 3689 2145 3692
rect 2179 3689 2191 3723
rect 2133 3683 2191 3689
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 2777 3723 2835 3729
rect 2777 3720 2789 3723
rect 2280 3692 2789 3720
rect 2280 3680 2286 3692
rect 2777 3689 2789 3692
rect 2823 3689 2835 3723
rect 2777 3683 2835 3689
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 4430 3720 4436 3732
rect 3283 3692 4436 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 4430 3680 4436 3692
rect 4488 3680 4494 3732
rect 4893 3723 4951 3729
rect 4893 3689 4905 3723
rect 4939 3720 4951 3723
rect 5074 3720 5080 3732
rect 4939 3692 5080 3720
rect 4939 3689 4951 3692
rect 4893 3683 4951 3689
rect 5074 3680 5080 3692
rect 5132 3720 5138 3732
rect 5810 3720 5816 3732
rect 5132 3692 5816 3720
rect 5132 3680 5138 3692
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 6549 3723 6607 3729
rect 5960 3692 6005 3720
rect 5960 3680 5966 3692
rect 6549 3689 6561 3723
rect 6595 3689 6607 3723
rect 6549 3683 6607 3689
rect 3786 3652 3792 3664
rect 2240 3624 3792 3652
rect 2240 3593 2268 3624
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 5442 3652 5448 3664
rect 5316 3624 5448 3652
rect 5316 3612 5322 3624
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 6564 3652 6592 3683
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 6917 3723 6975 3729
rect 6917 3720 6929 3723
rect 6788 3692 6929 3720
rect 6788 3680 6794 3692
rect 6917 3689 6929 3692
rect 6963 3720 6975 3723
rect 7190 3720 7196 3732
rect 6963 3692 7196 3720
rect 6963 3689 6975 3692
rect 6917 3683 6975 3689
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7561 3723 7619 3729
rect 7561 3689 7573 3723
rect 7607 3720 7619 3723
rect 7650 3720 7656 3732
rect 7607 3692 7656 3720
rect 7607 3689 7619 3692
rect 7561 3683 7619 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 9033 3723 9091 3729
rect 9033 3720 9045 3723
rect 8260 3692 9045 3720
rect 8260 3680 8266 3692
rect 9033 3689 9045 3692
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 10597 3723 10655 3729
rect 10597 3689 10609 3723
rect 10643 3689 10655 3723
rect 10962 3720 10968 3732
rect 10923 3692 10968 3720
rect 10597 3683 10655 3689
rect 7929 3655 7987 3661
rect 7929 3652 7941 3655
rect 6564 3624 7941 3652
rect 7929 3621 7941 3624
rect 7975 3621 7987 3655
rect 7929 3615 7987 3621
rect 8021 3655 8079 3661
rect 8021 3621 8033 3655
rect 8067 3652 8079 3655
rect 8386 3652 8392 3664
rect 8067 3624 8392 3652
rect 8067 3621 8079 3624
rect 8021 3615 8079 3621
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 10502 3652 10508 3664
rect 8956 3624 10508 3652
rect 8956 3596 8984 3624
rect 10502 3612 10508 3624
rect 10560 3612 10566 3664
rect 10612 3652 10640 3683
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12618 3720 12624 3732
rect 12579 3692 12624 3720
rect 12618 3680 12624 3692
rect 12676 3680 12682 3732
rect 14458 3680 14464 3732
rect 14516 3720 14522 3732
rect 14553 3723 14611 3729
rect 14553 3720 14565 3723
rect 14516 3692 14565 3720
rect 14516 3680 14522 3692
rect 14553 3689 14565 3692
rect 14599 3689 14611 3723
rect 15654 3720 15660 3732
rect 15615 3692 15660 3720
rect 14553 3683 14611 3689
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 15804 3692 15849 3720
rect 15804 3680 15810 3692
rect 12342 3652 12348 3664
rect 10612 3624 12348 3652
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12526 3652 12532 3664
rect 12487 3624 12532 3652
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 13440 3655 13498 3661
rect 13440 3621 13452 3655
rect 13486 3652 13498 3655
rect 13814 3652 13820 3664
rect 13486 3624 13820 3652
rect 13486 3621 13498 3624
rect 13440 3615 13498 3621
rect 13814 3612 13820 3624
rect 13872 3652 13878 3664
rect 14090 3652 14096 3664
rect 13872 3624 14096 3652
rect 13872 3612 13878 3624
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3553 2283 3587
rect 3145 3587 3203 3593
rect 3145 3584 3157 3587
rect 2225 3547 2283 3553
rect 2332 3556 3157 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2332 3516 2360 3556
rect 3145 3553 3157 3556
rect 3191 3584 3203 3587
rect 4706 3584 4712 3596
rect 3191 3556 4712 3584
rect 3191 3553 3203 3556
rect 3145 3547 3203 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 5810 3584 5816 3596
rect 5684 3556 5816 3584
rect 5684 3544 5690 3556
rect 5810 3544 5816 3556
rect 5868 3584 5874 3596
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5868 3556 6009 3584
rect 5868 3544 5874 3556
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7098 3584 7104 3596
rect 7055 3556 7104 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 8478 3584 8484 3596
rect 7208 3556 8484 3584
rect 1728 3488 2360 3516
rect 2409 3519 2467 3525
rect 1728 3476 1734 3488
rect 2409 3485 2421 3519
rect 2455 3516 2467 3519
rect 3050 3516 3056 3528
rect 2455 3488 3056 3516
rect 2455 3485 2467 3488
rect 2409 3479 2467 3485
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3326 3516 3332 3528
rect 3287 3488 3332 3516
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 4062 3516 4068 3528
rect 4023 3488 4068 3516
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5442 3516 5448 3528
rect 5215 3488 5448 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 1854 3408 1860 3460
rect 1912 3448 1918 3460
rect 5000 3448 5028 3479
rect 5442 3476 5448 3488
rect 5500 3516 5506 3528
rect 6181 3519 6239 3525
rect 6181 3516 6193 3519
rect 5500 3488 6193 3516
rect 5500 3476 5506 3488
rect 6181 3485 6193 3488
rect 6227 3516 6239 3519
rect 6454 3516 6460 3528
rect 6227 3488 6460 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 7208 3525 7236 3556
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 8938 3584 8944 3596
rect 8899 3556 8944 3584
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 9953 3587 10011 3593
rect 9953 3553 9965 3587
rect 9999 3584 10011 3587
rect 10870 3584 10876 3596
rect 9999 3556 10876 3584
rect 9999 3553 10011 3556
rect 9953 3547 10011 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11609 3587 11667 3593
rect 11609 3553 11621 3587
rect 11655 3584 11667 3587
rect 11974 3584 11980 3596
rect 11655 3556 11980 3584
rect 11655 3553 11667 3556
rect 11609 3547 11667 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 7742 3516 7748 3528
rect 7340 3488 7748 3516
rect 7340 3476 7346 3488
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9214 3476 9220 3488
rect 9272 3516 9278 3528
rect 9398 3516 9404 3528
rect 9272 3488 9404 3516
rect 9272 3476 9278 3488
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10468 3488 11069 3516
rect 10468 3476 10474 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3516 11299 3519
rect 11698 3516 11704 3528
rect 11287 3488 11704 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 12710 3516 12716 3528
rect 12671 3488 12716 3516
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13170 3516 13176 3528
rect 13131 3488 13176 3516
rect 13170 3476 13176 3488
rect 13228 3476 13234 3528
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 14976 3488 15853 3516
rect 14976 3476 14982 3488
rect 15841 3485 15853 3488
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 5994 3448 6000 3460
rect 1912 3420 4936 3448
rect 5000 3420 6000 3448
rect 1912 3408 1918 3420
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3380 1823 3383
rect 2222 3380 2228 3392
rect 1811 3352 2228 3380
rect 1811 3349 1823 3352
rect 1765 3343 1823 3349
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 3568 3352 4537 3380
rect 3568 3340 3574 3352
rect 4525 3349 4537 3352
rect 4571 3349 4583 3383
rect 4908 3380 4936 3420
rect 5994 3408 6000 3420
rect 6052 3408 6058 3460
rect 7834 3408 7840 3460
rect 7892 3448 7898 3460
rect 11146 3448 11152 3460
rect 7892 3420 11152 3448
rect 7892 3408 7898 3420
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 5074 3380 5080 3392
rect 4908 3352 5080 3380
rect 4525 3343 4583 3349
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5534 3380 5540 3392
rect 5495 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 8294 3380 8300 3392
rect 5684 3352 8300 3380
rect 5684 3340 5690 3352
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 8573 3383 8631 3389
rect 8573 3349 8585 3383
rect 8619 3380 8631 3383
rect 10686 3380 10692 3392
rect 8619 3352 10692 3380
rect 8619 3349 8631 3352
rect 8573 3343 8631 3349
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 11793 3383 11851 3389
rect 11793 3349 11805 3383
rect 11839 3380 11851 3383
rect 11974 3380 11980 3392
rect 11839 3352 11980 3380
rect 11839 3349 11851 3352
rect 11793 3343 11851 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12161 3383 12219 3389
rect 12161 3349 12173 3383
rect 12207 3380 12219 3383
rect 13538 3380 13544 3392
rect 12207 3352 13544 3380
rect 12207 3349 12219 3352
rect 12161 3343 12219 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 15102 3340 15108 3392
rect 15160 3380 15166 3392
rect 15289 3383 15347 3389
rect 15289 3380 15301 3383
rect 15160 3352 15301 3380
rect 15160 3340 15166 3352
rect 15289 3349 15301 3352
rect 15335 3349 15347 3383
rect 15289 3343 15347 3349
rect 1104 3290 16836 3312
rect 1104 3238 3614 3290
rect 3666 3238 3678 3290
rect 3730 3238 3742 3290
rect 3794 3238 3806 3290
rect 3858 3238 8878 3290
rect 8930 3238 8942 3290
rect 8994 3238 9006 3290
rect 9058 3238 9070 3290
rect 9122 3238 14142 3290
rect 14194 3238 14206 3290
rect 14258 3238 14270 3290
rect 14322 3238 14334 3290
rect 14386 3238 16836 3290
rect 1104 3216 16836 3238
rect 474 3136 480 3188
rect 532 3176 538 3188
rect 2777 3179 2835 3185
rect 532 3148 2360 3176
rect 532 3136 538 3148
rect 2332 3108 2360 3148
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 3326 3176 3332 3188
rect 2823 3148 3332 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 3326 3136 3332 3148
rect 3384 3136 3390 3188
rect 4154 3176 4160 3188
rect 4115 3148 4160 3176
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4632 3148 6500 3176
rect 4632 3108 4660 3148
rect 2332 3080 4660 3108
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 4764 3080 6377 3108
rect 4764 3068 4770 3080
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 6472 3108 6500 3148
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 7101 3179 7159 3185
rect 7101 3176 7113 3179
rect 6696 3148 7113 3176
rect 6696 3136 6702 3148
rect 7101 3145 7113 3148
rect 7147 3145 7159 3179
rect 7101 3139 7159 3145
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 7892 3148 8309 3176
rect 7892 3136 7898 3148
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 9582 3176 9588 3188
rect 8297 3139 8355 3145
rect 8404 3148 9588 3176
rect 7282 3108 7288 3120
rect 6472 3080 7288 3108
rect 6365 3071 6423 3077
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 7926 3068 7932 3120
rect 7984 3068 7990 3120
rect 8404 3108 8432 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10134 3176 10140 3188
rect 9916 3148 10140 3176
rect 9916 3136 9922 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 11698 3176 11704 3188
rect 10560 3148 11560 3176
rect 11659 3148 11704 3176
rect 10560 3136 10566 3148
rect 8036 3080 8432 3108
rect 9309 3111 9367 3117
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4246 3040 4252 3052
rect 3835 3012 4252 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4798 3040 4804 3052
rect 4759 3012 4804 3040
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5534 3040 5540 3052
rect 5224 3012 5540 3040
rect 5224 3000 5230 3012
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 5718 3040 5724 3052
rect 5679 3012 5724 3040
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 7745 3043 7803 3049
rect 5868 3012 7512 3040
rect 5868 3000 5874 3012
rect 3510 2972 3516 2984
rect 3471 2944 3516 2972
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 4982 2972 4988 2984
rect 3651 2944 4988 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5626 2972 5632 2984
rect 5587 2944 5632 2972
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 7374 2972 7380 2984
rect 6227 2944 7380 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7484 2972 7512 3012
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 7944 3040 7972 3068
rect 7791 3012 7972 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 7926 2972 7932 2984
rect 7484 2944 7932 2972
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 1642 2907 1700 2913
rect 1642 2904 1654 2907
rect 1412 2876 1654 2904
rect 1412 2848 1440 2876
rect 1642 2873 1654 2876
rect 1688 2873 1700 2907
rect 4617 2907 4675 2913
rect 4617 2904 4629 2907
rect 1642 2867 1700 2873
rect 3160 2876 4629 2904
rect 1394 2796 1400 2848
rect 1452 2796 1458 2848
rect 3160 2845 3188 2876
rect 4617 2873 4629 2876
rect 4663 2873 4675 2907
rect 4617 2867 4675 2873
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 5537 2907 5595 2913
rect 5537 2904 5549 2907
rect 5132 2876 5549 2904
rect 5132 2864 5138 2876
rect 5537 2873 5549 2876
rect 5583 2873 5595 2907
rect 5537 2867 5595 2873
rect 5994 2864 6000 2916
rect 6052 2904 6058 2916
rect 7561 2907 7619 2913
rect 7561 2904 7573 2907
rect 6052 2876 7573 2904
rect 6052 2864 6058 2876
rect 7561 2873 7573 2876
rect 7607 2904 7619 2907
rect 8036 2904 8064 3080
rect 9309 3077 9321 3111
rect 9355 3108 9367 3111
rect 10318 3108 10324 3120
rect 9355 3080 10324 3108
rect 9355 3077 9367 3080
rect 9309 3071 9367 3077
rect 10318 3068 10324 3080
rect 10376 3068 10382 3120
rect 11532 3108 11560 3148
rect 11698 3136 11704 3148
rect 11756 3176 11762 3188
rect 11756 3148 12480 3176
rect 11756 3136 11762 3148
rect 12250 3108 12256 3120
rect 11532 3080 12256 3108
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9953 3043 10011 3049
rect 9953 3040 9965 3043
rect 9272 3012 9965 3040
rect 9272 3000 9278 3012
rect 9953 3009 9965 3012
rect 9999 3009 10011 3043
rect 12452 3040 12480 3148
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 13814 3176 13820 3188
rect 13775 3148 13820 3176
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 13372 3108 13400 3136
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 13372 3080 14105 3108
rect 14093 3077 14105 3080
rect 14139 3077 14151 3111
rect 14093 3071 14151 3077
rect 14458 3068 14464 3120
rect 14516 3108 14522 3120
rect 14516 3080 14688 3108
rect 14516 3068 14522 3080
rect 12452 3012 12572 3040
rect 9953 3003 10011 3009
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 8628 2944 8677 2972
rect 8628 2932 8634 2944
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 9490 2972 9496 2984
rect 8665 2935 8723 2941
rect 9324 2944 9496 2972
rect 9324 2904 9352 2944
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 9677 2975 9735 2981
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 9766 2972 9772 2984
rect 9723 2944 9772 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 7607 2876 8064 2904
rect 8680 2876 9352 2904
rect 7607 2873 7619 2876
rect 7561 2867 7619 2873
rect 3145 2839 3203 2845
rect 3145 2805 3157 2839
rect 3191 2805 3203 2839
rect 4522 2836 4528 2848
rect 4483 2808 4528 2836
rect 3145 2799 3203 2805
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 5166 2836 5172 2848
rect 5127 2808 5172 2836
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 7469 2839 7527 2845
rect 7469 2805 7481 2839
rect 7515 2836 7527 2839
rect 8680 2836 8708 2876
rect 9398 2864 9404 2916
rect 9456 2904 9462 2916
rect 9968 2904 9996 3003
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10594 2981 10600 2984
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 10284 2944 10333 2972
rect 10284 2932 10290 2944
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 10588 2972 10600 2981
rect 10555 2944 10600 2972
rect 10321 2935 10379 2941
rect 10588 2935 10600 2944
rect 10594 2932 10600 2935
rect 10652 2932 10658 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2941 12495 2975
rect 12544 2972 12572 3012
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 14660 3049 14688 3080
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 13504 3012 14565 3040
rect 13504 3000 13510 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 15381 3043 15439 3049
rect 14792 3012 15332 3040
rect 14792 3000 14798 3012
rect 12693 2975 12751 2981
rect 12693 2972 12705 2975
rect 12544 2944 12705 2972
rect 12437 2935 12495 2941
rect 12693 2941 12705 2944
rect 12739 2941 12751 2975
rect 12693 2935 12751 2941
rect 11054 2904 11060 2916
rect 9456 2876 9904 2904
rect 9968 2876 11060 2904
rect 9456 2864 9462 2876
rect 7515 2808 8708 2836
rect 7515 2805 7527 2808
rect 7469 2799 7527 2805
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 9766 2836 9772 2848
rect 8812 2808 8857 2836
rect 9727 2808 9772 2836
rect 8812 2796 8818 2808
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 9876 2836 9904 2876
rect 11054 2864 11060 2876
rect 11112 2904 11118 2916
rect 12066 2904 12072 2916
rect 11112 2876 12072 2904
rect 11112 2864 11118 2876
rect 12066 2864 12072 2876
rect 12124 2864 12130 2916
rect 12452 2904 12480 2935
rect 13998 2932 14004 2984
rect 14056 2972 14062 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14056 2944 14473 2972
rect 14056 2932 14062 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 15102 2972 15108 2984
rect 15063 2944 15108 2972
rect 14461 2935 14519 2941
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 15304 2972 15332 3012
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 17494 3040 17500 3052
rect 15427 3012 17500 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 15841 2975 15899 2981
rect 15841 2972 15853 2975
rect 15304 2944 15853 2972
rect 15841 2941 15853 2944
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 13170 2904 13176 2916
rect 12452 2876 13176 2904
rect 13170 2864 13176 2876
rect 13228 2864 13234 2916
rect 13906 2864 13912 2916
rect 13964 2864 13970 2916
rect 14918 2904 14924 2916
rect 14375 2876 14924 2904
rect 13924 2836 13952 2864
rect 14375 2836 14403 2876
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 15654 2864 15660 2916
rect 15712 2904 15718 2916
rect 16117 2907 16175 2913
rect 16117 2904 16129 2907
rect 15712 2876 16129 2904
rect 15712 2864 15718 2876
rect 16117 2873 16129 2876
rect 16163 2873 16175 2907
rect 16117 2867 16175 2873
rect 9876 2808 14403 2836
rect 1104 2746 16836 2768
rect 1104 2694 6246 2746
rect 6298 2694 6310 2746
rect 6362 2694 6374 2746
rect 6426 2694 6438 2746
rect 6490 2694 11510 2746
rect 11562 2694 11574 2746
rect 11626 2694 11638 2746
rect 11690 2694 11702 2746
rect 11754 2694 16836 2746
rect 1104 2672 16836 2694
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 4062 2632 4068 2644
rect 3375 2604 4068 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4982 2632 4988 2644
rect 4943 2604 4988 2632
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5445 2635 5503 2641
rect 5445 2632 5457 2635
rect 5224 2604 5457 2632
rect 5224 2592 5230 2604
rect 5445 2601 5457 2604
rect 5491 2601 5503 2635
rect 7006 2632 7012 2644
rect 6967 2604 7012 2632
rect 5445 2595 5503 2601
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 8754 2632 8760 2644
rect 8711 2604 8760 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 9030 2632 9036 2644
rect 8991 2604 9036 2632
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9122 2592 9128 2644
rect 9180 2632 9186 2644
rect 10410 2632 10416 2644
rect 9180 2604 9225 2632
rect 10371 2604 10416 2632
rect 9180 2592 9186 2604
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10744 2604 10885 2632
rect 10744 2592 10750 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 11330 2592 11336 2644
rect 11388 2632 11394 2644
rect 11425 2635 11483 2641
rect 11425 2632 11437 2635
rect 11388 2604 11437 2632
rect 11388 2592 11394 2604
rect 11425 2601 11437 2604
rect 11471 2601 11483 2635
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11425 2595 11483 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 13538 2592 13544 2644
rect 13596 2632 13602 2644
rect 15289 2635 15347 2641
rect 15289 2632 15301 2635
rect 13596 2604 15301 2632
rect 13596 2592 13602 2604
rect 15289 2601 15301 2604
rect 15335 2601 15347 2635
rect 15289 2595 15347 2601
rect 3694 2524 3700 2576
rect 3752 2564 3758 2576
rect 4706 2564 4712 2576
rect 3752 2536 4712 2564
rect 3752 2524 3758 2536
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 5350 2564 5356 2576
rect 5311 2536 5356 2564
rect 5350 2524 5356 2536
rect 5408 2524 5414 2576
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 5592 2536 7481 2564
rect 5592 2524 5598 2536
rect 7469 2533 7481 2536
rect 7515 2533 7527 2567
rect 7469 2527 7527 2533
rect 10318 2524 10324 2576
rect 10376 2564 10382 2576
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 10376 2536 10793 2564
rect 10376 2524 10382 2536
rect 10781 2533 10793 2536
rect 10827 2533 10839 2567
rect 10781 2527 10839 2533
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 11793 2567 11851 2573
rect 11793 2564 11805 2567
rect 11204 2536 11805 2564
rect 11204 2524 11210 2536
rect 11793 2533 11805 2536
rect 11839 2533 11851 2567
rect 11793 2527 11851 2533
rect 12250 2524 12256 2576
rect 12308 2564 12314 2576
rect 12308 2536 12736 2564
rect 12308 2524 12314 2536
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 3421 2499 3479 2505
rect 3421 2465 3433 2499
rect 3467 2496 3479 2499
rect 4154 2496 4160 2508
rect 3467 2468 4160 2496
rect 3467 2465 3479 2468
rect 3421 2459 3479 2465
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4614 2496 4620 2508
rect 4295 2468 4620 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 6086 2496 6092 2508
rect 6047 2468 6092 2496
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7248 2468 8033 2496
rect 7248 2456 7254 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 8021 2459 8079 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12400 2468 12633 2496
rect 12400 2456 12406 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12708 2496 12736 2536
rect 12802 2524 12808 2576
rect 12860 2564 12866 2576
rect 15749 2567 15807 2573
rect 15749 2564 15761 2567
rect 12860 2536 15761 2564
rect 12860 2524 12866 2536
rect 15749 2533 15761 2536
rect 15795 2533 15807 2567
rect 15749 2527 15807 2533
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 12708 2468 13461 2496
rect 12621 2459 12679 2465
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 13909 2499 13967 2505
rect 13909 2465 13921 2499
rect 13955 2496 13967 2499
rect 14001 2499 14059 2505
rect 14001 2496 14013 2499
rect 13955 2468 14013 2496
rect 13955 2465 13967 2468
rect 13909 2459 13967 2465
rect 14001 2465 14013 2468
rect 14047 2465 14059 2499
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14001 2459 14059 2465
rect 14108 2468 14841 2496
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 3234 2428 3240 2440
rect 2547 2400 3240 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 4430 2428 4436 2440
rect 3651 2400 4436 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4571 2400 4660 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 4632 2360 4660 2400
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 5442 2428 5448 2440
rect 4764 2400 5448 2428
rect 4764 2388 4770 2400
rect 5442 2388 5448 2400
rect 5500 2428 5506 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 5500 2400 5549 2428
rect 5500 2388 5506 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 7098 2428 7104 2440
rect 6411 2400 7104 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7524 2400 7573 2428
rect 7524 2388 7530 2400
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 7984 2400 8432 2428
rect 7984 2388 7990 2400
rect 6086 2360 6092 2372
rect 4632 2332 6092 2360
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 8404 2360 8432 2400
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 8536 2400 9229 2428
rect 8536 2388 8542 2400
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10652 2400 10977 2428
rect 10652 2388 10658 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 12066 2428 12072 2440
rect 12027 2400 12072 2428
rect 10965 2391 11023 2397
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 11698 2360 11704 2372
rect 8404 2332 11704 2360
rect 11698 2320 11704 2332
rect 11756 2320 11762 2372
rect 11790 2320 11796 2372
rect 11848 2360 11854 2372
rect 12820 2360 12848 2391
rect 13354 2388 13360 2440
rect 13412 2428 13418 2440
rect 14108 2428 14136 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 15289 2499 15347 2505
rect 15289 2465 15301 2499
rect 15335 2496 15347 2499
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15335 2468 15485 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 13412 2400 14136 2428
rect 14277 2431 14335 2437
rect 13412 2388 13418 2400
rect 14277 2397 14289 2431
rect 14323 2428 14335 2431
rect 14642 2428 14648 2440
rect 14323 2400 14648 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 13814 2360 13820 2372
rect 11848 2332 12848 2360
rect 13556 2332 13820 2360
rect 11848 2320 11854 2332
rect 1857 2295 1915 2301
rect 1857 2261 1869 2295
rect 1903 2292 1915 2295
rect 2774 2292 2780 2304
rect 1903 2264 2780 2292
rect 1903 2261 1915 2264
rect 1857 2255 1915 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 2961 2295 3019 2301
rect 2961 2261 2973 2295
rect 3007 2292 3019 2295
rect 4890 2292 4896 2304
rect 3007 2264 4896 2292
rect 3007 2261 3019 2264
rect 2961 2255 3019 2261
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 8202 2292 8208 2304
rect 8163 2264 8208 2292
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 9953 2295 10011 2301
rect 9953 2261 9965 2295
rect 9999 2292 10011 2295
rect 13556 2292 13584 2332
rect 13814 2320 13820 2332
rect 13872 2320 13878 2372
rect 13909 2363 13967 2369
rect 13909 2329 13921 2363
rect 13955 2360 13967 2363
rect 14550 2360 14556 2372
rect 13955 2332 14556 2360
rect 13955 2329 13967 2332
rect 13909 2323 13967 2329
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 9999 2264 13584 2292
rect 13633 2295 13691 2301
rect 9999 2261 10011 2264
rect 9953 2255 10011 2261
rect 13633 2261 13645 2295
rect 13679 2292 13691 2295
rect 14918 2292 14924 2304
rect 13679 2264 14924 2292
rect 13679 2261 13691 2264
rect 13633 2255 13691 2261
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 15068 2264 15113 2292
rect 15068 2252 15074 2264
rect 1104 2202 16836 2224
rect 1104 2150 3614 2202
rect 3666 2150 3678 2202
rect 3730 2150 3742 2202
rect 3794 2150 3806 2202
rect 3858 2150 8878 2202
rect 8930 2150 8942 2202
rect 8994 2150 9006 2202
rect 9058 2150 9070 2202
rect 9122 2150 14142 2202
rect 14194 2150 14206 2202
rect 14258 2150 14270 2202
rect 14322 2150 14334 2202
rect 14386 2150 16836 2202
rect 1104 2128 16836 2150
rect 2498 2048 2504 2100
rect 2556 2088 2562 2100
rect 9766 2088 9772 2100
rect 2556 2060 9772 2088
rect 2556 2048 2562 2060
rect 9766 2048 9772 2060
rect 9824 2048 9830 2100
rect 2314 1436 2320 1488
rect 2372 1476 2378 1488
rect 9398 1476 9404 1488
rect 2372 1448 9404 1476
rect 2372 1436 2378 1448
rect 9398 1436 9404 1448
rect 9456 1436 9462 1488
rect 3694 1028 3700 1080
rect 3752 1068 3758 1080
rect 8202 1068 8208 1080
rect 3752 1040 8208 1068
rect 3752 1028 3758 1040
rect 8202 1028 8208 1040
rect 8260 1028 8266 1080
<< via1 >>
rect 4068 15172 4120 15224
rect 8944 15172 8996 15224
rect 9312 15172 9364 15224
rect 14924 15172 14976 15224
rect 6246 14662 6298 14714
rect 6310 14662 6362 14714
rect 6374 14662 6426 14714
rect 6438 14662 6490 14714
rect 11510 14662 11562 14714
rect 11574 14662 11626 14714
rect 11638 14662 11690 14714
rect 11702 14662 11754 14714
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 10324 14560 10376 14612
rect 11060 14492 11112 14544
rect 6644 14424 6696 14476
rect 8760 14424 8812 14476
rect 10416 14424 10468 14476
rect 10692 14424 10744 14476
rect 6092 14356 6144 14408
rect 7104 14356 7156 14408
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 9220 14399 9272 14408
rect 9220 14365 9229 14399
rect 9229 14365 9263 14399
rect 9263 14365 9272 14399
rect 9220 14356 9272 14365
rect 4068 14220 4120 14272
rect 5540 14220 5592 14272
rect 6184 14220 6236 14272
rect 7656 14220 7708 14272
rect 8576 14263 8628 14272
rect 8576 14229 8585 14263
rect 8585 14229 8619 14263
rect 8619 14229 8628 14263
rect 8576 14220 8628 14229
rect 16304 14220 16356 14272
rect 3614 14118 3666 14170
rect 3678 14118 3730 14170
rect 3742 14118 3794 14170
rect 3806 14118 3858 14170
rect 8878 14118 8930 14170
rect 8942 14118 8994 14170
rect 9006 14118 9058 14170
rect 9070 14118 9122 14170
rect 14142 14118 14194 14170
rect 14206 14118 14258 14170
rect 14270 14118 14322 14170
rect 14334 14118 14386 14170
rect 9496 14016 9548 14068
rect 14832 14016 14884 14068
rect 5540 13948 5592 14000
rect 13544 13948 13596 14000
rect 3148 13880 3200 13932
rect 5080 13880 5132 13932
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 6920 13880 6972 13932
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 9220 13923 9272 13932
rect 7840 13880 7892 13889
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 9864 13880 9916 13932
rect 15200 13880 15252 13932
rect 3976 13812 4028 13864
rect 8392 13812 8444 13864
rect 9312 13812 9364 13864
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 4896 13744 4948 13796
rect 7380 13744 7432 13796
rect 9680 13744 9732 13796
rect 2228 13719 2280 13728
rect 2228 13685 2237 13719
rect 2237 13685 2271 13719
rect 2271 13685 2280 13719
rect 2228 13676 2280 13685
rect 3332 13676 3384 13728
rect 4528 13676 4580 13728
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 7012 13676 7064 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7748 13676 7800 13728
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 8852 13676 8904 13728
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 10508 13719 10560 13728
rect 10508 13685 10517 13719
rect 10517 13685 10551 13719
rect 10551 13685 10560 13719
rect 10508 13676 10560 13685
rect 12532 13744 12584 13796
rect 13360 13744 13412 13796
rect 14924 13676 14976 13728
rect 15108 13719 15160 13728
rect 15108 13685 15117 13719
rect 15117 13685 15151 13719
rect 15151 13685 15160 13719
rect 15108 13676 15160 13685
rect 15476 13719 15528 13728
rect 15476 13685 15485 13719
rect 15485 13685 15519 13719
rect 15519 13685 15528 13719
rect 15476 13676 15528 13685
rect 15660 13676 15712 13728
rect 6246 13574 6298 13626
rect 6310 13574 6362 13626
rect 6374 13574 6426 13626
rect 6438 13574 6490 13626
rect 11510 13574 11562 13626
rect 11574 13574 11626 13626
rect 11638 13574 11690 13626
rect 11702 13574 11754 13626
rect 8668 13472 8720 13524
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 2504 13379 2556 13388
rect 2504 13345 2513 13379
rect 2513 13345 2547 13379
rect 2547 13345 2556 13379
rect 2504 13336 2556 13345
rect 5632 13336 5684 13388
rect 7564 13404 7616 13456
rect 8024 13404 8076 13456
rect 15476 13472 15528 13524
rect 12532 13404 12584 13456
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 5080 13311 5132 13320
rect 2688 13268 2740 13277
rect 5080 13277 5089 13311
rect 5089 13277 5123 13311
rect 5123 13277 5132 13311
rect 5080 13268 5132 13277
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 5816 13200 5868 13252
rect 5908 13200 5960 13252
rect 6828 13336 6880 13388
rect 7840 13336 7892 13388
rect 8208 13336 8260 13388
rect 8576 13336 8628 13388
rect 8852 13336 8904 13388
rect 10692 13336 10744 13388
rect 11888 13336 11940 13388
rect 7656 13268 7708 13320
rect 10876 13268 10928 13320
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 13452 13336 13504 13388
rect 13636 13379 13688 13388
rect 13636 13345 13670 13379
rect 13670 13345 13688 13379
rect 13636 13336 13688 13345
rect 12900 13311 12952 13320
rect 12900 13277 12909 13311
rect 12909 13277 12943 13311
rect 12943 13277 12952 13311
rect 15016 13404 15068 13456
rect 15936 13379 15988 13388
rect 15936 13345 15945 13379
rect 15945 13345 15979 13379
rect 15979 13345 15988 13379
rect 15936 13336 15988 13345
rect 16396 13336 16448 13388
rect 12900 13268 12952 13277
rect 13084 13200 13136 13252
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 4436 13175 4488 13184
rect 4436 13141 4445 13175
rect 4445 13141 4479 13175
rect 4479 13141 4488 13175
rect 4436 13132 4488 13141
rect 5172 13132 5224 13184
rect 7288 13132 7340 13184
rect 8300 13132 8352 13184
rect 9220 13132 9272 13184
rect 9496 13132 9548 13184
rect 9772 13132 9824 13184
rect 12256 13132 12308 13184
rect 13176 13132 13228 13184
rect 16028 13200 16080 13252
rect 14464 13132 14516 13184
rect 14832 13132 14884 13184
rect 3614 13030 3666 13082
rect 3678 13030 3730 13082
rect 3742 13030 3794 13082
rect 3806 13030 3858 13082
rect 8878 13030 8930 13082
rect 8942 13030 8994 13082
rect 9006 13030 9058 13082
rect 9070 13030 9122 13082
rect 14142 13030 14194 13082
rect 14206 13030 14258 13082
rect 14270 13030 14322 13082
rect 14334 13030 14386 13082
rect 4712 12928 4764 12980
rect 6828 12928 6880 12980
rect 2688 12792 2740 12844
rect 4160 12860 4212 12912
rect 5356 12860 5408 12912
rect 3976 12792 4028 12844
rect 5448 12835 5500 12844
rect 5448 12801 5457 12835
rect 5457 12801 5491 12835
rect 5491 12801 5500 12835
rect 5448 12792 5500 12801
rect 7196 12792 7248 12844
rect 7656 12792 7708 12844
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 2228 12724 2280 12776
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 7932 12724 7984 12776
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 9864 12792 9916 12844
rect 11888 12835 11940 12844
rect 9956 12724 10008 12776
rect 3424 12656 3476 12708
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 2780 12631 2832 12640
rect 2780 12597 2789 12631
rect 2789 12597 2823 12631
rect 2823 12597 2832 12631
rect 2780 12588 2832 12597
rect 4068 12588 4120 12640
rect 4252 12631 4304 12640
rect 4252 12597 4261 12631
rect 4261 12597 4295 12631
rect 4295 12597 4304 12631
rect 4252 12588 4304 12597
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 9496 12699 9548 12708
rect 9496 12665 9505 12699
rect 9505 12665 9539 12699
rect 9539 12665 9548 12699
rect 9496 12656 9548 12665
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 13452 12928 13504 12980
rect 13636 12860 13688 12912
rect 12072 12724 12124 12776
rect 13452 12724 13504 12776
rect 10416 12656 10468 12708
rect 5264 12588 5316 12597
rect 7932 12631 7984 12640
rect 7932 12597 7941 12631
rect 7941 12597 7975 12631
rect 7975 12597 7984 12631
rect 7932 12588 7984 12597
rect 9036 12631 9088 12640
rect 9036 12597 9045 12631
rect 9045 12597 9079 12631
rect 9079 12597 9088 12631
rect 9036 12588 9088 12597
rect 9128 12588 9180 12640
rect 11336 12588 11388 12640
rect 11980 12656 12032 12708
rect 12808 12656 12860 12708
rect 15200 12656 15252 12708
rect 14740 12588 14792 12640
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 6246 12486 6298 12538
rect 6310 12486 6362 12538
rect 6374 12486 6426 12538
rect 6438 12486 6490 12538
rect 11510 12486 11562 12538
rect 11574 12486 11626 12538
rect 11638 12486 11690 12538
rect 11702 12486 11754 12538
rect 1768 12384 1820 12436
rect 2136 12384 2188 12436
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 5816 12427 5868 12436
rect 5816 12393 5825 12427
rect 5825 12393 5859 12427
rect 5859 12393 5868 12427
rect 5816 12384 5868 12393
rect 7840 12384 7892 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 10508 12384 10560 12436
rect 11980 12384 12032 12436
rect 12256 12384 12308 12436
rect 14464 12384 14516 12436
rect 15568 12384 15620 12436
rect 4620 12316 4672 12368
rect 11336 12316 11388 12368
rect 12532 12316 12584 12368
rect 14648 12316 14700 12368
rect 2964 12291 3016 12300
rect 2964 12257 2973 12291
rect 2973 12257 3007 12291
rect 3007 12257 3016 12291
rect 2964 12248 3016 12257
rect 3056 12291 3108 12300
rect 3056 12257 3065 12291
rect 3065 12257 3099 12291
rect 3099 12257 3108 12291
rect 3056 12248 3108 12257
rect 5816 12248 5868 12300
rect 6000 12248 6052 12300
rect 8208 12248 8260 12300
rect 10324 12248 10376 12300
rect 2872 12180 2924 12232
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 2596 12112 2648 12164
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 4344 12044 4396 12096
rect 4804 12044 4856 12096
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 5632 12044 5684 12096
rect 6184 12044 6236 12096
rect 7748 12180 7800 12232
rect 9128 12180 9180 12232
rect 9956 12180 10008 12232
rect 12348 12248 12400 12300
rect 12624 12291 12676 12300
rect 12624 12257 12633 12291
rect 12633 12257 12667 12291
rect 12667 12257 12676 12291
rect 12624 12248 12676 12257
rect 14832 12248 14884 12300
rect 15476 12248 15528 12300
rect 7564 12112 7616 12164
rect 12440 12180 12492 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 13452 12180 13504 12232
rect 14924 12180 14976 12232
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 13084 12112 13136 12164
rect 6736 12044 6788 12096
rect 9312 12044 9364 12096
rect 10048 12044 10100 12096
rect 10876 12044 10928 12096
rect 13912 12044 13964 12096
rect 15200 12044 15252 12096
rect 15844 12044 15896 12096
rect 3614 11942 3666 11994
rect 3678 11942 3730 11994
rect 3742 11942 3794 11994
rect 3806 11942 3858 11994
rect 8878 11942 8930 11994
rect 8942 11942 8994 11994
rect 9006 11942 9058 11994
rect 9070 11942 9122 11994
rect 14142 11942 14194 11994
rect 14206 11942 14258 11994
rect 14270 11942 14322 11994
rect 14334 11942 14386 11994
rect 2780 11840 2832 11892
rect 3976 11840 4028 11892
rect 4252 11840 4304 11892
rect 4436 11840 4488 11892
rect 4804 11840 4856 11892
rect 5264 11840 5316 11892
rect 5540 11840 5592 11892
rect 6092 11772 6144 11824
rect 8484 11840 8536 11892
rect 9864 11840 9916 11892
rect 10324 11883 10376 11892
rect 10324 11849 10333 11883
rect 10333 11849 10367 11883
rect 10367 11849 10376 11883
rect 10324 11840 10376 11849
rect 11796 11840 11848 11892
rect 13084 11840 13136 11892
rect 13360 11840 13412 11892
rect 10600 11772 10652 11824
rect 10968 11772 11020 11824
rect 12532 11772 12584 11824
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 3516 11704 3568 11756
rect 4804 11747 4856 11756
rect 2596 11636 2648 11688
rect 4436 11636 4488 11688
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 5816 11704 5868 11756
rect 6552 11704 6604 11756
rect 6736 11636 6788 11688
rect 8484 11704 8536 11756
rect 6828 11568 6880 11620
rect 7840 11636 7892 11688
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 9864 11704 9916 11756
rect 11336 11704 11388 11756
rect 12808 11704 12860 11756
rect 13268 11704 13320 11756
rect 13912 11747 13964 11756
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 13912 11704 13964 11713
rect 15936 11704 15988 11756
rect 12532 11636 12584 11688
rect 13176 11636 13228 11688
rect 11244 11568 11296 11620
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 5632 11500 5684 11552
rect 7564 11500 7616 11552
rect 8392 11500 8444 11552
rect 10600 11500 10652 11552
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11336 11500 11388 11552
rect 13452 11568 13504 11620
rect 14740 11611 14792 11620
rect 14740 11577 14774 11611
rect 14774 11577 14792 11611
rect 14740 11568 14792 11577
rect 12532 11500 12584 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 15200 11500 15252 11552
rect 6246 11398 6298 11450
rect 6310 11398 6362 11450
rect 6374 11398 6426 11450
rect 6438 11398 6490 11450
rect 11510 11398 11562 11450
rect 11574 11398 11626 11450
rect 11638 11398 11690 11450
rect 11702 11398 11754 11450
rect 1400 11228 1452 11280
rect 2596 11296 2648 11348
rect 9312 11296 9364 11348
rect 10876 11296 10928 11348
rect 12900 11296 12952 11348
rect 13636 11296 13688 11348
rect 3976 11228 4028 11280
rect 4620 11228 4672 11280
rect 3884 11092 3936 11144
rect 5540 11228 5592 11280
rect 6092 11228 6144 11280
rect 9772 11228 9824 11280
rect 9864 11228 9916 11280
rect 5448 11203 5500 11212
rect 5448 11169 5482 11203
rect 5482 11169 5500 11203
rect 5448 11160 5500 11169
rect 6552 11160 6604 11212
rect 2044 10956 2096 11008
rect 2136 10956 2188 11008
rect 5080 11024 5132 11076
rect 3516 10999 3568 11008
rect 3516 10965 3525 10999
rect 3525 10965 3559 10999
rect 3559 10965 3568 10999
rect 3516 10956 3568 10965
rect 6736 11092 6788 11144
rect 7104 11160 7156 11212
rect 7748 11160 7800 11212
rect 9588 11160 9640 11212
rect 10600 11160 10652 11212
rect 12532 11160 12584 11212
rect 13176 11160 13228 11212
rect 13728 11228 13780 11280
rect 13912 11203 13964 11212
rect 13912 11169 13921 11203
rect 13921 11169 13955 11203
rect 13955 11169 13964 11203
rect 13912 11160 13964 11169
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 6552 11067 6604 11076
rect 6552 11033 6561 11067
rect 6561 11033 6595 11067
rect 6595 11033 6604 11067
rect 6552 11024 6604 11033
rect 6828 11067 6880 11076
rect 6828 11033 6837 11067
rect 6837 11033 6871 11067
rect 6871 11033 6880 11067
rect 6828 11024 6880 11033
rect 8668 11092 8720 11144
rect 9220 11135 9272 11144
rect 8760 11024 8812 11076
rect 8852 11024 8904 11076
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 9956 11135 10008 11144
rect 9956 11101 9965 11135
rect 9965 11101 9999 11135
rect 9999 11101 10008 11135
rect 9956 11092 10008 11101
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 9772 11024 9824 11076
rect 12256 11024 12308 11076
rect 12532 11024 12584 11076
rect 13084 11092 13136 11144
rect 13728 11092 13780 11144
rect 14004 11135 14056 11144
rect 14004 11101 14013 11135
rect 14013 11101 14047 11135
rect 14047 11101 14056 11135
rect 14004 11092 14056 11101
rect 15292 11160 15344 11212
rect 15936 11160 15988 11212
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 13452 11024 13504 11076
rect 14556 11024 14608 11076
rect 14648 11024 14700 11076
rect 8668 10956 8720 11008
rect 10600 10956 10652 11008
rect 12900 10956 12952 11008
rect 13360 10956 13412 11008
rect 15476 11024 15528 11076
rect 15384 10999 15436 11008
rect 15384 10965 15393 10999
rect 15393 10965 15427 10999
rect 15427 10965 15436 10999
rect 15384 10956 15436 10965
rect 3614 10854 3666 10906
rect 3678 10854 3730 10906
rect 3742 10854 3794 10906
rect 3806 10854 3858 10906
rect 8878 10854 8930 10906
rect 8942 10854 8994 10906
rect 9006 10854 9058 10906
rect 9070 10854 9122 10906
rect 14142 10854 14194 10906
rect 14206 10854 14258 10906
rect 14270 10854 14322 10906
rect 14334 10854 14386 10906
rect 2596 10752 2648 10804
rect 3148 10752 3200 10804
rect 2412 10684 2464 10736
rect 5540 10752 5592 10804
rect 5632 10752 5684 10804
rect 8208 10752 8260 10804
rect 9588 10795 9640 10804
rect 9588 10761 9597 10795
rect 9597 10761 9631 10795
rect 9631 10761 9640 10795
rect 9588 10752 9640 10761
rect 4068 10684 4120 10736
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 3516 10616 3568 10668
rect 3240 10548 3292 10600
rect 4252 10548 4304 10600
rect 2780 10480 2832 10532
rect 4620 10684 4672 10736
rect 5632 10659 5684 10668
rect 4988 10548 5040 10600
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6092 10548 6144 10600
rect 6828 10616 6880 10668
rect 6736 10548 6788 10600
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 2412 10412 2464 10464
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 3516 10412 3568 10421
rect 3884 10412 3936 10464
rect 4620 10412 4672 10464
rect 4988 10455 5040 10464
rect 4988 10421 4997 10455
rect 4997 10421 5031 10455
rect 5031 10421 5040 10455
rect 4988 10412 5040 10421
rect 8116 10591 8168 10600
rect 8116 10557 8150 10591
rect 8150 10557 8168 10591
rect 8116 10548 8168 10557
rect 9496 10548 9548 10600
rect 11152 10752 11204 10804
rect 11336 10795 11388 10804
rect 11336 10761 11345 10795
rect 11345 10761 11379 10795
rect 11379 10761 11388 10795
rect 11336 10752 11388 10761
rect 10600 10684 10652 10736
rect 15660 10752 15712 10804
rect 9128 10480 9180 10532
rect 9404 10480 9456 10532
rect 6828 10412 6880 10464
rect 6920 10412 6972 10464
rect 7104 10412 7156 10464
rect 7472 10412 7524 10464
rect 9588 10412 9640 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 10600 10412 10652 10464
rect 12072 10616 12124 10668
rect 13452 10548 13504 10600
rect 13820 10548 13872 10600
rect 12072 10412 12124 10464
rect 12624 10480 12676 10532
rect 13176 10480 13228 10532
rect 15200 10523 15252 10532
rect 12808 10412 12860 10464
rect 13268 10412 13320 10464
rect 14832 10412 14884 10464
rect 15200 10489 15234 10523
rect 15234 10489 15252 10523
rect 15200 10480 15252 10489
rect 6246 10310 6298 10362
rect 6310 10310 6362 10362
rect 6374 10310 6426 10362
rect 6438 10310 6490 10362
rect 11510 10310 11562 10362
rect 11574 10310 11626 10362
rect 11638 10310 11690 10362
rect 11702 10310 11754 10362
rect 2504 10208 2556 10260
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 3240 10208 3292 10260
rect 2320 10183 2372 10192
rect 2320 10149 2329 10183
rect 2329 10149 2363 10183
rect 2363 10149 2372 10183
rect 2320 10140 2372 10149
rect 2412 10183 2464 10192
rect 2412 10149 2421 10183
rect 2421 10149 2455 10183
rect 2455 10149 2464 10183
rect 2412 10140 2464 10149
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2504 10072 2556 10124
rect 4068 10140 4120 10192
rect 4436 10140 4488 10192
rect 5448 10208 5500 10260
rect 5632 10208 5684 10260
rect 6000 10208 6052 10260
rect 7472 10208 7524 10260
rect 8116 10208 8168 10260
rect 10416 10251 10468 10260
rect 10416 10217 10425 10251
rect 10425 10217 10459 10251
rect 10459 10217 10468 10251
rect 10416 10208 10468 10217
rect 11888 10208 11940 10260
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 4344 10115 4396 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 6000 10072 6052 10124
rect 7104 10115 7156 10124
rect 7104 10081 7138 10115
rect 7138 10081 7156 10115
rect 7104 10072 7156 10081
rect 6828 10047 6880 10056
rect 3608 10004 3660 10013
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 8484 10140 8536 10192
rect 8300 10072 8352 10124
rect 9588 10072 9640 10124
rect 11428 10115 11480 10124
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 10232 10004 10284 10056
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 12808 10208 12860 10260
rect 13728 10208 13780 10260
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 15384 10208 15436 10260
rect 1584 9979 1636 9988
rect 1584 9945 1593 9979
rect 1593 9945 1627 9979
rect 1627 9945 1636 9979
rect 1584 9936 1636 9945
rect 2044 9936 2096 9988
rect 3240 9936 3292 9988
rect 3332 9936 3384 9988
rect 5632 9936 5684 9988
rect 6736 9936 6788 9988
rect 3424 9868 3476 9920
rect 4252 9868 4304 9920
rect 4988 9868 5040 9920
rect 9404 9936 9456 9988
rect 11060 10004 11112 10056
rect 15200 10140 15252 10192
rect 15752 10183 15804 10192
rect 15752 10149 15761 10183
rect 15761 10149 15795 10183
rect 15795 10149 15804 10183
rect 15752 10140 15804 10149
rect 12532 10072 12584 10124
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 14188 10004 14240 10056
rect 14280 10004 14332 10056
rect 14556 10004 14608 10056
rect 16028 10072 16080 10124
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 8668 9868 8720 9920
rect 10784 9936 10836 9988
rect 15752 9936 15804 9988
rect 9680 9868 9732 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 14924 9868 14976 9920
rect 15200 9868 15252 9920
rect 3614 9766 3666 9818
rect 3678 9766 3730 9818
rect 3742 9766 3794 9818
rect 3806 9766 3858 9818
rect 8878 9766 8930 9818
rect 8942 9766 8994 9818
rect 9006 9766 9058 9818
rect 9070 9766 9122 9818
rect 14142 9766 14194 9818
rect 14206 9766 14258 9818
rect 14270 9766 14322 9818
rect 14334 9766 14386 9818
rect 2688 9596 2740 9648
rect 3056 9639 3108 9648
rect 3056 9605 3065 9639
rect 3065 9605 3099 9639
rect 3099 9605 3108 9639
rect 3056 9596 3108 9605
rect 3240 9596 3292 9648
rect 3516 9528 3568 9580
rect 1492 9460 1544 9512
rect 2596 9460 2648 9512
rect 3056 9460 3108 9512
rect 3240 9460 3292 9512
rect 5172 9664 5224 9716
rect 5540 9664 5592 9716
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 3792 9392 3844 9444
rect 2136 9324 2188 9376
rect 3884 9324 3936 9376
rect 4528 9596 4580 9648
rect 4712 9596 4764 9648
rect 5632 9596 5684 9648
rect 6736 9596 6788 9648
rect 7104 9664 7156 9716
rect 10600 9664 10652 9716
rect 9404 9596 9456 9648
rect 12532 9664 12584 9716
rect 14556 9664 14608 9716
rect 4252 9528 4304 9580
rect 4620 9528 4672 9580
rect 4528 9324 4580 9376
rect 4620 9324 4672 9376
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 14096 9596 14148 9648
rect 14372 9596 14424 9648
rect 14740 9596 14792 9648
rect 5080 9460 5132 9512
rect 5356 9460 5408 9512
rect 5908 9460 5960 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7840 9460 7892 9512
rect 9588 9503 9640 9512
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 7196 9392 7248 9444
rect 7472 9392 7524 9444
rect 9680 9392 9732 9444
rect 9864 9435 9916 9444
rect 9864 9401 9898 9435
rect 9898 9401 9916 9435
rect 9864 9392 9916 9401
rect 10048 9392 10100 9444
rect 11612 9460 11664 9512
rect 11704 9460 11756 9512
rect 14648 9528 14700 9580
rect 15016 9528 15068 9580
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 5080 9324 5132 9376
rect 5448 9324 5500 9376
rect 5908 9324 5960 9376
rect 10232 9324 10284 9376
rect 11428 9392 11480 9444
rect 12532 9392 12584 9444
rect 15108 9503 15160 9512
rect 15108 9469 15117 9503
rect 15117 9469 15151 9503
rect 15151 9469 15160 9503
rect 15108 9460 15160 9469
rect 13176 9435 13228 9444
rect 13176 9401 13210 9435
rect 13210 9401 13228 9435
rect 13176 9392 13228 9401
rect 14004 9392 14056 9444
rect 16580 9392 16632 9444
rect 12072 9324 12124 9376
rect 12348 9324 12400 9376
rect 12716 9324 12768 9376
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 13452 9324 13504 9376
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 14740 9367 14792 9376
rect 14740 9333 14749 9367
rect 14749 9333 14783 9367
rect 14783 9333 14792 9367
rect 14740 9324 14792 9333
rect 6246 9222 6298 9274
rect 6310 9222 6362 9274
rect 6374 9222 6426 9274
rect 6438 9222 6490 9274
rect 11510 9222 11562 9274
rect 11574 9222 11626 9274
rect 11638 9222 11690 9274
rect 11702 9222 11754 9274
rect 1492 9120 1544 9172
rect 1952 9120 2004 9172
rect 2412 9120 2464 9172
rect 2688 9052 2740 9104
rect 4068 9120 4120 9172
rect 4160 9052 4212 9104
rect 4344 9052 4396 9104
rect 4712 9052 4764 9104
rect 1952 8984 2004 9036
rect 2504 8984 2556 9036
rect 4068 8984 4120 9036
rect 5632 8984 5684 9036
rect 5816 8984 5868 9036
rect 6828 9052 6880 9104
rect 8668 9052 8720 9104
rect 12624 9120 12676 9172
rect 14004 9163 14056 9172
rect 14004 9129 14013 9163
rect 14013 9129 14047 9163
rect 14047 9129 14056 9163
rect 14004 9120 14056 9129
rect 3056 8916 3108 8968
rect 5264 8916 5316 8968
rect 7840 8984 7892 9036
rect 9220 8984 9272 9036
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10232 8984 10284 9036
rect 12072 8984 12124 9036
rect 12440 8984 12492 9036
rect 14280 8984 14332 9036
rect 2872 8848 2924 8900
rect 3424 8848 3476 8900
rect 4252 8780 4304 8832
rect 5540 8780 5592 8832
rect 7196 8848 7248 8900
rect 7472 8780 7524 8832
rect 8208 8780 8260 8832
rect 9864 8916 9916 8968
rect 9956 8916 10008 8968
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10600 8916 10652 8968
rect 9680 8848 9732 8900
rect 9312 8823 9364 8832
rect 9312 8789 9321 8823
rect 9321 8789 9355 8823
rect 9355 8789 9364 8823
rect 9312 8780 9364 8789
rect 12164 8780 12216 8832
rect 13820 8916 13872 8968
rect 14004 8916 14056 8968
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 13452 8848 13504 8900
rect 12716 8780 12768 8832
rect 12992 8780 13044 8832
rect 3614 8678 3666 8730
rect 3678 8678 3730 8730
rect 3742 8678 3794 8730
rect 3806 8678 3858 8730
rect 8878 8678 8930 8730
rect 8942 8678 8994 8730
rect 9006 8678 9058 8730
rect 9070 8678 9122 8730
rect 14142 8678 14194 8730
rect 14206 8678 14258 8730
rect 14270 8678 14322 8730
rect 14334 8678 14386 8730
rect 2228 8576 2280 8628
rect 4344 8576 4396 8628
rect 4896 8576 4948 8628
rect 2872 8508 2924 8560
rect 4160 8508 4212 8560
rect 5264 8508 5316 8560
rect 2596 8440 2648 8492
rect 2780 8440 2832 8492
rect 3056 8440 3108 8492
rect 4344 8440 4396 8492
rect 6920 8440 6972 8492
rect 11888 8576 11940 8628
rect 13820 8576 13872 8628
rect 14004 8576 14056 8628
rect 9588 8508 9640 8560
rect 1952 8372 2004 8424
rect 8116 8440 8168 8492
rect 9680 8440 9732 8492
rect 7748 8372 7800 8424
rect 9220 8372 9272 8424
rect 12532 8508 12584 8560
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12716 8440 12768 8492
rect 15568 8508 15620 8560
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 12164 8372 12216 8424
rect 12624 8372 12676 8424
rect 3424 8347 3476 8356
rect 3424 8313 3458 8347
rect 3458 8313 3476 8347
rect 3424 8304 3476 8313
rect 3608 8304 3660 8356
rect 7104 8304 7156 8356
rect 7288 8304 7340 8356
rect 2412 8236 2464 8288
rect 2596 8279 2648 8288
rect 2596 8245 2605 8279
rect 2605 8245 2639 8279
rect 2639 8245 2648 8279
rect 2596 8236 2648 8245
rect 3056 8236 3108 8288
rect 5080 8236 5132 8288
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 5632 8279 5684 8288
rect 5632 8245 5641 8279
rect 5641 8245 5675 8279
rect 5675 8245 5684 8279
rect 5632 8236 5684 8245
rect 6736 8236 6788 8288
rect 7380 8236 7432 8288
rect 8944 8304 8996 8356
rect 9128 8304 9180 8356
rect 9312 8304 9364 8356
rect 12900 8304 12952 8356
rect 13452 8372 13504 8424
rect 14924 8372 14976 8424
rect 15844 8440 15896 8492
rect 13360 8304 13412 8356
rect 12072 8236 12124 8288
rect 12716 8236 12768 8288
rect 13268 8236 13320 8288
rect 15292 8304 15344 8356
rect 16212 8372 16264 8424
rect 15476 8279 15528 8288
rect 15476 8245 15485 8279
rect 15485 8245 15519 8279
rect 15519 8245 15528 8279
rect 15476 8236 15528 8245
rect 6246 8134 6298 8186
rect 6310 8134 6362 8186
rect 6374 8134 6426 8186
rect 6438 8134 6490 8186
rect 11510 8134 11562 8186
rect 11574 8134 11626 8186
rect 11638 8134 11690 8186
rect 11702 8134 11754 8186
rect 5264 8032 5316 8084
rect 5632 8032 5684 8084
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 8300 8032 8352 8084
rect 8576 8032 8628 8084
rect 9404 8032 9456 8084
rect 9588 8032 9640 8084
rect 4344 8007 4396 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 3516 7896 3568 7948
rect 4344 7973 4378 8007
rect 4378 7973 4396 8007
rect 4344 7964 4396 7973
rect 5724 7964 5776 8016
rect 8392 7964 8444 8016
rect 8760 7964 8812 8016
rect 5908 7896 5960 7948
rect 2228 7828 2280 7880
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 4068 7871 4120 7880
rect 2780 7760 2832 7812
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 6000 7828 6052 7880
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 9772 7896 9824 7948
rect 10508 8032 10560 8084
rect 10784 8032 10836 8084
rect 10968 8032 11020 8084
rect 11980 8032 12032 8084
rect 6276 7828 6328 7837
rect 8024 7828 8076 7880
rect 5080 7760 5132 7812
rect 8116 7760 8168 7812
rect 8208 7760 8260 7812
rect 8484 7828 8536 7880
rect 8944 7828 8996 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 12624 7964 12676 8016
rect 12716 7964 12768 8016
rect 14648 7964 14700 8016
rect 11704 7896 11756 7948
rect 11796 7896 11848 7948
rect 13268 7896 13320 7948
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 10324 7828 10376 7880
rect 13360 7828 13412 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 4436 7692 4488 7744
rect 5724 7735 5776 7744
rect 5724 7701 5733 7735
rect 5733 7701 5767 7735
rect 5767 7701 5776 7735
rect 5724 7692 5776 7701
rect 6184 7692 6236 7744
rect 9496 7692 9548 7744
rect 12900 7760 12952 7812
rect 13176 7760 13228 7812
rect 14464 7828 14516 7880
rect 15016 7828 15068 7880
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 13728 7760 13780 7812
rect 14832 7760 14884 7812
rect 14924 7692 14976 7744
rect 15752 7692 15804 7744
rect 3614 7590 3666 7642
rect 3678 7590 3730 7642
rect 3742 7590 3794 7642
rect 3806 7590 3858 7642
rect 8878 7590 8930 7642
rect 8942 7590 8994 7642
rect 9006 7590 9058 7642
rect 9070 7590 9122 7642
rect 14142 7590 14194 7642
rect 14206 7590 14258 7642
rect 14270 7590 14322 7642
rect 14334 7590 14386 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 3516 7488 3568 7540
rect 4344 7488 4396 7540
rect 6736 7488 6788 7540
rect 12348 7488 12400 7540
rect 13544 7488 13596 7540
rect 14648 7488 14700 7540
rect 16212 7531 16264 7540
rect 16212 7497 16221 7531
rect 16221 7497 16255 7531
rect 16255 7497 16264 7531
rect 16212 7488 16264 7497
rect 10048 7463 10100 7472
rect 10048 7429 10057 7463
rect 10057 7429 10091 7463
rect 10091 7429 10100 7463
rect 10048 7420 10100 7429
rect 11704 7463 11756 7472
rect 11704 7429 11713 7463
rect 11713 7429 11747 7463
rect 11747 7429 11756 7463
rect 11704 7420 11756 7429
rect 13176 7420 13228 7472
rect 13728 7420 13780 7472
rect 2412 7352 2464 7404
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 2228 7284 2280 7336
rect 6276 7352 6328 7404
rect 6736 7352 6788 7404
rect 12808 7352 12860 7404
rect 13360 7352 13412 7404
rect 13544 7352 13596 7404
rect 1400 7216 1452 7268
rect 3056 7216 3108 7268
rect 5448 7284 5500 7336
rect 4068 7216 4120 7268
rect 4252 7216 4304 7268
rect 6184 7284 6236 7336
rect 6920 7284 6972 7336
rect 8024 7284 8076 7336
rect 10324 7327 10376 7336
rect 10324 7293 10333 7327
rect 10333 7293 10367 7327
rect 10367 7293 10376 7327
rect 10324 7284 10376 7293
rect 756 7148 808 7200
rect 3240 7148 3292 7200
rect 3516 7148 3568 7200
rect 4528 7148 4580 7200
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 5264 7148 5316 7200
rect 6000 7148 6052 7200
rect 7380 7148 7432 7200
rect 7564 7148 7616 7200
rect 9220 7216 9272 7268
rect 9404 7216 9456 7268
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 14464 7284 14516 7336
rect 15016 7284 15068 7336
rect 16028 7327 16080 7336
rect 16028 7293 16037 7327
rect 16037 7293 16071 7327
rect 16071 7293 16080 7327
rect 16028 7284 16080 7293
rect 10784 7216 10836 7268
rect 10968 7216 11020 7268
rect 14004 7216 14056 7268
rect 10508 7148 10560 7200
rect 11152 7148 11204 7200
rect 12072 7148 12124 7200
rect 13636 7148 13688 7200
rect 14280 7148 14332 7200
rect 15844 7148 15896 7200
rect 6246 7046 6298 7098
rect 6310 7046 6362 7098
rect 6374 7046 6426 7098
rect 6438 7046 6490 7098
rect 11510 7046 11562 7098
rect 11574 7046 11626 7098
rect 11638 7046 11690 7098
rect 11702 7046 11754 7098
rect 2320 6944 2372 6996
rect 3240 6944 3292 6996
rect 1768 6808 1820 6860
rect 2504 6876 2556 6928
rect 4160 6944 4212 6996
rect 4712 6987 4764 6996
rect 4712 6953 4721 6987
rect 4721 6953 4755 6987
rect 4755 6953 4764 6987
rect 4712 6944 4764 6953
rect 5080 6944 5132 6996
rect 6736 6987 6788 6996
rect 6736 6953 6745 6987
rect 6745 6953 6779 6987
rect 6779 6953 6788 6987
rect 6736 6944 6788 6953
rect 7288 6944 7340 6996
rect 8116 6944 8168 6996
rect 10048 6944 10100 6996
rect 10692 6944 10744 6996
rect 11888 6944 11940 6996
rect 13912 6944 13964 6996
rect 14280 6944 14332 6996
rect 4252 6876 4304 6928
rect 5632 6919 5684 6928
rect 5632 6885 5666 6919
rect 5666 6885 5684 6919
rect 5632 6876 5684 6885
rect 6828 6876 6880 6928
rect 2688 6808 2740 6860
rect 6920 6808 6972 6860
rect 7104 6808 7156 6860
rect 7288 6851 7340 6860
rect 7288 6817 7322 6851
rect 7322 6817 7340 6851
rect 7288 6808 7340 6817
rect 7564 6876 7616 6928
rect 10600 6876 10652 6928
rect 11980 6876 12032 6928
rect 16028 6876 16080 6928
rect 9588 6808 9640 6860
rect 9864 6808 9916 6860
rect 11796 6808 11848 6860
rect 2504 6783 2556 6792
rect 2504 6749 2513 6783
rect 2513 6749 2547 6783
rect 2547 6749 2556 6783
rect 2504 6740 2556 6749
rect 4252 6740 4304 6792
rect 4344 6740 4396 6792
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10784 6783 10836 6792
rect 3056 6672 3108 6724
rect 8668 6715 8720 6724
rect 8668 6681 8677 6715
rect 8677 6681 8711 6715
rect 8711 6681 8720 6715
rect 8668 6672 8720 6681
rect 10784 6749 10793 6783
rect 10793 6749 10827 6783
rect 10827 6749 10836 6783
rect 10784 6740 10836 6749
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 12900 6808 12952 6860
rect 13360 6808 13412 6860
rect 14372 6808 14424 6860
rect 14924 6808 14976 6860
rect 15568 6808 15620 6860
rect 6552 6604 6604 6656
rect 7196 6604 7248 6656
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 12164 6715 12216 6724
rect 12164 6681 12173 6715
rect 12173 6681 12207 6715
rect 12207 6681 12216 6715
rect 12164 6672 12216 6681
rect 12348 6672 12400 6724
rect 13176 6740 13228 6792
rect 14004 6740 14056 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 15660 6672 15712 6724
rect 15016 6604 15068 6656
rect 15292 6647 15344 6656
rect 15292 6613 15301 6647
rect 15301 6613 15335 6647
rect 15335 6613 15344 6647
rect 15292 6604 15344 6613
rect 3614 6502 3666 6554
rect 3678 6502 3730 6554
rect 3742 6502 3794 6554
rect 3806 6502 3858 6554
rect 8878 6502 8930 6554
rect 8942 6502 8994 6554
rect 9006 6502 9058 6554
rect 9070 6502 9122 6554
rect 14142 6502 14194 6554
rect 14206 6502 14258 6554
rect 14270 6502 14322 6554
rect 14334 6502 14386 6554
rect 2504 6400 2556 6452
rect 3148 6400 3200 6452
rect 3976 6400 4028 6452
rect 4528 6400 4580 6452
rect 5448 6443 5500 6452
rect 5448 6409 5457 6443
rect 5457 6409 5491 6443
rect 5491 6409 5500 6443
rect 5448 6400 5500 6409
rect 5632 6332 5684 6384
rect 5724 6264 5776 6316
rect 6092 6332 6144 6384
rect 6828 6332 6880 6384
rect 8392 6332 8444 6384
rect 12348 6400 12400 6452
rect 12440 6400 12492 6452
rect 9220 6332 9272 6384
rect 12624 6332 12676 6384
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 2320 6196 2372 6248
rect 3148 6239 3200 6248
rect 3148 6205 3157 6239
rect 3157 6205 3191 6239
rect 3191 6205 3200 6239
rect 3148 6196 3200 6205
rect 2412 6128 2464 6180
rect 2596 6060 2648 6112
rect 2964 6060 3016 6112
rect 3884 6196 3936 6248
rect 7196 6239 7248 6248
rect 7196 6205 7230 6239
rect 7230 6205 7248 6239
rect 3976 6128 4028 6180
rect 4712 6128 4764 6180
rect 6460 6128 6512 6180
rect 7196 6196 7248 6205
rect 8484 6264 8536 6316
rect 9312 6264 9364 6316
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 11152 6264 11204 6316
rect 11336 6264 11388 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 8760 6196 8812 6248
rect 13728 6264 13780 6316
rect 12440 6196 12492 6248
rect 12716 6196 12768 6248
rect 13820 6196 13872 6248
rect 15844 6196 15896 6248
rect 6736 6128 6788 6180
rect 4344 6060 4396 6112
rect 5724 6060 5776 6112
rect 8208 6060 8260 6112
rect 8392 6060 8444 6112
rect 9312 6060 9364 6112
rect 9772 6060 9824 6112
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 11336 6060 11388 6112
rect 12624 6060 12676 6112
rect 13452 6060 13504 6112
rect 13912 6060 13964 6112
rect 15844 6060 15896 6112
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 6246 5958 6298 6010
rect 6310 5958 6362 6010
rect 6374 5958 6426 6010
rect 6438 5958 6490 6010
rect 11510 5958 11562 6010
rect 11574 5958 11626 6010
rect 11638 5958 11690 6010
rect 11702 5958 11754 6010
rect 4068 5856 4120 5908
rect 7564 5856 7616 5908
rect 9772 5856 9824 5908
rect 10508 5856 10560 5908
rect 10692 5856 10744 5908
rect 10968 5856 11020 5908
rect 11152 5856 11204 5908
rect 12440 5856 12492 5908
rect 12624 5856 12676 5908
rect 15384 5856 15436 5908
rect 16396 5856 16448 5908
rect 4344 5788 4396 5840
rect 9680 5788 9732 5840
rect 13268 5831 13320 5840
rect 1676 5720 1728 5772
rect 2320 5763 2372 5772
rect 2320 5729 2329 5763
rect 2329 5729 2363 5763
rect 2363 5729 2372 5763
rect 2320 5720 2372 5729
rect 2596 5763 2648 5772
rect 2596 5729 2630 5763
rect 2630 5729 2648 5763
rect 2596 5720 2648 5729
rect 4252 5720 4304 5772
rect 4896 5695 4948 5704
rect 4896 5661 4905 5695
rect 4905 5661 4939 5695
rect 4939 5661 4948 5695
rect 4896 5652 4948 5661
rect 5724 5763 5776 5772
rect 5724 5729 5758 5763
rect 5758 5729 5776 5763
rect 5724 5720 5776 5729
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 7656 5720 7708 5772
rect 8024 5763 8076 5772
rect 8024 5729 8033 5763
rect 8033 5729 8067 5763
rect 8067 5729 8076 5763
rect 8024 5720 8076 5729
rect 10048 5763 10100 5772
rect 7196 5652 7248 5704
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 7932 5584 7984 5636
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10416 5720 10468 5772
rect 9312 5652 9364 5704
rect 10140 5652 10192 5704
rect 11060 5720 11112 5772
rect 11704 5720 11756 5772
rect 13268 5797 13277 5831
rect 13277 5797 13311 5831
rect 13311 5797 13320 5831
rect 13268 5788 13320 5797
rect 13360 5720 13412 5772
rect 11336 5652 11388 5704
rect 13544 5652 13596 5704
rect 14464 5652 14516 5704
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 9220 5584 9272 5636
rect 11428 5584 11480 5636
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 3240 5516 3292 5568
rect 3976 5516 4028 5568
rect 6736 5516 6788 5568
rect 6828 5559 6880 5568
rect 6828 5525 6837 5559
rect 6837 5525 6871 5559
rect 6871 5525 6880 5559
rect 6828 5516 6880 5525
rect 7104 5516 7156 5568
rect 9680 5516 9732 5568
rect 12348 5516 12400 5568
rect 13544 5516 13596 5568
rect 15384 5559 15436 5568
rect 15384 5525 15393 5559
rect 15393 5525 15427 5559
rect 15427 5525 15436 5559
rect 15384 5516 15436 5525
rect 3614 5414 3666 5466
rect 3678 5414 3730 5466
rect 3742 5414 3794 5466
rect 3806 5414 3858 5466
rect 8878 5414 8930 5466
rect 8942 5414 8994 5466
rect 9006 5414 9058 5466
rect 9070 5414 9122 5466
rect 14142 5414 14194 5466
rect 14206 5414 14258 5466
rect 14270 5414 14322 5466
rect 14334 5414 14386 5466
rect 4160 5312 4212 5364
rect 5632 5355 5684 5364
rect 2412 5176 2464 5228
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 4252 5219 4304 5228
rect 4252 5185 4261 5219
rect 4261 5185 4295 5219
rect 4295 5185 4304 5219
rect 4252 5176 4304 5185
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 8024 5312 8076 5364
rect 11704 5355 11756 5364
rect 11704 5321 11713 5355
rect 11713 5321 11747 5355
rect 11747 5321 11756 5355
rect 11704 5312 11756 5321
rect 12440 5312 12492 5364
rect 13360 5312 13412 5364
rect 13728 5312 13780 5364
rect 5540 5244 5592 5296
rect 6920 5244 6972 5296
rect 3332 5108 3384 5160
rect 2504 5040 2556 5092
rect 5632 5108 5684 5160
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 4804 5040 4856 5092
rect 5448 5040 5500 5092
rect 3424 4972 3476 5024
rect 4068 4972 4120 5024
rect 6000 4972 6052 5024
rect 7288 5176 7340 5228
rect 11428 5244 11480 5296
rect 14924 5312 14976 5364
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 12900 5176 12952 5228
rect 6736 5108 6788 5160
rect 9496 5151 9548 5160
rect 9496 5117 9505 5151
rect 9505 5117 9539 5151
rect 9539 5117 9548 5151
rect 9496 5108 9548 5117
rect 6552 5040 6604 5092
rect 8208 5040 8260 5092
rect 10048 5108 10100 5160
rect 12072 5108 12124 5160
rect 12532 5108 12584 5160
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 9956 5040 10008 5092
rect 12624 5040 12676 5092
rect 13728 5040 13780 5092
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 11980 5015 12032 5024
rect 11980 4981 11989 5015
rect 11989 4981 12023 5015
rect 12023 4981 12032 5015
rect 11980 4972 12032 4981
rect 12532 4972 12584 5024
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 14464 5151 14516 5160
rect 14464 5117 14498 5151
rect 14498 5117 14516 5151
rect 14464 5108 14516 5117
rect 15016 5040 15068 5092
rect 6246 4870 6298 4922
rect 6310 4870 6362 4922
rect 6374 4870 6426 4922
rect 6438 4870 6490 4922
rect 11510 4870 11562 4922
rect 11574 4870 11626 4922
rect 11638 4870 11690 4922
rect 11702 4870 11754 4922
rect 2412 4768 2464 4820
rect 2688 4700 2740 4752
rect 3240 4768 3292 4820
rect 6920 4768 6972 4820
rect 11888 4768 11940 4820
rect 11980 4768 12032 4820
rect 12624 4768 12676 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 15292 4768 15344 4820
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 8024 4700 8076 4752
rect 1400 4632 1452 4684
rect 2320 4632 2372 4684
rect 2872 4632 2924 4684
rect 3056 4632 3108 4684
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 4344 4675 4396 4684
rect 4344 4641 4378 4675
rect 4378 4641 4396 4675
rect 5816 4675 5868 4684
rect 4344 4632 4396 4641
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6828 4675 6880 4684
rect 6828 4641 6862 4675
rect 6862 4641 6880 4675
rect 6828 4632 6880 4641
rect 7104 4632 7156 4684
rect 9220 4700 9272 4752
rect 8668 4632 8720 4684
rect 9772 4632 9824 4684
rect 10324 4632 10376 4684
rect 8300 4564 8352 4616
rect 9128 4564 9180 4616
rect 9404 4564 9456 4616
rect 6552 4496 6604 4548
rect 8208 4539 8260 4548
rect 8208 4505 8217 4539
rect 8217 4505 8251 4539
rect 8251 4505 8260 4539
rect 8208 4496 8260 4505
rect 12900 4632 12952 4684
rect 14004 4632 14056 4684
rect 14832 4632 14884 4684
rect 11336 4564 11388 4616
rect 13084 4564 13136 4616
rect 14464 4564 14516 4616
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 3516 4471 3568 4480
rect 3516 4437 3525 4471
rect 3525 4437 3559 4471
rect 3559 4437 3568 4471
rect 3516 4428 3568 4437
rect 4804 4428 4856 4480
rect 6460 4428 6512 4480
rect 10876 4428 10928 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 12348 4428 12400 4480
rect 14924 4496 14976 4548
rect 14832 4471 14884 4480
rect 14832 4437 14841 4471
rect 14841 4437 14875 4471
rect 14875 4437 14884 4471
rect 14832 4428 14884 4437
rect 15752 4428 15804 4480
rect 3614 4326 3666 4378
rect 3678 4326 3730 4378
rect 3742 4326 3794 4378
rect 3806 4326 3858 4378
rect 8878 4326 8930 4378
rect 8942 4326 8994 4378
rect 9006 4326 9058 4378
rect 9070 4326 9122 4378
rect 14142 4326 14194 4378
rect 14206 4326 14258 4378
rect 14270 4326 14322 4378
rect 14334 4326 14386 4378
rect 6736 4224 6788 4276
rect 2412 4156 2464 4208
rect 2596 4156 2648 4208
rect 2688 4088 2740 4140
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 4988 4088 5040 4140
rect 6460 4156 6512 4208
rect 6920 4156 6972 4208
rect 7104 4156 7156 4208
rect 2228 3927 2280 3936
rect 2228 3893 2237 3927
rect 2237 3893 2271 3927
rect 2271 3893 2280 3927
rect 4160 4020 4212 4072
rect 4896 4020 4948 4072
rect 7288 4088 7340 4140
rect 9220 4156 9272 4208
rect 10600 4199 10652 4208
rect 10600 4165 10609 4199
rect 10609 4165 10643 4199
rect 10643 4165 10652 4199
rect 10600 4156 10652 4165
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12072 4088 12124 4140
rect 12900 4088 12952 4140
rect 15844 4156 15896 4208
rect 13268 4088 13320 4140
rect 14096 4131 14148 4140
rect 14096 4097 14105 4131
rect 14105 4097 14139 4131
rect 14139 4097 14148 4131
rect 14096 4088 14148 4097
rect 14464 4088 14516 4140
rect 15476 4088 15528 4140
rect 8760 4020 8812 4072
rect 9772 4020 9824 4072
rect 10232 4020 10284 4072
rect 10876 4020 10928 4072
rect 11336 4020 11388 4072
rect 11980 4020 12032 4072
rect 15200 4020 15252 4072
rect 15384 4020 15436 4072
rect 2228 3884 2280 3893
rect 3056 3884 3108 3936
rect 4344 3952 4396 4004
rect 5540 3952 5592 4004
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 4068 3884 4120 3936
rect 4528 3884 4580 3936
rect 5816 3884 5868 3936
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7564 3927 7616 3936
rect 7564 3893 7573 3927
rect 7573 3893 7607 3927
rect 7607 3893 7616 3927
rect 7564 3884 7616 3893
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 8208 3927 8260 3936
rect 7656 3884 7708 3893
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 8300 3884 8352 3936
rect 9404 3952 9456 4004
rect 11152 3952 11204 4004
rect 12072 3952 12124 4004
rect 9772 3884 9824 3936
rect 10968 3884 11020 3936
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 12624 3884 12676 3936
rect 13360 3884 13412 3936
rect 13452 3927 13504 3936
rect 13452 3893 13461 3927
rect 13461 3893 13495 3927
rect 13495 3893 13504 3927
rect 13820 3927 13872 3936
rect 13452 3884 13504 3893
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 15660 3884 15712 3936
rect 6246 3782 6298 3834
rect 6310 3782 6362 3834
rect 6374 3782 6426 3834
rect 6438 3782 6490 3834
rect 11510 3782 11562 3834
rect 11574 3782 11626 3834
rect 11638 3782 11690 3834
rect 11702 3782 11754 3834
rect 1952 3680 2004 3732
rect 2228 3680 2280 3732
rect 4436 3680 4488 3732
rect 5080 3680 5132 3732
rect 5816 3680 5868 3732
rect 5908 3723 5960 3732
rect 5908 3689 5917 3723
rect 5917 3689 5951 3723
rect 5951 3689 5960 3723
rect 5908 3680 5960 3689
rect 3792 3612 3844 3664
rect 5264 3612 5316 3664
rect 5448 3612 5500 3664
rect 6736 3680 6788 3732
rect 7196 3680 7248 3732
rect 7656 3680 7708 3732
rect 8208 3680 8260 3732
rect 10968 3723 11020 3732
rect 8392 3612 8444 3664
rect 10508 3612 10560 3664
rect 10968 3689 10977 3723
rect 10977 3689 11011 3723
rect 11011 3689 11020 3723
rect 10968 3680 11020 3689
rect 12624 3723 12676 3732
rect 12624 3689 12633 3723
rect 12633 3689 12667 3723
rect 12667 3689 12676 3723
rect 12624 3680 12676 3689
rect 14464 3680 14516 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 15752 3723 15804 3732
rect 15752 3689 15761 3723
rect 15761 3689 15795 3723
rect 15795 3689 15804 3723
rect 15752 3680 15804 3689
rect 12348 3612 12400 3664
rect 12532 3655 12584 3664
rect 12532 3621 12541 3655
rect 12541 3621 12575 3655
rect 12575 3621 12584 3655
rect 12532 3612 12584 3621
rect 13820 3612 13872 3664
rect 14096 3612 14148 3664
rect 1676 3476 1728 3528
rect 4712 3544 4764 3596
rect 5632 3544 5684 3596
rect 5816 3544 5868 3596
rect 7104 3544 7156 3596
rect 3056 3476 3108 3528
rect 3332 3519 3384 3528
rect 3332 3485 3341 3519
rect 3341 3485 3375 3519
rect 3375 3485 3384 3519
rect 3332 3476 3384 3485
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 1860 3408 1912 3460
rect 5448 3476 5500 3528
rect 6460 3476 6512 3528
rect 8484 3544 8536 3596
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10876 3544 10928 3596
rect 11980 3544 12032 3596
rect 7288 3476 7340 3528
rect 7748 3476 7800 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9404 3476 9456 3528
rect 10416 3476 10468 3528
rect 11704 3476 11756 3528
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 13176 3519 13228 3528
rect 13176 3485 13185 3519
rect 13185 3485 13219 3519
rect 13219 3485 13228 3519
rect 13176 3476 13228 3485
rect 14924 3476 14976 3528
rect 2228 3340 2280 3392
rect 3516 3340 3568 3392
rect 6000 3408 6052 3460
rect 7840 3408 7892 3460
rect 11152 3408 11204 3460
rect 5080 3340 5132 3392
rect 5540 3383 5592 3392
rect 5540 3349 5549 3383
rect 5549 3349 5583 3383
rect 5583 3349 5592 3383
rect 5540 3340 5592 3349
rect 5632 3340 5684 3392
rect 8300 3340 8352 3392
rect 10692 3340 10744 3392
rect 11980 3340 12032 3392
rect 13544 3340 13596 3392
rect 15108 3340 15160 3392
rect 3614 3238 3666 3290
rect 3678 3238 3730 3290
rect 3742 3238 3794 3290
rect 3806 3238 3858 3290
rect 8878 3238 8930 3290
rect 8942 3238 8994 3290
rect 9006 3238 9058 3290
rect 9070 3238 9122 3290
rect 14142 3238 14194 3290
rect 14206 3238 14258 3290
rect 14270 3238 14322 3290
rect 14334 3238 14386 3290
rect 480 3136 532 3188
rect 3332 3136 3384 3188
rect 4160 3179 4212 3188
rect 4160 3145 4169 3179
rect 4169 3145 4203 3179
rect 4203 3145 4212 3179
rect 4160 3136 4212 3145
rect 4712 3068 4764 3120
rect 6644 3136 6696 3188
rect 7840 3136 7892 3188
rect 7288 3068 7340 3120
rect 7932 3068 7984 3120
rect 9588 3136 9640 3188
rect 9864 3136 9916 3188
rect 10140 3136 10192 3188
rect 10508 3136 10560 3188
rect 11704 3179 11756 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 4252 3000 4304 3052
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 5172 3000 5224 3052
rect 5540 3000 5592 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 5816 3000 5868 3052
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 4988 2932 5040 2984
rect 5632 2975 5684 2984
rect 5632 2941 5641 2975
rect 5641 2941 5675 2975
rect 5675 2941 5684 2975
rect 5632 2932 5684 2941
rect 7380 2932 7432 2984
rect 7932 2932 7984 2984
rect 1400 2796 1452 2848
rect 5080 2864 5132 2916
rect 6000 2864 6052 2916
rect 10324 3068 10376 3120
rect 11704 3145 11713 3179
rect 11713 3145 11747 3179
rect 11747 3145 11756 3179
rect 11704 3136 11756 3145
rect 12256 3068 12308 3120
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 9220 3000 9272 3052
rect 13360 3136 13412 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 14464 3068 14516 3120
rect 8576 2932 8628 2984
rect 9496 2932 9548 2984
rect 9772 2932 9824 2984
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 9404 2864 9456 2916
rect 10232 2932 10284 2984
rect 10600 2975 10652 2984
rect 10600 2941 10634 2975
rect 10634 2941 10652 2975
rect 10600 2932 10652 2941
rect 13452 3000 13504 3052
rect 14740 3000 14792 3052
rect 8760 2839 8812 2848
rect 8760 2805 8769 2839
rect 8769 2805 8803 2839
rect 8803 2805 8812 2839
rect 9772 2839 9824 2848
rect 8760 2796 8812 2805
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 11060 2864 11112 2916
rect 12072 2864 12124 2916
rect 14004 2932 14056 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 17500 3000 17552 3052
rect 13176 2864 13228 2916
rect 13912 2864 13964 2916
rect 14924 2864 14976 2916
rect 15660 2864 15712 2916
rect 6246 2694 6298 2746
rect 6310 2694 6362 2746
rect 6374 2694 6426 2746
rect 6438 2694 6490 2746
rect 11510 2694 11562 2746
rect 11574 2694 11626 2746
rect 11638 2694 11690 2746
rect 11702 2694 11754 2746
rect 4068 2592 4120 2644
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 4988 2592 5040 2601
rect 5172 2592 5224 2644
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 8760 2592 8812 2644
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 10416 2635 10468 2644
rect 9128 2592 9180 2601
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 10692 2592 10744 2644
rect 11336 2592 11388 2644
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 13544 2592 13596 2644
rect 3700 2524 3752 2576
rect 4712 2524 4764 2576
rect 5356 2567 5408 2576
rect 5356 2533 5365 2567
rect 5365 2533 5399 2567
rect 5399 2533 5408 2567
rect 5356 2524 5408 2533
rect 5540 2524 5592 2576
rect 10324 2524 10376 2576
rect 11152 2524 11204 2576
rect 12256 2524 12308 2576
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 4160 2456 4212 2508
rect 4620 2456 4672 2508
rect 6092 2499 6144 2508
rect 6092 2465 6101 2499
rect 6101 2465 6135 2499
rect 6135 2465 6144 2499
rect 6092 2456 6144 2465
rect 7196 2456 7248 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 12348 2456 12400 2508
rect 12808 2524 12860 2576
rect 3240 2388 3292 2440
rect 4436 2388 4488 2440
rect 4712 2388 4764 2440
rect 5448 2388 5500 2440
rect 7104 2388 7156 2440
rect 7472 2388 7524 2440
rect 7932 2388 7984 2440
rect 6092 2320 6144 2372
rect 8484 2388 8536 2440
rect 10600 2388 10652 2440
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 11704 2320 11756 2372
rect 11796 2320 11848 2372
rect 13360 2388 13412 2440
rect 14648 2388 14700 2440
rect 2780 2252 2832 2304
rect 4896 2252 4948 2304
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 13820 2320 13872 2372
rect 14556 2320 14608 2372
rect 14924 2252 14976 2304
rect 15016 2295 15068 2304
rect 15016 2261 15025 2295
rect 15025 2261 15059 2295
rect 15059 2261 15068 2295
rect 15016 2252 15068 2261
rect 3614 2150 3666 2202
rect 3678 2150 3730 2202
rect 3742 2150 3794 2202
rect 3806 2150 3858 2202
rect 8878 2150 8930 2202
rect 8942 2150 8994 2202
rect 9006 2150 9058 2202
rect 9070 2150 9122 2202
rect 14142 2150 14194 2202
rect 14206 2150 14258 2202
rect 14270 2150 14322 2202
rect 14334 2150 14386 2202
rect 2504 2048 2556 2100
rect 9772 2048 9824 2100
rect 2320 1436 2372 1488
rect 9404 1436 9456 1488
rect 3700 1028 3752 1080
rect 8208 1028 8260 1080
<< metal2 >>
rect 3514 16688 3570 16697
rect 3514 16623 3570 16632
rect 16394 16688 16450 16697
rect 16394 16623 16450 16632
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1320 9353 1348 15399
rect 2042 14648 2098 14657
rect 2042 14583 2098 14592
rect 1858 12744 1914 12753
rect 1858 12679 1914 12688
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1780 12442 1808 12582
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1872 12288 1900 12679
rect 1780 12260 1900 12288
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1400 11280 1452 11286
rect 1400 11222 1452 11228
rect 1412 10674 1440 11222
rect 1400 10668 1452 10674
rect 1452 10628 1532 10656
rect 1400 10610 1452 10616
rect 1398 10160 1454 10169
rect 1398 10095 1400 10104
rect 1452 10095 1454 10104
rect 1400 10066 1452 10072
rect 1504 9518 1532 10628
rect 1596 10577 1624 12038
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1582 10024 1638 10033
rect 1582 9959 1584 9968
rect 1636 9959 1638 9968
rect 1584 9930 1636 9936
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1504 9178 1532 9454
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1674 8392 1730 8401
rect 1674 8327 1730 8336
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7274 1440 7890
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1400 7268 1452 7274
rect 1400 7210 1452 7216
rect 756 7200 808 7206
rect 1596 7177 1624 7278
rect 756 7142 808 7148
rect 1582 7168 1638 7177
rect 480 3188 532 3194
rect 480 3130 532 3136
rect 492 480 520 3130
rect 768 1465 796 7142
rect 1582 7103 1638 7112
rect 1688 5778 1716 8327
rect 1780 6866 1808 12260
rect 2056 12186 2084 14583
rect 3238 14240 3294 14249
rect 3238 14175 3294 14184
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2148 12442 2176 13126
rect 2240 12782 2268 13670
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 1964 12158 2084 12186
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 9897 1900 11494
rect 1858 9888 1914 9897
rect 1858 9823 1914 9832
rect 1964 9178 1992 12158
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2148 11014 2176 11698
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2056 9994 2084 10950
rect 2044 9988 2096 9994
rect 2044 9930 2096 9936
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1964 8430 1992 8978
rect 2148 8673 2176 9318
rect 2134 8664 2190 8673
rect 2240 8634 2268 12582
rect 2318 12064 2374 12073
rect 2318 11999 2374 12008
rect 2332 10724 2360 11999
rect 2412 10736 2464 10742
rect 2332 10696 2412 10724
rect 2332 10198 2360 10696
rect 2412 10678 2464 10684
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10198 2452 10406
rect 2516 10266 2544 13330
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2608 12442 2636 13262
rect 2700 12850 2728 13262
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2608 11694 2636 12106
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 11354 2636 11630
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9489 2544 10066
rect 2608 10062 2636 10746
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2608 9518 2636 9998
rect 2700 9654 2728 12786
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 11898 2820 12582
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2688 9648 2740 9654
rect 2688 9590 2740 9596
rect 2596 9512 2648 9518
rect 2502 9480 2558 9489
rect 2596 9454 2648 9460
rect 2502 9415 2558 9424
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2134 8599 2190 8608
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 2424 8294 2452 9114
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1768 6860 1820 6866
rect 1820 6820 1900 6848
rect 1768 6802 1820 6808
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 3058 1440 4626
rect 1780 3641 1808 5510
rect 1766 3632 1822 3641
rect 1766 3567 1822 3576
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 754 1456 810 1465
rect 754 1391 810 1400
rect 1412 480 1440 2790
rect 1688 2514 1716 3470
rect 1872 3466 1900 6820
rect 1964 3738 1992 7686
rect 2240 7546 2268 7822
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2240 6236 2268 7278
rect 2332 7002 2360 7890
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2424 6746 2452 7346
rect 2516 6934 2544 8978
rect 2608 8498 2636 9454
rect 2700 9110 2728 9590
rect 2688 9104 2740 9110
rect 2792 9081 2820 10474
rect 2688 9046 2740 9052
rect 2778 9072 2834 9081
rect 2778 9007 2834 9016
rect 2884 8906 2912 12174
rect 2976 10266 3004 12242
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2962 9752 3018 9761
rect 2962 9687 3018 9696
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2594 8392 2650 8401
rect 2594 8327 2650 8336
rect 2608 8294 2636 8327
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2792 7970 2820 8434
rect 2700 7942 2820 7970
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2504 6792 2556 6798
rect 2424 6740 2504 6746
rect 2424 6734 2556 6740
rect 2424 6718 2544 6734
rect 2320 6248 2372 6254
rect 2240 6208 2320 6236
rect 2320 6190 2372 6196
rect 2332 5778 2360 6190
rect 2424 6186 2452 6718
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2412 6180 2464 6186
rect 2412 6122 2464 6128
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2332 4690 2360 5714
rect 2424 5234 2452 6122
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2424 4826 2452 5170
rect 2516 5098 2544 6394
rect 2608 6118 2636 7822
rect 2700 6866 2728 7942
rect 2780 7812 2832 7818
rect 2780 7754 2832 7760
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2608 5778 2636 6054
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2424 4214 2452 4762
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3738 2268 3878
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 2514 2268 3334
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2516 2106 2544 5034
rect 2608 4214 2636 5714
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 2700 4146 2728 4694
rect 2792 4457 2820 7754
rect 2884 4865 2912 8502
rect 2976 6497 3004 9687
rect 3068 9654 3096 12242
rect 3160 12238 3188 13874
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3160 10810 3188 12174
rect 3252 11801 3280 14175
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3238 11792 3294 11801
rect 3238 11727 3294 11736
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3146 10432 3202 10441
rect 3146 10367 3202 10376
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3068 9217 3096 9454
rect 3054 9208 3110 9217
rect 3054 9143 3110 9152
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3068 8498 3096 8910
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 3068 7274 3096 8230
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2962 6488 3018 6497
rect 2962 6423 3018 6432
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2870 4856 2926 4865
rect 2870 4791 2926 4800
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2778 4448 2834 4457
rect 2778 4383 2834 4392
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2504 2100 2556 2106
rect 2504 2042 2556 2048
rect 2320 1488 2372 1494
rect 2320 1430 2372 1436
rect 2332 480 2360 1430
rect 478 0 534 480
rect 1398 0 1454 480
rect 2318 0 2374 480
rect 2792 241 2820 2246
rect 2884 649 2912 4626
rect 2976 1873 3004 6054
rect 3068 4690 3096 6666
rect 3160 6458 3188 10367
rect 3252 10305 3280 10542
rect 3238 10296 3294 10305
rect 3238 10231 3240 10240
rect 3292 10231 3294 10240
rect 3240 10202 3292 10208
rect 3252 10171 3280 10202
rect 3238 10024 3294 10033
rect 3344 9994 3372 13670
rect 3422 12744 3478 12753
rect 3422 12679 3424 12688
rect 3476 12679 3478 12688
rect 3424 12650 3476 12656
rect 3528 11762 3556 16623
rect 4066 16280 4122 16289
rect 4066 16215 4122 16224
rect 14922 16280 14978 16289
rect 14922 16215 14978 16224
rect 4080 15230 4108 16215
rect 4894 15872 4950 15881
rect 4894 15807 4950 15816
rect 4068 15224 4120 15230
rect 4068 15166 4120 15172
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4080 14278 4108 14991
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3588 14172 3884 14192
rect 3644 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3666 14118 3668 14170
rect 3730 14118 3742 14170
rect 3804 14118 3806 14170
rect 3644 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3588 14096 3884 14116
rect 3976 13864 4028 13870
rect 3974 13832 3976 13841
rect 4028 13832 4030 13841
rect 4908 13802 4936 15807
rect 14462 15464 14518 15473
rect 14462 15399 14518 15408
rect 8944 15224 8996 15230
rect 8944 15166 8996 15172
rect 9312 15224 9364 15230
rect 9312 15166 9364 15172
rect 6220 14716 6516 14736
rect 6276 14714 6300 14716
rect 6356 14714 6380 14716
rect 6436 14714 6460 14716
rect 6298 14662 6300 14714
rect 6362 14662 6374 14714
rect 6436 14662 6438 14714
rect 6276 14660 6300 14662
rect 6356 14660 6380 14662
rect 6436 14660 6460 14662
rect 6220 14640 6516 14660
rect 8956 14618 8984 15166
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 14006 5580 14214
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 3974 13767 4030 13776
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 3588 13084 3884 13104
rect 3644 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3666 13030 3668 13082
rect 3730 13030 3742 13082
rect 3804 13030 3806 13082
rect 3644 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3588 13008 3884 13028
rect 4160 12912 4212 12918
rect 4448 12889 4476 13126
rect 4160 12854 4212 12860
rect 4434 12880 4490 12889
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3588 11996 3884 12016
rect 3644 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3666 11942 3668 11994
rect 3730 11942 3742 11994
rect 3804 11942 3806 11994
rect 3644 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3588 11920 3884 11940
rect 3988 11898 4016 12786
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3882 11656 3938 11665
rect 3882 11591 3938 11600
rect 3896 11150 3924 11591
rect 3988 11286 4016 11834
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3528 10674 3556 10950
rect 3588 10908 3884 10928
rect 3644 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3666 10854 3668 10906
rect 3730 10854 3742 10906
rect 3804 10854 3806 10906
rect 3644 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3588 10832 3884 10852
rect 4080 10742 4108 12582
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3516 10668 3568 10674
rect 3568 10628 3648 10656
rect 3516 10610 3568 10616
rect 3516 10464 3568 10470
rect 3514 10432 3516 10441
rect 3568 10432 3570 10441
rect 3514 10367 3570 10376
rect 3620 10062 3648 10628
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 10112 3924 10406
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 3896 10084 4016 10112
rect 3608 10056 3660 10062
rect 3528 10016 3608 10044
rect 3238 9959 3240 9968
rect 3292 9959 3294 9968
rect 3332 9988 3384 9994
rect 3240 9930 3292 9936
rect 3332 9930 3384 9936
rect 3424 9920 3476 9926
rect 3330 9888 3386 9897
rect 3424 9862 3476 9868
rect 3330 9823 3386 9832
rect 3238 9752 3294 9761
rect 3238 9687 3294 9696
rect 3252 9654 3280 9687
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3252 9353 3280 9454
rect 3238 9344 3294 9353
rect 3238 9279 3294 9288
rect 3252 7206 3280 9279
rect 3344 7426 3372 9823
rect 3436 9024 3464 9862
rect 3528 9586 3556 10016
rect 3608 9998 3660 10004
rect 3588 9820 3884 9840
rect 3644 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3666 9766 3668 9818
rect 3730 9766 3742 9818
rect 3804 9766 3806 9818
rect 3644 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3588 9744 3884 9764
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3804 9353 3832 9386
rect 3884 9376 3936 9382
rect 3790 9344 3846 9353
rect 3884 9318 3936 9324
rect 3790 9279 3846 9288
rect 3436 8996 3556 9024
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3436 8362 3464 8842
rect 3424 8356 3476 8362
rect 3528 8344 3556 8996
rect 3896 8945 3924 9318
rect 3882 8936 3938 8945
rect 3882 8871 3938 8880
rect 3588 8732 3884 8752
rect 3644 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3666 8678 3668 8730
rect 3730 8678 3742 8730
rect 3804 8678 3806 8730
rect 3644 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3588 8656 3884 8676
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3608 8356 3660 8362
rect 3528 8316 3608 8344
rect 3424 8298 3476 8304
rect 3608 8298 3660 8304
rect 3514 7984 3570 7993
rect 3514 7919 3516 7928
rect 3568 7919 3570 7928
rect 3516 7890 3568 7896
rect 3896 7732 3924 8463
rect 3988 7857 4016 10084
rect 4080 9897 4108 10134
rect 4066 9888 4122 9897
rect 4066 9823 4122 9832
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 9178 4108 9454
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4172 9110 4200 12854
rect 4434 12815 4490 12824
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4264 11898 4292 12582
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4264 9926 4292 10542
rect 4356 10130 4384 12038
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4448 11694 4476 11834
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4080 8673 4108 8978
rect 4264 8838 4292 9522
rect 4356 9353 4384 10066
rect 4342 9344 4398 9353
rect 4342 9279 4398 9288
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4066 8664 4122 8673
rect 4356 8634 4384 9046
rect 4066 8599 4122 8608
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 4172 8106 4200 8502
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4172 8078 4292 8106
rect 4158 7984 4214 7993
rect 4158 7919 4214 7928
rect 4068 7880 4120 7886
rect 3974 7848 4030 7857
rect 4068 7822 4120 7828
rect 3974 7783 4030 7792
rect 3896 7704 4016 7732
rect 3588 7644 3884 7664
rect 3644 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3666 7590 3668 7642
rect 3730 7590 3742 7642
rect 3804 7590 3806 7642
rect 3644 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3588 7568 3884 7588
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3528 7449 3556 7482
rect 3514 7440 3570 7449
rect 3344 7398 3464 7426
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3252 6905 3280 6938
rect 3238 6896 3294 6905
rect 3238 6831 3294 6840
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3146 6352 3202 6361
rect 3146 6287 3202 6296
rect 3160 6254 3188 6287
rect 3148 6248 3200 6254
rect 3200 6208 3372 6236
rect 3148 6190 3200 6196
rect 3240 5568 3292 5574
rect 3160 5516 3240 5522
rect 3160 5510 3292 5516
rect 3160 5494 3280 5510
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3641 3096 3878
rect 3054 3632 3110 3641
rect 3054 3567 3110 3576
rect 3056 3528 3108 3534
rect 3160 3516 3188 5494
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3252 4826 3280 5170
rect 3344 5166 3372 6208
rect 3332 5160 3384 5166
rect 3436 5137 3464 7398
rect 3514 7375 3570 7384
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 7041 3556 7142
rect 3514 7032 3570 7041
rect 3514 6967 3570 6976
rect 3588 6556 3884 6576
rect 3644 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3666 6502 3668 6554
rect 3730 6502 3742 6554
rect 3804 6502 3806 6554
rect 3644 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3588 6480 3884 6500
rect 3988 6458 4016 7704
rect 4080 7274 4108 7822
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4172 7002 4200 7919
rect 4264 7449 4292 8078
rect 4356 8022 4384 8434
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4356 7546 4384 7958
rect 4448 7750 4476 10134
rect 4540 9654 4568 13670
rect 5092 13326 5120 13874
rect 5172 13728 5224 13734
rect 5170 13696 5172 13705
rect 5724 13728 5776 13734
rect 5224 13696 5226 13705
rect 5724 13670 5776 13676
rect 5170 13631 5226 13640
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4632 11286 4660 12310
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4632 10470 4660 10678
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4632 9586 4660 10406
rect 4724 9654 4752 12922
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4816 11898 4844 12038
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4816 11762 4844 11834
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 5092 11082 5120 13262
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12782 5212 13126
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5172 12776 5224 12782
rect 5368 12753 5396 12854
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5172 12718 5224 12724
rect 5354 12744 5410 12753
rect 5354 12679 5410 12688
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5276 11898 5304 12582
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5092 10792 5120 11018
rect 5092 10764 5304 10792
rect 5078 10704 5134 10713
rect 5078 10639 5134 10648
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 5000 10470 5028 10542
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4894 9752 4950 9761
rect 4894 9687 4950 9696
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4710 9344 4766 9353
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4250 7440 4306 7449
rect 4250 7375 4306 7384
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4264 6934 4292 7210
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4356 6798 4384 7482
rect 4540 7206 4568 9318
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4252 6792 4304 6798
rect 4250 6760 4252 6769
rect 4344 6792 4396 6798
rect 4304 6760 4306 6769
rect 4344 6734 4396 6740
rect 4250 6695 4306 6704
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3896 6089 3924 6190
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3882 6080 3938 6089
rect 3882 6015 3938 6024
rect 3988 5574 4016 6122
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4080 5681 4108 5850
rect 4264 5778 4292 6695
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5846 4384 6054
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4066 5672 4122 5681
rect 4356 5658 4384 5782
rect 4066 5607 4122 5616
rect 4264 5630 4384 5658
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3588 5468 3884 5488
rect 3644 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3666 5414 3668 5466
rect 3730 5414 3742 5466
rect 3804 5414 3806 5466
rect 3644 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3588 5392 3884 5412
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 3332 5102 3384 5108
rect 3422 5128 3478 5137
rect 3422 5063 3478 5072
rect 3974 5128 4030 5137
rect 3974 5063 4030 5072
rect 3424 5024 3476 5030
rect 3330 4992 3386 5001
rect 3424 4966 3476 4972
rect 3330 4927 3386 4936
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3344 4690 3372 4927
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3534 3372 4082
rect 3108 3488 3188 3516
rect 3332 3528 3384 3534
rect 3056 3470 3108 3476
rect 3332 3470 3384 3476
rect 3344 3194 3372 3470
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 2962 1864 3018 1873
rect 2962 1799 3018 1808
rect 2870 640 2926 649
rect 2870 575 2926 584
rect 3252 480 3280 2382
rect 3436 2281 3464 4966
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 4049 3556 4422
rect 3588 4380 3884 4400
rect 3644 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3666 4326 3668 4378
rect 3730 4326 3742 4378
rect 3804 4326 3806 4378
rect 3644 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3588 4304 3884 4324
rect 3514 4040 3570 4049
rect 3514 3975 3570 3984
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3670 3832 3878
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3528 2990 3556 3334
rect 3588 3292 3884 3312
rect 3644 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3666 3238 3668 3290
rect 3730 3238 3742 3290
rect 3804 3238 3806 3290
rect 3644 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3588 3216 3884 3236
rect 3988 3097 4016 5063
rect 4080 5030 4108 5199
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4068 4616 4120 4622
rect 4066 4584 4068 4593
rect 4120 4584 4122 4593
rect 4066 4519 4122 4528
rect 4172 4162 4200 5306
rect 4264 5234 4292 5630
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4264 4593 4292 5170
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4250 4584 4306 4593
rect 4250 4519 4306 4528
rect 4356 4162 4384 4626
rect 4080 4134 4200 4162
rect 4264 4134 4384 4162
rect 4080 3942 4108 4134
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3974 3088 4030 3097
rect 3974 3023 4030 3032
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3698 2680 3754 2689
rect 4080 2650 4108 3470
rect 4172 3194 4200 4014
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4264 3058 4292 4134
rect 4540 4026 4568 6394
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4448 3998 4568 4026
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 3698 2615 3754 2624
rect 4068 2644 4120 2650
rect 3712 2582 3740 2615
rect 4068 2586 4120 2592
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 4158 2544 4214 2553
rect 4158 2479 4160 2488
rect 4212 2479 4214 2488
rect 4160 2450 4212 2456
rect 3422 2272 3478 2281
rect 3422 2207 3478 2216
rect 3588 2204 3884 2224
rect 3644 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3666 2150 3668 2202
rect 3730 2150 3742 2202
rect 3804 2150 3806 2202
rect 3644 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3588 2128 3884 2148
rect 4356 2020 4384 3946
rect 4448 3738 4476 3998
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4540 2854 4568 3878
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4632 2514 4660 9318
rect 4710 9279 4766 9288
rect 4724 9110 4752 9279
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4908 8634 4936 9687
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5000 8480 5028 9862
rect 5092 9518 5120 10639
rect 5170 10024 5226 10033
rect 5170 9959 5226 9968
rect 5184 9722 5212 9959
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 4908 8452 5028 8480
rect 4710 7032 4766 7041
rect 4710 6967 4712 6976
rect 4764 6967 4766 6976
rect 4712 6938 4764 6944
rect 4710 6624 4766 6633
rect 4710 6559 4766 6568
rect 4724 6186 4752 6559
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4724 3602 4752 6122
rect 4908 5710 4936 8452
rect 5092 8378 5120 9318
rect 5276 8974 5304 10764
rect 5368 10606 5396 12679
rect 5460 12102 5488 12786
rect 5644 12102 5672 13330
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5552 11286 5580 11834
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5460 10266 5488 11154
rect 5644 10810 5672 11494
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5460 9602 5488 10202
rect 5552 9722 5580 10746
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 10266 5672 10610
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5644 9654 5672 9930
rect 5632 9648 5684 9654
rect 5460 9586 5580 9602
rect 5632 9590 5684 9596
rect 5460 9580 5592 9586
rect 5460 9574 5540 9580
rect 5540 9522 5592 9528
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5368 9217 5396 9454
rect 5448 9376 5500 9382
rect 5446 9344 5448 9353
rect 5500 9344 5502 9353
rect 5446 9279 5502 9288
rect 5354 9208 5410 9217
rect 5354 9143 5410 9152
rect 5264 8968 5316 8974
rect 5170 8936 5226 8945
rect 5264 8910 5316 8916
rect 5170 8871 5226 8880
rect 5000 8350 5120 8378
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4816 4486 4844 5034
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4724 2582 4752 3062
rect 4816 3058 4844 4422
rect 5000 4264 5028 8350
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7818 5120 8230
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 7002 5120 7142
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5000 4236 5120 4264
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4436 2440 4488 2446
rect 4712 2440 4764 2446
rect 4488 2388 4712 2394
rect 4436 2382 4764 2388
rect 4448 2366 4752 2382
rect 4908 2310 4936 4014
rect 5000 3380 5028 4082
rect 5092 3738 5120 4236
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5080 3392 5132 3398
rect 5000 3352 5080 3380
rect 5080 3334 5132 3340
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5000 2650 5028 2926
rect 5092 2922 5120 3334
rect 5184 3058 5212 8871
rect 5262 8664 5318 8673
rect 5262 8599 5318 8608
rect 5276 8566 5304 8599
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 8090 5304 8230
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5262 7304 5318 7313
rect 5262 7239 5318 7248
rect 5276 7206 5304 7239
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 3913 5304 7142
rect 5262 3904 5318 3913
rect 5262 3839 5318 3848
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5184 2650 5212 2790
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5276 2530 5304 3606
rect 5368 3505 5396 9143
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5460 6458 5488 7278
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5284 5488 5646
rect 5552 5545 5580 8774
rect 5644 8378 5672 8978
rect 5736 8548 5764 13670
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5828 12442 5856 13194
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5828 11762 5856 12242
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5814 11248 5870 11257
rect 5814 11183 5870 11192
rect 5828 9081 5856 11183
rect 5920 9518 5948 13194
rect 6012 12306 6040 13262
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6104 11830 6132 14350
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 13938 6224 14214
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6220 13628 6516 13648
rect 6276 13626 6300 13628
rect 6356 13626 6380 13628
rect 6436 13626 6460 13628
rect 6298 13574 6300 13626
rect 6362 13574 6374 13626
rect 6436 13574 6438 13626
rect 6276 13572 6300 13574
rect 6356 13572 6380 13574
rect 6436 13572 6460 13574
rect 6220 13552 6516 13572
rect 6220 12540 6516 12560
rect 6276 12538 6300 12540
rect 6356 12538 6380 12540
rect 6436 12538 6460 12540
rect 6298 12486 6300 12538
rect 6362 12486 6374 12538
rect 6436 12486 6438 12538
rect 6276 12484 6300 12486
rect 6356 12484 6380 12486
rect 6436 12484 6460 12486
rect 6220 12464 6516 12484
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6196 11642 6224 12038
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6104 11614 6224 11642
rect 6104 11286 6132 11614
rect 6220 11452 6516 11472
rect 6276 11450 6300 11452
rect 6356 11450 6380 11452
rect 6436 11450 6460 11452
rect 6298 11398 6300 11450
rect 6362 11398 6374 11450
rect 6436 11398 6438 11450
rect 6276 11396 6300 11398
rect 6356 11396 6380 11398
rect 6436 11396 6460 11398
rect 6220 11376 6516 11396
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6564 11218 6592 11698
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 11082 6592 11154
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6550 10568 6606 10577
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6012 10130 6040 10202
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5814 9072 5870 9081
rect 5814 9007 5816 9016
rect 5868 9007 5870 9016
rect 5816 8978 5868 8984
rect 5828 8947 5856 8978
rect 5736 8520 5856 8548
rect 5644 8350 5764 8378
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8090 5672 8230
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5736 8022 5764 8350
rect 5724 8016 5776 8022
rect 5724 7958 5776 7964
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7041 5764 7686
rect 5722 7032 5778 7041
rect 5722 6967 5778 6976
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5644 6390 5672 6870
rect 5722 6488 5778 6497
rect 5722 6423 5778 6432
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5538 5536 5594 5545
rect 5538 5471 5594 5480
rect 5644 5370 5672 6326
rect 5736 6322 5764 6423
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5778 5764 6054
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 5296 5592 5302
rect 5460 5256 5540 5284
rect 5540 5238 5592 5244
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5460 3670 5488 5034
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5448 3528 5500 3534
rect 5354 3496 5410 3505
rect 5448 3470 5500 3476
rect 5354 3431 5410 3440
rect 5368 2582 5396 3431
rect 5184 2502 5304 2530
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4264 1992 4384 2020
rect 3700 1080 3752 1086
rect 3698 1048 3700 1057
rect 3752 1048 3754 1057
rect 3698 983 3754 992
rect 4264 480 4292 1992
rect 5184 480 5212 2502
rect 5460 2446 5488 3470
rect 5552 3398 5580 3946
rect 5644 3602 5672 5102
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5552 2582 5580 2994
rect 5644 2990 5672 3334
rect 5736 3058 5764 5714
rect 5828 4690 5856 8520
rect 5920 8265 5948 9318
rect 5906 8256 5962 8265
rect 5906 8191 5962 8200
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5920 5166 5948 7890
rect 6012 7886 6040 10066
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6012 5030 6040 7142
rect 6104 6390 6132 10542
rect 6550 10503 6606 10512
rect 6220 10364 6516 10384
rect 6276 10362 6300 10364
rect 6356 10362 6380 10364
rect 6436 10362 6460 10364
rect 6298 10310 6300 10362
rect 6362 10310 6374 10362
rect 6436 10310 6438 10362
rect 6276 10308 6300 10310
rect 6356 10308 6380 10310
rect 6436 10308 6460 10310
rect 6220 10288 6516 10308
rect 6220 9276 6516 9296
rect 6276 9274 6300 9276
rect 6356 9274 6380 9276
rect 6436 9274 6460 9276
rect 6298 9222 6300 9274
rect 6362 9222 6374 9274
rect 6436 9222 6438 9274
rect 6276 9220 6300 9222
rect 6356 9220 6380 9222
rect 6436 9220 6460 9222
rect 6220 9200 6516 9220
rect 6220 8188 6516 8208
rect 6276 8186 6300 8188
rect 6356 8186 6380 8188
rect 6436 8186 6460 8188
rect 6298 8134 6300 8186
rect 6362 8134 6374 8186
rect 6436 8134 6438 8186
rect 6276 8132 6300 8134
rect 6356 8132 6380 8134
rect 6436 8132 6460 8134
rect 6220 8112 6516 8132
rect 6184 7880 6236 7886
rect 6182 7848 6184 7857
rect 6276 7880 6328 7886
rect 6236 7848 6238 7857
rect 6276 7822 6328 7828
rect 6182 7783 6238 7792
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7342 6224 7686
rect 6288 7410 6316 7822
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6220 7100 6516 7120
rect 6276 7098 6300 7100
rect 6356 7098 6380 7100
rect 6436 7098 6460 7100
rect 6298 7046 6300 7098
rect 6362 7046 6374 7098
rect 6436 7046 6438 7098
rect 6276 7044 6300 7046
rect 6356 7044 6380 7046
rect 6436 7044 6460 7046
rect 6220 7024 6516 7044
rect 6564 6746 6592 10503
rect 6380 6718 6592 6746
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6380 6168 6408 6718
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6104 6140 6408 6168
rect 6458 6216 6514 6225
rect 6458 6151 6460 6160
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5998 4856 6054 4865
rect 5998 4791 6054 4800
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5906 4040 5962 4049
rect 5906 3975 5962 3984
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3738 5856 3878
rect 5920 3738 5948 3975
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5828 3058 5856 3538
rect 6012 3466 6040 4791
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 6012 2922 6040 3402
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 6104 2514 6132 6140
rect 6512 6151 6514 6160
rect 6460 6122 6512 6128
rect 6220 6012 6516 6032
rect 6276 6010 6300 6012
rect 6356 6010 6380 6012
rect 6436 6010 6460 6012
rect 6298 5958 6300 6010
rect 6362 5958 6374 6010
rect 6436 5958 6438 6010
rect 6276 5956 6300 5958
rect 6356 5956 6380 5958
rect 6436 5956 6460 5958
rect 6220 5936 6516 5956
rect 6564 5098 6592 6598
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6220 4924 6516 4944
rect 6276 4922 6300 4924
rect 6356 4922 6380 4924
rect 6436 4922 6460 4924
rect 6298 4870 6300 4922
rect 6362 4870 6374 4922
rect 6436 4870 6438 4922
rect 6276 4868 6300 4870
rect 6356 4868 6380 4870
rect 6436 4868 6460 4870
rect 6220 4848 6516 4868
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6472 4214 6500 4422
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6220 3836 6516 3856
rect 6276 3834 6300 3836
rect 6356 3834 6380 3836
rect 6436 3834 6460 3836
rect 6298 3782 6300 3834
rect 6362 3782 6374 3834
rect 6436 3782 6438 3834
rect 6276 3780 6300 3782
rect 6356 3780 6380 3782
rect 6436 3780 6460 3782
rect 6220 3760 6516 3780
rect 6460 3528 6512 3534
rect 6564 3516 6592 4490
rect 6512 3488 6592 3516
rect 6460 3470 6512 3476
rect 6656 3194 6684 14418
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6840 13025 6868 13330
rect 6826 13016 6882 13025
rect 6826 12951 6828 12960
rect 6880 12951 6882 12960
rect 6828 12922 6880 12928
rect 6840 12891 6868 12922
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11694 6776 12038
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6748 11150 6776 11630
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10962 6776 11086
rect 6840 11082 6868 11562
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6748 10934 6868 10962
rect 6840 10674 6868 10934
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 9994 6776 10542
rect 6840 10470 6868 10610
rect 6932 10470 6960 13874
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6840 10062 6868 10406
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9988 6788 9994
rect 6736 9930 6788 9936
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6748 8956 6776 9590
rect 6840 9518 6868 9998
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9110 6868 9454
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6748 8928 6868 8956
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6748 7546 6776 8230
rect 6840 8129 6868 8928
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6826 8120 6882 8129
rect 6826 8055 6882 8064
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 7002 6776 7346
rect 6932 7342 6960 8434
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6840 6390 6868 6870
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6828 6384 6880 6390
rect 6734 6352 6790 6361
rect 6828 6326 6880 6332
rect 6932 6322 6960 6802
rect 6734 6287 6790 6296
rect 6920 6316 6972 6322
rect 6748 6186 6776 6287
rect 6920 6258 6972 6264
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6748 5166 6776 5510
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6734 4992 6790 5001
rect 6734 4927 6790 4936
rect 6748 4282 6776 4927
rect 6840 4690 6868 5510
rect 6932 5302 6960 6258
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 4826 6960 5238
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6748 3738 6776 4218
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6220 2748 6516 2768
rect 6276 2746 6300 2748
rect 6356 2746 6380 2748
rect 6436 2746 6460 2748
rect 6298 2694 6300 2746
rect 6362 2694 6374 2746
rect 6436 2694 6438 2746
rect 6276 2692 6300 2694
rect 6356 2692 6380 2694
rect 6436 2692 6460 2694
rect 6220 2672 6516 2692
rect 6932 2553 6960 4150
rect 7024 2650 7052 13670
rect 7116 12050 7144 14350
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 13938 7696 14214
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 12850 7236 13670
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7300 12782 7328 13126
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7392 12628 7420 13738
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7300 12600 7420 12628
rect 7116 12022 7236 12050
rect 7102 11792 7158 11801
rect 7102 11727 7158 11736
rect 7116 11218 7144 11727
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 10130 7144 10406
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7116 9722 7144 10066
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7208 9450 7236 12022
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7116 8090 7144 8298
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7104 6860 7156 6866
rect 7208 6848 7236 8842
rect 7300 8362 7328 12600
rect 7576 12288 7604 13398
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 12850 7696 13262
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7760 12322 7788 13670
rect 7852 13394 7880 13874
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7932 12776 7984 12782
rect 7852 12724 7932 12730
rect 7852 12718 7984 12724
rect 7852 12702 7972 12718
rect 7852 12442 7880 12702
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7484 12260 7604 12288
rect 7668 12294 7788 12322
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10674 7420 11086
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7484 10470 7512 12260
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7576 11558 7604 12106
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 10266 7512 10406
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7378 9888 7434 9897
rect 7378 9823 7434 9832
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7392 8294 7420 9823
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7484 8838 7512 9386
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7300 6866 7328 6938
rect 7156 6820 7236 6848
rect 7288 6860 7340 6866
rect 7104 6802 7156 6808
rect 7288 6802 7340 6808
rect 7300 6769 7328 6802
rect 7286 6760 7342 6769
rect 7286 6695 7342 6704
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6254 7236 6598
rect 7196 6248 7248 6254
rect 7248 6208 7328 6236
rect 7196 6190 7248 6196
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 4690 7144 5510
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7116 4214 7144 4626
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7208 3942 7236 5646
rect 7300 5234 7328 6208
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7300 4146 7328 5170
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7102 3632 7158 3641
rect 7102 3567 7104 3576
rect 7156 3567 7158 3576
rect 7104 3538 7156 3544
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6918 2544 6974 2553
rect 6092 2508 6144 2514
rect 7208 2514 7236 3674
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7300 3126 7328 3470
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7392 2990 7420 7142
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7378 2680 7434 2689
rect 7378 2615 7380 2624
rect 7432 2615 7434 2624
rect 7380 2586 7432 2592
rect 6918 2479 6974 2488
rect 7196 2508 7248 2514
rect 6092 2450 6144 2456
rect 7196 2450 7248 2456
rect 7484 2446 7512 8774
rect 7576 7290 7604 11494
rect 7668 9761 7696 12294
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 11218 7788 12174
rect 7852 11694 7880 12378
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7654 9752 7710 9761
rect 7654 9687 7710 9696
rect 7668 9489 7696 9687
rect 7654 9480 7710 9489
rect 7654 9415 7710 9424
rect 7760 8514 7788 11154
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 9042 7880 9454
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7760 8486 7880 8514
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7576 7262 7696 7290
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 6934 7604 7142
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7562 6488 7618 6497
rect 7562 6423 7618 6432
rect 7576 5914 7604 6423
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7668 5778 7696 7262
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7576 3074 7604 3878
rect 7668 3738 7696 3878
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7760 3534 7788 8366
rect 7852 4049 7880 8486
rect 7944 5642 7972 12582
rect 8036 7886 8064 13398
rect 8128 10606 8156 14350
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8220 12306 8248 13330
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12782 8340 13126
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8298 12336 8354 12345
rect 8208 12300 8260 12306
rect 8298 12271 8354 12280
rect 8208 12242 8260 12248
rect 8220 10810 8248 12242
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8128 10266 8156 10542
rect 8312 10305 8340 12271
rect 8404 11558 8432 13806
rect 8588 13394 8616 14214
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13530 8708 13670
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8496 11898 8524 12786
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8496 11762 8524 11834
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8298 10296 8354 10305
rect 8116 10260 8168 10266
rect 8298 10231 8354 10240
rect 8116 10202 8168 10208
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8116 8492 8168 8498
rect 8220 8480 8248 8774
rect 8168 8452 8248 8480
rect 8116 8434 8168 8440
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8114 7848 8170 7857
rect 8036 7342 8064 7822
rect 8220 7818 8248 8452
rect 8312 8090 8340 10066
rect 8404 9500 8432 11494
rect 8680 11150 8708 11630
rect 8772 11234 8800 14418
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8852 14172 9148 14192
rect 8908 14170 8932 14172
rect 8988 14170 9012 14172
rect 9068 14170 9092 14172
rect 8930 14118 8932 14170
rect 8994 14118 9006 14170
rect 9068 14118 9070 14170
rect 8908 14116 8932 14118
rect 8988 14116 9012 14118
rect 9068 14116 9092 14118
rect 8852 14096 9148 14116
rect 9232 13938 9260 14350
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9324 13870 9352 15166
rect 11484 14716 11780 14736
rect 11540 14714 11564 14716
rect 11620 14714 11644 14716
rect 11700 14714 11724 14716
rect 11562 14662 11564 14714
rect 11626 14662 11638 14714
rect 11700 14662 11702 14714
rect 11540 14660 11564 14662
rect 11620 14660 11644 14662
rect 11700 14660 11724 14662
rect 11484 14640 11780 14660
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9312 13864 9364 13870
rect 8850 13832 8906 13841
rect 9364 13824 9444 13852
rect 9312 13806 9364 13812
rect 8850 13767 8906 13776
rect 8864 13734 8892 13767
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8864 13297 8892 13330
rect 8850 13288 8906 13297
rect 8850 13223 8906 13232
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 8852 13084 9148 13104
rect 8908 13082 8932 13084
rect 8988 13082 9012 13084
rect 9068 13082 9092 13084
rect 8930 13030 8932 13082
rect 8994 13030 9006 13082
rect 9068 13030 9070 13082
rect 8908 13028 8932 13030
rect 8988 13028 9012 13030
rect 9068 13028 9092 13030
rect 8852 13008 9148 13028
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9048 12442 9076 12582
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9140 12238 9168 12582
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 8852 11996 9148 12016
rect 8908 11994 8932 11996
rect 8988 11994 9012 11996
rect 9068 11994 9092 11996
rect 8930 11942 8932 11994
rect 8994 11942 9006 11994
rect 9068 11942 9070 11994
rect 8908 11940 8932 11942
rect 8988 11940 9012 11942
rect 9068 11940 9092 11942
rect 8852 11920 9148 11940
rect 9232 11234 9260 13126
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9324 11354 9352 12038
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 8772 11206 8892 11234
rect 9232 11206 9352 11234
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8864 11082 8892 11206
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8496 9897 8524 10134
rect 8680 9926 8708 10950
rect 8576 9920 8628 9926
rect 8482 9888 8538 9897
rect 8576 9862 8628 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8482 9823 8538 9832
rect 8404 9472 8524 9500
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8496 7970 8524 9472
rect 8588 8090 8616 9862
rect 8680 9625 8708 9862
rect 8666 9616 8722 9625
rect 8666 9551 8722 9560
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8404 7868 8432 7958
rect 8496 7942 8616 7970
rect 8484 7880 8536 7886
rect 8404 7840 8484 7868
rect 8114 7783 8116 7792
rect 8168 7783 8170 7792
rect 8208 7812 8260 7818
rect 8116 7754 8168 7760
rect 8208 7754 8260 7760
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7930 5536 7986 5545
rect 7930 5471 7986 5480
rect 7838 4040 7894 4049
rect 7838 3975 7894 3984
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7852 3466 7880 3975
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7576 3046 7696 3074
rect 7668 2938 7696 3046
rect 7852 2938 7880 3130
rect 7944 3126 7972 5471
rect 8036 5370 8064 5714
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7668 2910 7880 2938
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7944 2446 7972 2926
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6104 480 6132 2314
rect 7116 480 7144 2382
rect 8036 480 8064 4694
rect 8128 3534 8156 6938
rect 8404 6390 8432 7840
rect 8484 7822 8536 7828
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8220 5710 8248 6054
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5098 8248 5646
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8300 4616 8352 4622
rect 8206 4584 8262 4593
rect 8300 4558 8352 4564
rect 8206 4519 8208 4528
rect 8260 4519 8262 4528
rect 8208 4490 8260 4496
rect 8312 3942 8340 4558
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8220 3738 8248 3878
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8128 3097 8156 3470
rect 8312 3398 8340 3878
rect 8404 3670 8432 6054
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8496 3602 8524 6258
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8114 3088 8170 3097
rect 8114 3023 8170 3032
rect 8496 2446 8524 3538
rect 8588 2990 8616 7942
rect 8680 6730 8708 9046
rect 8772 8022 8800 11018
rect 8852 10908 9148 10928
rect 8908 10906 8932 10908
rect 8988 10906 9012 10908
rect 9068 10906 9092 10908
rect 8930 10854 8932 10906
rect 8994 10854 9006 10906
rect 9068 10854 9070 10906
rect 8908 10852 8932 10854
rect 8988 10852 9012 10854
rect 9068 10852 9092 10854
rect 8852 10832 9148 10852
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9140 10441 9168 10474
rect 9126 10432 9182 10441
rect 9126 10367 9182 10376
rect 9232 10062 9260 11086
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 8852 9820 9148 9840
rect 8908 9818 8932 9820
rect 8988 9818 9012 9820
rect 9068 9818 9092 9820
rect 8930 9766 8932 9818
rect 8994 9766 9006 9818
rect 9068 9766 9070 9818
rect 8908 9764 8932 9766
rect 8988 9764 9012 9766
rect 9068 9764 9092 9766
rect 8852 9744 9148 9764
rect 9232 9042 9260 9998
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9324 8922 9352 11206
rect 9416 10538 9444 13824
rect 9508 13190 9536 14010
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9508 10606 9536 12650
rect 9692 12442 9720 13738
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9678 11792 9734 11801
rect 9678 11727 9734 11736
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9600 10810 9628 11154
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9416 9994 9444 10474
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9494 10296 9550 10305
rect 9494 10231 9550 10240
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9508 9761 9536 10231
rect 9600 10130 9628 10406
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9692 10010 9720 11727
rect 9784 11286 9812 13126
rect 9876 12850 9904 13874
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13530 10180 13670
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10138 12880 10194 12889
rect 9864 12844 9916 12850
rect 10336 12866 10364 14554
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10428 12889 10456 14418
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10138 12815 10194 12824
rect 10244 12838 10364 12866
rect 10414 12880 10470 12889
rect 9864 12786 9916 12792
rect 9876 11898 9904 12786
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9968 12238 9996 12718
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9876 11762 9904 11834
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 11286 9904 11698
rect 9772 11280 9824 11286
rect 9772 11222 9824 11228
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9968 11150 9996 12174
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9600 9982 9720 10010
rect 9494 9752 9550 9761
rect 9494 9687 9550 9696
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9416 8945 9444 9590
rect 9232 8894 9352 8922
rect 9402 8936 9458 8945
rect 8852 8732 9148 8752
rect 8908 8730 8932 8732
rect 8988 8730 9012 8732
rect 9068 8730 9092 8732
rect 8930 8678 8932 8730
rect 8994 8678 9006 8730
rect 9068 8678 9070 8730
rect 8908 8676 8932 8678
rect 8988 8676 9012 8678
rect 9068 8676 9092 8678
rect 8852 8656 9148 8676
rect 9232 8514 9260 8894
rect 9402 8871 9458 8880
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9140 8486 9260 8514
rect 9140 8362 9168 8486
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8956 7886 8984 8298
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8852 7644 9148 7664
rect 8908 7642 8932 7644
rect 8988 7642 9012 7644
rect 9068 7642 9092 7644
rect 8930 7590 8932 7642
rect 8994 7590 9006 7642
rect 9068 7590 9070 7642
rect 8908 7588 8932 7590
rect 8988 7588 9012 7590
rect 9068 7588 9092 7590
rect 8852 7568 9148 7588
rect 9232 7274 9260 8366
rect 9324 8362 9352 8774
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 7886 9352 8298
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9416 7274 9444 8026
rect 9508 7834 9536 9687
rect 9600 9625 9628 9982
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9586 9616 9642 9625
rect 9586 9551 9642 9560
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9600 9330 9628 9454
rect 9692 9450 9720 9862
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9784 9330 9812 11018
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10033 9904 10406
rect 9862 10024 9918 10033
rect 9862 9959 9918 9968
rect 10060 9450 10088 12038
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9600 9302 9812 9330
rect 9692 8906 9720 9302
rect 9876 8974 9904 9386
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9600 8090 9628 8502
rect 9692 8498 9720 8842
rect 9770 8664 9826 8673
rect 9770 8599 9826 8608
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9784 7954 9812 8599
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9968 7857 9996 8910
rect 9954 7848 10010 7857
rect 9508 7806 9628 7834
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9232 6746 9260 7210
rect 8668 6724 8720 6730
rect 9232 6718 9352 6746
rect 8668 6666 8720 6672
rect 8680 4690 8708 6666
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 8852 6556 9148 6576
rect 8908 6554 8932 6556
rect 8988 6554 9012 6556
rect 9068 6554 9092 6556
rect 8930 6502 8932 6554
rect 8994 6502 9006 6554
rect 9068 6502 9070 6554
rect 8908 6500 8932 6502
rect 8988 6500 9012 6502
rect 9068 6500 9092 6502
rect 8852 6480 9148 6500
rect 9232 6390 9260 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9324 6322 9352 6718
rect 9416 6361 9444 7210
rect 9402 6352 9458 6361
rect 9312 6316 9364 6322
rect 9402 6287 9458 6296
rect 9312 6258 9364 6264
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 9310 6216 9366 6225
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8772 4078 8800 6190
rect 9310 6151 9366 6160
rect 9324 6118 9352 6151
rect 9312 6112 9364 6118
rect 9218 6080 9274 6089
rect 9312 6054 9364 6060
rect 9218 6015 9274 6024
rect 9232 5642 9260 6015
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 8852 5468 9148 5488
rect 8908 5466 8932 5468
rect 8988 5466 9012 5468
rect 9068 5466 9092 5468
rect 8930 5414 8932 5466
rect 8994 5414 9006 5466
rect 9068 5414 9070 5466
rect 8908 5412 8932 5414
rect 8988 5412 9012 5414
rect 9068 5412 9092 5414
rect 8852 5392 9148 5412
rect 9232 5352 9260 5578
rect 9140 5324 9260 5352
rect 9140 4622 9168 5324
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9232 4758 9260 4966
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 8852 4380 9148 4400
rect 8908 4378 8932 4380
rect 8988 4378 9012 4380
rect 9068 4378 9092 4380
rect 8930 4326 8932 4378
rect 8994 4326 9006 4378
rect 9068 4326 9070 4378
rect 8908 4324 8932 4326
rect 8988 4324 9012 4326
rect 9068 4324 9092 4326
rect 8852 4304 9148 4324
rect 9232 4214 9260 4694
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8956 3505 8984 3538
rect 9220 3528 9272 3534
rect 8942 3496 8998 3505
rect 9220 3470 9272 3476
rect 8942 3431 8998 3440
rect 8852 3292 9148 3312
rect 8908 3290 8932 3292
rect 8988 3290 9012 3292
rect 9068 3290 9092 3292
rect 8930 3238 8932 3290
rect 8994 3238 9006 3290
rect 9068 3238 9070 3290
rect 8908 3236 8932 3238
rect 8988 3236 9012 3238
rect 9068 3236 9092 3238
rect 8852 3216 9148 3236
rect 8942 3088 8998 3097
rect 9232 3058 9260 3470
rect 8942 3023 8944 3032
rect 8996 3023 8998 3032
rect 9220 3052 9272 3058
rect 8944 2994 8996 3000
rect 9220 2994 9272 3000
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 9034 2952 9090 2961
rect 9034 2887 9090 2896
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2650 8800 2790
rect 9048 2650 9076 2887
rect 9126 2816 9182 2825
rect 9126 2751 9182 2760
rect 9140 2650 9168 2751
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 1086 8248 2246
rect 8852 2204 9148 2224
rect 8908 2202 8932 2204
rect 8988 2202 9012 2204
rect 9068 2202 9092 2204
rect 8930 2150 8932 2202
rect 8994 2150 9006 2202
rect 9068 2150 9070 2202
rect 8908 2148 8932 2150
rect 8988 2148 9012 2150
rect 9068 2148 9092 2150
rect 8852 2128 9148 2148
rect 9324 1850 9352 5646
rect 9508 5166 9536 7686
rect 9600 6866 9628 7806
rect 9954 7783 10010 7792
rect 10060 7698 10088 8978
rect 10152 8974 10180 12815
rect 10244 11778 10272 12838
rect 10414 12815 10470 12824
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10336 11898 10364 12242
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10244 11750 10364 11778
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10244 9382 10272 9998
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10232 9036 10284 9042
rect 10336 9024 10364 11750
rect 10428 10266 10456 12650
rect 10520 12442 10548 13670
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10520 11665 10548 12378
rect 10612 11830 10640 13806
rect 10704 13394 10732 14418
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10506 11656 10562 11665
rect 10506 11591 10562 11600
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 11218 10640 11494
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10612 10742 10640 10950
rect 10600 10736 10652 10742
rect 10506 10704 10562 10713
rect 10600 10678 10652 10684
rect 10506 10639 10562 10648
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10284 8996 10364 9024
rect 10232 8978 10284 8984
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 9968 7670 10088 7698
rect 9968 7313 9996 7670
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9954 7304 10010 7313
rect 9954 7239 10010 7248
rect 9968 7041 9996 7239
rect 9954 7032 10010 7041
rect 10060 7002 10088 7414
rect 10336 7342 10364 7822
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 9954 6967 10010 6976
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9600 5012 9628 6802
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 5846 9720 6734
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5914 9812 6054
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9508 4984 9628 5012
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9416 4010 9444 4558
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3534 9444 3946
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9508 2990 9536 4984
rect 9692 3602 9720 5510
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9784 4078 9812 4626
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9772 3936 9824 3942
rect 9876 3924 9904 6802
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10060 5166 10088 5714
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9824 3896 9904 3924
rect 9772 3878 9824 3884
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9600 2938 9628 3130
rect 9784 2990 9812 3878
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 2984 9824 2990
rect 9404 2916 9456 2922
rect 9600 2910 9720 2938
rect 9772 2926 9824 2932
rect 9404 2858 9456 2864
rect 8956 1822 9352 1850
rect 8208 1080 8260 1086
rect 8208 1022 8260 1028
rect 8956 480 8984 1822
rect 9416 1494 9444 2858
rect 9692 2836 9720 2910
rect 9772 2848 9824 2854
rect 9692 2808 9772 2836
rect 9876 2836 9904 3130
rect 9824 2808 9904 2836
rect 9772 2790 9824 2796
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9784 2106 9812 2450
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 9404 1488 9456 1494
rect 9404 1430 9456 1436
rect 9968 480 9996 5034
rect 10152 3194 10180 5646
rect 10336 5234 10364 7278
rect 10428 5778 10456 10202
rect 10520 9897 10548 10639
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10612 10062 10640 10406
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10506 9888 10562 9897
rect 10506 9823 10562 9832
rect 10520 8090 10548 9823
rect 10612 9722 10640 9998
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10612 8974 10640 9658
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 6225 10548 7142
rect 10704 7002 10732 13330
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10888 12102 10916 13262
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 9994 10824 11494
rect 10888 11354 10916 12038
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10980 11234 11008 11766
rect 10888 11206 11008 11234
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10796 8090 10824 9930
rect 10888 8537 10916 11206
rect 11072 10062 11100 14486
rect 14116 14172 14412 14192
rect 14172 14170 14196 14172
rect 14252 14170 14276 14172
rect 14332 14170 14356 14172
rect 14194 14118 14196 14170
rect 14258 14118 14270 14170
rect 14332 14118 14334 14170
rect 14172 14116 14196 14118
rect 14252 14116 14276 14118
rect 14332 14116 14356 14118
rect 14116 14096 14412 14116
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 11484 13628 11780 13648
rect 11540 13626 11564 13628
rect 11620 13626 11644 13628
rect 11700 13626 11724 13628
rect 11562 13574 11564 13626
rect 11626 13574 11638 13626
rect 11700 13574 11702 13626
rect 11540 13572 11564 13574
rect 11620 13572 11644 13574
rect 11700 13572 11724 13574
rect 11484 13552 11780 13572
rect 12544 13462 12572 13738
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11348 12374 11376 12582
rect 11484 12540 11780 12560
rect 11540 12538 11564 12540
rect 11620 12538 11644 12540
rect 11700 12538 11724 12540
rect 11562 12486 11564 12538
rect 11626 12486 11638 12538
rect 11700 12486 11702 12538
rect 11540 12484 11564 12486
rect 11620 12484 11644 12486
rect 11700 12484 11724 12486
rect 11484 12464 11780 12484
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11348 11762 11376 12310
rect 11808 11898 11836 13262
rect 11900 12850 11928 13330
rect 11980 13320 12032 13326
rect 12900 13320 12952 13326
rect 11980 13262 12032 13268
rect 12820 13280 12900 13308
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11992 12714 12020 13262
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11992 12442 12020 12650
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11256 11121 11284 11562
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11242 11112 11298 11121
rect 11242 11047 11298 11056
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10056 11112 10062
rect 10980 10016 11060 10044
rect 10980 9466 11008 10016
rect 11060 9998 11112 10004
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9625 11100 9862
rect 11058 9616 11114 9625
rect 11058 9551 11114 9560
rect 10980 9438 11100 9466
rect 10874 8528 10930 8537
rect 10874 8463 10930 8472
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10980 7274 11008 8026
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10600 6928 10652 6934
rect 10598 6896 10600 6905
rect 10652 6896 10654 6905
rect 10598 6831 10654 6840
rect 10796 6798 10824 7210
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6361 10824 6734
rect 10782 6352 10838 6361
rect 10782 6287 10784 6296
rect 10836 6287 10838 6296
rect 10784 6258 10836 6264
rect 10506 6216 10562 6225
rect 10506 6151 10562 6160
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5914 10548 6054
rect 10980 5914 11008 7210
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10336 4690 10364 5170
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10704 4298 10732 5850
rect 11072 5778 11100 9438
rect 11164 7206 11192 10746
rect 11256 9160 11284 11047
rect 11348 10810 11376 11494
rect 11484 11452 11780 11472
rect 11540 11450 11564 11452
rect 11620 11450 11644 11452
rect 11700 11450 11724 11452
rect 11562 11398 11564 11450
rect 11626 11398 11638 11450
rect 11700 11398 11702 11450
rect 11540 11396 11564 11398
rect 11620 11396 11644 11398
rect 11700 11396 11724 11398
rect 11484 11376 11780 11396
rect 11794 11248 11850 11257
rect 11794 11183 11850 11192
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11484 10364 11780 10384
rect 11540 10362 11564 10364
rect 11620 10362 11644 10364
rect 11700 10362 11724 10364
rect 11562 10310 11564 10362
rect 11626 10310 11638 10362
rect 11700 10310 11702 10362
rect 11540 10308 11564 10310
rect 11620 10308 11644 10310
rect 11700 10308 11724 10310
rect 11484 10288 11780 10308
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11440 9897 11468 10066
rect 11426 9888 11482 9897
rect 11426 9823 11482 9832
rect 11702 9616 11758 9625
rect 11702 9551 11758 9560
rect 11716 9518 11744 9551
rect 11612 9512 11664 9518
rect 11426 9480 11482 9489
rect 11426 9415 11428 9424
rect 11480 9415 11482 9424
rect 11610 9480 11612 9489
rect 11704 9512 11756 9518
rect 11664 9480 11666 9489
rect 11704 9454 11756 9460
rect 11610 9415 11666 9424
rect 11428 9386 11480 9392
rect 11484 9276 11780 9296
rect 11540 9274 11564 9276
rect 11620 9274 11644 9276
rect 11700 9274 11724 9276
rect 11562 9222 11564 9274
rect 11626 9222 11638 9274
rect 11700 9222 11702 9274
rect 11540 9220 11564 9222
rect 11620 9220 11644 9222
rect 11700 9220 11724 9222
rect 11484 9200 11780 9220
rect 11256 9132 11376 9160
rect 11242 9072 11298 9081
rect 11242 9007 11298 9016
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11164 5914 11192 6258
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11060 5772 11112 5778
rect 11112 5732 11192 5760
rect 11060 5714 11112 5720
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10520 4270 10732 4298
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10244 2990 10272 4014
rect 10520 3670 10548 4270
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10336 2582 10364 3062
rect 10428 2650 10456 3470
rect 10520 3194 10548 3606
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10612 2990 10640 4150
rect 10888 4078 10916 4422
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3738 11008 3878
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10612 2446 10640 2926
rect 10704 2650 10732 3334
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10888 480 10916 3538
rect 11072 2922 11100 4422
rect 11164 4010 11192 5732
rect 11256 4162 11284 9007
rect 11348 6322 11376 9132
rect 11484 8188 11780 8208
rect 11540 8186 11564 8188
rect 11620 8186 11644 8188
rect 11700 8186 11724 8188
rect 11562 8134 11564 8186
rect 11626 8134 11638 8186
rect 11700 8134 11702 8186
rect 11540 8132 11564 8134
rect 11620 8132 11644 8134
rect 11700 8132 11724 8134
rect 11484 8112 11780 8132
rect 11808 7954 11836 11183
rect 12084 10674 12112 12718
rect 12268 12442 12296 13126
rect 12820 12714 12848 13280
rect 12900 13262 12952 13268
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12360 12209 12388 12242
rect 12440 12232 12492 12238
rect 12346 12200 12402 12209
rect 12544 12209 12572 12310
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12440 12174 12492 12180
rect 12530 12200 12586 12209
rect 12346 12135 12402 12144
rect 12452 11257 12480 12174
rect 12530 12135 12586 12144
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12544 11694 12572 11766
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12438 11248 12494 11257
rect 12544 11218 12572 11494
rect 12438 11183 12494 11192
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12072 10464 12124 10470
rect 11886 10432 11942 10441
rect 12072 10406 12124 10412
rect 11886 10367 11942 10376
rect 11900 10266 11928 10367
rect 12084 10266 12112 10406
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12162 9616 12218 9625
rect 12162 9551 12218 9560
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9217 12112 9318
rect 12070 9208 12126 9217
rect 12070 9143 12126 9152
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11900 7993 11928 8570
rect 12084 8498 12112 8978
rect 12176 8838 12204 9551
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12072 8492 12124 8498
rect 11992 8452 12072 8480
rect 11992 8090 12020 8452
rect 12072 8434 12124 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12072 8288 12124 8294
rect 12070 8256 12072 8265
rect 12124 8256 12126 8265
rect 12070 8191 12126 8200
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11886 7984 11942 7993
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11796 7948 11848 7954
rect 11886 7919 11942 7928
rect 11796 7890 11848 7896
rect 11716 7478 11744 7890
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11978 7304 12034 7313
rect 11978 7239 12034 7248
rect 11484 7100 11780 7120
rect 11540 7098 11564 7100
rect 11620 7098 11644 7100
rect 11700 7098 11724 7100
rect 11562 7046 11564 7098
rect 11626 7046 11638 7098
rect 11700 7046 11702 7098
rect 11540 7044 11564 7046
rect 11620 7044 11644 7046
rect 11700 7044 11724 7046
rect 11484 7024 11780 7044
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11704 6792 11756 6798
rect 11808 6769 11836 6802
rect 11704 6734 11756 6740
rect 11794 6760 11850 6769
rect 11716 6322 11744 6734
rect 11794 6695 11850 6704
rect 11336 6316 11388 6322
rect 11336 6258 11388 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11336 6112 11388 6118
rect 11716 6100 11744 6258
rect 11716 6072 11836 6100
rect 11336 6054 11388 6060
rect 11348 5896 11376 6054
rect 11484 6012 11780 6032
rect 11540 6010 11564 6012
rect 11620 6010 11644 6012
rect 11700 6010 11724 6012
rect 11562 5958 11564 6010
rect 11626 5958 11638 6010
rect 11700 5958 11702 6010
rect 11540 5956 11564 5958
rect 11620 5956 11644 5958
rect 11700 5956 11724 5958
rect 11484 5936 11780 5956
rect 11348 5868 11468 5896
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11348 4622 11376 5646
rect 11440 5642 11468 5868
rect 11704 5772 11756 5778
rect 11808 5760 11836 6072
rect 11756 5732 11836 5760
rect 11704 5714 11756 5720
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11440 5302 11468 5578
rect 11716 5370 11744 5714
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11428 5296 11480 5302
rect 11900 5250 11928 6938
rect 11992 6934 12020 7239
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11428 5238 11480 5244
rect 11808 5222 11928 5250
rect 11484 4924 11780 4944
rect 11540 4922 11564 4924
rect 11620 4922 11644 4924
rect 11700 4922 11724 4924
rect 11562 4870 11564 4922
rect 11626 4870 11638 4922
rect 11700 4870 11702 4922
rect 11540 4868 11564 4870
rect 11620 4868 11644 4870
rect 11700 4868 11724 4870
rect 11484 4848 11780 4868
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11256 4134 11376 4162
rect 11348 4078 11376 4134
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11164 2582 11192 3402
rect 11348 2650 11376 3878
rect 11484 3836 11780 3856
rect 11540 3834 11564 3836
rect 11620 3834 11644 3836
rect 11700 3834 11724 3836
rect 11562 3782 11564 3834
rect 11626 3782 11638 3834
rect 11700 3782 11702 3834
rect 11540 3780 11564 3782
rect 11620 3780 11644 3782
rect 11700 3780 11724 3782
rect 11484 3760 11780 3780
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11716 3194 11744 3470
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11484 2748 11780 2768
rect 11540 2746 11564 2748
rect 11620 2746 11644 2748
rect 11700 2746 11724 2748
rect 11562 2694 11564 2746
rect 11626 2694 11638 2746
rect 11700 2694 11702 2746
rect 11540 2692 11564 2694
rect 11620 2692 11644 2694
rect 11700 2692 11724 2694
rect 11484 2672 11780 2692
rect 11336 2644 11388 2650
rect 11808 2632 11836 5222
rect 12084 5166 12112 7142
rect 12176 6730 12204 8366
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12268 5273 12296 11018
rect 12544 10520 12572 11018
rect 12636 10713 12664 12242
rect 12820 12238 12848 12650
rect 13096 12594 13124 13194
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13004 12566 13124 12594
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12820 11762 12848 12174
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11354 12940 11494
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12622 10704 12678 10713
rect 12622 10639 12678 10648
rect 12624 10532 12676 10538
rect 12544 10492 12624 10520
rect 12624 10474 12676 10480
rect 12346 10296 12402 10305
rect 12346 10231 12402 10240
rect 12360 9761 12388 10231
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12544 9897 12572 10066
rect 12636 10062 12664 10474
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12530 9888 12586 9897
rect 12530 9823 12586 9832
rect 12346 9752 12402 9761
rect 12544 9722 12572 9823
rect 12346 9687 12402 9696
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12532 9444 12584 9450
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 9081 12388 9318
rect 12346 9072 12402 9081
rect 12452 9042 12480 9415
rect 12532 9386 12584 9392
rect 12346 9007 12402 9016
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12544 8673 12572 9386
rect 12636 9178 12664 9998
rect 12728 9382 12756 11086
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10266 12848 10406
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12912 9500 12940 10950
rect 13004 9625 13032 12566
rect 13082 12200 13138 12209
rect 13082 12135 13084 12144
rect 13136 12135 13138 12144
rect 13084 12106 13136 12112
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13096 11150 13124 11834
rect 13188 11694 13216 13126
rect 13372 11898 13400 13738
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13464 12986 13492 13330
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13464 12782 13492 12922
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13556 12730 13584 13942
rect 14002 13832 14058 13841
rect 14002 13767 14058 13776
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12918 13676 13330
rect 13910 13288 13966 13297
rect 13910 13223 13966 13232
rect 13636 12912 13688 12918
rect 13688 12860 13768 12866
rect 13636 12854 13768 12860
rect 13648 12838 13768 12854
rect 13464 12238 13492 12718
rect 13556 12702 13676 12730
rect 13542 12608 13598 12617
rect 13542 12543 13598 12552
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13174 11248 13230 11257
rect 13174 11183 13176 11192
rect 13228 11183 13230 11192
rect 13176 11154 13228 11160
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13188 10690 13216 11154
rect 13096 10662 13216 10690
rect 12990 9616 13046 9625
rect 12990 9551 13046 9560
rect 12912 9472 13032 9500
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12820 8922 12848 9318
rect 12728 8894 12848 8922
rect 12728 8838 12756 8894
rect 13004 8838 13032 9472
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12530 8664 12586 8673
rect 12530 8599 12586 8608
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12360 7449 12388 7482
rect 12346 7440 12402 7449
rect 12346 7375 12402 7384
rect 12438 6760 12494 6769
rect 12348 6724 12400 6730
rect 12438 6695 12494 6704
rect 12348 6666 12400 6672
rect 12360 6458 12388 6666
rect 12452 6458 12480 6695
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5914 12480 6190
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12254 5264 12310 5273
rect 12254 5199 12310 5208
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4826 12020 4966
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11900 4146 11928 4762
rect 12360 4486 12388 5510
rect 12452 5370 12480 5850
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12544 5166 12572 8502
rect 12728 8498 12756 8774
rect 12990 8528 13046 8537
rect 12716 8492 12768 8498
rect 12990 8463 13046 8472
rect 12716 8434 12768 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 8265 12664 8366
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12716 8288 12768 8294
rect 12622 8256 12678 8265
rect 12716 8230 12768 8236
rect 12622 8191 12678 8200
rect 12728 8106 12756 8230
rect 12636 8078 12756 8106
rect 12636 8022 12664 8078
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12806 7984 12862 7993
rect 12728 7528 12756 7958
rect 12806 7919 12862 7928
rect 12636 7500 12756 7528
rect 12636 6390 12664 7500
rect 12714 7440 12770 7449
rect 12820 7410 12848 7919
rect 12912 7818 12940 8298
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 13004 7698 13032 8463
rect 12912 7670 13032 7698
rect 12714 7375 12770 7384
rect 12808 7404 12860 7410
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12728 6254 12756 7375
rect 12808 7346 12860 7352
rect 12912 6866 12940 7670
rect 13096 6905 13124 10662
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 9450 13216 10474
rect 13280 10470 13308 11698
rect 13464 11626 13492 12174
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13464 11082 13492 11562
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13266 10160 13322 10169
rect 13266 10095 13322 10104
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13280 8294 13308 10095
rect 13372 8362 13400 10950
rect 13464 10606 13492 11018
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13464 9382 13492 10542
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13464 8430 13492 8842
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13556 7993 13584 12543
rect 13648 11354 13676 12702
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13542 7984 13598 7993
rect 13268 7948 13320 7954
rect 13542 7919 13598 7928
rect 13268 7890 13320 7896
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13188 7478 13216 7754
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13082 6896 13138 6905
rect 12900 6860 12952 6866
rect 13082 6831 13138 6840
rect 12900 6802 12952 6808
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12636 5914 12664 6054
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11992 3602 12020 4014
rect 12084 4010 12112 4082
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 12544 3670 12572 4966
rect 12636 4826 12664 5034
rect 12624 4820 12676 4826
rect 12676 4780 12756 4808
rect 12624 4762 12676 4768
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3738 12664 3878
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 2689 12020 3334
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12072 2916 12124 2922
rect 12072 2858 12124 2864
rect 11978 2680 12034 2689
rect 11888 2644 11940 2650
rect 11336 2586 11388 2592
rect 11716 2604 11888 2632
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11716 2378 11744 2604
rect 11978 2615 12034 2624
rect 11888 2586 11940 2592
rect 12084 2446 12112 2858
rect 12268 2582 12296 3062
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 12360 2514 12388 3606
rect 12728 3534 12756 4780
rect 12912 4690 12940 5170
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12912 4146 12940 4626
rect 13096 4622 13124 6831
rect 13188 6798 13216 7414
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13280 5846 13308 7890
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13372 7410 13400 7822
rect 13556 7546 13584 7822
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13372 5778 13400 6802
rect 13556 6361 13584 7346
rect 13648 7206 13676 11290
rect 13740 11286 13768 12838
rect 13924 12617 13952 13223
rect 13910 12608 13966 12617
rect 13910 12543 13966 12552
rect 14016 12458 14044 13767
rect 14476 13190 14504 15399
rect 14936 15230 14964 16215
rect 15014 15872 15070 15881
rect 15014 15807 15070 15816
rect 14924 15224 14976 15230
rect 14924 15166 14976 15172
rect 14830 14648 14886 14657
rect 14830 14583 14886 14592
rect 14646 14240 14702 14249
rect 14646 14175 14702 14184
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14116 13084 14412 13104
rect 14172 13082 14196 13084
rect 14252 13082 14276 13084
rect 14332 13082 14356 13084
rect 14194 13030 14196 13082
rect 14258 13030 14270 13082
rect 14332 13030 14334 13082
rect 14172 13028 14196 13030
rect 14252 13028 14276 13030
rect 14332 13028 14356 13030
rect 14116 13008 14412 13028
rect 13924 12430 14044 12458
rect 14464 12436 14516 12442
rect 13924 12209 13952 12430
rect 14464 12378 14516 12384
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11762 13952 12038
rect 14116 11996 14412 12016
rect 14172 11994 14196 11996
rect 14252 11994 14276 11996
rect 14332 11994 14356 11996
rect 14194 11942 14196 11994
rect 14258 11942 14270 11994
rect 14332 11942 14334 11994
rect 14172 11940 14196 11942
rect 14252 11940 14276 11942
rect 14332 11940 14356 11942
rect 14116 11920 14412 11940
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10690 13768 11086
rect 13740 10662 13860 10690
rect 13832 10606 13860 10662
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13740 9217 13768 10202
rect 13726 9208 13782 9217
rect 13726 9143 13782 9152
rect 13740 7818 13768 9143
rect 13832 8974 13860 10542
rect 13924 9761 13952 11154
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14016 10792 14044 11086
rect 14116 10908 14412 10928
rect 14172 10906 14196 10908
rect 14252 10906 14276 10908
rect 14332 10906 14356 10908
rect 14194 10854 14196 10906
rect 14258 10854 14270 10906
rect 14332 10854 14334 10906
rect 14172 10852 14196 10854
rect 14252 10852 14276 10854
rect 14332 10852 14356 10854
rect 14116 10832 14412 10852
rect 14016 10764 14320 10792
rect 14002 10704 14058 10713
rect 14002 10639 14058 10648
rect 13910 9752 13966 9761
rect 13910 9687 13966 9696
rect 14016 9568 14044 10639
rect 14186 10432 14242 10441
rect 14186 10367 14242 10376
rect 14200 10062 14228 10367
rect 14292 10062 14320 10764
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14116 9820 14412 9840
rect 14172 9818 14196 9820
rect 14252 9818 14276 9820
rect 14332 9818 14356 9820
rect 14194 9766 14196 9818
rect 14258 9766 14270 9818
rect 14332 9766 14334 9818
rect 14172 9764 14196 9766
rect 14252 9764 14276 9766
rect 14332 9764 14356 9766
rect 14116 9744 14412 9764
rect 14096 9648 14148 9654
rect 13924 9540 14044 9568
rect 14094 9616 14096 9625
rect 14372 9648 14424 9654
rect 14148 9616 14150 9625
rect 14372 9590 14424 9596
rect 14476 9602 14504 12378
rect 14660 12374 14688 14175
rect 14844 14074 14872 14583
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14752 11626 14780 12582
rect 14844 12306 14872 13126
rect 14936 12481 14964 13670
rect 15028 13462 15056 15807
rect 16210 15056 16266 15065
rect 16210 14991 16266 15000
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 14922 12472 14978 12481
rect 14922 12407 14978 12416
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14936 12238 14964 12407
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14568 10266 14596 11018
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14568 9722 14596 9998
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14094 9551 14150 9560
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13728 7472 13780 7478
rect 13832 7449 13860 8570
rect 13728 7414 13780 7420
rect 13818 7440 13874 7449
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13542 6352 13598 6361
rect 13740 6322 13768 7414
rect 13818 7375 13874 7384
rect 13820 7336 13872 7342
rect 13818 7304 13820 7313
rect 13872 7304 13874 7313
rect 13818 7239 13874 7248
rect 13924 7002 13952 9540
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 9178 14044 9386
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14292 9042 14320 9318
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 14016 8634 14044 8910
rect 14384 8820 14412 9590
rect 14476 9574 14596 9602
rect 14660 9586 14688 11018
rect 14752 9654 14780 11562
rect 14936 10962 14964 12174
rect 14936 10934 15056 10962
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14922 10432 14978 10441
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14464 8968 14516 8974
rect 14462 8936 14464 8945
rect 14516 8936 14518 8945
rect 14462 8871 14518 8880
rect 14384 8792 14504 8820
rect 14116 8732 14412 8752
rect 14172 8730 14196 8732
rect 14252 8730 14276 8732
rect 14332 8730 14356 8732
rect 14194 8678 14196 8730
rect 14258 8678 14270 8730
rect 14332 8678 14334 8730
rect 14172 8676 14196 8678
rect 14252 8676 14276 8678
rect 14332 8676 14356 8678
rect 14116 8656 14412 8676
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14476 7886 14504 8792
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14116 7644 14412 7664
rect 14172 7642 14196 7644
rect 14252 7642 14276 7644
rect 14332 7642 14356 7644
rect 14194 7590 14196 7642
rect 14258 7590 14270 7642
rect 14332 7590 14334 7642
rect 14172 7588 14196 7590
rect 14252 7588 14276 7590
rect 14332 7588 14356 7590
rect 14116 7568 14412 7588
rect 14476 7528 14504 7822
rect 14384 7500 14504 7528
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 14016 6798 14044 7210
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 7002 14320 7142
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14384 6866 14412 7500
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14476 6798 14504 7278
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14116 6556 14412 6576
rect 14172 6554 14196 6556
rect 14252 6554 14276 6556
rect 14332 6554 14356 6556
rect 14194 6502 14196 6554
rect 14258 6502 14270 6554
rect 14332 6502 14334 6554
rect 14172 6500 14196 6502
rect 14252 6500 14276 6502
rect 14332 6500 14356 6502
rect 14116 6480 14412 6500
rect 13542 6287 13598 6296
rect 13728 6316 13780 6322
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13372 4826 13400 5306
rect 13360 4820 13412 4826
rect 13188 4780 13360 4808
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 13188 3534 13216 4780
rect 13360 4762 13412 4768
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13188 2922 13216 3470
rect 13280 3074 13308 4082
rect 13464 4049 13492 6054
rect 13556 5710 13584 6287
rect 13728 6258 13780 6264
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13556 5166 13584 5510
rect 13740 5370 13768 6258
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 14002 6216 14058 6225
rect 13832 6089 13860 6190
rect 14002 6151 14058 6160
rect 13912 6112 13964 6118
rect 13818 6080 13874 6089
rect 13912 6054 13964 6060
rect 13818 6015 13874 6024
rect 13818 5944 13874 5953
rect 13818 5879 13874 5888
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4826 13676 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13450 4040 13506 4049
rect 13450 3975 13506 3984
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13452 3936 13504 3942
rect 13740 3890 13768 5034
rect 13832 3942 13860 5879
rect 13452 3878 13504 3884
rect 13372 3194 13400 3878
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13280 3046 13400 3074
rect 13464 3058 13492 3878
rect 13648 3862 13768 3890
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 12808 2576 12860 2582
rect 12808 2518 12860 2524
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11808 480 11836 2314
rect 12820 480 12848 2518
rect 13372 2446 13400 3046
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13556 2650 13584 3334
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13648 2530 13676 3862
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13832 3194 13860 3606
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13924 2922 13952 6054
rect 14016 4826 14044 6151
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14116 5468 14412 5488
rect 14172 5466 14196 5468
rect 14252 5466 14276 5468
rect 14332 5466 14356 5468
rect 14194 5414 14196 5466
rect 14258 5414 14270 5466
rect 14332 5414 14334 5466
rect 14172 5412 14196 5414
rect 14252 5412 14276 5414
rect 14332 5412 14356 5414
rect 14116 5392 14412 5412
rect 14476 5166 14504 5646
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 2990 14044 4626
rect 14476 4622 14504 5102
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14116 4380 14412 4400
rect 14172 4378 14196 4380
rect 14252 4378 14276 4380
rect 14332 4378 14356 4380
rect 14194 4326 14196 4378
rect 14258 4326 14270 4378
rect 14332 4326 14334 4378
rect 14172 4324 14196 4326
rect 14252 4324 14276 4326
rect 14332 4324 14356 4326
rect 14116 4304 14412 4324
rect 14476 4146 14504 4558
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14108 3670 14136 4082
rect 14476 3738 14504 4082
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14116 3292 14412 3312
rect 14172 3290 14196 3292
rect 14252 3290 14276 3292
rect 14332 3290 14356 3292
rect 14194 3238 14196 3290
rect 14258 3238 14270 3290
rect 14332 3238 14334 3290
rect 14172 3236 14196 3238
rect 14252 3236 14276 3238
rect 14332 3236 14356 3238
rect 14116 3216 14412 3236
rect 14476 3126 14504 3674
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13648 2502 13768 2530
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13740 480 13768 2502
rect 14568 2378 14596 9574
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14740 9376 14792 9382
rect 14646 9344 14702 9353
rect 14740 9318 14792 9324
rect 14646 9279 14702 9288
rect 14660 9081 14688 9279
rect 14646 9072 14702 9081
rect 14646 9007 14702 9016
rect 14660 8022 14688 9007
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14660 3641 14688 7482
rect 14646 3632 14702 3641
rect 14646 3567 14702 3576
rect 14752 3058 14780 9318
rect 14844 8265 14872 10406
rect 14922 10367 14978 10376
rect 14936 9926 14964 10367
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 15028 9738 15056 10934
rect 14936 9710 15056 9738
rect 14936 8430 14964 9710
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15028 9364 15056 9522
rect 15120 9518 15148 13670
rect 15212 12714 15240 13874
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13530 15516 13670
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15212 12102 15240 12650
rect 15580 12442 15608 13806
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 10538 15240 11494
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15212 10198 15240 10474
rect 15304 10305 15332 11154
rect 15488 11082 15516 12242
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15290 10296 15346 10305
rect 15396 10266 15424 10950
rect 15672 10810 15700 13670
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15290 10231 15346 10240
rect 15384 10260 15436 10266
rect 15200 10192 15252 10198
rect 15200 10134 15252 10140
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15212 9586 15240 9862
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15198 9480 15254 9489
rect 15198 9415 15254 9424
rect 15028 9336 15148 9364
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14830 8256 14886 8265
rect 14830 8191 14886 8200
rect 15028 7886 15056 8434
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14844 4690 14872 7754
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 7041 14964 7686
rect 15028 7342 15056 7822
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14922 7032 14978 7041
rect 14922 6967 14978 6976
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14936 5370 14964 6802
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15028 6338 15056 6598
rect 15120 6497 15148 9336
rect 15106 6488 15162 6497
rect 15106 6423 15162 6432
rect 15028 6310 15148 6338
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14924 4548 14976 4554
rect 14924 4490 14976 4496
rect 14832 4480 14884 4486
rect 14936 4457 14964 4490
rect 14832 4422 14884 4428
rect 14922 4448 14978 4457
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 13832 1873 13860 2314
rect 14116 2204 14412 2224
rect 14172 2202 14196 2204
rect 14252 2202 14276 2204
rect 14332 2202 14356 2204
rect 14194 2150 14196 2202
rect 14258 2150 14270 2202
rect 14332 2150 14334 2202
rect 14172 2148 14196 2150
rect 14252 2148 14276 2150
rect 14332 2148 14356 2150
rect 14116 2128 14412 2148
rect 13818 1864 13874 1873
rect 13818 1799 13874 1808
rect 14660 480 14688 2382
rect 14844 1057 14872 4422
rect 14922 4383 14978 4392
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14936 2922 14964 3470
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 15028 2394 15056 5034
rect 15120 3505 15148 6310
rect 15212 4078 15240 9415
rect 15304 8362 15332 10231
rect 15384 10202 15436 10208
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15382 10024 15438 10033
rect 15764 9994 15792 10134
rect 15856 10062 15884 12038
rect 15948 11762 15976 13330
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16040 12238 16068 13194
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15948 11121 15976 11154
rect 16040 11150 16068 12174
rect 16028 11144 16080 11150
rect 15934 11112 15990 11121
rect 16028 11086 16080 11092
rect 15934 11047 15990 11056
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15382 9959 15438 9968
rect 15752 9988 15804 9994
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 4826 15332 6598
rect 15396 5914 15424 9959
rect 15752 9930 15804 9936
rect 15948 9897 15976 11047
rect 16040 10130 16068 11086
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 15934 9888 15990 9897
rect 15934 9823 15990 9832
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15396 4078 15424 5510
rect 15488 4146 15516 8230
rect 15580 6866 15608 8502
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15672 6730 15700 7890
rect 15856 7886 15884 8434
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15764 4826 15792 7686
rect 15856 7206 15884 7822
rect 16132 7426 16160 12582
rect 16224 10169 16252 14991
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16210 10160 16266 10169
rect 16210 10095 16266 10104
rect 16224 8430 16252 10095
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16210 7848 16266 7857
rect 16210 7783 16266 7792
rect 16224 7546 16252 7783
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16132 7398 16252 7426
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 6798 15884 7142
rect 16040 6934 16068 7278
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15856 6254 15884 6734
rect 15844 6248 15896 6254
rect 15896 6196 15976 6202
rect 15844 6190 15976 6196
rect 15856 6174 15976 6190
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15856 4622 15884 6054
rect 15948 5710 15976 6174
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3738 15700 3878
rect 15764 3738 15792 4422
rect 15856 4214 15884 4558
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15106 3496 15162 3505
rect 15106 3431 15162 3440
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15120 2990 15148 3334
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15028 2366 15148 2394
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 14936 1465 14964 2246
rect 14922 1456 14978 1465
rect 14922 1391 14978 1400
rect 14830 1048 14886 1057
rect 14830 983 14886 992
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3238 0 3294 480
rect 4250 0 4306 480
rect 5170 0 5226 480
rect 6090 0 6146 480
rect 7102 0 7158 480
rect 8022 0 8078 480
rect 8942 0 8998 480
rect 9954 0 10010 480
rect 10874 0 10930 480
rect 11794 0 11850 480
rect 12806 0 12862 480
rect 13726 0 13782 480
rect 14646 0 14702 480
rect 15028 241 15056 2246
rect 15120 649 15148 2366
rect 15106 640 15162 649
rect 15106 575 15162 584
rect 15672 480 15700 2858
rect 16132 2281 16160 6054
rect 16224 5681 16252 7398
rect 16210 5672 16266 5681
rect 16210 5607 16266 5616
rect 16316 4865 16344 14214
rect 16408 13394 16436 16623
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16408 5914 16436 13330
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16302 4856 16358 4865
rect 16302 4791 16358 4800
rect 16118 2272 16174 2281
rect 16118 2207 16174 2216
rect 16592 480 16620 9386
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17512 480 17540 2994
rect 15014 232 15070 241
rect 15014 167 15070 176
rect 15658 0 15714 480
rect 16578 0 16634 480
rect 17498 0 17554 480
<< via2 >>
rect 3514 16632 3570 16688
rect 16394 16632 16450 16688
rect 1306 15408 1362 15464
rect 2042 14592 2098 14648
rect 1858 12688 1914 12744
rect 1398 10124 1454 10160
rect 1398 10104 1400 10124
rect 1400 10104 1452 10124
rect 1452 10104 1454 10124
rect 1582 10512 1638 10568
rect 1582 9988 1638 10024
rect 1582 9968 1584 9988
rect 1584 9968 1636 9988
rect 1636 9968 1638 9988
rect 1306 9288 1362 9344
rect 1674 8336 1730 8392
rect 1582 7112 1638 7168
rect 3238 14184 3294 14240
rect 1858 9832 1914 9888
rect 2134 8608 2190 8664
rect 2318 12008 2374 12064
rect 2502 9424 2558 9480
rect 1766 3576 1822 3632
rect 754 1400 810 1456
rect 2778 9016 2834 9072
rect 2962 9696 3018 9752
rect 2594 8336 2650 8392
rect 3238 11736 3294 11792
rect 3146 10376 3202 10432
rect 3054 9152 3110 9208
rect 2962 6432 3018 6488
rect 2870 4800 2926 4856
rect 2778 4392 2834 4448
rect 3238 10260 3294 10296
rect 3238 10240 3240 10260
rect 3240 10240 3292 10260
rect 3292 10240 3294 10260
rect 3238 9988 3294 10024
rect 3422 12708 3478 12744
rect 3422 12688 3424 12708
rect 3424 12688 3476 12708
rect 3476 12688 3478 12708
rect 4066 16224 4122 16280
rect 14922 16224 14978 16280
rect 4894 15816 4950 15872
rect 4066 15000 4122 15056
rect 3588 14170 3644 14172
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3588 14118 3614 14170
rect 3614 14118 3644 14170
rect 3668 14118 3678 14170
rect 3678 14118 3724 14170
rect 3748 14118 3794 14170
rect 3794 14118 3804 14170
rect 3828 14118 3858 14170
rect 3858 14118 3884 14170
rect 3588 14116 3644 14118
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3974 13812 3976 13832
rect 3976 13812 4028 13832
rect 4028 13812 4030 13832
rect 3974 13776 4030 13812
rect 14462 15408 14518 15464
rect 6220 14714 6276 14716
rect 6300 14714 6356 14716
rect 6380 14714 6436 14716
rect 6460 14714 6516 14716
rect 6220 14662 6246 14714
rect 6246 14662 6276 14714
rect 6300 14662 6310 14714
rect 6310 14662 6356 14714
rect 6380 14662 6426 14714
rect 6426 14662 6436 14714
rect 6460 14662 6490 14714
rect 6490 14662 6516 14714
rect 6220 14660 6276 14662
rect 6300 14660 6356 14662
rect 6380 14660 6436 14662
rect 6460 14660 6516 14662
rect 3588 13082 3644 13084
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3588 13030 3614 13082
rect 3614 13030 3644 13082
rect 3668 13030 3678 13082
rect 3678 13030 3724 13082
rect 3748 13030 3794 13082
rect 3794 13030 3804 13082
rect 3828 13030 3858 13082
rect 3858 13030 3884 13082
rect 3588 13028 3644 13030
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3588 11994 3644 11996
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3588 11942 3614 11994
rect 3614 11942 3644 11994
rect 3668 11942 3678 11994
rect 3678 11942 3724 11994
rect 3748 11942 3794 11994
rect 3794 11942 3804 11994
rect 3828 11942 3858 11994
rect 3858 11942 3884 11994
rect 3588 11940 3644 11942
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3882 11600 3938 11656
rect 3588 10906 3644 10908
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3588 10854 3614 10906
rect 3614 10854 3644 10906
rect 3668 10854 3678 10906
rect 3678 10854 3724 10906
rect 3748 10854 3794 10906
rect 3794 10854 3804 10906
rect 3828 10854 3858 10906
rect 3858 10854 3884 10906
rect 3588 10852 3644 10854
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3514 10412 3516 10432
rect 3516 10412 3568 10432
rect 3568 10412 3570 10432
rect 3514 10376 3570 10412
rect 3238 9968 3240 9988
rect 3240 9968 3292 9988
rect 3292 9968 3294 9988
rect 3330 9832 3386 9888
rect 3238 9696 3294 9752
rect 3238 9288 3294 9344
rect 3588 9818 3644 9820
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3588 9766 3614 9818
rect 3614 9766 3644 9818
rect 3668 9766 3678 9818
rect 3678 9766 3724 9818
rect 3748 9766 3794 9818
rect 3794 9766 3804 9818
rect 3828 9766 3858 9818
rect 3858 9766 3884 9818
rect 3588 9764 3644 9766
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3790 9288 3846 9344
rect 3882 8880 3938 8936
rect 3588 8730 3644 8732
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3588 8678 3614 8730
rect 3614 8678 3644 8730
rect 3668 8678 3678 8730
rect 3678 8678 3724 8730
rect 3748 8678 3794 8730
rect 3794 8678 3804 8730
rect 3828 8678 3858 8730
rect 3858 8678 3884 8730
rect 3588 8676 3644 8678
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3882 8472 3938 8528
rect 3514 7948 3570 7984
rect 3514 7928 3516 7948
rect 3516 7928 3568 7948
rect 3568 7928 3570 7948
rect 4066 9832 4122 9888
rect 4434 12824 4490 12880
rect 4342 9288 4398 9344
rect 4066 8608 4122 8664
rect 4158 7928 4214 7984
rect 3974 7792 4030 7848
rect 3588 7642 3644 7644
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3588 7590 3614 7642
rect 3614 7590 3644 7642
rect 3668 7590 3678 7642
rect 3678 7590 3724 7642
rect 3748 7590 3794 7642
rect 3794 7590 3804 7642
rect 3828 7590 3858 7642
rect 3858 7590 3884 7642
rect 3588 7588 3644 7590
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3238 6840 3294 6896
rect 3146 6296 3202 6352
rect 3054 3576 3110 3632
rect 3514 7384 3570 7440
rect 3514 6976 3570 7032
rect 3588 6554 3644 6556
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3588 6502 3614 6554
rect 3614 6502 3644 6554
rect 3668 6502 3678 6554
rect 3678 6502 3724 6554
rect 3748 6502 3794 6554
rect 3794 6502 3804 6554
rect 3828 6502 3858 6554
rect 3858 6502 3884 6554
rect 3588 6500 3644 6502
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 5170 13676 5172 13696
rect 5172 13676 5224 13696
rect 5224 13676 5226 13696
rect 5170 13640 5226 13676
rect 5354 12688 5410 12744
rect 5078 10648 5134 10704
rect 4894 9696 4950 9752
rect 4250 7384 4306 7440
rect 4250 6740 4252 6760
rect 4252 6740 4304 6760
rect 4304 6740 4306 6760
rect 4250 6704 4306 6740
rect 3882 6024 3938 6080
rect 4066 5616 4122 5672
rect 3588 5466 3644 5468
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3588 5414 3614 5466
rect 3614 5414 3644 5466
rect 3668 5414 3678 5466
rect 3678 5414 3724 5466
rect 3748 5414 3794 5466
rect 3794 5414 3804 5466
rect 3828 5414 3858 5466
rect 3858 5414 3884 5466
rect 3588 5412 3644 5414
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 4066 5208 4122 5264
rect 3422 5072 3478 5128
rect 3974 5072 4030 5128
rect 3330 4936 3386 4992
rect 2962 1808 3018 1864
rect 2870 584 2926 640
rect 3588 4378 3644 4380
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3588 4326 3614 4378
rect 3614 4326 3644 4378
rect 3668 4326 3678 4378
rect 3678 4326 3724 4378
rect 3748 4326 3794 4378
rect 3794 4326 3804 4378
rect 3828 4326 3858 4378
rect 3858 4326 3884 4378
rect 3588 4324 3644 4326
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3514 3984 3570 4040
rect 3588 3290 3644 3292
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3588 3238 3614 3290
rect 3614 3238 3644 3290
rect 3668 3238 3678 3290
rect 3678 3238 3724 3290
rect 3748 3238 3794 3290
rect 3794 3238 3804 3290
rect 3828 3238 3858 3290
rect 3858 3238 3884 3290
rect 3588 3236 3644 3238
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 4066 4564 4068 4584
rect 4068 4564 4120 4584
rect 4120 4564 4122 4584
rect 4066 4528 4122 4564
rect 4250 4528 4306 4584
rect 3974 3032 4030 3088
rect 3698 2624 3754 2680
rect 4158 2508 4214 2544
rect 4158 2488 4160 2508
rect 4160 2488 4212 2508
rect 4212 2488 4214 2508
rect 3422 2216 3478 2272
rect 3588 2202 3644 2204
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3588 2150 3614 2202
rect 3614 2150 3644 2202
rect 3668 2150 3678 2202
rect 3678 2150 3724 2202
rect 3748 2150 3794 2202
rect 3794 2150 3804 2202
rect 3828 2150 3858 2202
rect 3858 2150 3884 2202
rect 3588 2148 3644 2150
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 4710 9288 4766 9344
rect 5170 9968 5226 10024
rect 4710 6996 4766 7032
rect 4710 6976 4712 6996
rect 4712 6976 4764 6996
rect 4764 6976 4766 6996
rect 4710 6568 4766 6624
rect 5446 9324 5448 9344
rect 5448 9324 5500 9344
rect 5500 9324 5502 9344
rect 5446 9288 5502 9324
rect 5354 9152 5410 9208
rect 5170 8880 5226 8936
rect 5262 8608 5318 8664
rect 5262 7248 5318 7304
rect 5262 3848 5318 3904
rect 5814 11192 5870 11248
rect 6220 13626 6276 13628
rect 6300 13626 6356 13628
rect 6380 13626 6436 13628
rect 6460 13626 6516 13628
rect 6220 13574 6246 13626
rect 6246 13574 6276 13626
rect 6300 13574 6310 13626
rect 6310 13574 6356 13626
rect 6380 13574 6426 13626
rect 6426 13574 6436 13626
rect 6460 13574 6490 13626
rect 6490 13574 6516 13626
rect 6220 13572 6276 13574
rect 6300 13572 6356 13574
rect 6380 13572 6436 13574
rect 6460 13572 6516 13574
rect 6220 12538 6276 12540
rect 6300 12538 6356 12540
rect 6380 12538 6436 12540
rect 6460 12538 6516 12540
rect 6220 12486 6246 12538
rect 6246 12486 6276 12538
rect 6300 12486 6310 12538
rect 6310 12486 6356 12538
rect 6380 12486 6426 12538
rect 6426 12486 6436 12538
rect 6460 12486 6490 12538
rect 6490 12486 6516 12538
rect 6220 12484 6276 12486
rect 6300 12484 6356 12486
rect 6380 12484 6436 12486
rect 6460 12484 6516 12486
rect 6220 11450 6276 11452
rect 6300 11450 6356 11452
rect 6380 11450 6436 11452
rect 6460 11450 6516 11452
rect 6220 11398 6246 11450
rect 6246 11398 6276 11450
rect 6300 11398 6310 11450
rect 6310 11398 6356 11450
rect 6380 11398 6426 11450
rect 6426 11398 6436 11450
rect 6460 11398 6490 11450
rect 6490 11398 6516 11450
rect 6220 11396 6276 11398
rect 6300 11396 6356 11398
rect 6380 11396 6436 11398
rect 6460 11396 6516 11398
rect 5814 9036 5870 9072
rect 5814 9016 5816 9036
rect 5816 9016 5868 9036
rect 5868 9016 5870 9036
rect 5722 6976 5778 7032
rect 5722 6432 5778 6488
rect 5538 5480 5594 5536
rect 5354 3440 5410 3496
rect 3698 1028 3700 1048
rect 3700 1028 3752 1048
rect 3752 1028 3754 1048
rect 3698 992 3754 1028
rect 5906 8200 5962 8256
rect 6550 10512 6606 10568
rect 6220 10362 6276 10364
rect 6300 10362 6356 10364
rect 6380 10362 6436 10364
rect 6460 10362 6516 10364
rect 6220 10310 6246 10362
rect 6246 10310 6276 10362
rect 6300 10310 6310 10362
rect 6310 10310 6356 10362
rect 6380 10310 6426 10362
rect 6426 10310 6436 10362
rect 6460 10310 6490 10362
rect 6490 10310 6516 10362
rect 6220 10308 6276 10310
rect 6300 10308 6356 10310
rect 6380 10308 6436 10310
rect 6460 10308 6516 10310
rect 6220 9274 6276 9276
rect 6300 9274 6356 9276
rect 6380 9274 6436 9276
rect 6460 9274 6516 9276
rect 6220 9222 6246 9274
rect 6246 9222 6276 9274
rect 6300 9222 6310 9274
rect 6310 9222 6356 9274
rect 6380 9222 6426 9274
rect 6426 9222 6436 9274
rect 6460 9222 6490 9274
rect 6490 9222 6516 9274
rect 6220 9220 6276 9222
rect 6300 9220 6356 9222
rect 6380 9220 6436 9222
rect 6460 9220 6516 9222
rect 6220 8186 6276 8188
rect 6300 8186 6356 8188
rect 6380 8186 6436 8188
rect 6460 8186 6516 8188
rect 6220 8134 6246 8186
rect 6246 8134 6276 8186
rect 6300 8134 6310 8186
rect 6310 8134 6356 8186
rect 6380 8134 6426 8186
rect 6426 8134 6436 8186
rect 6460 8134 6490 8186
rect 6490 8134 6516 8186
rect 6220 8132 6276 8134
rect 6300 8132 6356 8134
rect 6380 8132 6436 8134
rect 6460 8132 6516 8134
rect 6182 7828 6184 7848
rect 6184 7828 6236 7848
rect 6236 7828 6238 7848
rect 6182 7792 6238 7828
rect 6220 7098 6276 7100
rect 6300 7098 6356 7100
rect 6380 7098 6436 7100
rect 6460 7098 6516 7100
rect 6220 7046 6246 7098
rect 6246 7046 6276 7098
rect 6300 7046 6310 7098
rect 6310 7046 6356 7098
rect 6380 7046 6426 7098
rect 6426 7046 6436 7098
rect 6460 7046 6490 7098
rect 6490 7046 6516 7098
rect 6220 7044 6276 7046
rect 6300 7044 6356 7046
rect 6380 7044 6436 7046
rect 6460 7044 6516 7046
rect 6458 6180 6514 6216
rect 6458 6160 6460 6180
rect 6460 6160 6512 6180
rect 6512 6160 6514 6180
rect 5998 4800 6054 4856
rect 5906 3984 5962 4040
rect 6220 6010 6276 6012
rect 6300 6010 6356 6012
rect 6380 6010 6436 6012
rect 6460 6010 6516 6012
rect 6220 5958 6246 6010
rect 6246 5958 6276 6010
rect 6300 5958 6310 6010
rect 6310 5958 6356 6010
rect 6380 5958 6426 6010
rect 6426 5958 6436 6010
rect 6460 5958 6490 6010
rect 6490 5958 6516 6010
rect 6220 5956 6276 5958
rect 6300 5956 6356 5958
rect 6380 5956 6436 5958
rect 6460 5956 6516 5958
rect 6220 4922 6276 4924
rect 6300 4922 6356 4924
rect 6380 4922 6436 4924
rect 6460 4922 6516 4924
rect 6220 4870 6246 4922
rect 6246 4870 6276 4922
rect 6300 4870 6310 4922
rect 6310 4870 6356 4922
rect 6380 4870 6426 4922
rect 6426 4870 6436 4922
rect 6460 4870 6490 4922
rect 6490 4870 6516 4922
rect 6220 4868 6276 4870
rect 6300 4868 6356 4870
rect 6380 4868 6436 4870
rect 6460 4868 6516 4870
rect 6220 3834 6276 3836
rect 6300 3834 6356 3836
rect 6380 3834 6436 3836
rect 6460 3834 6516 3836
rect 6220 3782 6246 3834
rect 6246 3782 6276 3834
rect 6300 3782 6310 3834
rect 6310 3782 6356 3834
rect 6380 3782 6426 3834
rect 6426 3782 6436 3834
rect 6460 3782 6490 3834
rect 6490 3782 6516 3834
rect 6220 3780 6276 3782
rect 6300 3780 6356 3782
rect 6380 3780 6436 3782
rect 6460 3780 6516 3782
rect 6826 12980 6882 13016
rect 6826 12960 6828 12980
rect 6828 12960 6880 12980
rect 6880 12960 6882 12980
rect 6826 8064 6882 8120
rect 6734 6296 6790 6352
rect 6734 4936 6790 4992
rect 6220 2746 6276 2748
rect 6300 2746 6356 2748
rect 6380 2746 6436 2748
rect 6460 2746 6516 2748
rect 6220 2694 6246 2746
rect 6246 2694 6276 2746
rect 6300 2694 6310 2746
rect 6310 2694 6356 2746
rect 6380 2694 6426 2746
rect 6426 2694 6436 2746
rect 6460 2694 6490 2746
rect 6490 2694 6516 2746
rect 6220 2692 6276 2694
rect 6300 2692 6356 2694
rect 6380 2692 6436 2694
rect 6460 2692 6516 2694
rect 7102 11736 7158 11792
rect 7378 9832 7434 9888
rect 7286 6704 7342 6760
rect 7102 3596 7158 3632
rect 7102 3576 7104 3596
rect 7104 3576 7156 3596
rect 7156 3576 7158 3596
rect 6918 2488 6974 2544
rect 7378 2644 7434 2680
rect 7378 2624 7380 2644
rect 7380 2624 7432 2644
rect 7432 2624 7434 2644
rect 7654 9696 7710 9752
rect 7654 9424 7710 9480
rect 7562 6432 7618 6488
rect 8298 12280 8354 12336
rect 8298 10240 8354 10296
rect 8114 7812 8170 7848
rect 8852 14170 8908 14172
rect 8932 14170 8988 14172
rect 9012 14170 9068 14172
rect 9092 14170 9148 14172
rect 8852 14118 8878 14170
rect 8878 14118 8908 14170
rect 8932 14118 8942 14170
rect 8942 14118 8988 14170
rect 9012 14118 9058 14170
rect 9058 14118 9068 14170
rect 9092 14118 9122 14170
rect 9122 14118 9148 14170
rect 8852 14116 8908 14118
rect 8932 14116 8988 14118
rect 9012 14116 9068 14118
rect 9092 14116 9148 14118
rect 11484 14714 11540 14716
rect 11564 14714 11620 14716
rect 11644 14714 11700 14716
rect 11724 14714 11780 14716
rect 11484 14662 11510 14714
rect 11510 14662 11540 14714
rect 11564 14662 11574 14714
rect 11574 14662 11620 14714
rect 11644 14662 11690 14714
rect 11690 14662 11700 14714
rect 11724 14662 11754 14714
rect 11754 14662 11780 14714
rect 11484 14660 11540 14662
rect 11564 14660 11620 14662
rect 11644 14660 11700 14662
rect 11724 14660 11780 14662
rect 8850 13776 8906 13832
rect 8850 13232 8906 13288
rect 8852 13082 8908 13084
rect 8932 13082 8988 13084
rect 9012 13082 9068 13084
rect 9092 13082 9148 13084
rect 8852 13030 8878 13082
rect 8878 13030 8908 13082
rect 8932 13030 8942 13082
rect 8942 13030 8988 13082
rect 9012 13030 9058 13082
rect 9058 13030 9068 13082
rect 9092 13030 9122 13082
rect 9122 13030 9148 13082
rect 8852 13028 8908 13030
rect 8932 13028 8988 13030
rect 9012 13028 9068 13030
rect 9092 13028 9148 13030
rect 8852 11994 8908 11996
rect 8932 11994 8988 11996
rect 9012 11994 9068 11996
rect 9092 11994 9148 11996
rect 8852 11942 8878 11994
rect 8878 11942 8908 11994
rect 8932 11942 8942 11994
rect 8942 11942 8988 11994
rect 9012 11942 9058 11994
rect 9058 11942 9068 11994
rect 9092 11942 9122 11994
rect 9122 11942 9148 11994
rect 8852 11940 8908 11942
rect 8932 11940 8988 11942
rect 9012 11940 9068 11942
rect 9092 11940 9148 11942
rect 8482 9832 8538 9888
rect 8666 9560 8722 9616
rect 8114 7792 8116 7812
rect 8116 7792 8168 7812
rect 8168 7792 8170 7812
rect 7930 5480 7986 5536
rect 7838 3984 7894 4040
rect 8206 4548 8262 4584
rect 8206 4528 8208 4548
rect 8208 4528 8260 4548
rect 8260 4528 8262 4548
rect 8114 3032 8170 3088
rect 8852 10906 8908 10908
rect 8932 10906 8988 10908
rect 9012 10906 9068 10908
rect 9092 10906 9148 10908
rect 8852 10854 8878 10906
rect 8878 10854 8908 10906
rect 8932 10854 8942 10906
rect 8942 10854 8988 10906
rect 9012 10854 9058 10906
rect 9058 10854 9068 10906
rect 9092 10854 9122 10906
rect 9122 10854 9148 10906
rect 8852 10852 8908 10854
rect 8932 10852 8988 10854
rect 9012 10852 9068 10854
rect 9092 10852 9148 10854
rect 9126 10376 9182 10432
rect 8852 9818 8908 9820
rect 8932 9818 8988 9820
rect 9012 9818 9068 9820
rect 9092 9818 9148 9820
rect 8852 9766 8878 9818
rect 8878 9766 8908 9818
rect 8932 9766 8942 9818
rect 8942 9766 8988 9818
rect 9012 9766 9058 9818
rect 9058 9766 9068 9818
rect 9092 9766 9122 9818
rect 9122 9766 9148 9818
rect 8852 9764 8908 9766
rect 8932 9764 8988 9766
rect 9012 9764 9068 9766
rect 9092 9764 9148 9766
rect 9678 11736 9734 11792
rect 9494 10240 9550 10296
rect 10138 12824 10194 12880
rect 9494 9696 9550 9752
rect 8852 8730 8908 8732
rect 8932 8730 8988 8732
rect 9012 8730 9068 8732
rect 9092 8730 9148 8732
rect 8852 8678 8878 8730
rect 8878 8678 8908 8730
rect 8932 8678 8942 8730
rect 8942 8678 8988 8730
rect 9012 8678 9058 8730
rect 9058 8678 9068 8730
rect 9092 8678 9122 8730
rect 9122 8678 9148 8730
rect 8852 8676 8908 8678
rect 8932 8676 8988 8678
rect 9012 8676 9068 8678
rect 9092 8676 9148 8678
rect 9402 8880 9458 8936
rect 8852 7642 8908 7644
rect 8932 7642 8988 7644
rect 9012 7642 9068 7644
rect 9092 7642 9148 7644
rect 8852 7590 8878 7642
rect 8878 7590 8908 7642
rect 8932 7590 8942 7642
rect 8942 7590 8988 7642
rect 9012 7590 9058 7642
rect 9058 7590 9068 7642
rect 9092 7590 9122 7642
rect 9122 7590 9148 7642
rect 8852 7588 8908 7590
rect 8932 7588 8988 7590
rect 9012 7588 9068 7590
rect 9092 7588 9148 7590
rect 9586 9560 9642 9616
rect 9862 9968 9918 10024
rect 9770 8608 9826 8664
rect 8852 6554 8908 6556
rect 8932 6554 8988 6556
rect 9012 6554 9068 6556
rect 9092 6554 9148 6556
rect 8852 6502 8878 6554
rect 8878 6502 8908 6554
rect 8932 6502 8942 6554
rect 8942 6502 8988 6554
rect 9012 6502 9058 6554
rect 9058 6502 9068 6554
rect 9092 6502 9122 6554
rect 9122 6502 9148 6554
rect 8852 6500 8908 6502
rect 8932 6500 8988 6502
rect 9012 6500 9068 6502
rect 9092 6500 9148 6502
rect 9402 6296 9458 6352
rect 9310 6160 9366 6216
rect 9218 6024 9274 6080
rect 8852 5466 8908 5468
rect 8932 5466 8988 5468
rect 9012 5466 9068 5468
rect 9092 5466 9148 5468
rect 8852 5414 8878 5466
rect 8878 5414 8908 5466
rect 8932 5414 8942 5466
rect 8942 5414 8988 5466
rect 9012 5414 9058 5466
rect 9058 5414 9068 5466
rect 9092 5414 9122 5466
rect 9122 5414 9148 5466
rect 8852 5412 8908 5414
rect 8932 5412 8988 5414
rect 9012 5412 9068 5414
rect 9092 5412 9148 5414
rect 8852 4378 8908 4380
rect 8932 4378 8988 4380
rect 9012 4378 9068 4380
rect 9092 4378 9148 4380
rect 8852 4326 8878 4378
rect 8878 4326 8908 4378
rect 8932 4326 8942 4378
rect 8942 4326 8988 4378
rect 9012 4326 9058 4378
rect 9058 4326 9068 4378
rect 9092 4326 9122 4378
rect 9122 4326 9148 4378
rect 8852 4324 8908 4326
rect 8932 4324 8988 4326
rect 9012 4324 9068 4326
rect 9092 4324 9148 4326
rect 8942 3440 8998 3496
rect 8852 3290 8908 3292
rect 8932 3290 8988 3292
rect 9012 3290 9068 3292
rect 9092 3290 9148 3292
rect 8852 3238 8878 3290
rect 8878 3238 8908 3290
rect 8932 3238 8942 3290
rect 8942 3238 8988 3290
rect 9012 3238 9058 3290
rect 9058 3238 9068 3290
rect 9092 3238 9122 3290
rect 9122 3238 9148 3290
rect 8852 3236 8908 3238
rect 8932 3236 8988 3238
rect 9012 3236 9068 3238
rect 9092 3236 9148 3238
rect 8942 3052 8998 3088
rect 8942 3032 8944 3052
rect 8944 3032 8996 3052
rect 8996 3032 8998 3052
rect 9034 2896 9090 2952
rect 9126 2760 9182 2816
rect 8852 2202 8908 2204
rect 8932 2202 8988 2204
rect 9012 2202 9068 2204
rect 9092 2202 9148 2204
rect 8852 2150 8878 2202
rect 8878 2150 8908 2202
rect 8932 2150 8942 2202
rect 8942 2150 8988 2202
rect 9012 2150 9058 2202
rect 9058 2150 9068 2202
rect 9092 2150 9122 2202
rect 9122 2150 9148 2202
rect 8852 2148 8908 2150
rect 8932 2148 8988 2150
rect 9012 2148 9068 2150
rect 9092 2148 9148 2150
rect 9954 7792 10010 7848
rect 10414 12824 10470 12880
rect 10506 11600 10562 11656
rect 10506 10648 10562 10704
rect 9954 7248 10010 7304
rect 9954 6976 10010 7032
rect 10506 9832 10562 9888
rect 14116 14170 14172 14172
rect 14196 14170 14252 14172
rect 14276 14170 14332 14172
rect 14356 14170 14412 14172
rect 14116 14118 14142 14170
rect 14142 14118 14172 14170
rect 14196 14118 14206 14170
rect 14206 14118 14252 14170
rect 14276 14118 14322 14170
rect 14322 14118 14332 14170
rect 14356 14118 14386 14170
rect 14386 14118 14412 14170
rect 14116 14116 14172 14118
rect 14196 14116 14252 14118
rect 14276 14116 14332 14118
rect 14356 14116 14412 14118
rect 11484 13626 11540 13628
rect 11564 13626 11620 13628
rect 11644 13626 11700 13628
rect 11724 13626 11780 13628
rect 11484 13574 11510 13626
rect 11510 13574 11540 13626
rect 11564 13574 11574 13626
rect 11574 13574 11620 13626
rect 11644 13574 11690 13626
rect 11690 13574 11700 13626
rect 11724 13574 11754 13626
rect 11754 13574 11780 13626
rect 11484 13572 11540 13574
rect 11564 13572 11620 13574
rect 11644 13572 11700 13574
rect 11724 13572 11780 13574
rect 11484 12538 11540 12540
rect 11564 12538 11620 12540
rect 11644 12538 11700 12540
rect 11724 12538 11780 12540
rect 11484 12486 11510 12538
rect 11510 12486 11540 12538
rect 11564 12486 11574 12538
rect 11574 12486 11620 12538
rect 11644 12486 11690 12538
rect 11690 12486 11700 12538
rect 11724 12486 11754 12538
rect 11754 12486 11780 12538
rect 11484 12484 11540 12486
rect 11564 12484 11620 12486
rect 11644 12484 11700 12486
rect 11724 12484 11780 12486
rect 11242 11056 11298 11112
rect 11058 9560 11114 9616
rect 10874 8472 10930 8528
rect 10598 6876 10600 6896
rect 10600 6876 10652 6896
rect 10652 6876 10654 6896
rect 10598 6840 10654 6876
rect 10782 6316 10838 6352
rect 10782 6296 10784 6316
rect 10784 6296 10836 6316
rect 10836 6296 10838 6316
rect 10506 6160 10562 6216
rect 11484 11450 11540 11452
rect 11564 11450 11620 11452
rect 11644 11450 11700 11452
rect 11724 11450 11780 11452
rect 11484 11398 11510 11450
rect 11510 11398 11540 11450
rect 11564 11398 11574 11450
rect 11574 11398 11620 11450
rect 11644 11398 11690 11450
rect 11690 11398 11700 11450
rect 11724 11398 11754 11450
rect 11754 11398 11780 11450
rect 11484 11396 11540 11398
rect 11564 11396 11620 11398
rect 11644 11396 11700 11398
rect 11724 11396 11780 11398
rect 11794 11192 11850 11248
rect 11484 10362 11540 10364
rect 11564 10362 11620 10364
rect 11644 10362 11700 10364
rect 11724 10362 11780 10364
rect 11484 10310 11510 10362
rect 11510 10310 11540 10362
rect 11564 10310 11574 10362
rect 11574 10310 11620 10362
rect 11644 10310 11690 10362
rect 11690 10310 11700 10362
rect 11724 10310 11754 10362
rect 11754 10310 11780 10362
rect 11484 10308 11540 10310
rect 11564 10308 11620 10310
rect 11644 10308 11700 10310
rect 11724 10308 11780 10310
rect 11426 9832 11482 9888
rect 11702 9560 11758 9616
rect 11426 9444 11482 9480
rect 11426 9424 11428 9444
rect 11428 9424 11480 9444
rect 11480 9424 11482 9444
rect 11610 9460 11612 9480
rect 11612 9460 11664 9480
rect 11664 9460 11666 9480
rect 11610 9424 11666 9460
rect 11484 9274 11540 9276
rect 11564 9274 11620 9276
rect 11644 9274 11700 9276
rect 11724 9274 11780 9276
rect 11484 9222 11510 9274
rect 11510 9222 11540 9274
rect 11564 9222 11574 9274
rect 11574 9222 11620 9274
rect 11644 9222 11690 9274
rect 11690 9222 11700 9274
rect 11724 9222 11754 9274
rect 11754 9222 11780 9274
rect 11484 9220 11540 9222
rect 11564 9220 11620 9222
rect 11644 9220 11700 9222
rect 11724 9220 11780 9222
rect 11242 9016 11298 9072
rect 11484 8186 11540 8188
rect 11564 8186 11620 8188
rect 11644 8186 11700 8188
rect 11724 8186 11780 8188
rect 11484 8134 11510 8186
rect 11510 8134 11540 8186
rect 11564 8134 11574 8186
rect 11574 8134 11620 8186
rect 11644 8134 11690 8186
rect 11690 8134 11700 8186
rect 11724 8134 11754 8186
rect 11754 8134 11780 8186
rect 11484 8132 11540 8134
rect 11564 8132 11620 8134
rect 11644 8132 11700 8134
rect 11724 8132 11780 8134
rect 12346 12144 12402 12200
rect 12530 12144 12586 12200
rect 12438 11192 12494 11248
rect 11886 10376 11942 10432
rect 12162 9560 12218 9616
rect 12070 9152 12126 9208
rect 12070 8236 12072 8256
rect 12072 8236 12124 8256
rect 12124 8236 12126 8256
rect 12070 8200 12126 8236
rect 11886 7928 11942 7984
rect 11978 7248 12034 7304
rect 11484 7098 11540 7100
rect 11564 7098 11620 7100
rect 11644 7098 11700 7100
rect 11724 7098 11780 7100
rect 11484 7046 11510 7098
rect 11510 7046 11540 7098
rect 11564 7046 11574 7098
rect 11574 7046 11620 7098
rect 11644 7046 11690 7098
rect 11690 7046 11700 7098
rect 11724 7046 11754 7098
rect 11754 7046 11780 7098
rect 11484 7044 11540 7046
rect 11564 7044 11620 7046
rect 11644 7044 11700 7046
rect 11724 7044 11780 7046
rect 11794 6704 11850 6760
rect 11484 6010 11540 6012
rect 11564 6010 11620 6012
rect 11644 6010 11700 6012
rect 11724 6010 11780 6012
rect 11484 5958 11510 6010
rect 11510 5958 11540 6010
rect 11564 5958 11574 6010
rect 11574 5958 11620 6010
rect 11644 5958 11690 6010
rect 11690 5958 11700 6010
rect 11724 5958 11754 6010
rect 11754 5958 11780 6010
rect 11484 5956 11540 5958
rect 11564 5956 11620 5958
rect 11644 5956 11700 5958
rect 11724 5956 11780 5958
rect 11484 4922 11540 4924
rect 11564 4922 11620 4924
rect 11644 4922 11700 4924
rect 11724 4922 11780 4924
rect 11484 4870 11510 4922
rect 11510 4870 11540 4922
rect 11564 4870 11574 4922
rect 11574 4870 11620 4922
rect 11644 4870 11690 4922
rect 11690 4870 11700 4922
rect 11724 4870 11754 4922
rect 11754 4870 11780 4922
rect 11484 4868 11540 4870
rect 11564 4868 11620 4870
rect 11644 4868 11700 4870
rect 11724 4868 11780 4870
rect 11484 3834 11540 3836
rect 11564 3834 11620 3836
rect 11644 3834 11700 3836
rect 11724 3834 11780 3836
rect 11484 3782 11510 3834
rect 11510 3782 11540 3834
rect 11564 3782 11574 3834
rect 11574 3782 11620 3834
rect 11644 3782 11690 3834
rect 11690 3782 11700 3834
rect 11724 3782 11754 3834
rect 11754 3782 11780 3834
rect 11484 3780 11540 3782
rect 11564 3780 11620 3782
rect 11644 3780 11700 3782
rect 11724 3780 11780 3782
rect 11484 2746 11540 2748
rect 11564 2746 11620 2748
rect 11644 2746 11700 2748
rect 11724 2746 11780 2748
rect 11484 2694 11510 2746
rect 11510 2694 11540 2746
rect 11564 2694 11574 2746
rect 11574 2694 11620 2746
rect 11644 2694 11690 2746
rect 11690 2694 11700 2746
rect 11724 2694 11754 2746
rect 11754 2694 11780 2746
rect 11484 2692 11540 2694
rect 11564 2692 11620 2694
rect 11644 2692 11700 2694
rect 11724 2692 11780 2694
rect 12622 10648 12678 10704
rect 12346 10240 12402 10296
rect 12530 9832 12586 9888
rect 12346 9696 12402 9752
rect 12438 9424 12494 9480
rect 12346 9016 12402 9072
rect 13082 12164 13138 12200
rect 13082 12144 13084 12164
rect 13084 12144 13136 12164
rect 13136 12144 13138 12164
rect 14002 13776 14058 13832
rect 13910 13232 13966 13288
rect 13542 12552 13598 12608
rect 13174 11212 13230 11248
rect 13174 11192 13176 11212
rect 13176 11192 13228 11212
rect 13228 11192 13230 11212
rect 12990 9560 13046 9616
rect 12530 8608 12586 8664
rect 12346 7384 12402 7440
rect 12438 6704 12494 6760
rect 12254 5208 12310 5264
rect 12990 8472 13046 8528
rect 12622 8200 12678 8256
rect 12806 7928 12862 7984
rect 12714 7384 12770 7440
rect 13266 10104 13322 10160
rect 13542 7928 13598 7984
rect 13082 6840 13138 6896
rect 11978 2624 12034 2680
rect 13910 12552 13966 12608
rect 15014 15816 15070 15872
rect 14830 14592 14886 14648
rect 14646 14184 14702 14240
rect 14116 13082 14172 13084
rect 14196 13082 14252 13084
rect 14276 13082 14332 13084
rect 14356 13082 14412 13084
rect 14116 13030 14142 13082
rect 14142 13030 14172 13082
rect 14196 13030 14206 13082
rect 14206 13030 14252 13082
rect 14276 13030 14322 13082
rect 14322 13030 14332 13082
rect 14356 13030 14386 13082
rect 14386 13030 14412 13082
rect 14116 13028 14172 13030
rect 14196 13028 14252 13030
rect 14276 13028 14332 13030
rect 14356 13028 14412 13030
rect 13910 12144 13966 12200
rect 14116 11994 14172 11996
rect 14196 11994 14252 11996
rect 14276 11994 14332 11996
rect 14356 11994 14412 11996
rect 14116 11942 14142 11994
rect 14142 11942 14172 11994
rect 14196 11942 14206 11994
rect 14206 11942 14252 11994
rect 14276 11942 14322 11994
rect 14322 11942 14332 11994
rect 14356 11942 14386 11994
rect 14386 11942 14412 11994
rect 14116 11940 14172 11942
rect 14196 11940 14252 11942
rect 14276 11940 14332 11942
rect 14356 11940 14412 11942
rect 13726 9152 13782 9208
rect 14116 10906 14172 10908
rect 14196 10906 14252 10908
rect 14276 10906 14332 10908
rect 14356 10906 14412 10908
rect 14116 10854 14142 10906
rect 14142 10854 14172 10906
rect 14196 10854 14206 10906
rect 14206 10854 14252 10906
rect 14276 10854 14322 10906
rect 14322 10854 14332 10906
rect 14356 10854 14386 10906
rect 14386 10854 14412 10906
rect 14116 10852 14172 10854
rect 14196 10852 14252 10854
rect 14276 10852 14332 10854
rect 14356 10852 14412 10854
rect 14002 10648 14058 10704
rect 13910 9696 13966 9752
rect 14186 10376 14242 10432
rect 14116 9818 14172 9820
rect 14196 9818 14252 9820
rect 14276 9818 14332 9820
rect 14356 9818 14412 9820
rect 14116 9766 14142 9818
rect 14142 9766 14172 9818
rect 14196 9766 14206 9818
rect 14206 9766 14252 9818
rect 14276 9766 14322 9818
rect 14322 9766 14332 9818
rect 14356 9766 14386 9818
rect 14386 9766 14412 9818
rect 14116 9764 14172 9766
rect 14196 9764 14252 9766
rect 14276 9764 14332 9766
rect 14356 9764 14412 9766
rect 14094 9596 14096 9616
rect 14096 9596 14148 9616
rect 14148 9596 14150 9616
rect 14094 9560 14150 9596
rect 16210 15000 16266 15056
rect 14922 12416 14978 12472
rect 13542 6296 13598 6352
rect 13818 7384 13874 7440
rect 13818 7284 13820 7304
rect 13820 7284 13872 7304
rect 13872 7284 13874 7304
rect 13818 7248 13874 7284
rect 14462 8916 14464 8936
rect 14464 8916 14516 8936
rect 14516 8916 14518 8936
rect 14462 8880 14518 8916
rect 14116 8730 14172 8732
rect 14196 8730 14252 8732
rect 14276 8730 14332 8732
rect 14356 8730 14412 8732
rect 14116 8678 14142 8730
rect 14142 8678 14172 8730
rect 14196 8678 14206 8730
rect 14206 8678 14252 8730
rect 14276 8678 14322 8730
rect 14322 8678 14332 8730
rect 14356 8678 14386 8730
rect 14386 8678 14412 8730
rect 14116 8676 14172 8678
rect 14196 8676 14252 8678
rect 14276 8676 14332 8678
rect 14356 8676 14412 8678
rect 14116 7642 14172 7644
rect 14196 7642 14252 7644
rect 14276 7642 14332 7644
rect 14356 7642 14412 7644
rect 14116 7590 14142 7642
rect 14142 7590 14172 7642
rect 14196 7590 14206 7642
rect 14206 7590 14252 7642
rect 14276 7590 14322 7642
rect 14322 7590 14332 7642
rect 14356 7590 14386 7642
rect 14386 7590 14412 7642
rect 14116 7588 14172 7590
rect 14196 7588 14252 7590
rect 14276 7588 14332 7590
rect 14356 7588 14412 7590
rect 14116 6554 14172 6556
rect 14196 6554 14252 6556
rect 14276 6554 14332 6556
rect 14356 6554 14412 6556
rect 14116 6502 14142 6554
rect 14142 6502 14172 6554
rect 14196 6502 14206 6554
rect 14206 6502 14252 6554
rect 14276 6502 14322 6554
rect 14322 6502 14332 6554
rect 14356 6502 14386 6554
rect 14386 6502 14412 6554
rect 14116 6500 14172 6502
rect 14196 6500 14252 6502
rect 14276 6500 14332 6502
rect 14356 6500 14412 6502
rect 14002 6160 14058 6216
rect 13818 6024 13874 6080
rect 13818 5888 13874 5944
rect 13450 3984 13506 4040
rect 14116 5466 14172 5468
rect 14196 5466 14252 5468
rect 14276 5466 14332 5468
rect 14356 5466 14412 5468
rect 14116 5414 14142 5466
rect 14142 5414 14172 5466
rect 14196 5414 14206 5466
rect 14206 5414 14252 5466
rect 14276 5414 14322 5466
rect 14322 5414 14332 5466
rect 14356 5414 14386 5466
rect 14386 5414 14412 5466
rect 14116 5412 14172 5414
rect 14196 5412 14252 5414
rect 14276 5412 14332 5414
rect 14356 5412 14412 5414
rect 14116 4378 14172 4380
rect 14196 4378 14252 4380
rect 14276 4378 14332 4380
rect 14356 4378 14412 4380
rect 14116 4326 14142 4378
rect 14142 4326 14172 4378
rect 14196 4326 14206 4378
rect 14206 4326 14252 4378
rect 14276 4326 14322 4378
rect 14322 4326 14332 4378
rect 14356 4326 14386 4378
rect 14386 4326 14412 4378
rect 14116 4324 14172 4326
rect 14196 4324 14252 4326
rect 14276 4324 14332 4326
rect 14356 4324 14412 4326
rect 14116 3290 14172 3292
rect 14196 3290 14252 3292
rect 14276 3290 14332 3292
rect 14356 3290 14412 3292
rect 14116 3238 14142 3290
rect 14142 3238 14172 3290
rect 14196 3238 14206 3290
rect 14206 3238 14252 3290
rect 14276 3238 14322 3290
rect 14322 3238 14332 3290
rect 14356 3238 14386 3290
rect 14386 3238 14412 3290
rect 14116 3236 14172 3238
rect 14196 3236 14252 3238
rect 14276 3236 14332 3238
rect 14356 3236 14412 3238
rect 14646 9288 14702 9344
rect 14646 9016 14702 9072
rect 14646 3576 14702 3632
rect 14922 10376 14978 10432
rect 15290 10240 15346 10296
rect 15198 9424 15254 9480
rect 14830 8200 14886 8256
rect 14922 6976 14978 7032
rect 15106 6432 15162 6488
rect 14116 2202 14172 2204
rect 14196 2202 14252 2204
rect 14276 2202 14332 2204
rect 14356 2202 14412 2204
rect 14116 2150 14142 2202
rect 14142 2150 14172 2202
rect 14196 2150 14206 2202
rect 14206 2150 14252 2202
rect 14276 2150 14322 2202
rect 14322 2150 14332 2202
rect 14356 2150 14386 2202
rect 14386 2150 14412 2202
rect 14116 2148 14172 2150
rect 14196 2148 14252 2150
rect 14276 2148 14332 2150
rect 14356 2148 14412 2150
rect 13818 1808 13874 1864
rect 14922 4392 14978 4448
rect 15382 9968 15438 10024
rect 15934 11056 15990 11112
rect 15934 9832 15990 9888
rect 16210 10104 16266 10160
rect 16210 7792 16266 7848
rect 15106 3440 15162 3496
rect 14922 1400 14978 1456
rect 14830 992 14886 1048
rect 2778 176 2834 232
rect 15106 584 15162 640
rect 16210 5616 16266 5672
rect 16302 4800 16358 4856
rect 16118 2216 16174 2272
rect 15014 176 15070 232
<< metal3 >>
rect 0 16690 480 16720
rect 3509 16690 3575 16693
rect 0 16688 3575 16690
rect 0 16632 3514 16688
rect 3570 16632 3575 16688
rect 0 16630 3575 16632
rect 0 16600 480 16630
rect 3509 16627 3575 16630
rect 16389 16690 16455 16693
rect 17520 16690 18000 16720
rect 16389 16688 18000 16690
rect 16389 16632 16394 16688
rect 16450 16632 18000 16688
rect 16389 16630 18000 16632
rect 16389 16627 16455 16630
rect 17520 16600 18000 16630
rect 0 16282 480 16312
rect 4061 16282 4127 16285
rect 0 16280 4127 16282
rect 0 16224 4066 16280
rect 4122 16224 4127 16280
rect 0 16222 4127 16224
rect 0 16192 480 16222
rect 4061 16219 4127 16222
rect 14917 16282 14983 16285
rect 17520 16282 18000 16312
rect 14917 16280 18000 16282
rect 14917 16224 14922 16280
rect 14978 16224 18000 16280
rect 14917 16222 18000 16224
rect 14917 16219 14983 16222
rect 17520 16192 18000 16222
rect 0 15874 480 15904
rect 4889 15874 4955 15877
rect 0 15872 4955 15874
rect 0 15816 4894 15872
rect 4950 15816 4955 15872
rect 0 15814 4955 15816
rect 0 15784 480 15814
rect 4889 15811 4955 15814
rect 15009 15874 15075 15877
rect 17520 15874 18000 15904
rect 15009 15872 18000 15874
rect 15009 15816 15014 15872
rect 15070 15816 18000 15872
rect 15009 15814 18000 15816
rect 15009 15811 15075 15814
rect 17520 15784 18000 15814
rect 0 15466 480 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 480 15406
rect 1301 15403 1367 15406
rect 14457 15466 14523 15469
rect 17520 15466 18000 15496
rect 14457 15464 18000 15466
rect 14457 15408 14462 15464
rect 14518 15408 18000 15464
rect 14457 15406 18000 15408
rect 14457 15403 14523 15406
rect 17520 15376 18000 15406
rect 0 15058 480 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 480 14998
rect 4061 14995 4127 14998
rect 16205 15058 16271 15061
rect 17520 15058 18000 15088
rect 16205 15056 18000 15058
rect 16205 15000 16210 15056
rect 16266 15000 18000 15056
rect 16205 14998 18000 15000
rect 16205 14995 16271 14998
rect 17520 14968 18000 14998
rect 6208 14720 6528 14721
rect 0 14650 480 14680
rect 6208 14656 6216 14720
rect 6280 14656 6296 14720
rect 6360 14656 6376 14720
rect 6440 14656 6456 14720
rect 6520 14656 6528 14720
rect 6208 14655 6528 14656
rect 11472 14720 11792 14721
rect 11472 14656 11480 14720
rect 11544 14656 11560 14720
rect 11624 14656 11640 14720
rect 11704 14656 11720 14720
rect 11784 14656 11792 14720
rect 11472 14655 11792 14656
rect 2037 14650 2103 14653
rect 0 14648 2103 14650
rect 0 14592 2042 14648
rect 2098 14592 2103 14648
rect 0 14590 2103 14592
rect 0 14560 480 14590
rect 2037 14587 2103 14590
rect 14825 14650 14891 14653
rect 17520 14650 18000 14680
rect 14825 14648 18000 14650
rect 14825 14592 14830 14648
rect 14886 14592 18000 14648
rect 14825 14590 18000 14592
rect 14825 14587 14891 14590
rect 17520 14560 18000 14590
rect 0 14242 480 14272
rect 3233 14242 3299 14245
rect 0 14240 3299 14242
rect 0 14184 3238 14240
rect 3294 14184 3299 14240
rect 0 14182 3299 14184
rect 0 14152 480 14182
rect 3233 14179 3299 14182
rect 14641 14242 14707 14245
rect 17520 14242 18000 14272
rect 14641 14240 18000 14242
rect 14641 14184 14646 14240
rect 14702 14184 18000 14240
rect 14641 14182 18000 14184
rect 14641 14179 14707 14182
rect 3576 14176 3896 14177
rect 3576 14112 3584 14176
rect 3648 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3896 14176
rect 3576 14111 3896 14112
rect 8840 14176 9160 14177
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8840 14111 9160 14112
rect 14104 14176 14424 14177
rect 14104 14112 14112 14176
rect 14176 14112 14192 14176
rect 14256 14112 14272 14176
rect 14336 14112 14352 14176
rect 14416 14112 14424 14176
rect 17520 14152 18000 14182
rect 14104 14111 14424 14112
rect 0 13834 480 13864
rect 3969 13834 4035 13837
rect 8845 13834 8911 13837
rect 0 13832 4035 13834
rect 0 13776 3974 13832
rect 4030 13776 4035 13832
rect 0 13774 4035 13776
rect 0 13744 480 13774
rect 3969 13771 4035 13774
rect 5168 13832 8911 13834
rect 5168 13776 8850 13832
rect 8906 13776 8911 13832
rect 5168 13774 8911 13776
rect 5168 13701 5228 13774
rect 8845 13771 8911 13774
rect 13997 13834 14063 13837
rect 17520 13834 18000 13864
rect 13997 13832 18000 13834
rect 13997 13776 14002 13832
rect 14058 13776 18000 13832
rect 13997 13774 18000 13776
rect 13997 13771 14063 13774
rect 17520 13744 18000 13774
rect 4654 13636 4660 13700
rect 4724 13698 4730 13700
rect 5165 13698 5231 13701
rect 4724 13696 5231 13698
rect 4724 13640 5170 13696
rect 5226 13640 5231 13696
rect 4724 13638 5231 13640
rect 4724 13636 4730 13638
rect 5165 13635 5231 13638
rect 6208 13632 6528 13633
rect 6208 13568 6216 13632
rect 6280 13568 6296 13632
rect 6360 13568 6376 13632
rect 6440 13568 6456 13632
rect 6520 13568 6528 13632
rect 6208 13567 6528 13568
rect 11472 13632 11792 13633
rect 11472 13568 11480 13632
rect 11544 13568 11560 13632
rect 11624 13568 11640 13632
rect 11704 13568 11720 13632
rect 11784 13568 11792 13632
rect 11472 13567 11792 13568
rect 0 13290 480 13320
rect 8845 13290 8911 13293
rect 0 13288 8911 13290
rect 0 13232 8850 13288
rect 8906 13232 8911 13288
rect 0 13230 8911 13232
rect 0 13200 480 13230
rect 8845 13227 8911 13230
rect 13905 13290 13971 13293
rect 17520 13290 18000 13320
rect 13905 13288 18000 13290
rect 13905 13232 13910 13288
rect 13966 13232 18000 13288
rect 13905 13230 18000 13232
rect 13905 13227 13971 13230
rect 17520 13200 18000 13230
rect 3576 13088 3896 13089
rect 3576 13024 3584 13088
rect 3648 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3896 13088
rect 3576 13023 3896 13024
rect 8840 13088 9160 13089
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 8840 13023 9160 13024
rect 14104 13088 14424 13089
rect 14104 13024 14112 13088
rect 14176 13024 14192 13088
rect 14256 13024 14272 13088
rect 14336 13024 14352 13088
rect 14416 13024 14424 13088
rect 14104 13023 14424 13024
rect 6821 13018 6887 13021
rect 4294 13016 6887 13018
rect 4294 12960 6826 13016
rect 6882 12960 6887 13016
rect 4294 12958 6887 12960
rect 0 12882 480 12912
rect 4294 12882 4354 12958
rect 6821 12955 6887 12958
rect 0 12822 4354 12882
rect 4429 12882 4495 12885
rect 7414 12882 7420 12884
rect 4429 12880 7420 12882
rect 4429 12824 4434 12880
rect 4490 12824 7420 12880
rect 4429 12822 7420 12824
rect 0 12792 480 12822
rect 4429 12819 4495 12822
rect 7414 12820 7420 12822
rect 7484 12820 7490 12884
rect 10133 12882 10199 12885
rect 10409 12882 10475 12885
rect 17520 12882 18000 12912
rect 10133 12880 18000 12882
rect 10133 12824 10138 12880
rect 10194 12824 10414 12880
rect 10470 12824 18000 12880
rect 10133 12822 18000 12824
rect 10133 12819 10199 12822
rect 10409 12819 10475 12822
rect 17520 12792 18000 12822
rect 1853 12746 1919 12749
rect 3417 12746 3483 12749
rect 5349 12746 5415 12749
rect 1853 12744 5415 12746
rect 1853 12688 1858 12744
rect 1914 12688 3422 12744
rect 3478 12688 5354 12744
rect 5410 12688 5415 12744
rect 1853 12686 5415 12688
rect 1853 12683 1919 12686
rect 3417 12683 3483 12686
rect 5349 12683 5415 12686
rect 13537 12610 13603 12613
rect 13905 12610 13971 12613
rect 13537 12608 13971 12610
rect 13537 12552 13542 12608
rect 13598 12552 13910 12608
rect 13966 12552 13971 12608
rect 13537 12550 13971 12552
rect 13537 12547 13603 12550
rect 13905 12547 13971 12550
rect 6208 12544 6528 12545
rect 0 12474 480 12504
rect 6208 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6528 12544
rect 6208 12479 6528 12480
rect 11472 12544 11792 12545
rect 11472 12480 11480 12544
rect 11544 12480 11560 12544
rect 11624 12480 11640 12544
rect 11704 12480 11720 12544
rect 11784 12480 11792 12544
rect 11472 12479 11792 12480
rect 14917 12474 14983 12477
rect 17520 12474 18000 12504
rect 0 12414 4538 12474
rect 0 12384 480 12414
rect 4478 12338 4538 12414
rect 14917 12472 18000 12474
rect 14917 12416 14922 12472
rect 14978 12416 18000 12472
rect 14917 12414 18000 12416
rect 14917 12411 14983 12414
rect 17520 12384 18000 12414
rect 8293 12338 8359 12341
rect 4478 12336 8359 12338
rect 4478 12280 8298 12336
rect 8354 12280 8359 12336
rect 4478 12278 8359 12280
rect 8293 12275 8359 12278
rect 12341 12202 12407 12205
rect 12525 12202 12591 12205
rect 12341 12200 12591 12202
rect 12341 12144 12346 12200
rect 12402 12144 12530 12200
rect 12586 12144 12591 12200
rect 12341 12142 12591 12144
rect 12341 12139 12407 12142
rect 12525 12139 12591 12142
rect 13077 12202 13143 12205
rect 13905 12202 13971 12205
rect 13077 12200 13971 12202
rect 13077 12144 13082 12200
rect 13138 12144 13910 12200
rect 13966 12144 13971 12200
rect 13077 12142 13971 12144
rect 13077 12139 13143 12142
rect 13905 12139 13971 12142
rect 0 12066 480 12096
rect 2313 12066 2379 12069
rect 17520 12066 18000 12096
rect 0 12064 2379 12066
rect 0 12008 2318 12064
rect 2374 12008 2379 12064
rect 0 12006 2379 12008
rect 0 11976 480 12006
rect 2313 12003 2379 12006
rect 14782 12006 18000 12066
rect 3576 12000 3896 12001
rect 3576 11936 3584 12000
rect 3648 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3896 12000
rect 3576 11935 3896 11936
rect 8840 12000 9160 12001
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8840 11935 9160 11936
rect 14104 12000 14424 12001
rect 14104 11936 14112 12000
rect 14176 11936 14192 12000
rect 14256 11936 14272 12000
rect 14336 11936 14352 12000
rect 14416 11936 14424 12000
rect 14104 11935 14424 11936
rect 3233 11794 3299 11797
rect 7097 11794 7163 11797
rect 3233 11792 7163 11794
rect 3233 11736 3238 11792
rect 3294 11736 7102 11792
rect 7158 11736 7163 11792
rect 3233 11734 7163 11736
rect 3233 11731 3299 11734
rect 7097 11731 7163 11734
rect 9673 11794 9739 11797
rect 14782 11794 14842 12006
rect 17520 11976 18000 12006
rect 9673 11792 14842 11794
rect 9673 11736 9678 11792
rect 9734 11736 14842 11792
rect 9673 11734 14842 11736
rect 9673 11731 9739 11734
rect 0 11658 480 11688
rect 3877 11658 3943 11661
rect 0 11656 3943 11658
rect 0 11600 3882 11656
rect 3938 11600 3943 11656
rect 0 11598 3943 11600
rect 0 11568 480 11598
rect 3877 11595 3943 11598
rect 10501 11658 10567 11661
rect 17520 11658 18000 11688
rect 10501 11656 18000 11658
rect 10501 11600 10506 11656
rect 10562 11600 18000 11656
rect 10501 11598 18000 11600
rect 10501 11595 10567 11598
rect 17520 11568 18000 11598
rect 6208 11456 6528 11457
rect 6208 11392 6216 11456
rect 6280 11392 6296 11456
rect 6360 11392 6376 11456
rect 6440 11392 6456 11456
rect 6520 11392 6528 11456
rect 6208 11391 6528 11392
rect 11472 11456 11792 11457
rect 11472 11392 11480 11456
rect 11544 11392 11560 11456
rect 11624 11392 11640 11456
rect 11704 11392 11720 11456
rect 11784 11392 11792 11456
rect 11472 11391 11792 11392
rect 0 11250 480 11280
rect 5809 11250 5875 11253
rect 0 11248 5875 11250
rect 0 11192 5814 11248
rect 5870 11192 5875 11248
rect 0 11190 5875 11192
rect 0 11160 480 11190
rect 5809 11187 5875 11190
rect 11789 11250 11855 11253
rect 12433 11250 12499 11253
rect 11789 11248 12499 11250
rect 11789 11192 11794 11248
rect 11850 11192 12438 11248
rect 12494 11192 12499 11248
rect 11789 11190 12499 11192
rect 11789 11187 11855 11190
rect 12433 11187 12499 11190
rect 13169 11250 13235 11253
rect 17520 11250 18000 11280
rect 13169 11248 18000 11250
rect 13169 11192 13174 11248
rect 13230 11192 18000 11248
rect 13169 11190 18000 11192
rect 13169 11187 13235 11190
rect 17520 11160 18000 11190
rect 11237 11114 11303 11117
rect 15929 11114 15995 11117
rect 11237 11112 15995 11114
rect 11237 11056 11242 11112
rect 11298 11056 15934 11112
rect 15990 11056 15995 11112
rect 11237 11054 15995 11056
rect 11237 11051 11303 11054
rect 15929 11051 15995 11054
rect 3576 10912 3896 10913
rect 0 10842 480 10872
rect 3576 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3896 10912
rect 3576 10847 3896 10848
rect 8840 10912 9160 10913
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 10847 9160 10848
rect 14104 10912 14424 10913
rect 14104 10848 14112 10912
rect 14176 10848 14192 10912
rect 14256 10848 14272 10912
rect 14336 10848 14352 10912
rect 14416 10848 14424 10912
rect 14104 10847 14424 10848
rect 17520 10842 18000 10872
rect 0 10782 3480 10842
rect 0 10752 480 10782
rect 3420 10706 3480 10782
rect 14552 10782 18000 10842
rect 5073 10706 5139 10709
rect 3420 10704 5139 10706
rect 3420 10648 5078 10704
rect 5134 10648 5139 10704
rect 3420 10646 5139 10648
rect 5073 10643 5139 10646
rect 10501 10706 10567 10709
rect 12617 10706 12683 10709
rect 10501 10704 12683 10706
rect 10501 10648 10506 10704
rect 10562 10648 12622 10704
rect 12678 10648 12683 10704
rect 10501 10646 12683 10648
rect 10501 10643 10567 10646
rect 12617 10643 12683 10646
rect 13997 10706 14063 10709
rect 14552 10706 14612 10782
rect 17520 10752 18000 10782
rect 13997 10704 14612 10706
rect 13997 10648 14002 10704
rect 14058 10648 14612 10704
rect 13997 10646 14612 10648
rect 13997 10643 14063 10646
rect 1577 10570 1643 10573
rect 6545 10570 6611 10573
rect 1577 10568 6611 10570
rect 1577 10512 1582 10568
rect 1638 10512 6550 10568
rect 6606 10512 6611 10568
rect 1577 10510 6611 10512
rect 1577 10507 1643 10510
rect 6545 10507 6611 10510
rect 0 10434 480 10464
rect 3141 10434 3207 10437
rect 3509 10434 3575 10437
rect 0 10432 3575 10434
rect 0 10376 3146 10432
rect 3202 10376 3514 10432
rect 3570 10376 3575 10432
rect 0 10374 3575 10376
rect 0 10344 480 10374
rect 3141 10371 3207 10374
rect 3509 10371 3575 10374
rect 9121 10434 9187 10437
rect 9254 10434 9260 10436
rect 9121 10432 9260 10434
rect 9121 10376 9126 10432
rect 9182 10376 9260 10432
rect 9121 10374 9260 10376
rect 9121 10371 9187 10374
rect 9254 10372 9260 10374
rect 9324 10372 9330 10436
rect 11881 10434 11947 10437
rect 14181 10434 14247 10437
rect 14590 10434 14596 10436
rect 11881 10432 14596 10434
rect 11881 10376 11886 10432
rect 11942 10376 14186 10432
rect 14242 10376 14596 10432
rect 11881 10374 14596 10376
rect 11881 10371 11947 10374
rect 14181 10371 14247 10374
rect 14590 10372 14596 10374
rect 14660 10372 14666 10436
rect 14917 10434 14983 10437
rect 17520 10434 18000 10464
rect 14917 10432 18000 10434
rect 14917 10376 14922 10432
rect 14978 10376 18000 10432
rect 14917 10374 18000 10376
rect 14917 10371 14983 10374
rect 6208 10368 6528 10369
rect 6208 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6528 10368
rect 6208 10303 6528 10304
rect 11472 10368 11792 10369
rect 11472 10304 11480 10368
rect 11544 10304 11560 10368
rect 11624 10304 11640 10368
rect 11704 10304 11720 10368
rect 11784 10304 11792 10368
rect 17520 10344 18000 10374
rect 11472 10303 11792 10304
rect 3233 10300 3299 10301
rect 3182 10236 3188 10300
rect 3252 10298 3299 10300
rect 8293 10298 8359 10301
rect 9489 10298 9555 10301
rect 3252 10296 3344 10298
rect 3294 10240 3344 10296
rect 3252 10238 3344 10240
rect 8293 10296 9555 10298
rect 8293 10240 8298 10296
rect 8354 10240 9494 10296
rect 9550 10240 9555 10296
rect 8293 10238 9555 10240
rect 3252 10236 3299 10238
rect 3233 10235 3299 10236
rect 8293 10235 8359 10238
rect 9489 10235 9555 10238
rect 12341 10298 12407 10301
rect 15285 10298 15351 10301
rect 12341 10296 15351 10298
rect 12341 10240 12346 10296
rect 12402 10240 15290 10296
rect 15346 10240 15351 10296
rect 12341 10238 15351 10240
rect 12341 10235 12407 10238
rect 15285 10235 15351 10238
rect 1393 10162 1459 10165
rect 13261 10162 13327 10165
rect 16205 10162 16271 10165
rect 1393 10160 16271 10162
rect 1393 10104 1398 10160
rect 1454 10104 13266 10160
rect 13322 10104 16210 10160
rect 16266 10104 16271 10160
rect 1393 10102 16271 10104
rect 1393 10099 1459 10102
rect 13261 10099 13327 10102
rect 16205 10099 16271 10102
rect 1577 10026 1643 10029
rect 2814 10026 2820 10028
rect 1577 10024 2820 10026
rect 1577 9968 1582 10024
rect 1638 9968 2820 10024
rect 1577 9966 2820 9968
rect 1577 9963 1643 9966
rect 2814 9964 2820 9966
rect 2884 9964 2890 10028
rect 3233 10026 3299 10029
rect 5165 10026 5231 10029
rect 9857 10026 9923 10029
rect 15377 10026 15443 10029
rect 3233 10024 3434 10026
rect 3233 9968 3238 10024
rect 3294 9968 3434 10024
rect 3233 9966 3434 9968
rect 3233 9963 3299 9966
rect 0 9890 480 9920
rect 3374 9893 3434 9966
rect 5165 10024 9690 10026
rect 5165 9968 5170 10024
rect 5226 9968 9690 10024
rect 5165 9966 9690 9968
rect 5165 9963 5231 9966
rect 1853 9890 1919 9893
rect 0 9888 3250 9890
rect 0 9832 1858 9888
rect 1914 9832 3250 9888
rect 0 9830 3250 9832
rect 0 9800 480 9830
rect 1853 9827 1919 9830
rect 3190 9757 3250 9830
rect 3325 9888 3434 9893
rect 3325 9832 3330 9888
rect 3386 9832 3434 9888
rect 3325 9830 3434 9832
rect 4061 9890 4127 9893
rect 7373 9890 7439 9893
rect 8477 9890 8543 9893
rect 4061 9888 4170 9890
rect 4061 9832 4066 9888
rect 4122 9832 4170 9888
rect 3325 9827 3391 9830
rect 4061 9827 4170 9832
rect 7373 9888 8543 9890
rect 7373 9832 7378 9888
rect 7434 9832 8482 9888
rect 8538 9832 8543 9888
rect 7373 9830 8543 9832
rect 9630 9890 9690 9966
rect 9857 10024 15443 10026
rect 9857 9968 9862 10024
rect 9918 9968 15382 10024
rect 15438 9968 15443 10024
rect 9857 9966 15443 9968
rect 9857 9963 9923 9966
rect 15377 9963 15443 9966
rect 10501 9890 10567 9893
rect 9630 9888 10567 9890
rect 9630 9832 10506 9888
rect 10562 9832 10567 9888
rect 9630 9830 10567 9832
rect 7373 9827 7439 9830
rect 8477 9827 8543 9830
rect 10501 9827 10567 9830
rect 11421 9890 11487 9893
rect 12525 9890 12591 9893
rect 11421 9888 12591 9890
rect 11421 9832 11426 9888
rect 11482 9832 12530 9888
rect 12586 9832 12591 9888
rect 11421 9830 12591 9832
rect 11421 9827 11487 9830
rect 12525 9827 12591 9830
rect 15929 9890 15995 9893
rect 17520 9890 18000 9920
rect 15929 9888 18000 9890
rect 15929 9832 15934 9888
rect 15990 9832 18000 9888
rect 15929 9830 18000 9832
rect 15929 9827 15995 9830
rect 3576 9824 3896 9825
rect 3576 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3896 9824
rect 3576 9759 3896 9760
rect 2814 9692 2820 9756
rect 2884 9754 2890 9756
rect 2957 9754 3023 9757
rect 2884 9752 3023 9754
rect 2884 9696 2962 9752
rect 3018 9696 3023 9752
rect 2884 9694 3023 9696
rect 3190 9752 3299 9757
rect 3190 9696 3238 9752
rect 3294 9696 3299 9752
rect 3190 9694 3299 9696
rect 4110 9754 4170 9827
rect 8840 9824 9160 9825
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8840 9759 9160 9760
rect 14104 9824 14424 9825
rect 14104 9760 14112 9824
rect 14176 9760 14192 9824
rect 14256 9760 14272 9824
rect 14336 9760 14352 9824
rect 14416 9760 14424 9824
rect 17520 9800 18000 9830
rect 14104 9759 14424 9760
rect 4889 9754 4955 9757
rect 7649 9754 7715 9757
rect 4110 9752 7715 9754
rect 4110 9696 4894 9752
rect 4950 9696 7654 9752
rect 7710 9696 7715 9752
rect 4110 9694 7715 9696
rect 2884 9692 2890 9694
rect 2957 9691 3023 9694
rect 3233 9691 3299 9694
rect 4889 9691 4955 9694
rect 7649 9691 7715 9694
rect 9489 9754 9555 9757
rect 12341 9754 12407 9757
rect 13905 9754 13971 9757
rect 9489 9752 12407 9754
rect 9489 9696 9494 9752
rect 9550 9696 12346 9752
rect 12402 9696 12407 9752
rect 9489 9694 12407 9696
rect 9489 9691 9555 9694
rect 12341 9691 12407 9694
rect 13724 9752 13971 9754
rect 13724 9696 13910 9752
rect 13966 9696 13971 9752
rect 13724 9694 13971 9696
rect 8661 9618 8727 9621
rect 4110 9616 8727 9618
rect 4110 9560 8666 9616
rect 8722 9560 8727 9616
rect 4110 9558 8727 9560
rect 0 9482 480 9512
rect 2497 9482 2563 9485
rect 0 9480 2563 9482
rect 0 9424 2502 9480
rect 2558 9424 2563 9480
rect 0 9422 2563 9424
rect 0 9392 480 9422
rect 2497 9419 2563 9422
rect 1301 9346 1367 9349
rect 3233 9346 3299 9349
rect 1301 9344 3299 9346
rect 1301 9288 1306 9344
rect 1362 9288 3238 9344
rect 3294 9288 3299 9344
rect 1301 9286 3299 9288
rect 1301 9283 1367 9286
rect 3233 9283 3299 9286
rect 3785 9346 3851 9349
rect 4110 9348 4170 9558
rect 8661 9555 8727 9558
rect 9438 9556 9444 9620
rect 9508 9618 9514 9620
rect 9581 9618 9647 9621
rect 9508 9616 9647 9618
rect 9508 9560 9586 9616
rect 9642 9560 9647 9616
rect 9508 9558 9647 9560
rect 9508 9556 9514 9558
rect 9581 9555 9647 9558
rect 11053 9618 11119 9621
rect 11697 9618 11763 9621
rect 11053 9616 11763 9618
rect 11053 9560 11058 9616
rect 11114 9560 11702 9616
rect 11758 9560 11763 9616
rect 11053 9558 11763 9560
rect 11053 9555 11119 9558
rect 11697 9555 11763 9558
rect 12157 9618 12223 9621
rect 12985 9618 13051 9621
rect 12157 9616 13051 9618
rect 12157 9560 12162 9616
rect 12218 9560 12990 9616
rect 13046 9560 13051 9616
rect 12157 9558 13051 9560
rect 12157 9555 12223 9558
rect 12985 9555 13051 9558
rect 7649 9482 7715 9485
rect 11421 9482 11487 9485
rect 7649 9480 11487 9482
rect 7649 9424 7654 9480
rect 7710 9424 11426 9480
rect 11482 9424 11487 9480
rect 7649 9422 11487 9424
rect 7649 9419 7715 9422
rect 11421 9419 11487 9422
rect 11605 9482 11671 9485
rect 12433 9482 12499 9485
rect 11605 9480 12499 9482
rect 11605 9424 11610 9480
rect 11666 9424 12438 9480
rect 12494 9424 12499 9480
rect 11605 9422 12499 9424
rect 11605 9419 11671 9422
rect 12433 9419 12499 9422
rect 4102 9346 4108 9348
rect 3785 9344 4108 9346
rect 3785 9288 3790 9344
rect 3846 9288 4108 9344
rect 3785 9286 4108 9288
rect 3785 9283 3851 9286
rect 4102 9284 4108 9286
rect 4172 9284 4178 9348
rect 4337 9346 4403 9349
rect 4705 9346 4771 9349
rect 4337 9344 4771 9346
rect 4337 9288 4342 9344
rect 4398 9288 4710 9344
rect 4766 9288 4771 9344
rect 4337 9286 4771 9288
rect 4337 9283 4403 9286
rect 4705 9283 4771 9286
rect 5441 9346 5507 9349
rect 5574 9346 5580 9348
rect 5441 9344 5580 9346
rect 5441 9288 5446 9344
rect 5502 9288 5580 9344
rect 5441 9286 5580 9288
rect 5441 9283 5507 9286
rect 5574 9284 5580 9286
rect 5644 9284 5650 9348
rect 13724 9346 13784 9694
rect 13905 9691 13971 9694
rect 14590 9692 14596 9756
rect 14660 9692 14666 9756
rect 13854 9556 13860 9620
rect 13924 9618 13930 9620
rect 14089 9618 14155 9621
rect 13924 9616 14155 9618
rect 13924 9560 14094 9616
rect 14150 9560 14155 9616
rect 13924 9558 14155 9560
rect 13924 9556 13930 9558
rect 14089 9555 14155 9558
rect 14598 9482 14658 9692
rect 15193 9482 15259 9485
rect 17520 9482 18000 9512
rect 14598 9480 18000 9482
rect 14598 9424 15198 9480
rect 15254 9424 18000 9480
rect 14598 9422 18000 9424
rect 15193 9419 15259 9422
rect 17520 9392 18000 9422
rect 14641 9346 14707 9349
rect 13724 9344 14707 9346
rect 13724 9288 14646 9344
rect 14702 9288 14707 9344
rect 13724 9286 14707 9288
rect 14641 9283 14707 9286
rect 6208 9280 6528 9281
rect 6208 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6528 9280
rect 6208 9215 6528 9216
rect 11472 9280 11792 9281
rect 11472 9216 11480 9280
rect 11544 9216 11560 9280
rect 11624 9216 11640 9280
rect 11704 9216 11720 9280
rect 11784 9216 11792 9280
rect 11472 9215 11792 9216
rect 3049 9210 3115 9213
rect 5349 9210 5415 9213
rect 3049 9208 5415 9210
rect 3049 9152 3054 9208
rect 3110 9152 5354 9208
rect 5410 9152 5415 9208
rect 3049 9150 5415 9152
rect 3049 9147 3115 9150
rect 5349 9147 5415 9150
rect 12065 9210 12131 9213
rect 13721 9210 13787 9213
rect 12065 9208 13787 9210
rect 12065 9152 12070 9208
rect 12126 9152 13726 9208
rect 13782 9152 13787 9208
rect 12065 9150 13787 9152
rect 12065 9147 12131 9150
rect 13721 9147 13787 9150
rect 0 9074 480 9104
rect 2773 9074 2839 9077
rect 0 9072 2839 9074
rect 0 9016 2778 9072
rect 2834 9016 2839 9072
rect 0 9014 2839 9016
rect 0 8984 480 9014
rect 2773 9011 2839 9014
rect 5809 9074 5875 9077
rect 11237 9074 11303 9077
rect 12341 9074 12407 9077
rect 5809 9072 12407 9074
rect 5809 9016 5814 9072
rect 5870 9016 11242 9072
rect 11298 9016 12346 9072
rect 12402 9016 12407 9072
rect 5809 9014 12407 9016
rect 5809 9011 5875 9014
rect 11237 9011 11303 9014
rect 12341 9011 12407 9014
rect 14641 9074 14707 9077
rect 17520 9074 18000 9104
rect 14641 9072 18000 9074
rect 14641 9016 14646 9072
rect 14702 9016 18000 9072
rect 14641 9014 18000 9016
rect 14641 9011 14707 9014
rect 17520 8984 18000 9014
rect 3877 8938 3943 8941
rect 5165 8938 5231 8941
rect 3877 8936 5231 8938
rect 3877 8880 3882 8936
rect 3938 8880 5170 8936
rect 5226 8880 5231 8936
rect 3877 8878 5231 8880
rect 3877 8875 3943 8878
rect 5165 8875 5231 8878
rect 9397 8938 9463 8941
rect 14457 8938 14523 8941
rect 9397 8936 14523 8938
rect 9397 8880 9402 8936
rect 9458 8880 14462 8936
rect 14518 8880 14523 8936
rect 9397 8878 14523 8880
rect 9397 8875 9463 8878
rect 14457 8875 14523 8878
rect 3576 8736 3896 8737
rect 0 8666 480 8696
rect 3576 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3896 8736
rect 3576 8671 3896 8672
rect 8840 8736 9160 8737
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8840 8671 9160 8672
rect 14104 8736 14424 8737
rect 14104 8672 14112 8736
rect 14176 8672 14192 8736
rect 14256 8672 14272 8736
rect 14336 8672 14352 8736
rect 14416 8672 14424 8736
rect 14104 8671 14424 8672
rect 2129 8666 2195 8669
rect 4061 8666 4127 8669
rect 5257 8666 5323 8669
rect 0 8664 3480 8666
rect 0 8608 2134 8664
rect 2190 8608 3480 8664
rect 0 8606 3480 8608
rect 0 8576 480 8606
rect 2129 8603 2195 8606
rect 3420 8530 3480 8606
rect 4061 8664 5323 8666
rect 4061 8608 4066 8664
rect 4122 8608 5262 8664
rect 5318 8608 5323 8664
rect 4061 8606 5323 8608
rect 4061 8603 4127 8606
rect 5257 8603 5323 8606
rect 9765 8666 9831 8669
rect 12525 8666 12591 8669
rect 17520 8666 18000 8696
rect 9765 8664 12591 8666
rect 9765 8608 9770 8664
rect 9826 8608 12530 8664
rect 12586 8608 12591 8664
rect 9765 8606 12591 8608
rect 9765 8603 9831 8606
rect 12525 8603 12591 8606
rect 15104 8606 18000 8666
rect 3877 8530 3943 8533
rect 3420 8528 3943 8530
rect 3420 8472 3882 8528
rect 3938 8472 3943 8528
rect 3420 8470 3943 8472
rect 3877 8467 3943 8470
rect 10869 8530 10935 8533
rect 12985 8530 13051 8533
rect 10869 8528 13051 8530
rect 10869 8472 10874 8528
rect 10930 8472 12990 8528
rect 13046 8472 13051 8528
rect 10869 8470 13051 8472
rect 10869 8467 10935 8470
rect 12985 8467 13051 8470
rect 13854 8468 13860 8532
rect 13924 8530 13930 8532
rect 15104 8530 15164 8606
rect 17520 8576 18000 8606
rect 13924 8470 15164 8530
rect 13924 8468 13930 8470
rect 1669 8394 1735 8397
rect 2589 8394 2655 8397
rect 9438 8394 9444 8396
rect 1669 8392 9444 8394
rect 1669 8336 1674 8392
rect 1730 8336 2594 8392
rect 2650 8336 9444 8392
rect 1669 8334 9444 8336
rect 1669 8331 1735 8334
rect 2589 8331 2655 8334
rect 9438 8332 9444 8334
rect 9508 8332 9514 8396
rect 0 8258 480 8288
rect 5901 8258 5967 8261
rect 0 8256 5967 8258
rect 0 8200 5906 8256
rect 5962 8200 5967 8256
rect 0 8198 5967 8200
rect 0 8168 480 8198
rect 5901 8195 5967 8198
rect 12065 8258 12131 8261
rect 12617 8258 12683 8261
rect 12065 8256 12683 8258
rect 12065 8200 12070 8256
rect 12126 8200 12622 8256
rect 12678 8200 12683 8256
rect 12065 8198 12683 8200
rect 12065 8195 12131 8198
rect 12617 8195 12683 8198
rect 14825 8258 14891 8261
rect 17520 8258 18000 8288
rect 14825 8256 18000 8258
rect 14825 8200 14830 8256
rect 14886 8200 18000 8256
rect 14825 8198 18000 8200
rect 14825 8195 14891 8198
rect 6208 8192 6528 8193
rect 6208 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6528 8192
rect 6208 8127 6528 8128
rect 11472 8192 11792 8193
rect 11472 8128 11480 8192
rect 11544 8128 11560 8192
rect 11624 8128 11640 8192
rect 11704 8128 11720 8192
rect 11784 8128 11792 8192
rect 17520 8168 18000 8198
rect 11472 8127 11792 8128
rect 6821 8122 6887 8125
rect 8702 8122 8708 8124
rect 6821 8120 8708 8122
rect 6821 8064 6826 8120
rect 6882 8064 8708 8120
rect 6821 8062 8708 8064
rect 6821 8059 6887 8062
rect 8702 8060 8708 8062
rect 8772 8122 8778 8124
rect 8772 8062 11392 8122
rect 8772 8060 8778 8062
rect 3509 7986 3575 7989
rect 4153 7986 4219 7989
rect 3509 7984 4219 7986
rect 3509 7928 3514 7984
rect 3570 7928 4158 7984
rect 4214 7928 4219 7984
rect 3509 7926 4219 7928
rect 3509 7923 3575 7926
rect 4153 7923 4219 7926
rect 0 7850 480 7880
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 480 7790
rect 3969 7787 4035 7790
rect 6177 7850 6243 7853
rect 6678 7850 6684 7852
rect 6177 7848 6684 7850
rect 6177 7792 6182 7848
rect 6238 7792 6684 7848
rect 6177 7790 6684 7792
rect 6177 7787 6243 7790
rect 6678 7788 6684 7790
rect 6748 7788 6754 7852
rect 8109 7850 8175 7853
rect 9949 7850 10015 7853
rect 8109 7848 10015 7850
rect 8109 7792 8114 7848
rect 8170 7792 9954 7848
rect 10010 7792 10015 7848
rect 8109 7790 10015 7792
rect 8109 7787 8175 7790
rect 9949 7787 10015 7790
rect 3576 7648 3896 7649
rect 3576 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3896 7648
rect 3576 7583 3896 7584
rect 8840 7648 9160 7649
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 7583 9160 7584
rect 0 7442 480 7472
rect 3509 7442 3575 7445
rect 0 7440 3575 7442
rect 0 7384 3514 7440
rect 3570 7384 3575 7440
rect 0 7382 3575 7384
rect 0 7352 480 7382
rect 3509 7379 3575 7382
rect 4245 7442 4311 7445
rect 11332 7442 11392 8062
rect 11881 7986 11947 7989
rect 12801 7986 12867 7989
rect 13537 7986 13603 7989
rect 11881 7984 13603 7986
rect 11881 7928 11886 7984
rect 11942 7928 12806 7984
rect 12862 7928 13542 7984
rect 13598 7928 13603 7984
rect 11881 7926 13603 7928
rect 11881 7923 11947 7926
rect 12801 7923 12867 7926
rect 13537 7923 13603 7926
rect 16205 7850 16271 7853
rect 17520 7850 18000 7880
rect 16205 7848 18000 7850
rect 16205 7792 16210 7848
rect 16266 7792 18000 7848
rect 16205 7790 18000 7792
rect 16205 7787 16271 7790
rect 17520 7760 18000 7790
rect 14104 7648 14424 7649
rect 14104 7584 14112 7648
rect 14176 7584 14192 7648
rect 14256 7584 14272 7648
rect 14336 7584 14352 7648
rect 14416 7584 14424 7648
rect 14104 7583 14424 7584
rect 12341 7442 12407 7445
rect 12709 7442 12775 7445
rect 4245 7440 4906 7442
rect 4245 7384 4250 7440
rect 4306 7384 4906 7440
rect 4245 7382 4906 7384
rect 11332 7382 12266 7442
rect 4245 7379 4311 7382
rect 4846 7306 4906 7382
rect 5257 7306 5323 7309
rect 4846 7304 5323 7306
rect 4846 7248 5262 7304
rect 5318 7248 5323 7304
rect 4846 7246 5323 7248
rect 5257 7243 5323 7246
rect 9949 7306 10015 7309
rect 11973 7306 12039 7309
rect 9949 7304 12039 7306
rect 9949 7248 9954 7304
rect 10010 7248 11978 7304
rect 12034 7248 12039 7304
rect 9949 7246 12039 7248
rect 12206 7306 12266 7382
rect 12341 7440 12775 7442
rect 12341 7384 12346 7440
rect 12402 7384 12714 7440
rect 12770 7384 12775 7440
rect 12341 7382 12775 7384
rect 12341 7379 12407 7382
rect 12709 7379 12775 7382
rect 13813 7442 13879 7445
rect 17520 7442 18000 7472
rect 13813 7440 18000 7442
rect 13813 7384 13818 7440
rect 13874 7384 18000 7440
rect 13813 7382 18000 7384
rect 13813 7379 13879 7382
rect 17520 7352 18000 7382
rect 13813 7306 13879 7309
rect 12206 7304 13879 7306
rect 12206 7248 13818 7304
rect 13874 7248 13879 7304
rect 12206 7246 13879 7248
rect 9949 7243 10015 7246
rect 11973 7243 12039 7246
rect 13813 7243 13879 7246
rect 1577 7170 1643 7173
rect 5574 7170 5580 7172
rect 1577 7168 5580 7170
rect 1577 7112 1582 7168
rect 1638 7112 5580 7168
rect 1577 7110 5580 7112
rect 1577 7107 1643 7110
rect 5574 7108 5580 7110
rect 5644 7108 5650 7172
rect 6208 7104 6528 7105
rect 0 7034 480 7064
rect 6208 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6528 7104
rect 6208 7039 6528 7040
rect 11472 7104 11792 7105
rect 11472 7040 11480 7104
rect 11544 7040 11560 7104
rect 11624 7040 11640 7104
rect 11704 7040 11720 7104
rect 11784 7040 11792 7104
rect 11472 7039 11792 7040
rect 3509 7034 3575 7037
rect 0 7032 3575 7034
rect 0 6976 3514 7032
rect 3570 6976 3575 7032
rect 0 6974 3575 6976
rect 0 6944 480 6974
rect 3509 6971 3575 6974
rect 4705 7034 4771 7037
rect 5717 7034 5783 7037
rect 9949 7034 10015 7037
rect 4705 7032 5783 7034
rect 4705 6976 4710 7032
rect 4766 6976 5722 7032
rect 5778 6976 5783 7032
rect 4705 6974 5783 6976
rect 4705 6971 4771 6974
rect 5717 6971 5783 6974
rect 9814 7032 10015 7034
rect 9814 6976 9954 7032
rect 10010 6976 10015 7032
rect 9814 6974 10015 6976
rect 3233 6898 3299 6901
rect 9814 6898 9874 6974
rect 9949 6971 10015 6974
rect 14917 7034 14983 7037
rect 17520 7034 18000 7064
rect 14917 7032 18000 7034
rect 14917 6976 14922 7032
rect 14978 6976 18000 7032
rect 14917 6974 18000 6976
rect 14917 6971 14983 6974
rect 17520 6944 18000 6974
rect 3233 6896 9874 6898
rect 3233 6840 3238 6896
rect 3294 6840 9874 6896
rect 3233 6838 9874 6840
rect 10593 6898 10659 6901
rect 13077 6898 13143 6901
rect 10593 6896 13143 6898
rect 10593 6840 10598 6896
rect 10654 6840 13082 6896
rect 13138 6840 13143 6896
rect 10593 6838 13143 6840
rect 3233 6835 3299 6838
rect 10593 6835 10659 6838
rect 13077 6835 13143 6838
rect 4245 6762 4311 6765
rect 7281 6762 7347 6765
rect 4245 6760 7347 6762
rect 4245 6704 4250 6760
rect 4306 6704 7286 6760
rect 7342 6704 7347 6760
rect 4245 6702 7347 6704
rect 4245 6699 4311 6702
rect 7281 6699 7347 6702
rect 11789 6762 11855 6765
rect 12433 6762 12499 6765
rect 11789 6760 12499 6762
rect 11789 6704 11794 6760
rect 11850 6704 12438 6760
rect 12494 6704 12499 6760
rect 11789 6702 12499 6704
rect 11789 6699 11855 6702
rect 12433 6699 12499 6702
rect 4102 6564 4108 6628
rect 4172 6626 4178 6628
rect 4705 6626 4771 6629
rect 4172 6624 4771 6626
rect 4172 6568 4710 6624
rect 4766 6568 4771 6624
rect 4172 6566 4771 6568
rect 4172 6564 4178 6566
rect 4705 6563 4771 6566
rect 3576 6560 3896 6561
rect 0 6490 480 6520
rect 3576 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3896 6560
rect 3576 6495 3896 6496
rect 8840 6560 9160 6561
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8840 6495 9160 6496
rect 14104 6560 14424 6561
rect 14104 6496 14112 6560
rect 14176 6496 14192 6560
rect 14256 6496 14272 6560
rect 14336 6496 14352 6560
rect 14416 6496 14424 6560
rect 14104 6495 14424 6496
rect 2957 6490 3023 6493
rect 0 6488 3023 6490
rect 0 6432 2962 6488
rect 3018 6432 3023 6488
rect 0 6430 3023 6432
rect 0 6400 480 6430
rect 2957 6427 3023 6430
rect 5717 6490 5783 6493
rect 7557 6490 7623 6493
rect 5717 6488 7623 6490
rect 5717 6432 5722 6488
rect 5778 6432 7562 6488
rect 7618 6432 7623 6488
rect 5717 6430 7623 6432
rect 5717 6427 5783 6430
rect 7557 6427 7623 6430
rect 15101 6490 15167 6493
rect 17520 6490 18000 6520
rect 15101 6488 18000 6490
rect 15101 6432 15106 6488
rect 15162 6432 18000 6488
rect 15101 6430 18000 6432
rect 15101 6427 15167 6430
rect 17520 6400 18000 6430
rect 3141 6356 3207 6357
rect 3141 6354 3188 6356
rect 3096 6352 3188 6354
rect 3096 6296 3146 6352
rect 3096 6294 3188 6296
rect 3141 6292 3188 6294
rect 3252 6292 3258 6356
rect 6729 6354 6795 6357
rect 9397 6354 9463 6357
rect 6729 6352 9463 6354
rect 6729 6296 6734 6352
rect 6790 6296 9402 6352
rect 9458 6296 9463 6352
rect 6729 6294 9463 6296
rect 3141 6291 3207 6292
rect 6729 6291 6795 6294
rect 9397 6291 9463 6294
rect 10777 6354 10843 6357
rect 13537 6354 13603 6357
rect 10777 6352 13603 6354
rect 10777 6296 10782 6352
rect 10838 6296 13542 6352
rect 13598 6296 13603 6352
rect 10777 6294 13603 6296
rect 10777 6291 10843 6294
rect 13537 6291 13603 6294
rect 6453 6218 6519 6221
rect 9305 6218 9371 6221
rect 6453 6216 9371 6218
rect 6453 6160 6458 6216
rect 6514 6160 9310 6216
rect 9366 6160 9371 6216
rect 6453 6158 9371 6160
rect 6453 6155 6519 6158
rect 9305 6155 9371 6158
rect 10501 6218 10567 6221
rect 13997 6218 14063 6221
rect 10501 6216 14063 6218
rect 10501 6160 10506 6216
rect 10562 6160 14002 6216
rect 14058 6160 14063 6216
rect 10501 6158 14063 6160
rect 10501 6155 10567 6158
rect 13997 6155 14063 6158
rect 0 6082 480 6112
rect 3877 6082 3943 6085
rect 0 6080 3943 6082
rect 0 6024 3882 6080
rect 3938 6024 3943 6080
rect 0 6022 3943 6024
rect 0 5992 480 6022
rect 3877 6019 3943 6022
rect 9213 6084 9279 6085
rect 9213 6080 9260 6084
rect 9324 6082 9330 6084
rect 13813 6082 13879 6085
rect 17520 6082 18000 6112
rect 9213 6024 9218 6080
rect 9213 6020 9260 6024
rect 9324 6022 9370 6082
rect 13813 6080 18000 6082
rect 13813 6024 13818 6080
rect 13874 6024 18000 6080
rect 13813 6022 18000 6024
rect 9324 6020 9330 6022
rect 9213 6019 9279 6020
rect 13813 6019 13879 6022
rect 6208 6016 6528 6017
rect 6208 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6528 6016
rect 6208 5951 6528 5952
rect 11472 6016 11792 6017
rect 11472 5952 11480 6016
rect 11544 5952 11560 6016
rect 11624 5952 11640 6016
rect 11704 5952 11720 6016
rect 11784 5952 11792 6016
rect 17520 5992 18000 6022
rect 11472 5951 11792 5952
rect 13813 5948 13879 5949
rect 13813 5944 13860 5948
rect 13924 5946 13930 5948
rect 13813 5888 13818 5944
rect 13813 5884 13860 5888
rect 13924 5886 13970 5946
rect 13924 5884 13930 5886
rect 13813 5883 13879 5884
rect 0 5674 480 5704
rect 4061 5674 4127 5677
rect 0 5672 4127 5674
rect 0 5616 4066 5672
rect 4122 5616 4127 5672
rect 0 5614 4127 5616
rect 0 5584 480 5614
rect 4061 5611 4127 5614
rect 16205 5674 16271 5677
rect 17520 5674 18000 5704
rect 16205 5672 18000 5674
rect 16205 5616 16210 5672
rect 16266 5616 18000 5672
rect 16205 5614 18000 5616
rect 16205 5611 16271 5614
rect 17520 5584 18000 5614
rect 5533 5538 5599 5541
rect 7925 5538 7991 5541
rect 5533 5536 7991 5538
rect 5533 5480 5538 5536
rect 5594 5480 7930 5536
rect 7986 5480 7991 5536
rect 5533 5478 7991 5480
rect 5533 5475 5599 5478
rect 7925 5475 7991 5478
rect 3576 5472 3896 5473
rect 3576 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3896 5472
rect 3576 5407 3896 5408
rect 8840 5472 9160 5473
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8840 5407 9160 5408
rect 14104 5472 14424 5473
rect 14104 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 14424 5472
rect 14104 5407 14424 5408
rect 0 5266 480 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 480 5206
rect 4061 5203 4127 5206
rect 12249 5266 12315 5269
rect 17520 5266 18000 5296
rect 12249 5264 18000 5266
rect 12249 5208 12254 5264
rect 12310 5208 18000 5264
rect 12249 5206 18000 5208
rect 12249 5203 12315 5206
rect 17520 5176 18000 5206
rect 3417 5130 3483 5133
rect 3969 5130 4035 5133
rect 3417 5128 4035 5130
rect 3417 5072 3422 5128
rect 3478 5072 3974 5128
rect 4030 5072 4035 5128
rect 3417 5070 4035 5072
rect 3417 5067 3483 5070
rect 3969 5067 4035 5070
rect 3325 4994 3391 4997
rect 6729 4996 6795 4997
rect 4654 4994 4660 4996
rect 3325 4992 4660 4994
rect 3325 4936 3330 4992
rect 3386 4936 4660 4992
rect 3325 4934 4660 4936
rect 3325 4931 3391 4934
rect 4654 4932 4660 4934
rect 4724 4932 4730 4996
rect 6678 4994 6684 4996
rect 6638 4934 6684 4994
rect 6748 4992 6795 4996
rect 6790 4936 6795 4992
rect 6678 4932 6684 4934
rect 6748 4932 6795 4936
rect 6729 4931 6795 4932
rect 6208 4928 6528 4929
rect 0 4858 480 4888
rect 6208 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6528 4928
rect 6208 4863 6528 4864
rect 11472 4928 11792 4929
rect 11472 4864 11480 4928
rect 11544 4864 11560 4928
rect 11624 4864 11640 4928
rect 11704 4864 11720 4928
rect 11784 4864 11792 4928
rect 11472 4863 11792 4864
rect 2865 4858 2931 4861
rect 0 4856 2931 4858
rect 0 4800 2870 4856
rect 2926 4800 2931 4856
rect 0 4798 2931 4800
rect 0 4768 480 4798
rect 2865 4795 2931 4798
rect 5574 4796 5580 4860
rect 5644 4858 5650 4860
rect 5993 4858 6059 4861
rect 5644 4856 6059 4858
rect 5644 4800 5998 4856
rect 6054 4800 6059 4856
rect 5644 4798 6059 4800
rect 5644 4796 5650 4798
rect 5993 4795 6059 4798
rect 16297 4858 16363 4861
rect 17520 4858 18000 4888
rect 16297 4856 18000 4858
rect 16297 4800 16302 4856
rect 16358 4800 18000 4856
rect 16297 4798 18000 4800
rect 16297 4795 16363 4798
rect 17520 4768 18000 4798
rect 4061 4586 4127 4589
rect 4245 4586 4311 4589
rect 8201 4586 8267 4589
rect 4061 4584 8267 4586
rect 4061 4528 4066 4584
rect 4122 4528 4250 4584
rect 4306 4528 8206 4584
rect 8262 4528 8267 4584
rect 4061 4526 8267 4528
rect 4061 4523 4127 4526
rect 4245 4523 4311 4526
rect 8201 4523 8267 4526
rect 0 4450 480 4480
rect 2773 4450 2839 4453
rect 0 4448 2839 4450
rect 0 4392 2778 4448
rect 2834 4392 2839 4448
rect 0 4390 2839 4392
rect 0 4360 480 4390
rect 2773 4387 2839 4390
rect 14917 4450 14983 4453
rect 17520 4450 18000 4480
rect 14917 4448 18000 4450
rect 14917 4392 14922 4448
rect 14978 4392 18000 4448
rect 14917 4390 18000 4392
rect 14917 4387 14983 4390
rect 3576 4384 3896 4385
rect 3576 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3896 4384
rect 3576 4319 3896 4320
rect 8840 4384 9160 4385
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8840 4319 9160 4320
rect 14104 4384 14424 4385
rect 14104 4320 14112 4384
rect 14176 4320 14192 4384
rect 14256 4320 14272 4384
rect 14336 4320 14352 4384
rect 14416 4320 14424 4384
rect 17520 4360 18000 4390
rect 14104 4319 14424 4320
rect 0 4042 480 4072
rect 3509 4042 3575 4045
rect 0 4040 3575 4042
rect 0 3984 3514 4040
rect 3570 3984 3575 4040
rect 0 3982 3575 3984
rect 0 3952 480 3982
rect 3509 3979 3575 3982
rect 5901 4042 5967 4045
rect 7833 4042 7899 4045
rect 5901 4040 7899 4042
rect 5901 3984 5906 4040
rect 5962 3984 7838 4040
rect 7894 3984 7899 4040
rect 5901 3982 7899 3984
rect 5901 3979 5967 3982
rect 7833 3979 7899 3982
rect 13445 4042 13511 4045
rect 17520 4042 18000 4072
rect 13445 4040 18000 4042
rect 13445 3984 13450 4040
rect 13506 3984 18000 4040
rect 13445 3982 18000 3984
rect 13445 3979 13511 3982
rect 17520 3952 18000 3982
rect 5257 3906 5323 3909
rect 5214 3904 5323 3906
rect 5214 3848 5262 3904
rect 5318 3848 5323 3904
rect 5214 3843 5323 3848
rect 0 3634 480 3664
rect 1761 3634 1827 3637
rect 0 3632 1827 3634
rect 0 3576 1766 3632
rect 1822 3576 1827 3632
rect 0 3574 1827 3576
rect 0 3544 480 3574
rect 1761 3571 1827 3574
rect 3049 3634 3115 3637
rect 5214 3634 5274 3843
rect 6208 3840 6528 3841
rect 6208 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6528 3840
rect 6208 3775 6528 3776
rect 11472 3840 11792 3841
rect 11472 3776 11480 3840
rect 11544 3776 11560 3840
rect 11624 3776 11640 3840
rect 11704 3776 11720 3840
rect 11784 3776 11792 3840
rect 11472 3775 11792 3776
rect 7097 3634 7163 3637
rect 3049 3632 7163 3634
rect 3049 3576 3054 3632
rect 3110 3576 7102 3632
rect 7158 3576 7163 3632
rect 3049 3574 7163 3576
rect 3049 3571 3115 3574
rect 7097 3571 7163 3574
rect 14641 3634 14707 3637
rect 17520 3634 18000 3664
rect 14641 3632 18000 3634
rect 14641 3576 14646 3632
rect 14702 3576 18000 3632
rect 14641 3574 18000 3576
rect 14641 3571 14707 3574
rect 17520 3544 18000 3574
rect 5349 3498 5415 3501
rect 8937 3498 9003 3501
rect 5349 3496 9003 3498
rect 5349 3440 5354 3496
rect 5410 3440 8942 3496
rect 8998 3440 9003 3496
rect 5349 3438 9003 3440
rect 5349 3435 5415 3438
rect 8937 3435 9003 3438
rect 15101 3498 15167 3501
rect 15101 3496 15210 3498
rect 15101 3440 15106 3496
rect 15162 3440 15210 3496
rect 15101 3435 15210 3440
rect 3576 3296 3896 3297
rect 3576 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3896 3296
rect 3576 3231 3896 3232
rect 8840 3296 9160 3297
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 8840 3231 9160 3232
rect 14104 3296 14424 3297
rect 14104 3232 14112 3296
rect 14176 3232 14192 3296
rect 14256 3232 14272 3296
rect 14336 3232 14352 3296
rect 14416 3232 14424 3296
rect 14104 3231 14424 3232
rect 0 3090 480 3120
rect 3969 3090 4035 3093
rect 0 3088 4035 3090
rect 0 3032 3974 3088
rect 4030 3032 4035 3088
rect 0 3030 4035 3032
rect 0 3000 480 3030
rect 3969 3027 4035 3030
rect 8109 3090 8175 3093
rect 8937 3090 9003 3093
rect 8109 3088 9003 3090
rect 8109 3032 8114 3088
rect 8170 3032 8942 3088
rect 8998 3032 9003 3088
rect 8109 3030 9003 3032
rect 15150 3090 15210 3435
rect 17520 3090 18000 3120
rect 15150 3030 18000 3090
rect 8109 3027 8175 3030
rect 8937 3027 9003 3030
rect 17520 3000 18000 3030
rect 9029 2954 9095 2957
rect 9438 2954 9444 2956
rect 9029 2952 9444 2954
rect 9029 2896 9034 2952
rect 9090 2896 9444 2952
rect 9029 2894 9444 2896
rect 9029 2891 9095 2894
rect 9438 2892 9444 2894
rect 9508 2892 9514 2956
rect 8702 2756 8708 2820
rect 8772 2818 8778 2820
rect 9121 2818 9187 2821
rect 8772 2816 9187 2818
rect 8772 2760 9126 2816
rect 9182 2760 9187 2816
rect 8772 2758 9187 2760
rect 8772 2756 8778 2758
rect 9121 2755 9187 2758
rect 6208 2752 6528 2753
rect 0 2682 480 2712
rect 6208 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6528 2752
rect 6208 2687 6528 2688
rect 11472 2752 11792 2753
rect 11472 2688 11480 2752
rect 11544 2688 11560 2752
rect 11624 2688 11640 2752
rect 11704 2688 11720 2752
rect 11784 2688 11792 2752
rect 11472 2687 11792 2688
rect 3693 2682 3759 2685
rect 7373 2684 7439 2685
rect 7373 2682 7420 2684
rect 0 2680 3759 2682
rect 0 2624 3698 2680
rect 3754 2624 3759 2680
rect 0 2622 3759 2624
rect 7328 2680 7420 2682
rect 7328 2624 7378 2680
rect 7328 2622 7420 2624
rect 0 2592 480 2622
rect 3693 2619 3759 2622
rect 7373 2620 7420 2622
rect 7484 2620 7490 2684
rect 11973 2682 12039 2685
rect 17520 2682 18000 2712
rect 11973 2680 18000 2682
rect 11973 2624 11978 2680
rect 12034 2624 18000 2680
rect 11973 2622 18000 2624
rect 7373 2619 7439 2620
rect 11973 2619 12039 2622
rect 17520 2592 18000 2622
rect 4153 2546 4219 2549
rect 6913 2546 6979 2549
rect 4153 2544 6979 2546
rect 4153 2488 4158 2544
rect 4214 2488 6918 2544
rect 6974 2488 6979 2544
rect 4153 2486 6979 2488
rect 4153 2483 4219 2486
rect 6913 2483 6979 2486
rect 0 2274 480 2304
rect 3417 2274 3483 2277
rect 0 2272 3483 2274
rect 0 2216 3422 2272
rect 3478 2216 3483 2272
rect 0 2214 3483 2216
rect 0 2184 480 2214
rect 3417 2211 3483 2214
rect 16113 2274 16179 2277
rect 17520 2274 18000 2304
rect 16113 2272 18000 2274
rect 16113 2216 16118 2272
rect 16174 2216 18000 2272
rect 16113 2214 18000 2216
rect 16113 2211 16179 2214
rect 3576 2208 3896 2209
rect 3576 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3896 2208
rect 3576 2143 3896 2144
rect 8840 2208 9160 2209
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8840 2143 9160 2144
rect 14104 2208 14424 2209
rect 14104 2144 14112 2208
rect 14176 2144 14192 2208
rect 14256 2144 14272 2208
rect 14336 2144 14352 2208
rect 14416 2144 14424 2208
rect 17520 2184 18000 2214
rect 14104 2143 14424 2144
rect 0 1866 480 1896
rect 2957 1866 3023 1869
rect 0 1864 3023 1866
rect 0 1808 2962 1864
rect 3018 1808 3023 1864
rect 0 1806 3023 1808
rect 0 1776 480 1806
rect 2957 1803 3023 1806
rect 13813 1866 13879 1869
rect 17520 1866 18000 1896
rect 13813 1864 18000 1866
rect 13813 1808 13818 1864
rect 13874 1808 18000 1864
rect 13813 1806 18000 1808
rect 13813 1803 13879 1806
rect 17520 1776 18000 1806
rect 0 1458 480 1488
rect 749 1458 815 1461
rect 0 1456 815 1458
rect 0 1400 754 1456
rect 810 1400 815 1456
rect 0 1398 815 1400
rect 0 1368 480 1398
rect 749 1395 815 1398
rect 14917 1458 14983 1461
rect 17520 1458 18000 1488
rect 14917 1456 18000 1458
rect 14917 1400 14922 1456
rect 14978 1400 18000 1456
rect 14917 1398 18000 1400
rect 14917 1395 14983 1398
rect 17520 1368 18000 1398
rect 0 1050 480 1080
rect 3693 1050 3759 1053
rect 0 1048 3759 1050
rect 0 992 3698 1048
rect 3754 992 3759 1048
rect 0 990 3759 992
rect 0 960 480 990
rect 3693 987 3759 990
rect 14825 1050 14891 1053
rect 17520 1050 18000 1080
rect 14825 1048 18000 1050
rect 14825 992 14830 1048
rect 14886 992 18000 1048
rect 14825 990 18000 992
rect 14825 987 14891 990
rect 17520 960 18000 990
rect 0 642 480 672
rect 2865 642 2931 645
rect 0 640 2931 642
rect 0 584 2870 640
rect 2926 584 2931 640
rect 0 582 2931 584
rect 0 552 480 582
rect 2865 579 2931 582
rect 15101 642 15167 645
rect 17520 642 18000 672
rect 15101 640 18000 642
rect 15101 584 15106 640
rect 15162 584 18000 640
rect 15101 582 18000 584
rect 15101 579 15167 582
rect 17520 552 18000 582
rect 0 234 480 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 480 174
rect 2773 171 2839 174
rect 15009 234 15075 237
rect 17520 234 18000 264
rect 15009 232 18000 234
rect 15009 176 15014 232
rect 15070 176 18000 232
rect 15009 174 18000 176
rect 15009 171 15075 174
rect 17520 144 18000 174
<< via3 >>
rect 6216 14716 6280 14720
rect 6216 14660 6220 14716
rect 6220 14660 6276 14716
rect 6276 14660 6280 14716
rect 6216 14656 6280 14660
rect 6296 14716 6360 14720
rect 6296 14660 6300 14716
rect 6300 14660 6356 14716
rect 6356 14660 6360 14716
rect 6296 14656 6360 14660
rect 6376 14716 6440 14720
rect 6376 14660 6380 14716
rect 6380 14660 6436 14716
rect 6436 14660 6440 14716
rect 6376 14656 6440 14660
rect 6456 14716 6520 14720
rect 6456 14660 6460 14716
rect 6460 14660 6516 14716
rect 6516 14660 6520 14716
rect 6456 14656 6520 14660
rect 11480 14716 11544 14720
rect 11480 14660 11484 14716
rect 11484 14660 11540 14716
rect 11540 14660 11544 14716
rect 11480 14656 11544 14660
rect 11560 14716 11624 14720
rect 11560 14660 11564 14716
rect 11564 14660 11620 14716
rect 11620 14660 11624 14716
rect 11560 14656 11624 14660
rect 11640 14716 11704 14720
rect 11640 14660 11644 14716
rect 11644 14660 11700 14716
rect 11700 14660 11704 14716
rect 11640 14656 11704 14660
rect 11720 14716 11784 14720
rect 11720 14660 11724 14716
rect 11724 14660 11780 14716
rect 11780 14660 11784 14716
rect 11720 14656 11784 14660
rect 3584 14172 3648 14176
rect 3584 14116 3588 14172
rect 3588 14116 3644 14172
rect 3644 14116 3648 14172
rect 3584 14112 3648 14116
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 8848 14172 8912 14176
rect 8848 14116 8852 14172
rect 8852 14116 8908 14172
rect 8908 14116 8912 14172
rect 8848 14112 8912 14116
rect 8928 14172 8992 14176
rect 8928 14116 8932 14172
rect 8932 14116 8988 14172
rect 8988 14116 8992 14172
rect 8928 14112 8992 14116
rect 9008 14172 9072 14176
rect 9008 14116 9012 14172
rect 9012 14116 9068 14172
rect 9068 14116 9072 14172
rect 9008 14112 9072 14116
rect 9088 14172 9152 14176
rect 9088 14116 9092 14172
rect 9092 14116 9148 14172
rect 9148 14116 9152 14172
rect 9088 14112 9152 14116
rect 14112 14172 14176 14176
rect 14112 14116 14116 14172
rect 14116 14116 14172 14172
rect 14172 14116 14176 14172
rect 14112 14112 14176 14116
rect 14192 14172 14256 14176
rect 14192 14116 14196 14172
rect 14196 14116 14252 14172
rect 14252 14116 14256 14172
rect 14192 14112 14256 14116
rect 14272 14172 14336 14176
rect 14272 14116 14276 14172
rect 14276 14116 14332 14172
rect 14332 14116 14336 14172
rect 14272 14112 14336 14116
rect 14352 14172 14416 14176
rect 14352 14116 14356 14172
rect 14356 14116 14412 14172
rect 14412 14116 14416 14172
rect 14352 14112 14416 14116
rect 4660 13636 4724 13700
rect 6216 13628 6280 13632
rect 6216 13572 6220 13628
rect 6220 13572 6276 13628
rect 6276 13572 6280 13628
rect 6216 13568 6280 13572
rect 6296 13628 6360 13632
rect 6296 13572 6300 13628
rect 6300 13572 6356 13628
rect 6356 13572 6360 13628
rect 6296 13568 6360 13572
rect 6376 13628 6440 13632
rect 6376 13572 6380 13628
rect 6380 13572 6436 13628
rect 6436 13572 6440 13628
rect 6376 13568 6440 13572
rect 6456 13628 6520 13632
rect 6456 13572 6460 13628
rect 6460 13572 6516 13628
rect 6516 13572 6520 13628
rect 6456 13568 6520 13572
rect 11480 13628 11544 13632
rect 11480 13572 11484 13628
rect 11484 13572 11540 13628
rect 11540 13572 11544 13628
rect 11480 13568 11544 13572
rect 11560 13628 11624 13632
rect 11560 13572 11564 13628
rect 11564 13572 11620 13628
rect 11620 13572 11624 13628
rect 11560 13568 11624 13572
rect 11640 13628 11704 13632
rect 11640 13572 11644 13628
rect 11644 13572 11700 13628
rect 11700 13572 11704 13628
rect 11640 13568 11704 13572
rect 11720 13628 11784 13632
rect 11720 13572 11724 13628
rect 11724 13572 11780 13628
rect 11780 13572 11784 13628
rect 11720 13568 11784 13572
rect 3584 13084 3648 13088
rect 3584 13028 3588 13084
rect 3588 13028 3644 13084
rect 3644 13028 3648 13084
rect 3584 13024 3648 13028
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 8848 13084 8912 13088
rect 8848 13028 8852 13084
rect 8852 13028 8908 13084
rect 8908 13028 8912 13084
rect 8848 13024 8912 13028
rect 8928 13084 8992 13088
rect 8928 13028 8932 13084
rect 8932 13028 8988 13084
rect 8988 13028 8992 13084
rect 8928 13024 8992 13028
rect 9008 13084 9072 13088
rect 9008 13028 9012 13084
rect 9012 13028 9068 13084
rect 9068 13028 9072 13084
rect 9008 13024 9072 13028
rect 9088 13084 9152 13088
rect 9088 13028 9092 13084
rect 9092 13028 9148 13084
rect 9148 13028 9152 13084
rect 9088 13024 9152 13028
rect 14112 13084 14176 13088
rect 14112 13028 14116 13084
rect 14116 13028 14172 13084
rect 14172 13028 14176 13084
rect 14112 13024 14176 13028
rect 14192 13084 14256 13088
rect 14192 13028 14196 13084
rect 14196 13028 14252 13084
rect 14252 13028 14256 13084
rect 14192 13024 14256 13028
rect 14272 13084 14336 13088
rect 14272 13028 14276 13084
rect 14276 13028 14332 13084
rect 14332 13028 14336 13084
rect 14272 13024 14336 13028
rect 14352 13084 14416 13088
rect 14352 13028 14356 13084
rect 14356 13028 14412 13084
rect 14412 13028 14416 13084
rect 14352 13024 14416 13028
rect 7420 12820 7484 12884
rect 6216 12540 6280 12544
rect 6216 12484 6220 12540
rect 6220 12484 6276 12540
rect 6276 12484 6280 12540
rect 6216 12480 6280 12484
rect 6296 12540 6360 12544
rect 6296 12484 6300 12540
rect 6300 12484 6356 12540
rect 6356 12484 6360 12540
rect 6296 12480 6360 12484
rect 6376 12540 6440 12544
rect 6376 12484 6380 12540
rect 6380 12484 6436 12540
rect 6436 12484 6440 12540
rect 6376 12480 6440 12484
rect 6456 12540 6520 12544
rect 6456 12484 6460 12540
rect 6460 12484 6516 12540
rect 6516 12484 6520 12540
rect 6456 12480 6520 12484
rect 11480 12540 11544 12544
rect 11480 12484 11484 12540
rect 11484 12484 11540 12540
rect 11540 12484 11544 12540
rect 11480 12480 11544 12484
rect 11560 12540 11624 12544
rect 11560 12484 11564 12540
rect 11564 12484 11620 12540
rect 11620 12484 11624 12540
rect 11560 12480 11624 12484
rect 11640 12540 11704 12544
rect 11640 12484 11644 12540
rect 11644 12484 11700 12540
rect 11700 12484 11704 12540
rect 11640 12480 11704 12484
rect 11720 12540 11784 12544
rect 11720 12484 11724 12540
rect 11724 12484 11780 12540
rect 11780 12484 11784 12540
rect 11720 12480 11784 12484
rect 3584 11996 3648 12000
rect 3584 11940 3588 11996
rect 3588 11940 3644 11996
rect 3644 11940 3648 11996
rect 3584 11936 3648 11940
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 8848 11996 8912 12000
rect 8848 11940 8852 11996
rect 8852 11940 8908 11996
rect 8908 11940 8912 11996
rect 8848 11936 8912 11940
rect 8928 11996 8992 12000
rect 8928 11940 8932 11996
rect 8932 11940 8988 11996
rect 8988 11940 8992 11996
rect 8928 11936 8992 11940
rect 9008 11996 9072 12000
rect 9008 11940 9012 11996
rect 9012 11940 9068 11996
rect 9068 11940 9072 11996
rect 9008 11936 9072 11940
rect 9088 11996 9152 12000
rect 9088 11940 9092 11996
rect 9092 11940 9148 11996
rect 9148 11940 9152 11996
rect 9088 11936 9152 11940
rect 14112 11996 14176 12000
rect 14112 11940 14116 11996
rect 14116 11940 14172 11996
rect 14172 11940 14176 11996
rect 14112 11936 14176 11940
rect 14192 11996 14256 12000
rect 14192 11940 14196 11996
rect 14196 11940 14252 11996
rect 14252 11940 14256 11996
rect 14192 11936 14256 11940
rect 14272 11996 14336 12000
rect 14272 11940 14276 11996
rect 14276 11940 14332 11996
rect 14332 11940 14336 11996
rect 14272 11936 14336 11940
rect 14352 11996 14416 12000
rect 14352 11940 14356 11996
rect 14356 11940 14412 11996
rect 14412 11940 14416 11996
rect 14352 11936 14416 11940
rect 6216 11452 6280 11456
rect 6216 11396 6220 11452
rect 6220 11396 6276 11452
rect 6276 11396 6280 11452
rect 6216 11392 6280 11396
rect 6296 11452 6360 11456
rect 6296 11396 6300 11452
rect 6300 11396 6356 11452
rect 6356 11396 6360 11452
rect 6296 11392 6360 11396
rect 6376 11452 6440 11456
rect 6376 11396 6380 11452
rect 6380 11396 6436 11452
rect 6436 11396 6440 11452
rect 6376 11392 6440 11396
rect 6456 11452 6520 11456
rect 6456 11396 6460 11452
rect 6460 11396 6516 11452
rect 6516 11396 6520 11452
rect 6456 11392 6520 11396
rect 11480 11452 11544 11456
rect 11480 11396 11484 11452
rect 11484 11396 11540 11452
rect 11540 11396 11544 11452
rect 11480 11392 11544 11396
rect 11560 11452 11624 11456
rect 11560 11396 11564 11452
rect 11564 11396 11620 11452
rect 11620 11396 11624 11452
rect 11560 11392 11624 11396
rect 11640 11452 11704 11456
rect 11640 11396 11644 11452
rect 11644 11396 11700 11452
rect 11700 11396 11704 11452
rect 11640 11392 11704 11396
rect 11720 11452 11784 11456
rect 11720 11396 11724 11452
rect 11724 11396 11780 11452
rect 11780 11396 11784 11452
rect 11720 11392 11784 11396
rect 3584 10908 3648 10912
rect 3584 10852 3588 10908
rect 3588 10852 3644 10908
rect 3644 10852 3648 10908
rect 3584 10848 3648 10852
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 8848 10908 8912 10912
rect 8848 10852 8852 10908
rect 8852 10852 8908 10908
rect 8908 10852 8912 10908
rect 8848 10848 8912 10852
rect 8928 10908 8992 10912
rect 8928 10852 8932 10908
rect 8932 10852 8988 10908
rect 8988 10852 8992 10908
rect 8928 10848 8992 10852
rect 9008 10908 9072 10912
rect 9008 10852 9012 10908
rect 9012 10852 9068 10908
rect 9068 10852 9072 10908
rect 9008 10848 9072 10852
rect 9088 10908 9152 10912
rect 9088 10852 9092 10908
rect 9092 10852 9148 10908
rect 9148 10852 9152 10908
rect 9088 10848 9152 10852
rect 14112 10908 14176 10912
rect 14112 10852 14116 10908
rect 14116 10852 14172 10908
rect 14172 10852 14176 10908
rect 14112 10848 14176 10852
rect 14192 10908 14256 10912
rect 14192 10852 14196 10908
rect 14196 10852 14252 10908
rect 14252 10852 14256 10908
rect 14192 10848 14256 10852
rect 14272 10908 14336 10912
rect 14272 10852 14276 10908
rect 14276 10852 14332 10908
rect 14332 10852 14336 10908
rect 14272 10848 14336 10852
rect 14352 10908 14416 10912
rect 14352 10852 14356 10908
rect 14356 10852 14412 10908
rect 14412 10852 14416 10908
rect 14352 10848 14416 10852
rect 9260 10372 9324 10436
rect 14596 10372 14660 10436
rect 6216 10364 6280 10368
rect 6216 10308 6220 10364
rect 6220 10308 6276 10364
rect 6276 10308 6280 10364
rect 6216 10304 6280 10308
rect 6296 10364 6360 10368
rect 6296 10308 6300 10364
rect 6300 10308 6356 10364
rect 6356 10308 6360 10364
rect 6296 10304 6360 10308
rect 6376 10364 6440 10368
rect 6376 10308 6380 10364
rect 6380 10308 6436 10364
rect 6436 10308 6440 10364
rect 6376 10304 6440 10308
rect 6456 10364 6520 10368
rect 6456 10308 6460 10364
rect 6460 10308 6516 10364
rect 6516 10308 6520 10364
rect 6456 10304 6520 10308
rect 11480 10364 11544 10368
rect 11480 10308 11484 10364
rect 11484 10308 11540 10364
rect 11540 10308 11544 10364
rect 11480 10304 11544 10308
rect 11560 10364 11624 10368
rect 11560 10308 11564 10364
rect 11564 10308 11620 10364
rect 11620 10308 11624 10364
rect 11560 10304 11624 10308
rect 11640 10364 11704 10368
rect 11640 10308 11644 10364
rect 11644 10308 11700 10364
rect 11700 10308 11704 10364
rect 11640 10304 11704 10308
rect 11720 10364 11784 10368
rect 11720 10308 11724 10364
rect 11724 10308 11780 10364
rect 11780 10308 11784 10364
rect 11720 10304 11784 10308
rect 3188 10296 3252 10300
rect 3188 10240 3238 10296
rect 3238 10240 3252 10296
rect 3188 10236 3252 10240
rect 2820 9964 2884 10028
rect 3584 9820 3648 9824
rect 3584 9764 3588 9820
rect 3588 9764 3644 9820
rect 3644 9764 3648 9820
rect 3584 9760 3648 9764
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 2820 9692 2884 9756
rect 8848 9820 8912 9824
rect 8848 9764 8852 9820
rect 8852 9764 8908 9820
rect 8908 9764 8912 9820
rect 8848 9760 8912 9764
rect 8928 9820 8992 9824
rect 8928 9764 8932 9820
rect 8932 9764 8988 9820
rect 8988 9764 8992 9820
rect 8928 9760 8992 9764
rect 9008 9820 9072 9824
rect 9008 9764 9012 9820
rect 9012 9764 9068 9820
rect 9068 9764 9072 9820
rect 9008 9760 9072 9764
rect 9088 9820 9152 9824
rect 9088 9764 9092 9820
rect 9092 9764 9148 9820
rect 9148 9764 9152 9820
rect 9088 9760 9152 9764
rect 14112 9820 14176 9824
rect 14112 9764 14116 9820
rect 14116 9764 14172 9820
rect 14172 9764 14176 9820
rect 14112 9760 14176 9764
rect 14192 9820 14256 9824
rect 14192 9764 14196 9820
rect 14196 9764 14252 9820
rect 14252 9764 14256 9820
rect 14192 9760 14256 9764
rect 14272 9820 14336 9824
rect 14272 9764 14276 9820
rect 14276 9764 14332 9820
rect 14332 9764 14336 9820
rect 14272 9760 14336 9764
rect 14352 9820 14416 9824
rect 14352 9764 14356 9820
rect 14356 9764 14412 9820
rect 14412 9764 14416 9820
rect 14352 9760 14416 9764
rect 9444 9556 9508 9620
rect 4108 9284 4172 9348
rect 5580 9284 5644 9348
rect 14596 9692 14660 9756
rect 13860 9556 13924 9620
rect 6216 9276 6280 9280
rect 6216 9220 6220 9276
rect 6220 9220 6276 9276
rect 6276 9220 6280 9276
rect 6216 9216 6280 9220
rect 6296 9276 6360 9280
rect 6296 9220 6300 9276
rect 6300 9220 6356 9276
rect 6356 9220 6360 9276
rect 6296 9216 6360 9220
rect 6376 9276 6440 9280
rect 6376 9220 6380 9276
rect 6380 9220 6436 9276
rect 6436 9220 6440 9276
rect 6376 9216 6440 9220
rect 6456 9276 6520 9280
rect 6456 9220 6460 9276
rect 6460 9220 6516 9276
rect 6516 9220 6520 9276
rect 6456 9216 6520 9220
rect 11480 9276 11544 9280
rect 11480 9220 11484 9276
rect 11484 9220 11540 9276
rect 11540 9220 11544 9276
rect 11480 9216 11544 9220
rect 11560 9276 11624 9280
rect 11560 9220 11564 9276
rect 11564 9220 11620 9276
rect 11620 9220 11624 9276
rect 11560 9216 11624 9220
rect 11640 9276 11704 9280
rect 11640 9220 11644 9276
rect 11644 9220 11700 9276
rect 11700 9220 11704 9276
rect 11640 9216 11704 9220
rect 11720 9276 11784 9280
rect 11720 9220 11724 9276
rect 11724 9220 11780 9276
rect 11780 9220 11784 9276
rect 11720 9216 11784 9220
rect 3584 8732 3648 8736
rect 3584 8676 3588 8732
rect 3588 8676 3644 8732
rect 3644 8676 3648 8732
rect 3584 8672 3648 8676
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 8848 8732 8912 8736
rect 8848 8676 8852 8732
rect 8852 8676 8908 8732
rect 8908 8676 8912 8732
rect 8848 8672 8912 8676
rect 8928 8732 8992 8736
rect 8928 8676 8932 8732
rect 8932 8676 8988 8732
rect 8988 8676 8992 8732
rect 8928 8672 8992 8676
rect 9008 8732 9072 8736
rect 9008 8676 9012 8732
rect 9012 8676 9068 8732
rect 9068 8676 9072 8732
rect 9008 8672 9072 8676
rect 9088 8732 9152 8736
rect 9088 8676 9092 8732
rect 9092 8676 9148 8732
rect 9148 8676 9152 8732
rect 9088 8672 9152 8676
rect 14112 8732 14176 8736
rect 14112 8676 14116 8732
rect 14116 8676 14172 8732
rect 14172 8676 14176 8732
rect 14112 8672 14176 8676
rect 14192 8732 14256 8736
rect 14192 8676 14196 8732
rect 14196 8676 14252 8732
rect 14252 8676 14256 8732
rect 14192 8672 14256 8676
rect 14272 8732 14336 8736
rect 14272 8676 14276 8732
rect 14276 8676 14332 8732
rect 14332 8676 14336 8732
rect 14272 8672 14336 8676
rect 14352 8732 14416 8736
rect 14352 8676 14356 8732
rect 14356 8676 14412 8732
rect 14412 8676 14416 8732
rect 14352 8672 14416 8676
rect 13860 8468 13924 8532
rect 9444 8332 9508 8396
rect 6216 8188 6280 8192
rect 6216 8132 6220 8188
rect 6220 8132 6276 8188
rect 6276 8132 6280 8188
rect 6216 8128 6280 8132
rect 6296 8188 6360 8192
rect 6296 8132 6300 8188
rect 6300 8132 6356 8188
rect 6356 8132 6360 8188
rect 6296 8128 6360 8132
rect 6376 8188 6440 8192
rect 6376 8132 6380 8188
rect 6380 8132 6436 8188
rect 6436 8132 6440 8188
rect 6376 8128 6440 8132
rect 6456 8188 6520 8192
rect 6456 8132 6460 8188
rect 6460 8132 6516 8188
rect 6516 8132 6520 8188
rect 6456 8128 6520 8132
rect 11480 8188 11544 8192
rect 11480 8132 11484 8188
rect 11484 8132 11540 8188
rect 11540 8132 11544 8188
rect 11480 8128 11544 8132
rect 11560 8188 11624 8192
rect 11560 8132 11564 8188
rect 11564 8132 11620 8188
rect 11620 8132 11624 8188
rect 11560 8128 11624 8132
rect 11640 8188 11704 8192
rect 11640 8132 11644 8188
rect 11644 8132 11700 8188
rect 11700 8132 11704 8188
rect 11640 8128 11704 8132
rect 11720 8188 11784 8192
rect 11720 8132 11724 8188
rect 11724 8132 11780 8188
rect 11780 8132 11784 8188
rect 11720 8128 11784 8132
rect 8708 8060 8772 8124
rect 6684 7788 6748 7852
rect 3584 7644 3648 7648
rect 3584 7588 3588 7644
rect 3588 7588 3644 7644
rect 3644 7588 3648 7644
rect 3584 7584 3648 7588
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 8848 7644 8912 7648
rect 8848 7588 8852 7644
rect 8852 7588 8908 7644
rect 8908 7588 8912 7644
rect 8848 7584 8912 7588
rect 8928 7644 8992 7648
rect 8928 7588 8932 7644
rect 8932 7588 8988 7644
rect 8988 7588 8992 7644
rect 8928 7584 8992 7588
rect 9008 7644 9072 7648
rect 9008 7588 9012 7644
rect 9012 7588 9068 7644
rect 9068 7588 9072 7644
rect 9008 7584 9072 7588
rect 9088 7644 9152 7648
rect 9088 7588 9092 7644
rect 9092 7588 9148 7644
rect 9148 7588 9152 7644
rect 9088 7584 9152 7588
rect 14112 7644 14176 7648
rect 14112 7588 14116 7644
rect 14116 7588 14172 7644
rect 14172 7588 14176 7644
rect 14112 7584 14176 7588
rect 14192 7644 14256 7648
rect 14192 7588 14196 7644
rect 14196 7588 14252 7644
rect 14252 7588 14256 7644
rect 14192 7584 14256 7588
rect 14272 7644 14336 7648
rect 14272 7588 14276 7644
rect 14276 7588 14332 7644
rect 14332 7588 14336 7644
rect 14272 7584 14336 7588
rect 14352 7644 14416 7648
rect 14352 7588 14356 7644
rect 14356 7588 14412 7644
rect 14412 7588 14416 7644
rect 14352 7584 14416 7588
rect 5580 7108 5644 7172
rect 6216 7100 6280 7104
rect 6216 7044 6220 7100
rect 6220 7044 6276 7100
rect 6276 7044 6280 7100
rect 6216 7040 6280 7044
rect 6296 7100 6360 7104
rect 6296 7044 6300 7100
rect 6300 7044 6356 7100
rect 6356 7044 6360 7100
rect 6296 7040 6360 7044
rect 6376 7100 6440 7104
rect 6376 7044 6380 7100
rect 6380 7044 6436 7100
rect 6436 7044 6440 7100
rect 6376 7040 6440 7044
rect 6456 7100 6520 7104
rect 6456 7044 6460 7100
rect 6460 7044 6516 7100
rect 6516 7044 6520 7100
rect 6456 7040 6520 7044
rect 11480 7100 11544 7104
rect 11480 7044 11484 7100
rect 11484 7044 11540 7100
rect 11540 7044 11544 7100
rect 11480 7040 11544 7044
rect 11560 7100 11624 7104
rect 11560 7044 11564 7100
rect 11564 7044 11620 7100
rect 11620 7044 11624 7100
rect 11560 7040 11624 7044
rect 11640 7100 11704 7104
rect 11640 7044 11644 7100
rect 11644 7044 11700 7100
rect 11700 7044 11704 7100
rect 11640 7040 11704 7044
rect 11720 7100 11784 7104
rect 11720 7044 11724 7100
rect 11724 7044 11780 7100
rect 11780 7044 11784 7100
rect 11720 7040 11784 7044
rect 4108 6564 4172 6628
rect 3584 6556 3648 6560
rect 3584 6500 3588 6556
rect 3588 6500 3644 6556
rect 3644 6500 3648 6556
rect 3584 6496 3648 6500
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 8848 6556 8912 6560
rect 8848 6500 8852 6556
rect 8852 6500 8908 6556
rect 8908 6500 8912 6556
rect 8848 6496 8912 6500
rect 8928 6556 8992 6560
rect 8928 6500 8932 6556
rect 8932 6500 8988 6556
rect 8988 6500 8992 6556
rect 8928 6496 8992 6500
rect 9008 6556 9072 6560
rect 9008 6500 9012 6556
rect 9012 6500 9068 6556
rect 9068 6500 9072 6556
rect 9008 6496 9072 6500
rect 9088 6556 9152 6560
rect 9088 6500 9092 6556
rect 9092 6500 9148 6556
rect 9148 6500 9152 6556
rect 9088 6496 9152 6500
rect 14112 6556 14176 6560
rect 14112 6500 14116 6556
rect 14116 6500 14172 6556
rect 14172 6500 14176 6556
rect 14112 6496 14176 6500
rect 14192 6556 14256 6560
rect 14192 6500 14196 6556
rect 14196 6500 14252 6556
rect 14252 6500 14256 6556
rect 14192 6496 14256 6500
rect 14272 6556 14336 6560
rect 14272 6500 14276 6556
rect 14276 6500 14332 6556
rect 14332 6500 14336 6556
rect 14272 6496 14336 6500
rect 14352 6556 14416 6560
rect 14352 6500 14356 6556
rect 14356 6500 14412 6556
rect 14412 6500 14416 6556
rect 14352 6496 14416 6500
rect 3188 6352 3252 6356
rect 3188 6296 3202 6352
rect 3202 6296 3252 6352
rect 3188 6292 3252 6296
rect 9260 6080 9324 6084
rect 9260 6024 9274 6080
rect 9274 6024 9324 6080
rect 9260 6020 9324 6024
rect 6216 6012 6280 6016
rect 6216 5956 6220 6012
rect 6220 5956 6276 6012
rect 6276 5956 6280 6012
rect 6216 5952 6280 5956
rect 6296 6012 6360 6016
rect 6296 5956 6300 6012
rect 6300 5956 6356 6012
rect 6356 5956 6360 6012
rect 6296 5952 6360 5956
rect 6376 6012 6440 6016
rect 6376 5956 6380 6012
rect 6380 5956 6436 6012
rect 6436 5956 6440 6012
rect 6376 5952 6440 5956
rect 6456 6012 6520 6016
rect 6456 5956 6460 6012
rect 6460 5956 6516 6012
rect 6516 5956 6520 6012
rect 6456 5952 6520 5956
rect 11480 6012 11544 6016
rect 11480 5956 11484 6012
rect 11484 5956 11540 6012
rect 11540 5956 11544 6012
rect 11480 5952 11544 5956
rect 11560 6012 11624 6016
rect 11560 5956 11564 6012
rect 11564 5956 11620 6012
rect 11620 5956 11624 6012
rect 11560 5952 11624 5956
rect 11640 6012 11704 6016
rect 11640 5956 11644 6012
rect 11644 5956 11700 6012
rect 11700 5956 11704 6012
rect 11640 5952 11704 5956
rect 11720 6012 11784 6016
rect 11720 5956 11724 6012
rect 11724 5956 11780 6012
rect 11780 5956 11784 6012
rect 11720 5952 11784 5956
rect 13860 5944 13924 5948
rect 13860 5888 13874 5944
rect 13874 5888 13924 5944
rect 13860 5884 13924 5888
rect 3584 5468 3648 5472
rect 3584 5412 3588 5468
rect 3588 5412 3644 5468
rect 3644 5412 3648 5468
rect 3584 5408 3648 5412
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 8848 5468 8912 5472
rect 8848 5412 8852 5468
rect 8852 5412 8908 5468
rect 8908 5412 8912 5468
rect 8848 5408 8912 5412
rect 8928 5468 8992 5472
rect 8928 5412 8932 5468
rect 8932 5412 8988 5468
rect 8988 5412 8992 5468
rect 8928 5408 8992 5412
rect 9008 5468 9072 5472
rect 9008 5412 9012 5468
rect 9012 5412 9068 5468
rect 9068 5412 9072 5468
rect 9008 5408 9072 5412
rect 9088 5468 9152 5472
rect 9088 5412 9092 5468
rect 9092 5412 9148 5468
rect 9148 5412 9152 5468
rect 9088 5408 9152 5412
rect 14112 5468 14176 5472
rect 14112 5412 14116 5468
rect 14116 5412 14172 5468
rect 14172 5412 14176 5468
rect 14112 5408 14176 5412
rect 14192 5468 14256 5472
rect 14192 5412 14196 5468
rect 14196 5412 14252 5468
rect 14252 5412 14256 5468
rect 14192 5408 14256 5412
rect 14272 5468 14336 5472
rect 14272 5412 14276 5468
rect 14276 5412 14332 5468
rect 14332 5412 14336 5468
rect 14272 5408 14336 5412
rect 14352 5468 14416 5472
rect 14352 5412 14356 5468
rect 14356 5412 14412 5468
rect 14412 5412 14416 5468
rect 14352 5408 14416 5412
rect 4660 4932 4724 4996
rect 6684 4992 6748 4996
rect 6684 4936 6734 4992
rect 6734 4936 6748 4992
rect 6684 4932 6748 4936
rect 6216 4924 6280 4928
rect 6216 4868 6220 4924
rect 6220 4868 6276 4924
rect 6276 4868 6280 4924
rect 6216 4864 6280 4868
rect 6296 4924 6360 4928
rect 6296 4868 6300 4924
rect 6300 4868 6356 4924
rect 6356 4868 6360 4924
rect 6296 4864 6360 4868
rect 6376 4924 6440 4928
rect 6376 4868 6380 4924
rect 6380 4868 6436 4924
rect 6436 4868 6440 4924
rect 6376 4864 6440 4868
rect 6456 4924 6520 4928
rect 6456 4868 6460 4924
rect 6460 4868 6516 4924
rect 6516 4868 6520 4924
rect 6456 4864 6520 4868
rect 11480 4924 11544 4928
rect 11480 4868 11484 4924
rect 11484 4868 11540 4924
rect 11540 4868 11544 4924
rect 11480 4864 11544 4868
rect 11560 4924 11624 4928
rect 11560 4868 11564 4924
rect 11564 4868 11620 4924
rect 11620 4868 11624 4924
rect 11560 4864 11624 4868
rect 11640 4924 11704 4928
rect 11640 4868 11644 4924
rect 11644 4868 11700 4924
rect 11700 4868 11704 4924
rect 11640 4864 11704 4868
rect 11720 4924 11784 4928
rect 11720 4868 11724 4924
rect 11724 4868 11780 4924
rect 11780 4868 11784 4924
rect 11720 4864 11784 4868
rect 5580 4796 5644 4860
rect 3584 4380 3648 4384
rect 3584 4324 3588 4380
rect 3588 4324 3644 4380
rect 3644 4324 3648 4380
rect 3584 4320 3648 4324
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 8848 4380 8912 4384
rect 8848 4324 8852 4380
rect 8852 4324 8908 4380
rect 8908 4324 8912 4380
rect 8848 4320 8912 4324
rect 8928 4380 8992 4384
rect 8928 4324 8932 4380
rect 8932 4324 8988 4380
rect 8988 4324 8992 4380
rect 8928 4320 8992 4324
rect 9008 4380 9072 4384
rect 9008 4324 9012 4380
rect 9012 4324 9068 4380
rect 9068 4324 9072 4380
rect 9008 4320 9072 4324
rect 9088 4380 9152 4384
rect 9088 4324 9092 4380
rect 9092 4324 9148 4380
rect 9148 4324 9152 4380
rect 9088 4320 9152 4324
rect 14112 4380 14176 4384
rect 14112 4324 14116 4380
rect 14116 4324 14172 4380
rect 14172 4324 14176 4380
rect 14112 4320 14176 4324
rect 14192 4380 14256 4384
rect 14192 4324 14196 4380
rect 14196 4324 14252 4380
rect 14252 4324 14256 4380
rect 14192 4320 14256 4324
rect 14272 4380 14336 4384
rect 14272 4324 14276 4380
rect 14276 4324 14332 4380
rect 14332 4324 14336 4380
rect 14272 4320 14336 4324
rect 14352 4380 14416 4384
rect 14352 4324 14356 4380
rect 14356 4324 14412 4380
rect 14412 4324 14416 4380
rect 14352 4320 14416 4324
rect 6216 3836 6280 3840
rect 6216 3780 6220 3836
rect 6220 3780 6276 3836
rect 6276 3780 6280 3836
rect 6216 3776 6280 3780
rect 6296 3836 6360 3840
rect 6296 3780 6300 3836
rect 6300 3780 6356 3836
rect 6356 3780 6360 3836
rect 6296 3776 6360 3780
rect 6376 3836 6440 3840
rect 6376 3780 6380 3836
rect 6380 3780 6436 3836
rect 6436 3780 6440 3836
rect 6376 3776 6440 3780
rect 6456 3836 6520 3840
rect 6456 3780 6460 3836
rect 6460 3780 6516 3836
rect 6516 3780 6520 3836
rect 6456 3776 6520 3780
rect 11480 3836 11544 3840
rect 11480 3780 11484 3836
rect 11484 3780 11540 3836
rect 11540 3780 11544 3836
rect 11480 3776 11544 3780
rect 11560 3836 11624 3840
rect 11560 3780 11564 3836
rect 11564 3780 11620 3836
rect 11620 3780 11624 3836
rect 11560 3776 11624 3780
rect 11640 3836 11704 3840
rect 11640 3780 11644 3836
rect 11644 3780 11700 3836
rect 11700 3780 11704 3836
rect 11640 3776 11704 3780
rect 11720 3836 11784 3840
rect 11720 3780 11724 3836
rect 11724 3780 11780 3836
rect 11780 3780 11784 3836
rect 11720 3776 11784 3780
rect 3584 3292 3648 3296
rect 3584 3236 3588 3292
rect 3588 3236 3644 3292
rect 3644 3236 3648 3292
rect 3584 3232 3648 3236
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 8848 3292 8912 3296
rect 8848 3236 8852 3292
rect 8852 3236 8908 3292
rect 8908 3236 8912 3292
rect 8848 3232 8912 3236
rect 8928 3292 8992 3296
rect 8928 3236 8932 3292
rect 8932 3236 8988 3292
rect 8988 3236 8992 3292
rect 8928 3232 8992 3236
rect 9008 3292 9072 3296
rect 9008 3236 9012 3292
rect 9012 3236 9068 3292
rect 9068 3236 9072 3292
rect 9008 3232 9072 3236
rect 9088 3292 9152 3296
rect 9088 3236 9092 3292
rect 9092 3236 9148 3292
rect 9148 3236 9152 3292
rect 9088 3232 9152 3236
rect 14112 3292 14176 3296
rect 14112 3236 14116 3292
rect 14116 3236 14172 3292
rect 14172 3236 14176 3292
rect 14112 3232 14176 3236
rect 14192 3292 14256 3296
rect 14192 3236 14196 3292
rect 14196 3236 14252 3292
rect 14252 3236 14256 3292
rect 14192 3232 14256 3236
rect 14272 3292 14336 3296
rect 14272 3236 14276 3292
rect 14276 3236 14332 3292
rect 14332 3236 14336 3292
rect 14272 3232 14336 3236
rect 14352 3292 14416 3296
rect 14352 3236 14356 3292
rect 14356 3236 14412 3292
rect 14412 3236 14416 3292
rect 14352 3232 14416 3236
rect 9444 2892 9508 2956
rect 8708 2756 8772 2820
rect 6216 2748 6280 2752
rect 6216 2692 6220 2748
rect 6220 2692 6276 2748
rect 6276 2692 6280 2748
rect 6216 2688 6280 2692
rect 6296 2748 6360 2752
rect 6296 2692 6300 2748
rect 6300 2692 6356 2748
rect 6356 2692 6360 2748
rect 6296 2688 6360 2692
rect 6376 2748 6440 2752
rect 6376 2692 6380 2748
rect 6380 2692 6436 2748
rect 6436 2692 6440 2748
rect 6376 2688 6440 2692
rect 6456 2748 6520 2752
rect 6456 2692 6460 2748
rect 6460 2692 6516 2748
rect 6516 2692 6520 2748
rect 6456 2688 6520 2692
rect 11480 2748 11544 2752
rect 11480 2692 11484 2748
rect 11484 2692 11540 2748
rect 11540 2692 11544 2748
rect 11480 2688 11544 2692
rect 11560 2748 11624 2752
rect 11560 2692 11564 2748
rect 11564 2692 11620 2748
rect 11620 2692 11624 2748
rect 11560 2688 11624 2692
rect 11640 2748 11704 2752
rect 11640 2692 11644 2748
rect 11644 2692 11700 2748
rect 11700 2692 11704 2748
rect 11640 2688 11704 2692
rect 11720 2748 11784 2752
rect 11720 2692 11724 2748
rect 11724 2692 11780 2748
rect 11780 2692 11784 2748
rect 11720 2688 11784 2692
rect 7420 2680 7484 2684
rect 7420 2624 7434 2680
rect 7434 2624 7484 2680
rect 7420 2620 7484 2624
rect 3584 2204 3648 2208
rect 3584 2148 3588 2204
rect 3588 2148 3644 2204
rect 3644 2148 3648 2204
rect 3584 2144 3648 2148
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 8848 2204 8912 2208
rect 8848 2148 8852 2204
rect 8852 2148 8908 2204
rect 8908 2148 8912 2204
rect 8848 2144 8912 2148
rect 8928 2204 8992 2208
rect 8928 2148 8932 2204
rect 8932 2148 8988 2204
rect 8988 2148 8992 2204
rect 8928 2144 8992 2148
rect 9008 2204 9072 2208
rect 9008 2148 9012 2204
rect 9012 2148 9068 2204
rect 9068 2148 9072 2204
rect 9008 2144 9072 2148
rect 9088 2204 9152 2208
rect 9088 2148 9092 2204
rect 9092 2148 9148 2204
rect 9148 2148 9152 2204
rect 9088 2144 9152 2148
rect 14112 2204 14176 2208
rect 14112 2148 14116 2204
rect 14116 2148 14172 2204
rect 14172 2148 14176 2204
rect 14112 2144 14176 2148
rect 14192 2204 14256 2208
rect 14192 2148 14196 2204
rect 14196 2148 14252 2204
rect 14252 2148 14256 2204
rect 14192 2144 14256 2148
rect 14272 2204 14336 2208
rect 14272 2148 14276 2204
rect 14276 2148 14332 2204
rect 14332 2148 14336 2204
rect 14272 2144 14336 2148
rect 14352 2204 14416 2208
rect 14352 2148 14356 2204
rect 14356 2148 14412 2204
rect 14412 2148 14416 2204
rect 14352 2144 14416 2148
<< metal4 >>
rect 3576 14176 3896 14736
rect 3576 14112 3584 14176
rect 3648 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3896 14176
rect 3576 13088 3896 14112
rect 6208 14720 6528 14736
rect 6208 14656 6216 14720
rect 6280 14656 6296 14720
rect 6360 14656 6376 14720
rect 6440 14656 6456 14720
rect 6520 14656 6528 14720
rect 4659 13700 4725 13701
rect 4659 13636 4660 13700
rect 4724 13636 4725 13700
rect 4659 13635 4725 13636
rect 3576 13024 3584 13088
rect 3648 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3896 13088
rect 3576 12000 3896 13024
rect 3576 11936 3584 12000
rect 3648 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3896 12000
rect 3576 10912 3896 11936
rect 3576 10848 3584 10912
rect 3648 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3896 10912
rect 3187 10300 3253 10301
rect 3187 10236 3188 10300
rect 3252 10236 3253 10300
rect 3187 10235 3253 10236
rect 2819 10028 2885 10029
rect 2819 9964 2820 10028
rect 2884 9964 2885 10028
rect 2819 9963 2885 9964
rect 2822 9757 2882 9963
rect 2819 9756 2885 9757
rect 2819 9692 2820 9756
rect 2884 9692 2885 9756
rect 2819 9691 2885 9692
rect 3190 6357 3250 10235
rect 3576 9824 3896 10848
rect 3576 9760 3584 9824
rect 3648 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3896 9824
rect 3576 8736 3896 9760
rect 4107 9348 4173 9349
rect 4107 9284 4108 9348
rect 4172 9284 4173 9348
rect 4107 9283 4173 9284
rect 3576 8672 3584 8736
rect 3648 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3896 8736
rect 3576 7648 3896 8672
rect 3576 7584 3584 7648
rect 3648 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3896 7648
rect 3576 6560 3896 7584
rect 4110 6629 4170 9283
rect 4107 6628 4173 6629
rect 4107 6564 4108 6628
rect 4172 6564 4173 6628
rect 4107 6563 4173 6564
rect 3576 6496 3584 6560
rect 3648 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3896 6560
rect 3187 6356 3253 6357
rect 3187 6292 3188 6356
rect 3252 6292 3253 6356
rect 3187 6291 3253 6292
rect 3576 5472 3896 6496
rect 3576 5408 3584 5472
rect 3648 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3896 5472
rect 3576 4384 3896 5408
rect 4662 4997 4722 13635
rect 6208 13632 6528 14656
rect 6208 13568 6216 13632
rect 6280 13568 6296 13632
rect 6360 13568 6376 13632
rect 6440 13568 6456 13632
rect 6520 13568 6528 13632
rect 6208 12544 6528 13568
rect 8840 14176 9160 14736
rect 8840 14112 8848 14176
rect 8912 14112 8928 14176
rect 8992 14112 9008 14176
rect 9072 14112 9088 14176
rect 9152 14112 9160 14176
rect 8840 13088 9160 14112
rect 8840 13024 8848 13088
rect 8912 13024 8928 13088
rect 8992 13024 9008 13088
rect 9072 13024 9088 13088
rect 9152 13024 9160 13088
rect 7419 12884 7485 12885
rect 7419 12820 7420 12884
rect 7484 12820 7485 12884
rect 7419 12819 7485 12820
rect 6208 12480 6216 12544
rect 6280 12480 6296 12544
rect 6360 12480 6376 12544
rect 6440 12480 6456 12544
rect 6520 12480 6528 12544
rect 6208 11456 6528 12480
rect 6208 11392 6216 11456
rect 6280 11392 6296 11456
rect 6360 11392 6376 11456
rect 6440 11392 6456 11456
rect 6520 11392 6528 11456
rect 6208 10368 6528 11392
rect 6208 10304 6216 10368
rect 6280 10304 6296 10368
rect 6360 10304 6376 10368
rect 6440 10304 6456 10368
rect 6520 10304 6528 10368
rect 5579 9348 5645 9349
rect 5579 9284 5580 9348
rect 5644 9284 5645 9348
rect 5579 9283 5645 9284
rect 5582 7173 5642 9283
rect 6208 9280 6528 10304
rect 6208 9216 6216 9280
rect 6280 9216 6296 9280
rect 6360 9216 6376 9280
rect 6440 9216 6456 9280
rect 6520 9216 6528 9280
rect 6208 8192 6528 9216
rect 6208 8128 6216 8192
rect 6280 8128 6296 8192
rect 6360 8128 6376 8192
rect 6440 8128 6456 8192
rect 6520 8128 6528 8192
rect 5579 7172 5645 7173
rect 5579 7108 5580 7172
rect 5644 7108 5645 7172
rect 5579 7107 5645 7108
rect 4659 4996 4725 4997
rect 4659 4932 4660 4996
rect 4724 4932 4725 4996
rect 4659 4931 4725 4932
rect 5582 4861 5642 7107
rect 6208 7104 6528 8128
rect 6683 7852 6749 7853
rect 6683 7788 6684 7852
rect 6748 7788 6749 7852
rect 6683 7787 6749 7788
rect 6208 7040 6216 7104
rect 6280 7040 6296 7104
rect 6360 7040 6376 7104
rect 6440 7040 6456 7104
rect 6520 7040 6528 7104
rect 6208 6016 6528 7040
rect 6208 5952 6216 6016
rect 6280 5952 6296 6016
rect 6360 5952 6376 6016
rect 6440 5952 6456 6016
rect 6520 5952 6528 6016
rect 6208 4928 6528 5952
rect 6686 4997 6746 7787
rect 6683 4996 6749 4997
rect 6683 4932 6684 4996
rect 6748 4932 6749 4996
rect 6683 4931 6749 4932
rect 6208 4864 6216 4928
rect 6280 4864 6296 4928
rect 6360 4864 6376 4928
rect 6440 4864 6456 4928
rect 6520 4864 6528 4928
rect 5579 4860 5645 4861
rect 5579 4796 5580 4860
rect 5644 4796 5645 4860
rect 5579 4795 5645 4796
rect 3576 4320 3584 4384
rect 3648 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3896 4384
rect 3576 3296 3896 4320
rect 3576 3232 3584 3296
rect 3648 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3896 3296
rect 3576 2208 3896 3232
rect 3576 2144 3584 2208
rect 3648 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3896 2208
rect 3576 2128 3896 2144
rect 6208 3840 6528 4864
rect 6208 3776 6216 3840
rect 6280 3776 6296 3840
rect 6360 3776 6376 3840
rect 6440 3776 6456 3840
rect 6520 3776 6528 3840
rect 6208 2752 6528 3776
rect 6208 2688 6216 2752
rect 6280 2688 6296 2752
rect 6360 2688 6376 2752
rect 6440 2688 6456 2752
rect 6520 2688 6528 2752
rect 6208 2128 6528 2688
rect 7422 2685 7482 12819
rect 8840 12000 9160 13024
rect 8840 11936 8848 12000
rect 8912 11936 8928 12000
rect 8992 11936 9008 12000
rect 9072 11936 9088 12000
rect 9152 11936 9160 12000
rect 8840 10912 9160 11936
rect 8840 10848 8848 10912
rect 8912 10848 8928 10912
rect 8992 10848 9008 10912
rect 9072 10848 9088 10912
rect 9152 10848 9160 10912
rect 8840 9824 9160 10848
rect 11472 14720 11792 14736
rect 11472 14656 11480 14720
rect 11544 14656 11560 14720
rect 11624 14656 11640 14720
rect 11704 14656 11720 14720
rect 11784 14656 11792 14720
rect 11472 13632 11792 14656
rect 11472 13568 11480 13632
rect 11544 13568 11560 13632
rect 11624 13568 11640 13632
rect 11704 13568 11720 13632
rect 11784 13568 11792 13632
rect 11472 12544 11792 13568
rect 11472 12480 11480 12544
rect 11544 12480 11560 12544
rect 11624 12480 11640 12544
rect 11704 12480 11720 12544
rect 11784 12480 11792 12544
rect 11472 11456 11792 12480
rect 11472 11392 11480 11456
rect 11544 11392 11560 11456
rect 11624 11392 11640 11456
rect 11704 11392 11720 11456
rect 11784 11392 11792 11456
rect 9259 10436 9325 10437
rect 9259 10372 9260 10436
rect 9324 10372 9325 10436
rect 9259 10371 9325 10372
rect 8840 9760 8848 9824
rect 8912 9760 8928 9824
rect 8992 9760 9008 9824
rect 9072 9760 9088 9824
rect 9152 9760 9160 9824
rect 8840 8736 9160 9760
rect 8840 8672 8848 8736
rect 8912 8672 8928 8736
rect 8992 8672 9008 8736
rect 9072 8672 9088 8736
rect 9152 8672 9160 8736
rect 8707 8124 8773 8125
rect 8707 8060 8708 8124
rect 8772 8060 8773 8124
rect 8707 8059 8773 8060
rect 8710 2821 8770 8059
rect 8840 7648 9160 8672
rect 8840 7584 8848 7648
rect 8912 7584 8928 7648
rect 8992 7584 9008 7648
rect 9072 7584 9088 7648
rect 9152 7584 9160 7648
rect 8840 6560 9160 7584
rect 8840 6496 8848 6560
rect 8912 6496 8928 6560
rect 8992 6496 9008 6560
rect 9072 6496 9088 6560
rect 9152 6496 9160 6560
rect 8840 5472 9160 6496
rect 9262 6085 9322 10371
rect 11472 10368 11792 11392
rect 11472 10304 11480 10368
rect 11544 10304 11560 10368
rect 11624 10304 11640 10368
rect 11704 10304 11720 10368
rect 11784 10304 11792 10368
rect 9443 9620 9509 9621
rect 9443 9556 9444 9620
rect 9508 9556 9509 9620
rect 9443 9555 9509 9556
rect 9446 8397 9506 9555
rect 11472 9280 11792 10304
rect 14104 14176 14424 14736
rect 14104 14112 14112 14176
rect 14176 14112 14192 14176
rect 14256 14112 14272 14176
rect 14336 14112 14352 14176
rect 14416 14112 14424 14176
rect 14104 13088 14424 14112
rect 14104 13024 14112 13088
rect 14176 13024 14192 13088
rect 14256 13024 14272 13088
rect 14336 13024 14352 13088
rect 14416 13024 14424 13088
rect 14104 12000 14424 13024
rect 14104 11936 14112 12000
rect 14176 11936 14192 12000
rect 14256 11936 14272 12000
rect 14336 11936 14352 12000
rect 14416 11936 14424 12000
rect 14104 10912 14424 11936
rect 14104 10848 14112 10912
rect 14176 10848 14192 10912
rect 14256 10848 14272 10912
rect 14336 10848 14352 10912
rect 14416 10848 14424 10912
rect 14104 9824 14424 10848
rect 14595 10436 14661 10437
rect 14595 10372 14596 10436
rect 14660 10372 14661 10436
rect 14595 10371 14661 10372
rect 14104 9760 14112 9824
rect 14176 9760 14192 9824
rect 14256 9760 14272 9824
rect 14336 9760 14352 9824
rect 14416 9760 14424 9824
rect 13859 9620 13925 9621
rect 13859 9556 13860 9620
rect 13924 9556 13925 9620
rect 13859 9555 13925 9556
rect 11472 9216 11480 9280
rect 11544 9216 11560 9280
rect 11624 9216 11640 9280
rect 11704 9216 11720 9280
rect 11784 9216 11792 9280
rect 9443 8396 9509 8397
rect 9443 8332 9444 8396
rect 9508 8332 9509 8396
rect 9443 8331 9509 8332
rect 9259 6084 9325 6085
rect 9259 6020 9260 6084
rect 9324 6020 9325 6084
rect 9259 6019 9325 6020
rect 8840 5408 8848 5472
rect 8912 5408 8928 5472
rect 8992 5408 9008 5472
rect 9072 5408 9088 5472
rect 9152 5408 9160 5472
rect 8840 4384 9160 5408
rect 8840 4320 8848 4384
rect 8912 4320 8928 4384
rect 8992 4320 9008 4384
rect 9072 4320 9088 4384
rect 9152 4320 9160 4384
rect 8840 3296 9160 4320
rect 8840 3232 8848 3296
rect 8912 3232 8928 3296
rect 8992 3232 9008 3296
rect 9072 3232 9088 3296
rect 9152 3232 9160 3296
rect 8707 2820 8773 2821
rect 8707 2756 8708 2820
rect 8772 2756 8773 2820
rect 8707 2755 8773 2756
rect 7419 2684 7485 2685
rect 7419 2620 7420 2684
rect 7484 2620 7485 2684
rect 7419 2619 7485 2620
rect 8840 2208 9160 3232
rect 9446 2957 9506 8331
rect 11472 8192 11792 9216
rect 13862 8533 13922 9555
rect 14104 8736 14424 9760
rect 14598 9757 14658 10371
rect 14595 9756 14661 9757
rect 14595 9692 14596 9756
rect 14660 9692 14661 9756
rect 14595 9691 14661 9692
rect 14104 8672 14112 8736
rect 14176 8672 14192 8736
rect 14256 8672 14272 8736
rect 14336 8672 14352 8736
rect 14416 8672 14424 8736
rect 13859 8532 13925 8533
rect 13859 8468 13860 8532
rect 13924 8468 13925 8532
rect 13859 8467 13925 8468
rect 11472 8128 11480 8192
rect 11544 8128 11560 8192
rect 11624 8128 11640 8192
rect 11704 8128 11720 8192
rect 11784 8128 11792 8192
rect 11472 7104 11792 8128
rect 11472 7040 11480 7104
rect 11544 7040 11560 7104
rect 11624 7040 11640 7104
rect 11704 7040 11720 7104
rect 11784 7040 11792 7104
rect 11472 6016 11792 7040
rect 11472 5952 11480 6016
rect 11544 5952 11560 6016
rect 11624 5952 11640 6016
rect 11704 5952 11720 6016
rect 11784 5952 11792 6016
rect 11472 4928 11792 5952
rect 13862 5949 13922 8467
rect 14104 7648 14424 8672
rect 14104 7584 14112 7648
rect 14176 7584 14192 7648
rect 14256 7584 14272 7648
rect 14336 7584 14352 7648
rect 14416 7584 14424 7648
rect 14104 6560 14424 7584
rect 14104 6496 14112 6560
rect 14176 6496 14192 6560
rect 14256 6496 14272 6560
rect 14336 6496 14352 6560
rect 14416 6496 14424 6560
rect 13859 5948 13925 5949
rect 13859 5884 13860 5948
rect 13924 5884 13925 5948
rect 13859 5883 13925 5884
rect 11472 4864 11480 4928
rect 11544 4864 11560 4928
rect 11624 4864 11640 4928
rect 11704 4864 11720 4928
rect 11784 4864 11792 4928
rect 11472 3840 11792 4864
rect 11472 3776 11480 3840
rect 11544 3776 11560 3840
rect 11624 3776 11640 3840
rect 11704 3776 11720 3840
rect 11784 3776 11792 3840
rect 9443 2956 9509 2957
rect 9443 2892 9444 2956
rect 9508 2892 9509 2956
rect 9443 2891 9509 2892
rect 8840 2144 8848 2208
rect 8912 2144 8928 2208
rect 8992 2144 9008 2208
rect 9072 2144 9088 2208
rect 9152 2144 9160 2208
rect 8840 2128 9160 2144
rect 11472 2752 11792 3776
rect 11472 2688 11480 2752
rect 11544 2688 11560 2752
rect 11624 2688 11640 2752
rect 11704 2688 11720 2752
rect 11784 2688 11792 2752
rect 11472 2128 11792 2688
rect 14104 5472 14424 6496
rect 14104 5408 14112 5472
rect 14176 5408 14192 5472
rect 14256 5408 14272 5472
rect 14336 5408 14352 5472
rect 14416 5408 14424 5472
rect 14104 4384 14424 5408
rect 14104 4320 14112 4384
rect 14176 4320 14192 4384
rect 14256 4320 14272 4384
rect 14336 4320 14352 4384
rect 14416 4320 14424 4384
rect 14104 3296 14424 4320
rect 14104 3232 14112 3296
rect 14176 3232 14192 3296
rect 14256 3232 14272 3296
rect 14336 3232 14352 3296
rect 14416 3232 14424 3296
rect 14104 2208 14424 3232
rect 14104 2144 14112 2208
rect 14176 2144 14192 2208
rect 14256 2144 14272 2208
rect 14336 2144 14352 2208
rect 14416 2144 14424 2208
rect 14104 2128 14424 2144
use sky130_fd_sc_hd__fill_2  FILLER_0_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_19
timestamp 1605641404
transform 1 0 2852 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1605641404
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2208 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3128 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4140 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4232 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 1605641404
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_31
timestamp 1605641404
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1605641404
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51
timestamp 1605641404
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4968 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1605641404
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1605641404
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 6072 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1605641404
transform 1 0 6164 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1605641404
transform 1 0 8004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7084 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6992 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8280 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73
timestamp 1605641404
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79
timestamp 1605641404
transform 1 0 8372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_74 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10304 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9292 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 10396 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1605641404
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98
timestamp 1605641404
transform 1 0 10120 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1605641404
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_98
timestamp 1605641404
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11408 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1605641404
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1605641404
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1605641404
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14076 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13984 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_131
timestamp 1605641404
transform 1 0 13156 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1605641404
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1605641404
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_150
timestamp 1605641404
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_146
timestamp 1605641404
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15088 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp 1605641404
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1605641404
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1605641404
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1605641404
transform 1 0 16008 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15824 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 16836 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 16836 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2760 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1748 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_16
timestamp 1605641404
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 4508 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1605641404
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 5520 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6532 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_46
timestamp 1605641404
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1605641404
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_68
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_79
timestamp 1605641404
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10580 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1605641404
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1605641404
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1605641404
transform 1 0 11592 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12144 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1605641404
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1605641404
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13156 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1605641404
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_147
timestamp 1605641404
transform 1 0 14628 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1605641404
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_167
timestamp 1605641404
transform 1 0 16468 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2760 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1748 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_16
timestamp 1605641404
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3772 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4784 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_38
timestamp 1605641404
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 5704 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_46
timestamp 1605641404
transform 1 0 5336 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7176 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8188 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1605641404
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9200 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1605641404
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_104
timestamp 1605641404
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1605641404
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10856 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1605641404
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1605641404
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13432 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1605641404
transform 1 0 14444 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1605641404
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1605641404
transform 1 0 15456 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1605641404
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1605641404
transform 1 0 16284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 16836 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1656 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1605641404
transform 1 0 3312 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1605641404
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1605641404
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6532 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 5796 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_48
timestamp 1605641404
transform 1 0 5520 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 1605641404
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8556 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8188 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1605641404
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_80
timestamp 1605641404
transform 1 0 8464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1605641404
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 11684 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 11316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_109
timestamp 1605641404
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_114
timestamp 1605641404
transform 1 0 11592 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_131
timestamp 1605641404
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1605641404
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1605641404
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1605641404
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_163
timestamp 1605641404
transform 1 0 16100 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 16836 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 1605641404
transform 1 0 16468 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 2668 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1656 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1605641404
transform 1 0 3680 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4232 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 1605641404
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_32
timestamp 1605641404
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 5888 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_50
timestamp 1605641404
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_58
timestamp 1605641404
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7820 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1605641404
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10304 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9476 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1605641404
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_97
timestamp 1605641404
transform 1 0 10028 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_116
timestamp 1605641404
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1605641404
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14168 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13156 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1605641404
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1605641404
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1605641404
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1605641404
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1605641404
transform 1 0 16192 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 16836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1605641404
transform 1 0 1564 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1472 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2300 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1605641404
transform 1 0 1932 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_20
timestamp 1605641404
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1605641404
transform 1 0 3128 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3772 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 4416 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1605641404
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_26
timestamp 1605641404
transform 1 0 3496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5428 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5428 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1605641404
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1605641404
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_56
timestamp 1605641404
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1605641404
transform 1 0 8556 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1605641404
transform 1 0 7084 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 6900 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8648 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1605641404
transform 1 0 6900 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_69
timestamp 1605641404
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_80
timestamp 1605641404
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_79
timestamp 1605641404
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1605641404
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1605641404
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9108 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1605641404
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1605641404
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1605641404
transform 1 0 10028 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11592 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12604 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1605641404
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1605641404
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1605641404
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1605641404
transform 1 0 13248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14260 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13708 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_130
timestamp 1605641404
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_135
timestamp 1605641404
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp 1605641404
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1605641404
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15364 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1605641404
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1605641404
transform 1 0 16284 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1605641404
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1605641404
transform 1 0 16192 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1605641404
transform 1 0 15916 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 16836 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 1932 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2944 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1605641404
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_18
timestamp 1605641404
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1605641404
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5336 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_44
timestamp 1605641404
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp 1605641404
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6992 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 8648 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_80
timestamp 1605641404
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1605641404
transform 1 0 9016 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10120 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1605641404
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1605641404
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_96
timestamp 1605641404
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_107
timestamp 1605641404
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_118
timestamp 1605641404
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1605641404
transform 1 0 13248 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13800 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_136
timestamp 1605641404
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_147
timestamp 1605641404
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1605641404
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 16836 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1605641404
transform 1 0 16468 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1605641404
transform 1 0 1564 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp 1605641404
transform 1 0 1932 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 3220 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1605641404
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_39
timestamp 1605641404
transform 1 0 4692 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1605641404
transform 1 0 6072 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5060 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_52
timestamp 1605641404
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1605641404
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1605641404
transform 1 0 7728 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1605641404
transform 1 0 8096 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8648 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_71
timestamp 1605641404
transform 1 0 7636 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_80
timestamp 1605641404
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10304 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_98
timestamp 1605641404
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1605641404
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1605641404
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1605641404
transform 1 0 13800 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14352 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_132
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_142
timestamp 1605641404
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1605641404
transform 1 0 16008 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_160
timestamp 1605641404
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1605641404
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 16836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1605641404
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1605641404
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1605641404
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5704 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 6716 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1605641404
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1605641404
transform 1 0 6532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1605641404
transform 1 0 7820 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1605641404
transform 1 0 8648 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_70
timestamp 1605641404
transform 1 0 7544 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1605641404
transform 1 0 9844 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10396 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1605641404
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_99
timestamp 1605641404
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 1605641404
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13064 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14076 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1605641404
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_139
timestamp 1605641404
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1605641404
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1605641404
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_167
timestamp 1605641404
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1605641404
transform 1 0 1564 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1605641404
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_20
timestamp 1605641404
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1605641404
transform 1 0 4784 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3128 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_38
timestamp 1605641404
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1605641404
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 5244 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp 1605641404
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1605641404
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8188 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_11_71
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10028 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1605641404
transform 1 0 11500 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12788 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1605641404
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1605641404
transform 1 0 15456 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1605641404
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1605641404
transform 1 0 16284 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 16836 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1840 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 1564 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1605641404
transform 1 0 3496 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_24
timestamp 1605641404
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1605641404
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5888 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1605641404
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 7912 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 7544 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp 1605641404
transform 1 0 7820 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10672 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1605641404
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1605641404
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12328 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1605641404
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1605641404
transform 1 0 13984 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1605641404
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1605641404
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1605641404
transform 1 0 16100 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 16836 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1605641404
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1605641404
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1605641404
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1605641404
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1605641404
transform 1 0 4048 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4324 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1605641404
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_36
timestamp 1605641404
transform 1 0 4416 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1605641404
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1605641404
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4968 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1605641404
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1605641404
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_59
timestamp 1605641404
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8556 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_78
timestamp 1605641404
transform 1 0 8280 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_78
timestamp 1605641404
transform 1 0 8280 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9568 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10028 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1605641404
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1605641404
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11040 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_108
timestamp 1605641404
transform 1 0 11040 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1605641404
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_106
timestamp 1605641404
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1605641404
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12880 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13064 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14076 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1605641404
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_144
timestamp 1605641404
transform 1 0 14352 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_128
timestamp 1605641404
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_139
timestamp 1605641404
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1605641404
transform 1 0 14720 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15824 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_157
timestamp 1605641404
transform 1 0 15548 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1605641404
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1605641404
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_163
timestamp 1605641404
transform 1 0 16100 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1605641404
transform 1 0 16468 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1605641404
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1605641404
transform 1 0 4048 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1605641404
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_36
timestamp 1605641404
transform 1 0 4416 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4968 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1605641404
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1605641404
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7820 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1605641404
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1605641404
transform 1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 9568 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_89
timestamp 1605641404
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1605641404
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1605641404
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1605641404
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1605641404
transform 1 0 14352 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1605641404
transform 1 0 13892 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1605641404
transform 1 0 14260 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14904 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1605641404
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1605641404
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1605641404
transform 1 0 1564 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2116 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1605641404
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4140 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1605641404
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5152 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6808 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_42
timestamp 1605641404
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1605641404
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1605641404
transform 1 0 7820 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1605641404
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_76
timestamp 1605641404
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9936 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1605641404
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1605641404
transform 1 0 11684 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_112
timestamp 1605641404
transform 1 0 11408 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_119
timestamp 1605641404
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13524 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 13248 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1605641404
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_144
timestamp 1605641404
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1605641404
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15364 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1605641404
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1605641404
transform 1 0 16192 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2484 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1472 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_13
timestamp 1605641404
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4140 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1605641404
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 5336 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_42
timestamp 1605641404
transform 1 0 4968 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_55
timestamp 1605641404
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 6992 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8648 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1605641404
transform 1 0 8464 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10304 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_98
timestamp 1605641404
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1605641404
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1605641404
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14444 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1605641404
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1605641404
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1605641404
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1605641404
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1605641404
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 16836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2576 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_14
timestamp 1605641404
transform 1 0 2392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_25
timestamp 1605641404
transform 1 0 3404 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1605641404
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6532 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_48
timestamp 1605641404
transform 1 0 5520 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_54
timestamp 1605641404
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_58
timestamp 1605641404
transform 1 0 6440 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_18_75
timestamp 1605641404
transform 1 0 8004 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10488 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1605641404
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_96
timestamp 1605641404
transform 1 0 9936 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_118
timestamp 1605641404
transform 1 0 11960 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 13524 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_130
timestamp 1605641404
transform 1 0 13064 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp 1605641404
transform 1 0 13432 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1605641404
transform 1 0 15456 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1605641404
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_165
timestamp 1605641404
transform 1 0 16284 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 16836 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2760 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1605641404
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1605641404
transform 1 0 2944 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp 1605641404
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1605641404
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1605641404
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 5428 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_49 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5612 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1605641404
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_56
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6992 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8188 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1605641404
transform 1 0 7912 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1605641404
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_83
timestamp 1605641404
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1605641404
transform 1 0 7820 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10028 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1605641404
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_86
timestamp 1605641404
transform 1 0 9016 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1605641404
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1605641404
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12328 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1605641404
transform 1 0 11316 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1605641404
transform 1 0 11500 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1605641404
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1605641404
transform 1 0 11224 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1605641404
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13340 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 14076 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1605641404
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1605641404
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1605641404
transform 1 0 15916 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15548 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_157
timestamp 1605641404
transform 1 0 15548 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1605641404
transform 1 0 16284 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1605641404
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1605641404
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 16836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2208 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_11
timestamp 1605641404
transform 1 0 2116 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 4692 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_21
timestamp 1605641404
transform 1 0 3036 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_33
timestamp 1605641404
transform 1 0 4140 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1605641404
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7176 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8648 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_75
timestamp 1605641404
transform 1 0 8004 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_81
timestamp 1605641404
transform 1 0 8556 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10120 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_91
timestamp 1605641404
transform 1 0 9476 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 1605641404
transform 1 0 10028 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_107
timestamp 1605641404
transform 1 0 10948 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1605641404
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1605641404
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1605641404
transform 1 0 16100 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1605641404
transform 1 0 15088 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_151
timestamp 1605641404
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1605641404
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1605641404
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 16836 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_50
timestamp 1605641404
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1605641404
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1605641404
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_22_63
timestamp 1605641404
transform 1 0 6900 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1605641404
transform 1 0 7452 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1605641404
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_90
timestamp 1605641404
transform 1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1605641404
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1605641404
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1605641404
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1605641404
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1605641404
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1605641404
transform 1 0 15916 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1605641404
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1605641404
transform 1 0 15456 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_160
timestamp 1605641404
transform 1 0 15824 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1605641404
transform 1 0 16284 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 16836 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal2 s 3238 0 3294 480 6 bottom_grid_pin_0_
port 0 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 bottom_grid_pin_10_
port 1 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 bottom_grid_pin_11_
port 2 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 bottom_grid_pin_12_
port 3 nsew default tristate
rlabel metal2 s 15658 0 15714 480 6 bottom_grid_pin_13_
port 4 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 bottom_grid_pin_14_
port 5 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 bottom_grid_pin_15_
port 6 nsew default tristate
rlabel metal2 s 4250 0 4306 480 6 bottom_grid_pin_1_
port 7 nsew default tristate
rlabel metal2 s 5170 0 5226 480 6 bottom_grid_pin_2_
port 8 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 bottom_grid_pin_3_
port 9 nsew default tristate
rlabel metal2 s 7102 0 7158 480 6 bottom_grid_pin_4_
port 10 nsew default tristate
rlabel metal2 s 8022 0 8078 480 6 bottom_grid_pin_5_
port 11 nsew default tristate
rlabel metal2 s 8942 0 8998 480 6 bottom_grid_pin_6_
port 12 nsew default tristate
rlabel metal2 s 9954 0 10010 480 6 bottom_grid_pin_7_
port 13 nsew default tristate
rlabel metal2 s 10874 0 10930 480 6 bottom_grid_pin_8_
port 14 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 bottom_grid_pin_9_
port 15 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 ccff_head
port 16 nsew default input
rlabel metal2 s 2318 0 2374 480 6 ccff_tail
port 17 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[0]
port 18 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[10]
port 19 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[11]
port 20 nsew default input
rlabel metal3 s 0 13744 480 13864 6 chanx_left_in[12]
port 21 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chanx_left_in[13]
port 22 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[14]
port 23 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chanx_left_in[15]
port 24 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[16]
port 25 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[17]
port 26 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chanx_left_in[18]
port 27 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[19]
port 28 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[1]
port 29 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[2]
port 30 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[3]
port 31 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[4]
port 32 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[5]
port 33 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[6]
port 34 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[7]
port 35 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[8]
port 36 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[9]
port 37 nsew default input
rlabel metal3 s 0 144 480 264 6 chanx_left_out[0]
port 38 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[10]
port 39 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[11]
port 40 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 chanx_left_out[12]
port 41 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[13]
port 42 nsew default tristate
rlabel metal3 s 0 5992 480 6112 6 chanx_left_out[14]
port 43 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 chanx_left_out[15]
port 44 nsew default tristate
rlabel metal3 s 0 6944 480 7064 6 chanx_left_out[16]
port 45 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[17]
port 46 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 chanx_left_out[18]
port 47 nsew default tristate
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[19]
port 48 nsew default tristate
rlabel metal3 s 0 552 480 672 6 chanx_left_out[1]
port 49 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[2]
port 50 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[3]
port 51 nsew default tristate
rlabel metal3 s 0 1776 480 1896 6 chanx_left_out[4]
port 52 nsew default tristate
rlabel metal3 s 0 2184 480 2304 6 chanx_left_out[5]
port 53 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[6]
port 54 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[7]
port 55 nsew default tristate
rlabel metal3 s 0 3544 480 3664 6 chanx_left_out[8]
port 56 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_out[9]
port 57 nsew default tristate
rlabel metal3 s 17520 8576 18000 8696 6 chanx_right_in[0]
port 58 nsew default input
rlabel metal3 s 17520 12792 18000 12912 6 chanx_right_in[10]
port 59 nsew default input
rlabel metal3 s 17520 13200 18000 13320 6 chanx_right_in[11]
port 60 nsew default input
rlabel metal3 s 17520 13744 18000 13864 6 chanx_right_in[12]
port 61 nsew default input
rlabel metal3 s 17520 14152 18000 14272 6 chanx_right_in[13]
port 62 nsew default input
rlabel metal3 s 17520 14560 18000 14680 6 chanx_right_in[14]
port 63 nsew default input
rlabel metal3 s 17520 14968 18000 15088 6 chanx_right_in[15]
port 64 nsew default input
rlabel metal3 s 17520 15376 18000 15496 6 chanx_right_in[16]
port 65 nsew default input
rlabel metal3 s 17520 15784 18000 15904 6 chanx_right_in[17]
port 66 nsew default input
rlabel metal3 s 17520 16192 18000 16312 6 chanx_right_in[18]
port 67 nsew default input
rlabel metal3 s 17520 16600 18000 16720 6 chanx_right_in[19]
port 68 nsew default input
rlabel metal3 s 17520 8984 18000 9104 6 chanx_right_in[1]
port 69 nsew default input
rlabel metal3 s 17520 9392 18000 9512 6 chanx_right_in[2]
port 70 nsew default input
rlabel metal3 s 17520 9800 18000 9920 6 chanx_right_in[3]
port 71 nsew default input
rlabel metal3 s 17520 10344 18000 10464 6 chanx_right_in[4]
port 72 nsew default input
rlabel metal3 s 17520 10752 18000 10872 6 chanx_right_in[5]
port 73 nsew default input
rlabel metal3 s 17520 11160 18000 11280 6 chanx_right_in[6]
port 74 nsew default input
rlabel metal3 s 17520 11568 18000 11688 6 chanx_right_in[7]
port 75 nsew default input
rlabel metal3 s 17520 11976 18000 12096 6 chanx_right_in[8]
port 76 nsew default input
rlabel metal3 s 17520 12384 18000 12504 6 chanx_right_in[9]
port 77 nsew default input
rlabel metal3 s 17520 144 18000 264 6 chanx_right_out[0]
port 78 nsew default tristate
rlabel metal3 s 17520 4360 18000 4480 6 chanx_right_out[10]
port 79 nsew default tristate
rlabel metal3 s 17520 4768 18000 4888 6 chanx_right_out[11]
port 80 nsew default tristate
rlabel metal3 s 17520 5176 18000 5296 6 chanx_right_out[12]
port 81 nsew default tristate
rlabel metal3 s 17520 5584 18000 5704 6 chanx_right_out[13]
port 82 nsew default tristate
rlabel metal3 s 17520 5992 18000 6112 6 chanx_right_out[14]
port 83 nsew default tristate
rlabel metal3 s 17520 6400 18000 6520 6 chanx_right_out[15]
port 84 nsew default tristate
rlabel metal3 s 17520 6944 18000 7064 6 chanx_right_out[16]
port 85 nsew default tristate
rlabel metal3 s 17520 7352 18000 7472 6 chanx_right_out[17]
port 86 nsew default tristate
rlabel metal3 s 17520 7760 18000 7880 6 chanx_right_out[18]
port 87 nsew default tristate
rlabel metal3 s 17520 8168 18000 8288 6 chanx_right_out[19]
port 88 nsew default tristate
rlabel metal3 s 17520 552 18000 672 6 chanx_right_out[1]
port 89 nsew default tristate
rlabel metal3 s 17520 960 18000 1080 6 chanx_right_out[2]
port 90 nsew default tristate
rlabel metal3 s 17520 1368 18000 1488 6 chanx_right_out[3]
port 91 nsew default tristate
rlabel metal3 s 17520 1776 18000 1896 6 chanx_right_out[4]
port 92 nsew default tristate
rlabel metal3 s 17520 2184 18000 2304 6 chanx_right_out[5]
port 93 nsew default tristate
rlabel metal3 s 17520 2592 18000 2712 6 chanx_right_out[6]
port 94 nsew default tristate
rlabel metal3 s 17520 3000 18000 3120 6 chanx_right_out[7]
port 95 nsew default tristate
rlabel metal3 s 17520 3544 18000 3664 6 chanx_right_out[8]
port 96 nsew default tristate
rlabel metal3 s 17520 3952 18000 4072 6 chanx_right_out[9]
port 97 nsew default tristate
rlabel metal2 s 478 0 534 480 6 prog_clk
port 98 nsew default input
rlabel metal4 s 3576 2128 3896 14736 6 VPWR
port 99 nsew default input
rlabel metal4 s 6208 2128 6528 14736 6 VGND
port 100 nsew default input
<< properties >>
string FIXED_BBOX 0 0 18000 16720
<< end >>
